module fake_jpeg_24248_n_343 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_343);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_343;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx8_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_21),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_39),
.B(n_23),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx4_ASAP7_75t_SL g43 ( 
.A(n_17),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_47),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx6_ASAP7_75t_SL g47 ( 
.A(n_18),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx6_ASAP7_75t_SL g62 ( 
.A(n_48),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_20),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_50),
.B(n_51),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_40),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_54),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_20),
.Y(n_56)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

NAND3xp33_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_11),
.C(n_15),
.Y(n_59)
);

A2O1A1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_59),
.A2(n_70),
.B(n_36),
.C(n_17),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_48),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_60),
.Y(n_88)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_61),
.B(n_67),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_20),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_63),
.B(n_71),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_38),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_64),
.Y(n_89)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_69),
.B(n_34),
.Y(n_93)
);

NAND2xp33_ASAP7_75t_SL g70 ( 
.A(n_47),
.B(n_34),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_44),
.B(n_23),
.Y(n_71)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_72),
.Y(n_117)
);

INVx5_ASAP7_75t_SL g73 ( 
.A(n_58),
.Y(n_73)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_73),
.Y(n_105)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_75),
.B(n_77),
.Y(n_110)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_51),
.B(n_22),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_78),
.B(n_99),
.Y(n_106)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_79),
.Y(n_127)
);

OA22x2_ASAP7_75t_L g80 ( 
.A1(n_70),
.A2(n_28),
.B1(n_33),
.B2(n_46),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_80),
.A2(n_85),
.B1(n_24),
.B2(n_63),
.Y(n_107)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_81),
.B(n_83),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_54),
.B(n_28),
.C(n_33),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_82),
.B(n_96),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_84),
.B(n_90),
.Y(n_112)
);

O2A1O1Ixp33_ASAP7_75t_L g85 ( 
.A1(n_59),
.A2(n_28),
.B(n_32),
.C(n_29),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_68),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_91),
.B(n_92),
.Y(n_115)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_94),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_68),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_95),
.B(n_97),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_60),
.B(n_22),
.C(n_26),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_56),
.Y(n_98)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_98),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_50),
.B(n_22),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_53),
.Y(n_100)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_100),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_64),
.B(n_0),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_102),
.B(n_71),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_66),
.A2(n_19),
.B1(n_34),
.B2(n_32),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_103),
.A2(n_35),
.B1(n_24),
.B2(n_19),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_104),
.A2(n_109),
.B1(n_111),
.B2(n_120),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_107),
.A2(n_132),
.B1(n_65),
.B2(n_88),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_108),
.B(n_22),
.Y(n_157)
);

OA22x2_ASAP7_75t_L g109 ( 
.A1(n_80),
.A2(n_66),
.B1(n_53),
.B2(n_62),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_94),
.A2(n_66),
.B1(n_67),
.B2(n_69),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_101),
.B(n_29),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_118),
.B(n_126),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_83),
.A2(n_24),
.B1(n_35),
.B2(n_19),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_119),
.A2(n_19),
.B1(n_65),
.B2(n_35),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_80),
.A2(n_55),
.B1(n_57),
.B2(n_52),
.Y(n_120)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_76),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_123),
.B(n_125),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_80),
.A2(n_78),
.B1(n_90),
.B2(n_99),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_124),
.A2(n_62),
.B1(n_65),
.B2(n_61),
.Y(n_140)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_102),
.Y(n_126)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_102),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_129),
.B(n_130),
.Y(n_137)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_87),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_96),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_134),
.A2(n_146),
.B1(n_150),
.B2(n_152),
.Y(n_165)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_131),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_135),
.B(n_141),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_106),
.B(n_86),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_136),
.B(n_151),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_132),
.B(n_82),
.C(n_86),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_138),
.B(n_154),
.C(n_124),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_113),
.A2(n_62),
.B1(n_85),
.B2(n_74),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_139),
.A2(n_153),
.B(n_158),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_140),
.B(n_157),
.Y(n_167)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_117),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_110),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_142),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_126),
.A2(n_74),
.B(n_88),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_143),
.A2(n_159),
.B(n_161),
.Y(n_170)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_117),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_144),
.B(n_147),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_107),
.A2(n_55),
.B1(n_97),
.B2(n_100),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_127),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_131),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_148),
.A2(n_160),
.B1(n_105),
.B2(n_127),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_115),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_149),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_106),
.B(n_89),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_109),
.A2(n_52),
.B1(n_57),
.B2(n_89),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_120),
.A2(n_73),
.B(n_95),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_116),
.B(n_81),
.C(n_75),
.Y(n_154)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_121),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_156),
.B(n_162),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_129),
.A2(n_72),
.B1(n_23),
.B2(n_26),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_125),
.A2(n_21),
.B(n_31),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_109),
.A2(n_26),
.B1(n_91),
.B2(n_84),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_116),
.A2(n_21),
.B(n_31),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_121),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g163 ( 
.A(n_112),
.B(n_30),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_163),
.B(n_118),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_164),
.A2(n_191),
.B(n_194),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_145),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_166),
.B(n_176),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_169),
.B(n_173),
.C(n_190),
.Y(n_199)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_151),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_172),
.B(n_177),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_154),
.B(n_108),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_157),
.B(n_111),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_175),
.B(n_181),
.Y(n_212)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_141),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_136),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_179),
.B(n_184),
.Y(n_221)
);

XNOR2x2_ASAP7_75t_SL g181 ( 
.A(n_139),
.B(n_119),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_149),
.B(n_130),
.Y(n_182)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_182),
.Y(n_200)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_145),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_152),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_185),
.B(n_186),
.Y(n_223)
);

OR2x2_ASAP7_75t_L g186 ( 
.A(n_137),
.B(n_112),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_146),
.Y(n_187)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_187),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_138),
.B(n_109),
.Y(n_188)
);

OAI21xp33_ASAP7_75t_L g201 ( 
.A1(n_188),
.A2(n_193),
.B(n_148),
.Y(n_201)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_160),
.Y(n_189)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_189),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_161),
.B(n_128),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_153),
.Y(n_191)
);

OR2x2_ASAP7_75t_L g193 ( 
.A(n_142),
.B(n_109),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_143),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_156),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_195),
.Y(n_208)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_158),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_196),
.A2(n_134),
.B1(n_122),
.B2(n_104),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_162),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_197),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_201),
.A2(n_203),
.B(n_170),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_173),
.B(n_135),
.C(n_140),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_204),
.B(n_217),
.C(n_219),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_180),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_205),
.B(n_179),
.Y(n_245)
);

INVxp33_ASAP7_75t_SL g206 ( 
.A(n_176),
.Y(n_206)
);

A2O1A1Ixp33_ASAP7_75t_SL g243 ( 
.A1(n_206),
.A2(n_226),
.B(n_30),
.C(n_25),
.Y(n_243)
);

MAJx2_ASAP7_75t_L g207 ( 
.A(n_190),
.B(n_155),
.C(n_159),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_207),
.B(n_25),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_185),
.A2(n_133),
.B1(n_155),
.B2(n_122),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_209),
.A2(n_214),
.B1(n_215),
.B2(n_216),
.Y(n_242)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_174),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_211),
.B(n_225),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_169),
.B(n_133),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_213),
.B(n_167),
.Y(n_233)
);

AOI22x1_ASAP7_75t_L g214 ( 
.A1(n_181),
.A2(n_163),
.B1(n_105),
.B2(n_144),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_187),
.A2(n_114),
.B1(n_123),
.B2(n_163),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_191),
.A2(n_114),
.B1(n_147),
.B2(n_115),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_172),
.B(n_77),
.C(n_92),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_189),
.A2(n_31),
.B1(n_29),
.B2(n_32),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_218),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_177),
.B(n_79),
.C(n_22),
.Y(n_219)
);

BUFx24_ASAP7_75t_L g222 ( 
.A(n_192),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g229 ( 
.A(n_222),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_196),
.A2(n_30),
.B1(n_25),
.B2(n_17),
.Y(n_225)
);

AO22x2_ASAP7_75t_L g226 ( 
.A1(n_194),
.A2(n_17),
.B1(n_25),
.B2(n_2),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_202),
.A2(n_174),
.B1(n_188),
.B2(n_168),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_228),
.A2(n_230),
.B1(n_239),
.B2(n_240),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_211),
.A2(n_188),
.B1(n_168),
.B2(n_183),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_206),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_231),
.B(n_252),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_232),
.A2(n_237),
.B(n_247),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_233),
.B(n_235),
.C(n_250),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_199),
.B(n_175),
.C(n_167),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_200),
.B(n_182),
.Y(n_236)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_236),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_198),
.A2(n_171),
.B(n_170),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_224),
.A2(n_165),
.B1(n_178),
.B2(n_193),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_223),
.A2(n_214),
.B1(n_204),
.B2(n_220),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_221),
.B(n_184),
.Y(n_241)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_241),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_243),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_208),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_244),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_245),
.B(n_1),
.Y(n_274)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_222),
.Y(n_246)
);

INVx6_ASAP7_75t_L g260 ( 
.A(n_246),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_201),
.A2(n_186),
.B(n_165),
.Y(n_247)
);

HAxp5_ASAP7_75t_SL g248 ( 
.A(n_226),
.B(n_0),
.CON(n_248),
.SN(n_248)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_248),
.B(n_249),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_199),
.B(n_15),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_227),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_210),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_253),
.B(n_13),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_242),
.A2(n_226),
.B1(n_205),
.B2(n_217),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_257),
.A2(n_261),
.B1(n_262),
.B2(n_243),
.Y(n_288)
);

INVx13_ASAP7_75t_L g258 ( 
.A(n_229),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_258),
.B(n_9),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_238),
.A2(n_226),
.B1(n_213),
.B2(n_212),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_247),
.A2(n_212),
.B1(n_222),
.B2(n_207),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_235),
.B(n_219),
.C(n_36),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_264),
.B(n_265),
.C(n_266),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_233),
.B(n_36),
.C(n_2),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_234),
.B(n_1),
.C(n_3),
.Y(n_266)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_267),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_239),
.A2(n_230),
.B1(n_228),
.B2(n_240),
.Y(n_268)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_268),
.Y(n_292)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_270),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_249),
.B(n_13),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_272),
.B(n_250),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_229),
.B(n_246),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_273),
.B(n_274),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_259),
.B(n_251),
.Y(n_278)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_278),
.Y(n_298)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_279),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_256),
.B(n_234),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_281),
.B(n_282),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_256),
.B(n_232),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_264),
.B(n_241),
.C(n_236),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_283),
.B(n_266),
.C(n_265),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_261),
.B(n_237),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_284),
.B(n_275),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_257),
.A2(n_251),
.B1(n_243),
.B2(n_248),
.Y(n_285)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_285),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_269),
.B(n_243),
.Y(n_287)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_287),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_288),
.A2(n_263),
.B1(n_255),
.B2(n_254),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_289),
.B(n_291),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_275),
.A2(n_243),
.B(n_9),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_290),
.A2(n_274),
.B(n_277),
.Y(n_300)
);

FAx1_ASAP7_75t_SL g291 ( 
.A(n_262),
.B(n_3),
.CI(n_4),
.CON(n_291),
.SN(n_291)
);

AO221x1_ASAP7_75t_L g295 ( 
.A1(n_276),
.A2(n_260),
.B1(n_258),
.B2(n_255),
.C(n_254),
.Y(n_295)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_295),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_296),
.A2(n_306),
.B1(n_307),
.B2(n_288),
.Y(n_308)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_283),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_297),
.B(n_294),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_299),
.B(n_280),
.C(n_279),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_300),
.A2(n_12),
.B(n_6),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_301),
.B(n_302),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_282),
.B(n_263),
.Y(n_302)
);

MAJx2_ASAP7_75t_L g304 ( 
.A(n_284),
.B(n_271),
.C(n_272),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_304),
.B(n_281),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_292),
.A2(n_260),
.B1(n_271),
.B2(n_10),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_305),
.A2(n_286),
.B1(n_280),
.B2(n_291),
.Y(n_311)
);

AOI322xp5_ASAP7_75t_L g329 ( 
.A1(n_308),
.A2(n_5),
.A3(n_8),
.B1(n_315),
.B2(n_313),
.C1(n_314),
.C2(n_309),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_309),
.A2(n_318),
.B(n_319),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_310),
.B(n_311),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_298),
.B(n_290),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_312),
.A2(n_294),
.B1(n_6),
.B2(n_7),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_314),
.B(n_317),
.Y(n_324)
);

OR2x2_ASAP7_75t_L g315 ( 
.A(n_293),
.B(n_291),
.Y(n_315)
);

AOI221xp5_ASAP7_75t_L g322 ( 
.A1(n_315),
.A2(n_320),
.B1(n_5),
.B2(n_6),
.C(n_7),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_296),
.A2(n_13),
.B1(n_12),
.B2(n_11),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_299),
.B(n_3),
.C(n_5),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_302),
.B(n_12),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_316),
.A2(n_303),
.B(n_301),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_321),
.B(n_325),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_322),
.Y(n_334)
);

NAND4xp25_ASAP7_75t_SL g325 ( 
.A(n_320),
.B(n_304),
.C(n_6),
.D(n_7),
.Y(n_325)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_327),
.Y(n_335)
);

OAI21x1_ASAP7_75t_L g328 ( 
.A1(n_313),
.A2(n_5),
.B(n_8),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_328),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_329),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_324),
.B(n_318),
.Y(n_330)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_330),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_323),
.B(n_326),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_332),
.B(n_329),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_337),
.B(n_338),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_336),
.A2(n_322),
.B(n_333),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_340),
.B(n_339),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_341),
.A2(n_336),
.B1(n_331),
.B2(n_334),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_342),
.B(n_335),
.Y(n_343)
);


endmodule