module real_jpeg_11671_n_6 (n_5, n_4, n_36, n_0, n_37, n_1, n_2, n_33, n_34, n_35, n_3, n_6);

input n_5;
input n_4;
input n_36;
input n_0;
input n_37;
input n_1;
input n_2;
input n_33;
input n_34;
input n_35;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_21;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_7;
wire n_22;
wire n_18;
wire n_26;
wire n_27;
wire n_20;
wire n_19;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_0),
.B(n_20),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_1),
.B(n_18),
.C(n_29),
.Y(n_17)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

XOR2xp5_ASAP7_75t_L g7 ( 
.A(n_4),
.B(n_8),
.Y(n_7)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_5),
.B(n_14),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_L g6 ( 
.A(n_7),
.B(n_11),
.Y(n_6)
);

NOR2xp33_ASAP7_75t_L g8 ( 
.A(n_9),
.B(n_10),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_10),
.B(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_10),
.B(n_30),
.Y(n_29)
);

HB1xp67_ASAP7_75t_L g11 ( 
.A(n_12),
.Y(n_11)
);

A2O1A1Ixp33_ASAP7_75t_SL g12 ( 
.A1(n_13),
.A2(n_16),
.B(n_17),
.C(n_31),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_24),
.C(n_25),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_22),
.Y(n_20)
);

INVx4_ASAP7_75t_SL g22 ( 
.A(n_23),
.Y(n_22)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NOR2xp67_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_28),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_33),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_34),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_35),
.Y(n_21)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_36),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_37),
.Y(n_30)
);


endmodule