module fake_jpeg_24143_n_340 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_340);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_340;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx11_ASAP7_75t_SL g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_18),
.B(n_0),
.Y(n_36)
);

A2O1A1Ixp33_ASAP7_75t_L g64 ( 
.A1(n_36),
.A2(n_37),
.B(n_31),
.C(n_22),
.Y(n_64)
);

NAND2xp33_ASAP7_75t_SL g37 ( 
.A(n_31),
.B(n_34),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_47),
.Y(n_57)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_0),
.C(n_1),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_48),
.Y(n_61)
);

INVx3_ASAP7_75t_SL g42 ( 
.A(n_20),
.Y(n_42)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

BUFx8_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_26),
.B(n_6),
.Y(n_47)
);

CKINVDCx14_ASAP7_75t_R g48 ( 
.A(n_23),
.Y(n_48)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_50),
.B(n_56),
.Y(n_79)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_55),
.Y(n_114)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx4_ASAP7_75t_SL g96 ( 
.A(n_58),
.Y(n_96)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_60),
.Y(n_95)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_62),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_28),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_63),
.B(n_28),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_64),
.A2(n_24),
.B(n_17),
.Y(n_105)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx4_ASAP7_75t_SL g101 ( 
.A(n_65),
.Y(n_101)
);

BUFx16f_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_33),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_67),
.A2(n_73),
.B1(n_74),
.B2(n_76),
.Y(n_80)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_41),
.B(n_17),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_70),
.Y(n_86)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_71),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_39),
.A2(n_35),
.B1(n_21),
.B2(n_26),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_41),
.B(n_33),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_38),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_39),
.B(n_33),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_72),
.A2(n_35),
.B1(n_32),
.B2(n_21),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_77),
.A2(n_84),
.B(n_88),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_64),
.A2(n_40),
.B1(n_35),
.B2(n_39),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_78),
.A2(n_82),
.B1(n_100),
.B2(n_113),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_61),
.A2(n_35),
.B1(n_27),
.B2(n_42),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_72),
.A2(n_32),
.B1(n_27),
.B2(n_23),
.Y(n_84)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_85),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_58),
.A2(n_32),
.B1(n_27),
.B2(n_42),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_66),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_89),
.B(n_97),
.Y(n_122)
);

A2O1A1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_57),
.A2(n_31),
.B(n_25),
.C(n_30),
.Y(n_91)
);

A2O1A1Ixp33_ASAP7_75t_L g128 ( 
.A1(n_91),
.A2(n_22),
.B(n_19),
.C(n_44),
.Y(n_128)
);

AND2x2_ASAP7_75t_SL g92 ( 
.A(n_51),
.B(n_48),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_93),
.Y(n_118)
);

AND2x2_ASAP7_75t_SL g93 ( 
.A(n_51),
.B(n_48),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_75),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_53),
.A2(n_26),
.B1(n_29),
.B2(n_24),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_98),
.A2(n_22),
.B1(n_44),
.B2(n_18),
.Y(n_137)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_66),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_99),
.B(n_102),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_54),
.A2(n_42),
.B1(n_40),
.B2(n_29),
.Y(n_100)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_52),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_52),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_103),
.B(n_108),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_104),
.B(n_9),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_105),
.A2(n_18),
.B(n_9),
.Y(n_142)
);

AND2x6_ASAP7_75t_L g106 ( 
.A(n_63),
.B(n_14),
.Y(n_106)
);

FAx1_ASAP7_75t_SL g140 ( 
.A(n_106),
.B(n_10),
.CI(n_9),
.CON(n_140),
.SN(n_140)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_68),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_71),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_109),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_68),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_110),
.Y(n_131)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_53),
.Y(n_111)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_111),
.Y(n_126)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_55),
.Y(n_112)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_112),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_59),
.A2(n_42),
.B1(n_19),
.B2(n_43),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_86),
.B(n_42),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_115),
.A2(n_128),
.B(n_91),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_117),
.B(n_129),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_80),
.B(n_65),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_119),
.B(n_123),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_88),
.A2(n_69),
.B1(n_60),
.B2(n_43),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_120),
.A2(n_141),
.B1(n_96),
.B2(n_101),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_105),
.B(n_31),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_78),
.A2(n_44),
.B1(n_43),
.B2(n_49),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_124),
.A2(n_45),
.B1(n_16),
.B2(n_18),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_94),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_127),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_94),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_79),
.B(n_43),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_130),
.B(n_132),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_44),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_85),
.A2(n_49),
.B1(n_1),
.B2(n_2),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_134),
.A2(n_110),
.B(n_16),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_84),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_136),
.B(n_140),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_137),
.A2(n_142),
.B1(n_102),
.B2(n_96),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_77),
.A2(n_22),
.B1(n_45),
.B2(n_16),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_112),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_143),
.B(n_16),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_144),
.B(n_104),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_145),
.A2(n_159),
.B(n_164),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_118),
.B(n_93),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_147),
.B(n_156),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_148),
.A2(n_150),
.B1(n_178),
.B2(n_135),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_125),
.A2(n_114),
.B1(n_87),
.B2(n_95),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_152),
.A2(n_170),
.B1(n_137),
.B2(n_139),
.Y(n_201)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_127),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_153),
.B(n_173),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_154),
.B(n_161),
.Y(n_189)
);

MAJx2_ASAP7_75t_L g155 ( 
.A(n_115),
.B(n_106),
.C(n_93),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_SL g180 ( 
.A(n_155),
.B(n_128),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_118),
.B(n_119),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_123),
.A2(n_116),
.B(n_128),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_157),
.A2(n_169),
.B(n_140),
.Y(n_209)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_138),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_158),
.B(n_171),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_116),
.A2(n_92),
.B(n_83),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_121),
.B(n_90),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_121),
.B(n_133),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_162),
.B(n_126),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_131),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_163),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_130),
.B(n_92),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_120),
.B(n_101),
.C(n_45),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_165),
.B(n_166),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_115),
.B(n_114),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_115),
.B(n_97),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_168),
.B(n_172),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_125),
.B(n_132),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_141),
.A2(n_89),
.B1(n_81),
.B2(n_45),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_142),
.B(n_16),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_122),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_122),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_174),
.B(n_175),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_138),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_133),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_176),
.B(n_143),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_177),
.A2(n_124),
.B1(n_134),
.B2(n_135),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_180),
.B(n_196),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_181),
.B(n_182),
.Y(n_215)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_163),
.Y(n_182)
);

BUFx12_ASAP7_75t_L g183 ( 
.A(n_153),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_183),
.B(n_185),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_167),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_184),
.Y(n_213)
);

CKINVDCx14_ASAP7_75t_R g185 ( 
.A(n_146),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_160),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_187),
.B(n_188),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_177),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_190),
.A2(n_170),
.B1(n_149),
.B2(n_158),
.Y(n_226)
);

INVx13_ASAP7_75t_L g192 ( 
.A(n_173),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_192),
.Y(n_223)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_160),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_193),
.B(n_194),
.Y(n_228)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_166),
.Y(n_194)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_195),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_156),
.B(n_124),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_196),
.B(n_197),
.Y(n_233)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_152),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_164),
.B(n_126),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_198),
.A2(n_199),
.B(n_200),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_164),
.B(n_126),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_174),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_201),
.A2(n_165),
.B1(n_178),
.B2(n_151),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_176),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_202),
.Y(n_237)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_169),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_203),
.A2(n_207),
.B1(n_0),
.B2(n_2),
.Y(n_239)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_169),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_208),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_209),
.A2(n_145),
.B(n_172),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_151),
.B(n_139),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_212),
.B(n_150),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_211),
.B(n_168),
.C(n_159),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_214),
.B(n_217),
.C(n_179),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_216),
.A2(n_230),
.B1(n_232),
.B2(n_234),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_211),
.B(n_147),
.C(n_157),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_218),
.A2(n_226),
.B(n_239),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_220),
.B(n_229),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_184),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_222),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_180),
.B(n_155),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_224),
.B(n_236),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_195),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_203),
.A2(n_140),
.B1(n_131),
.B2(n_144),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_207),
.A2(n_140),
.B1(n_45),
.B2(n_18),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_205),
.A2(n_45),
.B1(n_1),
.B2(n_2),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_204),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_235),
.B(n_210),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_205),
.B(n_45),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_238),
.B(n_217),
.Y(n_251)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_183),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_240),
.B(n_183),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_241),
.B(n_244),
.C(n_254),
.Y(n_265)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_219),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_243),
.B(n_245),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_214),
.B(n_179),
.C(n_198),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_228),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_215),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_246),
.B(n_256),
.Y(n_275)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_247),
.Y(n_271)
);

AO21x1_ASAP7_75t_L g248 ( 
.A1(n_225),
.A2(n_194),
.B(n_209),
.Y(n_248)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_248),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_213),
.B(n_182),
.Y(n_249)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_249),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_251),
.B(n_253),
.Y(n_267)
);

AO22x1_ASAP7_75t_L g252 ( 
.A1(n_231),
.A2(n_188),
.B1(n_199),
.B2(n_186),
.Y(n_252)
);

OAI31xp33_ASAP7_75t_L g268 ( 
.A1(n_252),
.A2(n_220),
.A3(n_218),
.B(n_239),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_238),
.B(n_186),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_224),
.B(n_231),
.Y(n_254)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_228),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_227),
.B(n_187),
.C(n_193),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_257),
.B(n_264),
.C(n_226),
.Y(n_279)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_233),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_258),
.B(n_221),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_L g260 ( 
.A1(n_237),
.A2(n_197),
.B1(n_192),
.B2(n_200),
.Y(n_260)
);

CKINVDCx14_ASAP7_75t_R g278 ( 
.A(n_260),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_233),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_262),
.A2(n_261),
.B1(n_223),
.B2(n_206),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_263),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_216),
.B(n_212),
.C(n_181),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_252),
.A2(n_262),
.B1(n_264),
.B2(n_242),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_266),
.A2(n_255),
.B1(n_242),
.B2(n_257),
.Y(n_288)
);

XNOR2x2_ASAP7_75t_L g291 ( 
.A(n_268),
.B(n_234),
.Y(n_291)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_269),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_241),
.B(n_236),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_270),
.B(n_280),
.Y(n_298)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_252),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_276),
.A2(n_0),
.B(n_3),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_259),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_277),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_279),
.B(n_244),
.C(n_253),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_254),
.B(n_232),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_246),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_281),
.Y(n_295)
);

BUFx24_ASAP7_75t_SL g283 ( 
.A(n_248),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_283),
.B(n_230),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_284),
.A2(n_5),
.B1(n_11),
.B2(n_14),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_285),
.B(n_289),
.C(n_292),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_287),
.B(n_293),
.Y(n_313)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_288),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_265),
.B(n_251),
.C(n_250),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_291),
.A2(n_296),
.B1(n_276),
.B2(n_278),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_272),
.A2(n_255),
.B(n_191),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_265),
.B(n_250),
.C(n_240),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_266),
.A2(n_201),
.B1(n_189),
.B2(n_4),
.Y(n_294)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_294),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_268),
.B(n_8),
.Y(n_296)
);

INVx1_ASAP7_75t_SL g309 ( 
.A(n_297),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_267),
.B(n_279),
.C(n_275),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_299),
.B(n_293),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_300),
.B(n_274),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g301 ( 
.A(n_295),
.Y(n_301)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_301),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_303),
.B(n_306),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_304),
.B(n_310),
.Y(n_318)
);

INVxp33_ASAP7_75t_L g306 ( 
.A(n_291),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_308),
.B(n_285),
.C(n_289),
.Y(n_319)
);

FAx1_ASAP7_75t_SL g310 ( 
.A(n_288),
.B(n_273),
.CI(n_280),
.CON(n_310),
.SN(n_310)
);

A2O1A1Ixp33_ASAP7_75t_SL g311 ( 
.A1(n_292),
.A2(n_284),
.B(n_270),
.C(n_271),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_311),
.A2(n_294),
.B1(n_286),
.B2(n_298),
.Y(n_320)
);

OA21x2_ASAP7_75t_SL g312 ( 
.A1(n_296),
.A2(n_267),
.B(n_282),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_312),
.A2(n_290),
.B(n_299),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_314),
.A2(n_321),
.B(n_15),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_302),
.A2(n_307),
.B1(n_309),
.B2(n_306),
.Y(n_315)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_315),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_311),
.B(n_298),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_316),
.B(n_310),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_319),
.B(n_313),
.C(n_301),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_320),
.B(n_309),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_305),
.A2(n_5),
.B(n_11),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_311),
.B(n_11),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_323),
.B(n_15),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_317),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_324),
.B(n_325),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_326),
.A2(n_328),
.B(n_330),
.Y(n_331)
);

AO21x1_ASAP7_75t_L g333 ( 
.A1(n_327),
.A2(n_318),
.B(n_323),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_333),
.B(n_326),
.C(n_319),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_329),
.A2(n_322),
.B(n_316),
.Y(n_334)
);

INVxp33_ASAP7_75t_L g336 ( 
.A(n_334),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_335),
.B(n_331),
.C(n_332),
.Y(n_337)
);

AOI322xp5_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_3),
.A3(n_4),
.B1(n_15),
.B2(n_320),
.C1(n_336),
.C2(n_326),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_3),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_3),
.Y(n_340)
);


endmodule