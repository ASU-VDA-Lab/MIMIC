module fake_jpeg_22547_n_177 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_177);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_177;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_14),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx8_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_40),
.Y(n_46)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_0),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_36),
.B(n_25),
.Y(n_63)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_27),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_42),
.A2(n_16),
.B1(n_19),
.B2(n_31),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_24),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_43),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_25),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_32),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_29),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_48),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_29),
.Y(n_48)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_28),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_51),
.Y(n_83)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_55),
.B(n_58),
.Y(n_80)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

NAND2xp33_ASAP7_75t_SL g59 ( 
.A(n_37),
.B(n_27),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_35),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

AOI21xp33_ASAP7_75t_L g61 ( 
.A1(n_44),
.A2(n_17),
.B(n_22),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_61),
.Y(n_72)
);

A2O1A1Ixp33_ASAP7_75t_L g62 ( 
.A1(n_37),
.A2(n_26),
.B(n_27),
.C(n_32),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_62),
.B(n_65),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_20),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_35),
.B(n_15),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_47),
.A2(n_42),
.B1(n_38),
.B2(n_34),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_67),
.A2(n_68),
.B1(n_81),
.B2(n_84),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_62),
.A2(n_42),
.B1(n_29),
.B2(n_39),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_69),
.B(n_90),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_45),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_70),
.B(n_75),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_46),
.Y(n_71)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_71),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_50),
.A2(n_30),
.B1(n_16),
.B2(n_31),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_73),
.A2(n_40),
.B1(n_57),
.B2(n_56),
.Y(n_105)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_60),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_54),
.Y(n_91)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

A2O1A1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_76),
.A2(n_59),
.B(n_37),
.C(n_60),
.Y(n_94)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_50),
.A2(n_39),
.B1(n_30),
.B2(n_40),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_48),
.A2(n_30),
.B1(n_31),
.B2(n_28),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_54),
.A2(n_23),
.B1(n_15),
.B2(n_22),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_85),
.B(n_0),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_53),
.B(n_23),
.Y(n_86)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_86),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_63),
.B(n_37),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_89),
.B(n_63),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_45),
.B(n_22),
.Y(n_90)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_17),
.Y(n_93)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_94),
.A2(n_68),
.B(n_76),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_96),
.B(n_85),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_69),
.B(n_17),
.Y(n_99)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_99),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_66),
.B(n_13),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_100),
.B(n_106),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_77),
.B(n_58),
.Y(n_101)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_57),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_104),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_66),
.B(n_55),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_105),
.A2(n_107),
.B1(n_74),
.B2(n_82),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_72),
.B(n_6),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_89),
.B(n_52),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_109),
.B(n_84),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_113),
.B(n_123),
.Y(n_129)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_115),
.B(n_93),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_108),
.Y(n_117)
);

HB1xp67_ASAP7_75t_L g128 ( 
.A(n_117),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_104),
.B(n_67),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_118),
.A2(n_124),
.B(n_125),
.Y(n_131)
);

MAJx2_ASAP7_75t_L g119 ( 
.A(n_94),
.B(n_87),
.C(n_78),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_119),
.B(n_96),
.C(n_100),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_92),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_120),
.A2(n_122),
.B1(n_110),
.B2(n_98),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_101),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_80),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_109),
.A2(n_78),
.B(n_81),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_127),
.A2(n_105),
.B1(n_95),
.B2(n_99),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_130),
.A2(n_118),
.B1(n_121),
.B2(n_127),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_134),
.C(n_140),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_133),
.B(n_136),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_113),
.B(n_98),
.C(n_97),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_117),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_135),
.B(n_139),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_124),
.A2(n_106),
.B(n_102),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_137),
.A2(n_138),
.B1(n_141),
.B2(n_126),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_111),
.A2(n_74),
.B1(n_79),
.B2(n_103),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_116),
.A2(n_119),
.B(n_121),
.Y(n_139)
);

A2O1A1O1Ixp25_ASAP7_75t_L g140 ( 
.A1(n_125),
.A2(n_97),
.B(n_91),
.C(n_107),
.D(n_87),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_116),
.A2(n_108),
.B(n_110),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_142),
.A2(n_144),
.B1(n_147),
.B2(n_151),
.Y(n_158)
);

INVx13_ASAP7_75t_L g143 ( 
.A(n_128),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_143),
.B(n_146),
.Y(n_159)
);

INVx8_ASAP7_75t_L g144 ( 
.A(n_135),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_131),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_132),
.B(n_123),
.C(n_111),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_148),
.B(n_140),
.C(n_129),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_131),
.B(n_126),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_150),
.B(n_146),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_149),
.A2(n_134),
.B(n_114),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_152),
.A2(n_155),
.B(n_145),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_153),
.B(n_156),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_154),
.B(n_148),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_149),
.A2(n_114),
.B(n_129),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g156 ( 
.A(n_142),
.B(n_136),
.Y(n_156)
);

AOI321xp33_ASAP7_75t_L g157 ( 
.A1(n_150),
.A2(n_112),
.A3(n_18),
.B1(n_20),
.B2(n_12),
.C(n_6),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_157),
.A2(n_158),
.B(n_144),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_160),
.B(n_161),
.C(n_162),
.Y(n_169)
);

AOI221xp5_ASAP7_75t_L g161 ( 
.A1(n_159),
.A2(n_147),
.B1(n_145),
.B2(n_144),
.C(n_103),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_163),
.B(n_11),
.Y(n_166)
);

NOR2xp67_ASAP7_75t_SL g164 ( 
.A(n_153),
.B(n_143),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g168 ( 
.A(n_164),
.B(n_143),
.Y(n_168)
);

AOI322xp5_ASAP7_75t_L g173 ( 
.A1(n_166),
.A2(n_168),
.A3(n_75),
.B1(n_3),
.B2(n_4),
.C1(n_5),
.C2(n_2),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_165),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_167),
.B(n_169),
.Y(n_172)
);

OR2x2_ASAP7_75t_L g170 ( 
.A(n_164),
.B(n_13),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_170),
.B(n_1),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_171),
.B(n_172),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_173),
.A2(n_167),
.B(n_20),
.Y(n_174)
);

A2O1A1O1Ixp25_ASAP7_75t_L g176 ( 
.A1(n_174),
.A2(n_18),
.B(n_4),
.C(n_5),
.D(n_3),
.Y(n_176)
);

AOI221xp5_ASAP7_75t_L g177 ( 
.A1(n_176),
.A2(n_175),
.B1(n_4),
.B2(n_3),
.C(n_18),
.Y(n_177)
);


endmodule