module real_jpeg_2232_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_0),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_1),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_2),
.Y(n_74)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_4),
.A2(n_65),
.B1(n_66),
.B2(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_4),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_4),
.A2(n_38),
.B1(n_41),
.B2(n_104),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_4),
.A2(n_33),
.B1(n_34),
.B2(n_104),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_4),
.A2(n_54),
.B1(n_55),
.B2(n_104),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_5),
.A2(n_65),
.B1(n_66),
.B2(n_68),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_5),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_5),
.A2(n_38),
.B1(n_41),
.B2(n_68),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_5),
.A2(n_33),
.B1(n_34),
.B2(n_68),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_5),
.A2(n_54),
.B1(n_55),
.B2(n_68),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_6),
.A2(n_33),
.B1(n_34),
.B2(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_6),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_6),
.A2(n_38),
.B1(n_41),
.B2(n_58),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_6),
.A2(n_54),
.B1(n_55),
.B2(n_58),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_6),
.A2(n_58),
.B1(n_65),
.B2(n_66),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_7),
.A2(n_65),
.B1(n_66),
.B2(n_126),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_7),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_7),
.A2(n_33),
.B1(n_34),
.B2(n_126),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_7),
.A2(n_38),
.B1(n_41),
.B2(n_126),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_7),
.A2(n_54),
.B1(n_55),
.B2(n_126),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_8),
.A2(n_38),
.B1(n_41),
.B2(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_8),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_8),
.A2(n_33),
.B1(n_34),
.B2(n_46),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_8),
.A2(n_46),
.B1(n_65),
.B2(n_66),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_8),
.A2(n_46),
.B1(n_54),
.B2(n_55),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_9),
.A2(n_65),
.B1(n_66),
.B2(n_165),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_9),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_9),
.A2(n_38),
.B1(n_41),
.B2(n_165),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_9),
.A2(n_33),
.B1(n_34),
.B2(n_165),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_9),
.A2(n_54),
.B1(n_55),
.B2(n_165),
.Y(n_251)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_10),
.Y(n_67)
);

BUFx16f_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_13),
.A2(n_20),
.B(n_344),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_13),
.B(n_345),
.Y(n_344)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_14),
.A2(n_38),
.B1(n_41),
.B2(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_14),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_14),
.A2(n_43),
.B1(n_65),
.B2(n_66),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_14),
.A2(n_33),
.B1(n_34),
.B2(n_43),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_14),
.A2(n_43),
.B1(n_54),
.B2(n_55),
.Y(n_181)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_16),
.B(n_166),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_16),
.B(n_32),
.C(n_34),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_16),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_16),
.B(n_31),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_16),
.B(n_51),
.C(n_54),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_L g242 ( 
.A1(n_16),
.A2(n_33),
.B1(n_34),
.B2(n_201),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_16),
.B(n_97),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_16),
.B(n_83),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_16),
.A2(n_38),
.B1(n_41),
.B2(n_201),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_17),
.A2(n_33),
.B1(n_34),
.B2(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_17),
.A2(n_54),
.B1(n_55),
.B2(n_60),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_17),
.A2(n_38),
.B1(n_41),
.B2(n_60),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_17),
.A2(n_60),
.B1(n_65),
.B2(n_66),
.Y(n_333)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

AOI21xp33_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_339),
.B(n_342),
.Y(n_20)
);

OAI21x1_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_331),
.B(n_335),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_318),
.B(n_330),
.Y(n_22)
);

AO21x1_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_141),
.B(n_315),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_129),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_105),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_26),
.B(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_26),
.B(n_105),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_26),
.B(n_130),
.Y(n_317)
);

FAx1_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_61),
.CI(n_86),
.CON(n_26),
.SN(n_26)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_27),
.A2(n_28),
.B(n_47),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_47),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_29),
.A2(n_42),
.B1(n_44),
.B2(n_45),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_29),
.A2(n_44),
.B1(n_45),
.B2(n_80),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_29),
.A2(n_42),
.B1(n_44),
.B2(n_122),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_29),
.A2(n_44),
.B1(n_80),
.B2(n_139),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_29),
.A2(n_44),
.B1(n_174),
.B2(n_205),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_29),
.A2(n_266),
.B(n_267),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_29),
.A2(n_205),
.B(n_267),
.Y(n_285)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_30),
.B(n_162),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_30),
.A2(n_31),
.B(n_322),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_37),
.Y(n_30)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_31),
.B(n_162),
.Y(n_267)
);

AO22x1_ASAP7_75t_SL g31 ( 
.A1(n_32),
.A2(n_33),
.B1(n_34),
.B2(n_36),
.Y(n_31)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_32),
.A2(n_36),
.B1(n_38),
.B2(n_41),
.Y(n_37)
);

OAI22xp33_ASAP7_75t_L g50 ( 
.A1(n_33),
.A2(n_34),
.B1(n_51),
.B2(n_52),
.Y(n_50)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_34),
.B(n_240),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

OA22x2_ASAP7_75t_L g71 ( 
.A1(n_38),
.A2(n_41),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_38),
.B(n_191),
.Y(n_190)
);

NAND2xp33_ASAP7_75t_SL g215 ( 
.A(n_38),
.B(n_73),
.Y(n_215)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

AOI32xp33_ASAP7_75t_L g213 ( 
.A1(n_41),
.A2(n_66),
.A3(n_72),
.B1(n_214),
.B2(n_215),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_44),
.A2(n_122),
.B(n_161),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_44),
.A2(n_161),
.B(n_174),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_48),
.A2(n_53),
.B1(n_57),
.B2(n_59),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_48),
.A2(n_53),
.B1(n_57),
.B2(n_90),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_48),
.A2(n_186),
.B(n_242),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_48),
.A2(n_53),
.B1(n_184),
.B2(n_234),
.Y(n_268)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_49),
.A2(n_83),
.B(n_84),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_49),
.A2(n_83),
.B1(n_91),
.B2(n_120),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_49),
.A2(n_83),
.B1(n_120),
.B2(n_156),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_49),
.A2(n_183),
.B(n_185),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_49),
.B(n_187),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_53),
.Y(n_49)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_51),
.Y(n_52)
);

OA22x2_ASAP7_75t_L g53 ( 
.A1(n_51),
.A2(n_52),
.B1(n_54),
.B2(n_55),
.Y(n_53)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_53),
.A2(n_207),
.B(n_208),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_53),
.A2(n_208),
.B(n_234),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_54),
.B(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_54),
.B(n_247),
.Y(n_246)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_63),
.B1(n_77),
.B2(n_85),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_62),
.A2(n_63),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_SL g140 ( 
.A(n_63),
.B(n_78),
.C(n_82),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_63),
.B(n_133),
.C(n_140),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_69),
.B1(n_71),
.B2(n_76),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_64),
.A2(n_71),
.B(n_101),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_65),
.A2(n_66),
.B1(n_72),
.B2(n_73),
.Y(n_75)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

O2A1O1Ixp33_ASAP7_75t_L g200 ( 
.A1(n_66),
.A2(n_69),
.B(n_201),
.C(n_202),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_66),
.B(n_201),
.Y(n_202)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_69),
.A2(n_124),
.B(n_127),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_69),
.A2(n_71),
.B1(n_76),
.B2(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_70),
.B(n_102),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_70),
.A2(n_125),
.B1(n_164),
.B2(n_166),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_70),
.A2(n_166),
.B1(n_324),
.B2(n_325),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_70),
.A2(n_166),
.B1(n_325),
.B2(n_333),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_70),
.A2(n_166),
.B(n_333),
.Y(n_341)
);

AND2x2_ASAP7_75t_SL g70 ( 
.A(n_71),
.B(n_75),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_71),
.B(n_103),
.Y(n_128)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_71),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_71),
.A2(n_101),
.B(n_287),
.Y(n_286)
);

INVx4_ASAP7_75t_SL g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_77),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_79),
.B1(n_81),
.B2(n_82),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_81),
.A2(n_82),
.B1(n_137),
.B2(n_138),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_82),
.B(n_134),
.C(n_138),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_83),
.B(n_187),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_93),
.B(n_100),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_87),
.A2(n_88),
.B1(n_108),
.B2(n_109),
.Y(n_107)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_92),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_89),
.A2(n_92),
.B1(n_93),
.B2(n_151),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_89),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_92),
.A2(n_93),
.B1(n_100),
.B2(n_110),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_94),
.A2(n_97),
.B(n_98),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_94),
.A2(n_97),
.B1(n_117),
.B2(n_158),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_94),
.A2(n_201),
.B(n_228),
.Y(n_248)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_95),
.A2(n_96),
.B1(n_99),
.B2(n_116),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_95),
.A2(n_96),
.B1(n_180),
.B2(n_181),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_95),
.B(n_195),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_95),
.A2(n_96),
.B1(n_181),
.B2(n_218),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_95),
.A2(n_226),
.B(n_227),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_95),
.A2(n_96),
.B1(n_226),
.B2(n_256),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_96),
.A2(n_180),
.B(n_193),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_96),
.B(n_195),
.Y(n_228)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_97),
.A2(n_194),
.B(n_251),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_100),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_111),
.C(n_112),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_106),
.A2(n_107),
.B1(n_111),
.B2(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_111),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_112),
.B(n_144),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_121),
.C(n_123),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_113),
.A2(n_114),
.B1(n_148),
.B2(n_149),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_118),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_115),
.A2(n_118),
.B1(n_119),
.B2(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_115),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_SL g149 ( 
.A(n_121),
.B(n_123),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_128),
.B(n_200),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_129),
.A2(n_316),
.B(n_317),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_140),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_136),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_135),
.Y(n_324)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_139),
.Y(n_322)
);

AO21x1_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_167),
.B(n_314),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_143),
.B(n_146),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_143),
.B(n_146),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_150),
.C(n_152),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_147),
.B(n_150),
.Y(n_312)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_152),
.B(n_312),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_159),
.C(n_163),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_153),
.A2(n_154),
.B1(n_302),
.B2(n_304),
.Y(n_301)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_155),
.B(n_157),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_155),
.B(n_157),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_156),
.Y(n_207)
);

CKINVDCx14_ASAP7_75t_R g218 ( 
.A(n_158),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_159),
.A2(n_160),
.B1(n_163),
.B2(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_163),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_164),
.Y(n_287)
);

OAI21x1_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_309),
.B(n_313),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_169),
.A2(n_278),
.B(n_306),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_220),
.B(n_277),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_196),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_171),
.B(n_196),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_182),
.C(n_188),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_172),
.B(n_274),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_175),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_173),
.B(n_176),
.C(n_179),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_177),
.B1(n_178),
.B2(n_179),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_182),
.B(n_188),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_192),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_189),
.A2(n_190),
.B1(n_192),
.B2(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_192),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_210),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_197),
.B(n_211),
.C(n_219),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_199),
.B1(n_203),
.B2(n_209),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_198),
.B(n_204),
.C(n_206),
.Y(n_291)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_202),
.Y(n_214)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_203),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_204),
.B(n_206),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_219),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_213),
.B1(n_216),
.B2(n_217),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_212),
.B(n_217),
.Y(n_282)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_272),
.B(n_276),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_222),
.A2(n_261),
.B(n_271),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_243),
.B(n_260),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_224),
.B(n_237),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_224),
.B(n_237),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_229),
.B1(n_235),
.B2(n_236),
.Y(n_224)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_225),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_229),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_231),
.B1(n_232),
.B2(n_233),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_231),
.B(n_232),
.C(n_235),
.Y(n_262)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_241),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_238),
.A2(n_239),
.B1(n_241),
.B2(n_258),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_241),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_254),
.B(n_259),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_249),
.B(n_253),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_248),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_250),
.B(n_252),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_250),
.B(n_252),
.Y(n_253)
);

CKINVDCx14_ASAP7_75t_R g256 ( 
.A(n_251),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_257),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_255),
.B(n_257),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_262),
.B(n_263),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_269),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_268),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_265),
.B(n_268),
.C(n_269),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_273),
.B(n_275),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_273),
.B(n_275),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_293),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_280),
.B(n_292),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_280),
.B(n_292),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_289),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_281),
.B(n_290),
.C(n_291),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_SL g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_282),
.B(n_284),
.C(n_288),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_285),
.B1(n_286),
.B2(n_288),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_286),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_293),
.A2(n_307),
.B(n_308),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_294),
.B(n_305),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_294),
.B(n_305),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_295),
.A2(n_296),
.B1(n_297),
.B2(n_298),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_295),
.B(n_299),
.C(n_301),
.Y(n_310)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_SL g298 ( 
.A(n_299),
.B(n_301),
.Y(n_298)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_302),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_310),
.B(n_311),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_329),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_319),
.B(n_329),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_328),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_321),
.A2(n_323),
.B1(n_326),
.B2(n_327),
.Y(n_320)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_321),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_323),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_323),
.B(n_326),
.C(n_328),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_334),
.Y(n_331)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_332),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_332),
.B(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_334),
.Y(n_338)
);

CKINVDCx14_ASAP7_75t_R g335 ( 
.A(n_336),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_338),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_337),
.B(n_341),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_341),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_343),
.Y(n_342)
);


endmodule