module fake_jpeg_9019_n_227 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_227);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_227;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx11_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_29),
.B(n_32),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g30 ( 
.A(n_17),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_30),
.B(n_37),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_34),
.Y(n_46)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_15),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_36),
.Y(n_50)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_43),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_37),
.A2(n_20),
.B1(n_25),
.B2(n_24),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_41),
.A2(n_51),
.B1(n_54),
.B2(n_16),
.Y(n_65)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_37),
.A2(n_20),
.B1(n_25),
.B2(n_18),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_47),
.A2(n_49),
.B1(n_24),
.B2(n_22),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_33),
.A2(n_20),
.B1(n_36),
.B2(n_34),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_30),
.A2(n_25),
.B1(n_22),
.B2(n_21),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_52),
.B(n_57),
.Y(n_64)
);

BUFx8_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_53),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_30),
.A2(n_22),
.B1(n_16),
.B2(n_19),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_28),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_55),
.B(n_57),
.Y(n_76)
);

NAND2xp33_ASAP7_75t_SL g56 ( 
.A(n_30),
.B(n_23),
.Y(n_56)
);

A2O1A1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_56),
.A2(n_32),
.B(n_39),
.C(n_38),
.Y(n_59)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_59),
.A2(n_41),
.B(n_49),
.Y(n_79)
);

OR2x4_ASAP7_75t_L g60 ( 
.A(n_56),
.B(n_50),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_SL g95 ( 
.A(n_60),
.B(n_76),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_42),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_61),
.B(n_62),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_52),
.B(n_15),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_65),
.A2(n_69),
.B1(n_19),
.B2(n_44),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_27),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_67),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_39),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_28),
.Y(n_68)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_44),
.A2(n_28),
.B1(n_16),
.B2(n_19),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_39),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_70),
.B(n_48),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_71),
.A2(n_48),
.B1(n_27),
.B2(n_26),
.Y(n_87)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_73),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_24),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_21),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_74),
.B(n_75),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_21),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_63),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_85),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_79),
.A2(n_81),
.B1(n_86),
.B2(n_87),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_60),
.B(n_47),
.C(n_40),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_72),
.C(n_67),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_61),
.A2(n_44),
.B1(n_48),
.B2(n_45),
.Y(n_86)
);

INVx13_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_88),
.B(n_93),
.Y(n_110)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_91),
.B(n_70),
.Y(n_100)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_92),
.Y(n_112)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_59),
.A2(n_45),
.B1(n_26),
.B2(n_43),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_94),
.A2(n_93),
.B1(n_90),
.B2(n_82),
.Y(n_109)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_97),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_73),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_98),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_SL g122 ( 
.A(n_100),
.B(n_84),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_103),
.C(n_107),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_95),
.B(n_64),
.C(n_59),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_91),
.A2(n_45),
.B1(n_64),
.B2(n_68),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_105),
.A2(n_115),
.B1(n_92),
.B2(n_88),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_95),
.B(n_75),
.C(n_74),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_109),
.A2(n_111),
.B1(n_83),
.B2(n_90),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_94),
.A2(n_66),
.B1(n_62),
.B2(n_53),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_82),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_113),
.B(n_114),
.Y(n_121)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_80),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_79),
.A2(n_66),
.B1(n_53),
.B2(n_23),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_84),
.B(n_23),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_0),
.C(n_1),
.Y(n_137)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_80),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_13),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_96),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_118),
.A2(n_78),
.B(n_88),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_97),
.Y(n_119)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_119),
.Y(n_152)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_120),
.B(n_127),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_131),
.C(n_137),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_96),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_123),
.B(n_126),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_125),
.A2(n_106),
.B1(n_99),
.B2(n_111),
.Y(n_146)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_110),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_87),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_128),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_129),
.B(n_112),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_115),
.A2(n_92),
.B1(n_89),
.B2(n_53),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_130),
.A2(n_104),
.B1(n_4),
.B2(n_5),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_116),
.B(n_23),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_108),
.A2(n_23),
.B(n_53),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_132),
.A2(n_138),
.B1(n_2),
.B2(n_5),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_109),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_133),
.B(n_135),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_134),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_105),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_118),
.A2(n_0),
.B(n_1),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_136),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_99),
.A2(n_2),
.B(n_4),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_143),
.A2(n_149),
.B1(n_6),
.B2(n_7),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_122),
.B(n_107),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_144),
.B(n_119),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_146),
.B(n_147),
.Y(n_167)
);

INVx13_ASAP7_75t_L g147 ( 
.A(n_127),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_121),
.B(n_104),
.Y(n_148)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_148),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_133),
.B(n_120),
.Y(n_150)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_150),
.Y(n_168)
);

CKINVDCx14_ASAP7_75t_R g174 ( 
.A(n_151),
.Y(n_174)
);

INVxp67_ASAP7_75t_SL g153 ( 
.A(n_121),
.Y(n_153)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_153),
.Y(n_169)
);

INVx13_ASAP7_75t_L g154 ( 
.A(n_126),
.Y(n_154)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_154),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_134),
.B(n_5),
.Y(n_156)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_156),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_141),
.B(n_124),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_158),
.B(n_162),
.C(n_165),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_160),
.B(n_144),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_140),
.B(n_124),
.C(n_123),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_154),
.A2(n_132),
.B1(n_135),
.B2(n_129),
.Y(n_163)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_163),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_141),
.A2(n_138),
.B(n_128),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_164),
.A2(n_171),
.B1(n_139),
.B2(n_157),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_140),
.B(n_131),
.C(n_125),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_155),
.B(n_137),
.C(n_130),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_166),
.B(n_152),
.C(n_145),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_148),
.B(n_136),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_170),
.B(n_156),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_147),
.Y(n_173)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_173),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_173),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_175),
.B(n_183),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_176),
.A2(n_185),
.B1(n_167),
.B2(n_174),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_159),
.B(n_155),
.Y(n_177)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_177),
.Y(n_196)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_178),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_179),
.B(n_182),
.Y(n_195)
);

BUFx24_ASAP7_75t_SL g181 ( 
.A(n_158),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_181),
.B(n_184),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_160),
.B(n_146),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_168),
.B(n_142),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_172),
.A2(n_154),
.B1(n_145),
.B2(n_152),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_159),
.B(n_147),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_186),
.B(n_161),
.Y(n_190)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_190),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_188),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_191),
.B(n_157),
.Y(n_201)
);

AOI21x1_ASAP7_75t_L g192 ( 
.A1(n_185),
.A2(n_164),
.B(n_169),
.Y(n_192)
);

AO22x1_ASAP7_75t_L g207 ( 
.A1(n_192),
.A2(n_198),
.B1(n_199),
.B2(n_149),
.Y(n_207)
);

INVxp33_ASAP7_75t_L g193 ( 
.A(n_187),
.Y(n_193)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_193),
.Y(n_204)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_194),
.Y(n_208)
);

AO21x1_ASAP7_75t_L g198 ( 
.A1(n_182),
.A2(n_142),
.B(n_151),
.Y(n_198)
);

NOR2x1_ASAP7_75t_L g199 ( 
.A(n_183),
.B(n_166),
.Y(n_199)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_201),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_196),
.B(n_171),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_203),
.B(n_209),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_200),
.A2(n_165),
.B1(n_162),
.B2(n_180),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_205),
.B(n_206),
.C(n_9),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_195),
.B(n_179),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_199),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_204),
.A2(n_197),
.B(n_189),
.Y(n_210)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_210),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_203),
.B(n_198),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_211),
.B(n_207),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_202),
.A2(n_195),
.B(n_8),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_213),
.B(n_215),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_208),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_214),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_217),
.B(n_219),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_220),
.A2(n_216),
.B(n_212),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_222),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_218),
.B(n_220),
.C(n_215),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_224),
.B(n_221),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_225),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_226),
.B(n_223),
.Y(n_227)
);


endmodule