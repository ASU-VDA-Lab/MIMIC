module fake_jpeg_6118_n_279 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_279);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_279;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx14_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_33),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_37),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_38),
.A2(n_24),
.B1(n_30),
.B2(n_18),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_40),
.Y(n_44)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_38),
.A2(n_24),
.B1(n_22),
.B2(n_18),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_42),
.A2(n_25),
.B1(n_28),
.B2(n_27),
.Y(n_80)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_45),
.Y(n_62)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_46),
.A2(n_30),
.B1(n_17),
.B2(n_38),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_47),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_L g48 ( 
.A1(n_35),
.A2(n_21),
.B1(n_30),
.B2(n_32),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_48),
.A2(n_60),
.B1(n_31),
.B2(n_23),
.Y(n_86)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_49),
.B(n_51),
.Y(n_65)
);

OAI21xp33_ASAP7_75t_L g50 ( 
.A1(n_40),
.A2(n_22),
.B(n_27),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_50),
.A2(n_52),
.B1(n_17),
.B2(n_19),
.Y(n_75)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

NAND2xp33_ASAP7_75t_SL g52 ( 
.A(n_40),
.B(n_28),
.Y(n_52)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_54),
.B(n_58),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_55),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_36),
.B(n_23),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_57),
.B(n_31),
.Y(n_81)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_38),
.A2(n_32),
.B1(n_16),
.B2(n_25),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_59),
.B(n_34),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_61),
.B(n_71),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_60),
.B(n_16),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_63),
.B(n_81),
.Y(n_100)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_64),
.B(n_67),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_L g68 ( 
.A1(n_52),
.A2(n_35),
.B1(n_33),
.B2(n_34),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_68),
.A2(n_80),
.B1(n_86),
.B2(n_26),
.Y(n_107)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_69),
.B(n_77),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_70),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_34),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_44),
.B(n_34),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_72),
.B(n_73),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_41),
.B(n_33),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_33),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_74),
.B(n_82),
.Y(n_96)
);

A2O1A1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_75),
.A2(n_26),
.B(n_20),
.C(n_15),
.Y(n_110)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_78),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_53),
.B(n_33),
.Y(n_82)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_53),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_55),
.Y(n_90)
);

OA22x2_ASAP7_75t_L g87 ( 
.A1(n_53),
.A2(n_35),
.B1(n_33),
.B2(n_39),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_87),
.A2(n_43),
.B1(n_49),
.B2(n_45),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_55),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_88),
.Y(n_99)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_87),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_89),
.B(n_102),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_90),
.B(n_62),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_61),
.B(n_55),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_103),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_101),
.A2(n_106),
.B1(n_107),
.B2(n_87),
.Y(n_117)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_71),
.B(n_39),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_76),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_104),
.B(n_109),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_68),
.A2(n_21),
.B1(n_26),
.B2(n_20),
.Y(n_106)
);

OAI21xp33_ASAP7_75t_L g108 ( 
.A1(n_75),
.A2(n_0),
.B(n_2),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_108),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_65),
.B(n_2),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_110),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_74),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_112),
.B(n_69),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_72),
.B(n_26),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_113),
.B(n_114),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_73),
.A2(n_86),
.B(n_82),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_105),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_115),
.B(n_121),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_117),
.A2(n_98),
.B1(n_90),
.B2(n_7),
.Y(n_171)
);

INVx6_ASAP7_75t_SL g118 ( 
.A(n_111),
.Y(n_118)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_118),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_122),
.Y(n_145)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_91),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_123),
.B(n_125),
.Y(n_146)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_91),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_126),
.B(n_90),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_96),
.B(n_83),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_129),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_96),
.B(n_84),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_112),
.B(n_78),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_133),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_89),
.A2(n_70),
.B1(n_77),
.B2(n_64),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_131),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_99),
.B(n_67),
.Y(n_132)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_132),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_103),
.B(n_85),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_93),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_134),
.B(n_136),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_92),
.B(n_79),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_135),
.B(n_139),
.Y(n_170)
);

BUFx2_ASAP7_75t_SL g136 ( 
.A(n_94),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_99),
.B(n_3),
.Y(n_138)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_138),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_114),
.B(n_3),
.Y(n_139)
);

INVx13_ASAP7_75t_L g140 ( 
.A(n_104),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_140),
.B(n_142),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_92),
.B(n_79),
.Y(n_141)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_141),
.Y(n_152)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_97),
.Y(n_142)
);

OA21x2_ASAP7_75t_L g143 ( 
.A1(n_137),
.A2(n_101),
.B(n_102),
.Y(n_143)
);

OA21x2_ASAP7_75t_L g177 ( 
.A1(n_143),
.A2(n_133),
.B(n_117),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_124),
.B(n_113),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_144),
.B(n_140),
.C(n_121),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_132),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_150),
.B(n_164),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_118),
.Y(n_151)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_151),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_124),
.A2(n_95),
.B(n_110),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_153),
.A2(n_159),
.B(n_8),
.Y(n_194)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_129),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_155),
.B(n_157),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_127),
.A2(n_95),
.B1(n_107),
.B2(n_106),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_156),
.Y(n_187)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_130),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_135),
.A2(n_141),
.B(n_119),
.Y(n_159)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_122),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_161),
.B(n_163),
.Y(n_185)
);

CKINVDCx12_ASAP7_75t_R g163 ( 
.A(n_140),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_128),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_165),
.B(n_126),
.Y(n_172)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_119),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_167),
.B(n_14),
.Y(n_191)
);

OR2x2_ASAP7_75t_L g168 ( 
.A(n_139),
.B(n_100),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_168),
.A2(n_123),
.B1(n_125),
.B2(n_120),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_171),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_172),
.A2(n_177),
.B(n_192),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_173),
.B(n_152),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_160),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_174),
.Y(n_203)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_166),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_178),
.B(n_180),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_160),
.A2(n_115),
.B1(n_142),
.B2(n_98),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_179),
.A2(n_194),
.B(n_148),
.Y(n_215)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_147),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g181 ( 
.A(n_147),
.B(n_116),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_181),
.B(n_186),
.C(n_189),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_151),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_182),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_154),
.B(n_116),
.Y(n_183)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_183),
.Y(n_197)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_188),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_144),
.B(n_121),
.C(n_6),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_159),
.B(n_15),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_190),
.B(n_193),
.Y(n_205)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_191),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_153),
.A2(n_4),
.B(n_7),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_154),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_156),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_195),
.A2(n_171),
.B1(n_170),
.B2(n_149),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_152),
.B(n_9),
.Y(n_196)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_196),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_185),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_199),
.A2(n_212),
.B(n_215),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_206),
.A2(n_211),
.B1(n_195),
.B2(n_176),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_183),
.B(n_170),
.Y(n_207)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_207),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_180),
.B(n_155),
.Y(n_208)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_208),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_196),
.B(n_146),
.Y(n_210)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_210),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_186),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_187),
.A2(n_165),
.B1(n_157),
.B2(n_149),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_213),
.A2(n_214),
.B1(n_172),
.B2(n_175),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_187),
.A2(n_165),
.B1(n_143),
.B2(n_145),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_184),
.B(n_169),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_216),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_209),
.B(n_194),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_218),
.B(n_223),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_219),
.A2(n_221),
.B1(n_206),
.B2(n_207),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_198),
.A2(n_177),
.B1(n_181),
.B2(n_188),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_209),
.B(n_190),
.C(n_189),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_222),
.B(n_226),
.C(n_228),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_198),
.B(n_192),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_204),
.Y(n_224)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_224),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_205),
.B(n_177),
.C(n_176),
.Y(n_226)
);

FAx1_ASAP7_75t_SL g239 ( 
.A(n_227),
.B(n_215),
.CI(n_204),
.CON(n_239),
.SN(n_239)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_205),
.B(n_162),
.C(n_182),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_214),
.B(n_143),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_230),
.B(n_233),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_208),
.B(n_168),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_234),
.A2(n_239),
.B(n_240),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_226),
.A2(n_211),
.B1(n_213),
.B2(n_201),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_236),
.Y(n_253)
);

OA21x2_ASAP7_75t_SL g240 ( 
.A1(n_218),
.A2(n_197),
.B(n_216),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_221),
.B(n_219),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_241),
.B(n_242),
.C(n_234),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_232),
.A2(n_201),
.B1(n_197),
.B2(n_217),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_228),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_243),
.A2(n_244),
.B(n_225),
.Y(n_250)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_223),
.Y(n_244)
);

AO221x1_ASAP7_75t_L g246 ( 
.A1(n_238),
.A2(n_200),
.B1(n_203),
.B2(n_229),
.C(n_231),
.Y(n_246)
);

INVx11_ASAP7_75t_L g261 ( 
.A(n_246),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_235),
.B(n_237),
.C(n_241),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_248),
.B(n_249),
.C(n_255),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_250),
.B(n_254),
.Y(n_259)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_239),
.Y(n_251)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_251),
.Y(n_262)
);

OAI321xp33_ASAP7_75t_L g252 ( 
.A1(n_239),
.A2(n_233),
.A3(n_220),
.B1(n_230),
.B2(n_210),
.C(n_217),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_252),
.B(n_202),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_245),
.B(n_235),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_237),
.B(n_222),
.C(n_199),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_253),
.A2(n_203),
.B(n_245),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_256),
.A2(n_260),
.B(n_10),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_247),
.A2(n_200),
.B1(n_158),
.B2(n_202),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_257),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_258),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_251),
.B(n_10),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_262),
.B(n_255),
.Y(n_264)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_264),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_256),
.B(n_248),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_265),
.A2(n_266),
.B(n_268),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_267),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_261),
.B(n_12),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_269),
.B(n_261),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_273),
.B(n_257),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_274),
.B(n_275),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_270),
.A2(n_263),
.B(n_259),
.Y(n_275)
);

AOI211xp5_ASAP7_75t_L g277 ( 
.A1(n_276),
.A2(n_271),
.B(n_272),
.C(n_263),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_277),
.B(n_12),
.C(n_13),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_278),
.B(n_13),
.Y(n_279)
);


endmodule