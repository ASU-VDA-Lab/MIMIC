module fake_jpeg_24652_n_344 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_344);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_344;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_17),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_37),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_40),
.Y(n_63)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_17),
.B(n_21),
.Y(n_42)
);

NAND2xp33_ASAP7_75t_SL g57 ( 
.A(n_42),
.B(n_20),
.Y(n_57)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_43),
.B(n_44),
.Y(n_70)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_46),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_25),
.B(n_0),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_30),
.Y(n_66)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_50),
.B(n_58),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_46),
.A2(n_23),
.B1(n_32),
.B2(n_21),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_51),
.A2(n_54),
.B1(n_60),
.B2(n_62),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_21),
.C(n_26),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_52),
.B(n_57),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_46),
.A2(n_23),
.B1(n_32),
.B2(n_26),
.Y(n_54)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_59),
.A2(n_27),
.B1(n_35),
.B2(n_40),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_46),
.A2(n_25),
.B1(n_35),
.B2(n_22),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_42),
.A2(n_22),
.B1(n_27),
.B2(n_30),
.Y(n_62)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_66),
.B(n_67),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_48),
.A2(n_35),
.B1(n_30),
.B2(n_27),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_67),
.A2(n_31),
.B1(n_24),
.B2(n_18),
.Y(n_89)
);

BUFx16f_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_69),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_63),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_71),
.B(n_73),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_66),
.B(n_47),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_74),
.A2(n_91),
.B(n_102),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_51),
.A2(n_39),
.B1(n_44),
.B2(n_40),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_75),
.A2(n_89),
.B1(n_90),
.B2(n_100),
.Y(n_103)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_76),
.B(n_77),
.Y(n_132)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_52),
.A2(n_40),
.B1(n_44),
.B2(n_39),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_80),
.A2(n_88),
.B1(n_55),
.B2(n_65),
.Y(n_106)
);

BUFx8_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_82),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_83),
.B(n_84),
.Y(n_118)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

A2O1A1Ixp33_ASAP7_75t_L g86 ( 
.A1(n_57),
.A2(n_52),
.B(n_62),
.C(n_70),
.Y(n_86)
);

A2O1A1Ixp33_ASAP7_75t_L g109 ( 
.A1(n_86),
.A2(n_20),
.B(n_36),
.C(n_29),
.Y(n_109)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_87),
.B(n_92),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_55),
.A2(n_43),
.B1(n_41),
.B2(n_37),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_54),
.A2(n_43),
.B1(n_41),
.B2(n_42),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_69),
.A2(n_31),
.B1(n_19),
.B2(n_28),
.Y(n_91)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_94),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_63),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_95),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_97),
.B(n_36),
.Y(n_112)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_98),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_59),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_99),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_60),
.A2(n_43),
.B1(n_41),
.B2(n_42),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_61),
.B(n_18),
.Y(n_101)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_101),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_64),
.A2(n_42),
.B(n_24),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_106),
.A2(n_126),
.B1(n_87),
.B2(n_82),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_80),
.B(n_61),
.C(n_64),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_107),
.B(n_125),
.C(n_127),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_71),
.A2(n_95),
.B1(n_81),
.B2(n_89),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_108),
.A2(n_115),
.B1(n_122),
.B2(n_72),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_109),
.A2(n_112),
.B(n_84),
.Y(n_147)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_96),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_128),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_L g115 ( 
.A1(n_97),
.A2(n_64),
.B1(n_65),
.B2(n_58),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_69),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_117),
.B(n_119),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_85),
.B(n_58),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_99),
.A2(n_55),
.B1(n_53),
.B2(n_19),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_121),
.A2(n_94),
.B1(n_92),
.B2(n_98),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_81),
.A2(n_53),
.B1(n_69),
.B2(n_49),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_85),
.B(n_38),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_124),
.B(n_34),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_85),
.B(n_45),
.C(n_49),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_86),
.A2(n_50),
.B1(n_34),
.B2(n_45),
.Y(n_126)
);

MAJx2_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_83),
.C(n_90),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_88),
.Y(n_128)
);

AOI32xp33_ASAP7_75t_L g129 ( 
.A1(n_93),
.A2(n_45),
.A3(n_36),
.B1(n_29),
.B2(n_34),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g157 ( 
.A(n_129),
.B(n_122),
.Y(n_157)
);

AOI21xp33_ASAP7_75t_L g130 ( 
.A1(n_93),
.A2(n_28),
.B(n_20),
.Y(n_130)
);

AOI21xp33_ASAP7_75t_L g159 ( 
.A1(n_130),
.A2(n_9),
.B(n_16),
.Y(n_159)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_123),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_133),
.B(n_139),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_123),
.Y(n_136)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_136),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_137),
.A2(n_152),
.B1(n_128),
.B2(n_109),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_131),
.Y(n_138)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_138),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_113),
.B(n_72),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_114),
.B(n_75),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_141),
.B(n_148),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_113),
.B(n_105),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_142),
.B(n_149),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_143),
.A2(n_146),
.B(n_147),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_103),
.A2(n_79),
.B1(n_78),
.B2(n_76),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_144),
.A2(n_145),
.B1(n_109),
.B2(n_121),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_103),
.A2(n_79),
.B1(n_78),
.B2(n_77),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_119),
.B(n_20),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_118),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_118),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_150),
.B(n_151),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_110),
.B(n_82),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_105),
.B(n_82),
.Y(n_153)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_153),
.Y(n_165)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_114),
.B(n_20),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_154),
.B(n_155),
.Y(n_195)
);

OR2x2_ASAP7_75t_L g155 ( 
.A(n_117),
.B(n_34),
.Y(n_155)
);

AND2x2_ASAP7_75t_SL g156 ( 
.A(n_124),
.B(n_33),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_156),
.B(n_0),
.C(n_1),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_157),
.B(n_120),
.Y(n_170)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_132),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_158),
.A2(n_159),
.B(n_15),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_131),
.Y(n_160)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_160),
.Y(n_185)
);

INVx8_ASAP7_75t_L g161 ( 
.A(n_110),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_161),
.A2(n_116),
.B1(n_131),
.B2(n_129),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_112),
.B(n_33),
.Y(n_162)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_162),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_132),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_163),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_166),
.A2(n_169),
.B1(n_175),
.B2(n_177),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_170),
.B(n_173),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_134),
.B(n_125),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_152),
.A2(n_120),
.B1(n_104),
.B2(n_107),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_139),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_176),
.B(n_188),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_147),
.A2(n_127),
.B1(n_106),
.B2(n_117),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_134),
.B(n_140),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_178),
.B(n_183),
.Y(n_225)
);

NAND3xp33_ASAP7_75t_L g179 ( 
.A(n_149),
.B(n_111),
.C(n_127),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_179),
.B(n_192),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_181),
.A2(n_184),
.B1(n_133),
.B2(n_158),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_140),
.B(n_126),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_135),
.A2(n_116),
.B1(n_36),
.B2(n_29),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_148),
.B(n_33),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_186),
.B(n_190),
.C(n_196),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_141),
.A2(n_29),
.B1(n_33),
.B2(n_2),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_187),
.A2(n_193),
.B1(n_145),
.B2(n_144),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_163),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_156),
.B(n_33),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_142),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_191),
.B(n_192),
.Y(n_216)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_135),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_137),
.A2(n_16),
.B1(n_15),
.B2(n_14),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_194),
.A2(n_153),
.B(n_150),
.Y(n_200)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_168),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_197),
.B(n_211),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_199),
.A2(n_200),
.B(n_208),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_181),
.A2(n_157),
.B1(n_143),
.B2(n_146),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_201),
.A2(n_204),
.B1(n_207),
.B2(n_215),
.Y(n_240)
);

AO21x1_ASAP7_75t_L g251 ( 
.A1(n_203),
.A2(n_209),
.B(n_185),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_191),
.B(n_154),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_205),
.B(n_219),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_174),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_206),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_182),
.A2(n_161),
.B1(n_160),
.B2(n_138),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_195),
.A2(n_155),
.B(n_156),
.Y(n_208)
);

AND2x4_ASAP7_75t_SL g209 ( 
.A(n_195),
.B(n_155),
.Y(n_209)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_171),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_184),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_212),
.B(n_218),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_180),
.A2(n_162),
.B1(n_156),
.B2(n_154),
.Y(n_213)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_213),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_180),
.A2(n_160),
.B(n_138),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_172),
.B(n_189),
.Y(n_217)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_217),
.Y(n_236)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_182),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_172),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_187),
.Y(n_220)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_220),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_196),
.Y(n_221)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_221),
.Y(n_249)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_164),
.Y(n_222)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_222),
.Y(n_241)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_183),
.Y(n_223)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_223),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_189),
.B(n_161),
.Y(n_224)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_224),
.Y(n_252)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_169),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_226),
.A2(n_165),
.B1(n_185),
.B2(n_3),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_225),
.B(n_178),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_229),
.B(n_234),
.Y(n_256)
);

CKINVDCx14_ASAP7_75t_R g232 ( 
.A(n_215),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_232),
.B(n_238),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_210),
.B(n_173),
.C(n_190),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_233),
.B(n_235),
.C(n_245),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_225),
.B(n_170),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_210),
.B(n_186),
.C(n_177),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_202),
.B(n_167),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_237),
.B(n_221),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_224),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_214),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_239),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_216),
.Y(n_243)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_243),
.Y(n_258)
);

AND2x6_ASAP7_75t_L g244 ( 
.A(n_209),
.B(n_165),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_244),
.A2(n_251),
.B(n_212),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_202),
.B(n_194),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_246),
.A2(n_220),
.B1(n_206),
.B2(n_218),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_253),
.B(n_269),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_257),
.A2(n_274),
.B1(n_231),
.B2(n_236),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_242),
.B(n_197),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_259),
.B(n_268),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_228),
.A2(n_204),
.B1(n_230),
.B2(n_226),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_261),
.A2(n_264),
.B1(n_272),
.B2(n_4),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_233),
.B(n_223),
.C(n_198),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_262),
.B(n_263),
.C(n_266),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_249),
.B(n_198),
.C(n_217),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_250),
.A2(n_222),
.B1(n_201),
.B2(n_200),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_238),
.B(n_208),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_267),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_249),
.B(n_213),
.C(n_209),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_242),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_250),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_247),
.B(n_211),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_270),
.Y(n_285)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_251),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_271),
.B(n_227),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_231),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_235),
.B(n_229),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_273),
.B(n_245),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_240),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_254),
.B(n_241),
.Y(n_275)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_275),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_256),
.B(n_234),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_276),
.B(n_282),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_258),
.B(n_248),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_279),
.B(n_284),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_255),
.Y(n_281)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_281),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_256),
.B(n_237),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_286),
.B(n_289),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_263),
.B(n_252),
.C(n_236),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_287),
.B(n_266),
.C(n_255),
.Y(n_295)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_288),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_273),
.B(n_227),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_265),
.A2(n_244),
.B1(n_252),
.B2(n_9),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_290),
.B(n_291),
.Y(n_297)
);

NOR3xp33_ASAP7_75t_SL g292 ( 
.A(n_278),
.B(n_253),
.C(n_272),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_292),
.B(n_7),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_295),
.A2(n_299),
.B(n_302),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_287),
.B(n_283),
.C(n_277),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_291),
.B(n_257),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_301),
.B(n_306),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_283),
.B(n_277),
.C(n_282),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_285),
.A2(n_274),
.B1(n_270),
.B2(n_269),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_304),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_280),
.A2(n_260),
.B(n_262),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_305),
.B(n_14),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_286),
.B(n_260),
.Y(n_306)
);

BUFx24_ASAP7_75t_SL g307 ( 
.A(n_293),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_307),
.B(n_309),
.Y(n_328)
);

INVx11_ASAP7_75t_L g309 ( 
.A(n_298),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_292),
.B(n_289),
.Y(n_311)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_311),
.Y(n_321)
);

A2O1A1Ixp33_ASAP7_75t_L g312 ( 
.A1(n_297),
.A2(n_276),
.B(n_9),
.C(n_10),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_312),
.A2(n_316),
.B(n_300),
.Y(n_324)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_313),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_303),
.A2(n_8),
.B1(n_10),
.B2(n_12),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_314),
.A2(n_318),
.B1(n_319),
.B2(n_7),
.Y(n_322)
);

NOR2xp67_ASAP7_75t_L g315 ( 
.A(n_300),
.B(n_8),
.Y(n_315)
);

NOR2xp67_ASAP7_75t_SL g325 ( 
.A(n_315),
.B(n_296),
.Y(n_325)
);

OAI321xp33_ASAP7_75t_L g316 ( 
.A1(n_294),
.A2(n_14),
.A3(n_10),
.B1(n_7),
.B2(n_6),
.C(n_5),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_317),
.B(n_310),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_303),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_318)
);

A2O1A1Ixp33_ASAP7_75t_SL g320 ( 
.A1(n_309),
.A2(n_298),
.B(n_295),
.C(n_299),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_320),
.A2(n_323),
.B(n_326),
.Y(n_330)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_322),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_308),
.A2(n_302),
.B(n_305),
.Y(n_323)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_324),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_325),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_312),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_329),
.B(n_317),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_331),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_329),
.B(n_318),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_333),
.B(n_334),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_SL g334 ( 
.A(n_321),
.B(n_296),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_333),
.B(n_327),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_338),
.A2(n_339),
.B(n_332),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_330),
.A2(n_335),
.B(n_336),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_341),
.B(n_337),
.C(n_340),
.Y(n_342)
);

AO21x2_ASAP7_75t_L g343 ( 
.A1(n_342),
.A2(n_320),
.B(n_328),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_343),
.B(n_320),
.Y(n_344)
);


endmodule