module real_aes_1932_n_105 (n_17, n_28, n_76, n_56, n_34, n_98, n_832, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_104, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_833, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_105);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_832;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_104;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_833;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_105;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_785;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_L g234 ( .A(n_0), .B(n_156), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_1), .B(n_116), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g830 ( .A(n_2), .Y(n_830) );
INVx1_ASAP7_75t_L g149 ( .A(n_3), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_4), .B(n_162), .Y(n_175) );
NAND2xp33_ASAP7_75t_SL g226 ( .A(n_5), .B(n_160), .Y(n_226) );
INVx1_ASAP7_75t_L g207 ( .A(n_6), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g553 ( .A(n_7), .B(n_180), .Y(n_553) );
OAI22xp5_ASAP7_75t_SL g122 ( .A1(n_8), .A2(n_123), .B1(n_124), .B2(n_126), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_8), .Y(n_123) );
INVx1_ASAP7_75t_L g533 ( .A(n_9), .Y(n_533) );
CKINVDCx16_ASAP7_75t_R g116 ( .A(n_10), .Y(n_116) );
AND2x2_ASAP7_75t_L g173 ( .A(n_11), .B(n_166), .Y(n_173) );
CKINVDCx5p33_ASAP7_75t_R g500 ( .A(n_12), .Y(n_500) );
INVx2_ASAP7_75t_L g167 ( .A(n_13), .Y(n_167) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_14), .Y(n_125) );
NOR3xp33_ASAP7_75t_L g114 ( .A(n_15), .B(n_115), .C(n_117), .Y(n_114) );
CKINVDCx16_ASAP7_75t_R g132 ( .A(n_15), .Y(n_132) );
NOR2xp33_ASAP7_75t_L g729 ( .A(n_15), .B(n_28), .Y(n_729) );
INVx1_ASAP7_75t_L g561 ( .A(n_16), .Y(n_561) );
OAI22xp5_ASAP7_75t_SL g817 ( .A1(n_17), .A2(n_28), .B1(n_783), .B2(n_818), .Y(n_817) );
CKINVDCx20_ASAP7_75t_R g818 ( .A(n_17), .Y(n_818) );
AOI221x1_ASAP7_75t_L g220 ( .A1(n_18), .A2(n_144), .B1(n_221), .B2(n_223), .C(n_225), .Y(n_220) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_19), .B(n_162), .Y(n_195) );
INVx1_ASAP7_75t_L g112 ( .A(n_20), .Y(n_112) );
INVx1_ASAP7_75t_L g559 ( .A(n_21), .Y(n_559) );
INVx1_ASAP7_75t_SL g482 ( .A(n_22), .Y(n_482) );
NAND2xp5_ASAP7_75t_SL g549 ( .A(n_23), .B(n_163), .Y(n_549) );
AOI21xp5_ASAP7_75t_L g176 ( .A1(n_24), .A2(n_144), .B(n_177), .Y(n_176) );
AOI221xp5_ASAP7_75t_SL g187 ( .A1(n_25), .A2(n_41), .B1(n_144), .B2(n_162), .C(n_188), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_26), .B(n_156), .Y(n_178) );
AOI33xp33_ASAP7_75t_L g519 ( .A1(n_27), .A2(n_54), .A3(n_210), .B1(n_216), .B2(n_520), .B3(n_521), .Y(n_519) );
INVx1_ASAP7_75t_L g783 ( .A(n_28), .Y(n_783) );
INVx1_ASAP7_75t_L g493 ( .A(n_29), .Y(n_493) );
OR2x2_ASAP7_75t_L g168 ( .A(n_30), .B(n_94), .Y(n_168) );
OA21x2_ASAP7_75t_L g201 ( .A1(n_30), .A2(n_94), .B(n_167), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_31), .B(n_152), .Y(n_199) );
INVxp67_ASAP7_75t_L g219 ( .A(n_32), .Y(n_219) );
AND2x2_ASAP7_75t_L g250 ( .A(n_33), .B(n_165), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_34), .B(n_208), .Y(n_479) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_35), .A2(n_144), .B(n_233), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_36), .B(n_152), .Y(n_189) );
AND2x2_ASAP7_75t_L g145 ( .A(n_37), .B(n_146), .Y(n_145) );
AND2x2_ASAP7_75t_L g160 ( .A(n_37), .B(n_149), .Y(n_160) );
INVx1_ASAP7_75t_L g215 ( .A(n_37), .Y(n_215) );
INVxp67_ASAP7_75t_L g117 ( .A(n_38), .Y(n_117) );
OR2x6_ASAP7_75t_L g793 ( .A(n_38), .B(n_111), .Y(n_793) );
CKINVDCx20_ASAP7_75t_R g495 ( .A(n_39), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_40), .B(n_208), .Y(n_507) );
AOI22xp5_ASAP7_75t_L g542 ( .A1(n_42), .A2(n_180), .B1(n_224), .B2(n_543), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_43), .B(n_551), .Y(n_550) );
AOI22xp5_ASAP7_75t_L g286 ( .A1(n_44), .A2(n_84), .B1(n_144), .B2(n_213), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_45), .B(n_163), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_46), .B(n_156), .Y(n_248) );
INVx1_ASAP7_75t_L g791 ( .A(n_47), .Y(n_791) );
XNOR2xp5_ASAP7_75t_L g820 ( .A(n_48), .B(n_88), .Y(n_820) );
NAND2xp5_ASAP7_75t_SL g535 ( .A(n_49), .B(n_200), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_50), .B(n_163), .Y(n_534) );
CKINVDCx5p33_ASAP7_75t_R g546 ( .A(n_51), .Y(n_546) );
AND2x2_ASAP7_75t_L g237 ( .A(n_52), .B(n_165), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_53), .B(n_165), .Y(n_191) );
XOR2xp5_ASAP7_75t_L g812 ( .A(n_53), .B(n_813), .Y(n_812) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_55), .B(n_163), .Y(n_511) );
INVx1_ASAP7_75t_L g148 ( .A(n_56), .Y(n_148) );
INVx1_ASAP7_75t_L g158 ( .A(n_56), .Y(n_158) );
AND2x2_ASAP7_75t_L g512 ( .A(n_57), .B(n_165), .Y(n_512) );
AOI221xp5_ASAP7_75t_L g531 ( .A1(n_58), .A2(n_77), .B1(n_208), .B2(n_213), .C(n_532), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_59), .B(n_208), .Y(n_476) );
NAND2xp5_ASAP7_75t_SL g249 ( .A(n_60), .B(n_162), .Y(n_249) );
OAI22xp5_ASAP7_75t_SL g121 ( .A1(n_61), .A2(n_122), .B1(n_127), .B2(n_128), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_61), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_62), .B(n_224), .Y(n_502) );
AOI21xp5_ASAP7_75t_SL g471 ( .A1(n_63), .A2(n_213), .B(n_472), .Y(n_471) );
AND2x2_ASAP7_75t_L g169 ( .A(n_64), .B(n_165), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_65), .B(n_152), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_66), .B(n_156), .Y(n_155) );
AND2x2_ASAP7_75t_SL g202 ( .A(n_67), .B(n_166), .Y(n_202) );
INVx1_ASAP7_75t_L g556 ( .A(n_68), .Y(n_556) );
XNOR2xp5_ASAP7_75t_L g124 ( .A(n_69), .B(n_125), .Y(n_124) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_70), .A2(n_144), .B(n_246), .Y(n_245) );
INVx1_ASAP7_75t_L g510 ( .A(n_71), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_72), .B(n_152), .Y(n_179) );
AND2x2_ASAP7_75t_SL g287 ( .A(n_73), .B(n_200), .Y(n_287) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_74), .A2(n_213), .B(n_509), .Y(n_508) );
INVx1_ASAP7_75t_L g146 ( .A(n_75), .Y(n_146) );
INVx1_ASAP7_75t_L g154 ( .A(n_75), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_76), .B(n_208), .Y(n_522) );
AND2x2_ASAP7_75t_L g484 ( .A(n_78), .B(n_223), .Y(n_484) );
INVx1_ASAP7_75t_L g557 ( .A(n_79), .Y(n_557) );
AOI21xp5_ASAP7_75t_L g480 ( .A1(n_80), .A2(n_213), .B(n_481), .Y(n_480) );
A2O1A1Ixp33_ASAP7_75t_L g547 ( .A1(n_81), .A2(n_213), .B(n_283), .C(n_548), .Y(n_547) );
NAND2xp5_ASAP7_75t_SL g161 ( .A(n_82), .B(n_162), .Y(n_161) );
AOI22xp5_ASAP7_75t_L g285 ( .A1(n_83), .A2(n_87), .B1(n_162), .B2(n_208), .Y(n_285) );
INVx1_ASAP7_75t_L g113 ( .A(n_85), .Y(n_113) );
AND2x2_ASAP7_75t_SL g469 ( .A(n_86), .B(n_223), .Y(n_469) );
AOI22xp5_ASAP7_75t_L g516 ( .A1(n_89), .A2(n_213), .B1(n_517), .B2(n_518), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_90), .B(n_156), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_91), .B(n_156), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g794 ( .A(n_92), .B(n_795), .Y(n_794) );
AOI21xp5_ASAP7_75t_L g143 ( .A1(n_93), .A2(n_144), .B(n_150), .Y(n_143) );
INVx1_ASAP7_75t_L g473 ( .A(n_95), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_96), .B(n_152), .Y(n_151) );
AND2x2_ASAP7_75t_L g523 ( .A(n_97), .B(n_223), .Y(n_523) );
A2O1A1Ixp33_ASAP7_75t_L g490 ( .A1(n_98), .A2(n_491), .B(n_492), .C(n_494), .Y(n_490) );
INVxp67_ASAP7_75t_L g222 ( .A(n_99), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_100), .B(n_162), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_101), .B(n_152), .Y(n_247) );
AOI21xp5_ASAP7_75t_L g196 ( .A1(n_102), .A2(n_144), .B(n_197), .Y(n_196) );
BUFx2_ASAP7_75t_SL g789 ( .A(n_103), .Y(n_789) );
BUFx2_ASAP7_75t_L g804 ( .A(n_103), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_104), .B(n_163), .Y(n_475) );
AOI21xp5_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_118), .B(n_829), .Y(n_105) );
BUFx3_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_SL g107 ( .A(n_108), .Y(n_107) );
INVx2_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
NOR2xp33_ASAP7_75t_L g829 ( .A(n_109), .B(n_830), .Y(n_829) );
AND2x2_ASAP7_75t_SL g109 ( .A(n_110), .B(n_114), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_112), .B(n_113), .Y(n_111) );
AND2x4_ASAP7_75t_L g118 ( .A(n_119), .B(n_805), .Y(n_118) );
AOI21xp5_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_785), .B(n_799), .Y(n_119) );
NOR2xp33_ASAP7_75t_L g120 ( .A(n_121), .B(n_129), .Y(n_120) );
CKINVDCx16_ASAP7_75t_R g828 ( .A(n_121), .Y(n_828) );
INVxp33_ASAP7_75t_L g128 ( .A(n_122), .Y(n_128) );
INVx1_ASAP7_75t_L g126 ( .A(n_124), .Y(n_126) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
HB1xp67_ASAP7_75t_L g827 ( .A(n_130), .Y(n_827) );
OAI21x1_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_133), .B(n_459), .Y(n_130) );
HB1xp67_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
CKINVDCx16_ASAP7_75t_R g784 ( .A(n_132), .Y(n_784) );
OR2x2_ASAP7_75t_L g792 ( .A(n_132), .B(n_793), .Y(n_792) );
NAND2xp5_ASAP7_75t_L g797 ( .A(n_132), .B(n_798), .Y(n_797) );
AND2x4_ASAP7_75t_L g133 ( .A(n_134), .B(n_398), .Y(n_133) );
NOR3xp33_ASAP7_75t_L g134 ( .A(n_135), .B(n_291), .C(n_342), .Y(n_134) );
OAI211xp5_ASAP7_75t_SL g135 ( .A1(n_136), .A2(n_181), .B(n_238), .C(n_269), .Y(n_135) );
INVxp67_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
NOR2xp33_ASAP7_75t_L g137 ( .A(n_138), .B(n_170), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
HB1xp67_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_140), .B(n_243), .Y(n_406) );
INVx1_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
AND2x2_ASAP7_75t_L g251 ( .A(n_141), .B(n_172), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_141), .B(n_258), .Y(n_257) );
OR2x2_ASAP7_75t_L g268 ( .A(n_141), .B(n_258), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_141), .B(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g305 ( .A(n_141), .B(n_281), .Y(n_305) );
INVx2_ASAP7_75t_L g331 ( .A(n_141), .Y(n_331) );
AND2x4_ASAP7_75t_L g340 ( .A(n_141), .B(n_341), .Y(n_340) );
AND2x2_ASAP7_75t_L g445 ( .A(n_141), .B(n_312), .Y(n_445) );
AO21x2_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_164), .B(n_169), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_143), .B(n_161), .Y(n_142) );
AND2x6_ASAP7_75t_L g144 ( .A(n_145), .B(n_147), .Y(n_144) );
BUFx3_ASAP7_75t_L g212 ( .A(n_145), .Y(n_212) );
AND2x6_ASAP7_75t_L g156 ( .A(n_146), .B(n_157), .Y(n_156) );
INVx2_ASAP7_75t_L g217 ( .A(n_146), .Y(n_217) );
AND2x4_ASAP7_75t_L g213 ( .A(n_147), .B(n_214), .Y(n_213) );
AND2x2_ASAP7_75t_L g147 ( .A(n_148), .B(n_149), .Y(n_147) );
AND2x4_ASAP7_75t_L g152 ( .A(n_148), .B(n_153), .Y(n_152) );
INVx2_ASAP7_75t_L g210 ( .A(n_148), .Y(n_210) );
HB1xp67_ASAP7_75t_L g211 ( .A(n_149), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_155), .B(n_159), .Y(n_150) );
INVxp67_ASAP7_75t_L g562 ( .A(n_152), .Y(n_562) );
AND2x4_ASAP7_75t_L g163 ( .A(n_153), .B(n_157), .Y(n_163) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVxp67_ASAP7_75t_L g560 ( .A(n_156), .Y(n_560) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
AOI21xp5_ASAP7_75t_L g177 ( .A1(n_159), .A2(n_178), .B(n_179), .Y(n_177) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_159), .A2(n_189), .B(n_190), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g197 ( .A1(n_159), .A2(n_198), .B(n_199), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g233 ( .A1(n_159), .A2(n_234), .B(n_235), .Y(n_233) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_159), .A2(n_247), .B(n_248), .Y(n_246) );
O2A1O1Ixp33_ASAP7_75t_L g472 ( .A1(n_159), .A2(n_473), .B(n_474), .C(n_475), .Y(n_472) );
O2A1O1Ixp33_ASAP7_75t_SL g481 ( .A1(n_159), .A2(n_474), .B(n_482), .C(n_483), .Y(n_481) );
O2A1O1Ixp33_ASAP7_75t_L g509 ( .A1(n_159), .A2(n_474), .B(n_510), .C(n_511), .Y(n_509) );
INVx1_ASAP7_75t_L g517 ( .A(n_159), .Y(n_517) );
O2A1O1Ixp33_ASAP7_75t_SL g532 ( .A1(n_159), .A2(n_474), .B(n_533), .C(n_534), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g548 ( .A1(n_159), .A2(n_549), .B(n_550), .Y(n_548) );
NOR2xp33_ASAP7_75t_L g563 ( .A(n_159), .B(n_180), .Y(n_563) );
INVx5_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
AND2x4_ASAP7_75t_L g162 ( .A(n_160), .B(n_163), .Y(n_162) );
HB1xp67_ASAP7_75t_L g494 ( .A(n_160), .Y(n_494) );
INVx1_ASAP7_75t_L g227 ( .A(n_163), .Y(n_227) );
AO21x2_ASAP7_75t_L g243 ( .A1(n_164), .A2(n_244), .B(n_250), .Y(n_243) );
AO21x2_ASAP7_75t_L g258 ( .A1(n_164), .A2(n_244), .B(n_250), .Y(n_258) );
AO21x2_ASAP7_75t_L g477 ( .A1(n_164), .A2(n_478), .B(n_484), .Y(n_477) );
CKINVDCx5p33_ASAP7_75t_R g164 ( .A(n_165), .Y(n_164) );
OA21x2_ASAP7_75t_L g186 ( .A1(n_165), .A2(n_187), .B(n_191), .Y(n_186) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
AND2x2_ASAP7_75t_SL g166 ( .A(n_167), .B(n_168), .Y(n_166) );
AND2x4_ASAP7_75t_L g180 ( .A(n_167), .B(n_168), .Y(n_180) );
AND2x2_ASAP7_75t_L g329 ( .A(n_170), .B(n_330), .Y(n_329) );
OAI32xp33_ASAP7_75t_L g412 ( .A1(n_170), .A2(n_334), .A3(n_338), .B1(n_345), .B2(n_413), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_170), .B(n_445), .Y(n_444) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
AND2x2_ASAP7_75t_L g266 ( .A(n_171), .B(n_267), .Y(n_266) );
NAND3xp33_ASAP7_75t_L g339 ( .A(n_171), .B(n_261), .C(n_340), .Y(n_339) );
OR2x2_ASAP7_75t_L g365 ( .A(n_171), .B(n_268), .Y(n_365) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
HB1xp67_ASAP7_75t_L g255 ( .A(n_172), .Y(n_255) );
INVx5_ASAP7_75t_L g290 ( .A(n_172), .Y(n_290) );
AND2x4_ASAP7_75t_L g346 ( .A(n_172), .B(n_258), .Y(n_346) );
OR2x2_ASAP7_75t_L g361 ( .A(n_172), .B(n_281), .Y(n_361) );
OR2x2_ASAP7_75t_L g387 ( .A(n_172), .B(n_243), .Y(n_387) );
AND2x2_ASAP7_75t_L g395 ( .A(n_172), .B(n_341), .Y(n_395) );
AND2x4_ASAP7_75t_SL g420 ( .A(n_172), .B(n_340), .Y(n_420) );
OR2x6_ASAP7_75t_L g172 ( .A(n_173), .B(n_174), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g174 ( .A1(n_175), .A2(n_176), .B(n_180), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g206 ( .A(n_180), .B(n_207), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_180), .B(n_219), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_180), .B(n_222), .Y(n_221) );
NOR3xp33_ASAP7_75t_L g225 ( .A(n_180), .B(n_226), .C(n_227), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_180), .A2(n_471), .B(n_476), .Y(n_470) );
INVx1_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_182), .B(n_340), .Y(n_416) );
AND2x2_ASAP7_75t_L g182 ( .A(n_183), .B(n_192), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_183), .B(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
OR2x6_ASAP7_75t_SL g240 ( .A(n_184), .B(n_241), .Y(n_240) );
INVxp67_ASAP7_75t_SL g184 ( .A(n_185), .Y(n_184) );
INVx1_ASAP7_75t_L g265 ( .A(n_185), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_185), .B(n_300), .Y(n_318) );
HB1xp67_ASAP7_75t_L g456 ( .A(n_185), .Y(n_456) );
INVx1_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
INVx2_ASAP7_75t_L g273 ( .A(n_186), .Y(n_273) );
AND2x2_ASAP7_75t_L g298 ( .A(n_186), .B(n_229), .Y(n_298) );
INVx2_ASAP7_75t_L g326 ( .A(n_186), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_186), .B(n_193), .Y(n_367) );
BUFx3_ASAP7_75t_L g391 ( .A(n_186), .Y(n_391) );
OR2x2_ASAP7_75t_L g403 ( .A(n_186), .B(n_193), .Y(n_403) );
HB1xp67_ASAP7_75t_L g411 ( .A(n_186), .Y(n_411) );
AOI22xp5_ASAP7_75t_L g433 ( .A1(n_192), .A2(n_434), .B1(n_437), .B2(n_438), .Y(n_433) );
AND2x2_ASAP7_75t_L g192 ( .A(n_193), .B(n_203), .Y(n_192) );
INVx1_ASAP7_75t_L g261 ( .A(n_193), .Y(n_261) );
OR2x2_ASAP7_75t_L g272 ( .A(n_193), .B(n_273), .Y(n_272) );
INVx2_ASAP7_75t_L g279 ( .A(n_193), .Y(n_279) );
AND2x4_ASAP7_75t_SL g296 ( .A(n_193), .B(n_204), .Y(n_296) );
AND2x4_ASAP7_75t_L g301 ( .A(n_193), .B(n_302), .Y(n_301) );
INVx2_ASAP7_75t_L g310 ( .A(n_193), .Y(n_310) );
OR2x2_ASAP7_75t_L g316 ( .A(n_193), .B(n_204), .Y(n_316) );
OR2x2_ASAP7_75t_L g317 ( .A(n_193), .B(n_318), .Y(n_317) );
HB1xp67_ASAP7_75t_L g428 ( .A(n_193), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_193), .B(n_298), .Y(n_432) );
OR2x2_ASAP7_75t_L g448 ( .A(n_193), .B(n_351), .Y(n_448) );
OR2x6_ASAP7_75t_L g193 ( .A(n_194), .B(n_202), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_195), .A2(n_196), .B(n_200), .Y(n_194) );
INVx2_ASAP7_75t_SL g283 ( .A(n_200), .Y(n_283) );
OA21x2_ASAP7_75t_L g530 ( .A1(n_200), .A2(n_531), .B(n_535), .Y(n_530) );
BUFx4f_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
INVx3_ASAP7_75t_L g224 ( .A(n_201), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_203), .B(n_261), .Y(n_260) );
INVx1_ASAP7_75t_L g274 ( .A(n_203), .Y(n_274) );
AND2x2_ASAP7_75t_SL g381 ( .A(n_203), .B(n_265), .Y(n_381) );
AND2x4_ASAP7_75t_L g203 ( .A(n_204), .B(n_228), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_204), .B(n_229), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g262 ( .A(n_204), .B(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_204), .B(n_273), .Y(n_277) );
INVx3_ASAP7_75t_L g302 ( .A(n_204), .Y(n_302) );
INVx1_ASAP7_75t_L g335 ( .A(n_204), .Y(n_335) );
AND2x2_ASAP7_75t_L g415 ( .A(n_204), .B(n_279), .Y(n_415) );
AND2x4_ASAP7_75t_L g204 ( .A(n_205), .B(n_220), .Y(n_204) );
AOI22xp5_ASAP7_75t_L g205 ( .A1(n_206), .A2(n_208), .B1(n_213), .B2(n_218), .Y(n_205) );
INVx1_ASAP7_75t_L g503 ( .A(n_208), .Y(n_503) );
AND2x4_ASAP7_75t_L g208 ( .A(n_209), .B(n_212), .Y(n_208) );
INVx1_ASAP7_75t_L g544 ( .A(n_209), .Y(n_544) );
AND2x2_ASAP7_75t_L g209 ( .A(n_210), .B(n_211), .Y(n_209) );
OR2x6_ASAP7_75t_L g474 ( .A(n_210), .B(n_217), .Y(n_474) );
INVxp33_ASAP7_75t_L g520 ( .A(n_210), .Y(n_520) );
INVx1_ASAP7_75t_L g545 ( .A(n_212), .Y(n_545) );
INVxp67_ASAP7_75t_L g501 ( .A(n_213), .Y(n_501) );
NOR2x1p5_ASAP7_75t_L g214 ( .A(n_215), .B(n_216), .Y(n_214) );
INVx1_ASAP7_75t_L g521 ( .A(n_216), .Y(n_521) );
INVx3_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
OAI22xp5_ASAP7_75t_L g489 ( .A1(n_223), .A2(n_490), .B1(n_495), .B2(n_496), .Y(n_489) );
INVx3_ASAP7_75t_L g496 ( .A(n_223), .Y(n_496) );
INVx4_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
AOI21x1_ASAP7_75t_L g230 ( .A1(n_224), .A2(n_231), .B(n_237), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_224), .B(n_499), .Y(n_498) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_227), .B(n_493), .Y(n_492) );
OAI22xp5_ASAP7_75t_L g555 ( .A1(n_227), .A2(n_474), .B1(n_556), .B2(n_557), .Y(n_555) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_229), .B(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g300 ( .A(n_229), .Y(n_300) );
AND2x2_ASAP7_75t_L g325 ( .A(n_229), .B(n_326), .Y(n_325) );
OR2x2_ASAP7_75t_L g351 ( .A(n_229), .B(n_273), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_229), .B(n_302), .Y(n_368) );
INVx1_ASAP7_75t_L g374 ( .A(n_229), .Y(n_374) );
INVx3_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_232), .B(n_236), .Y(n_231) );
AOI222xp33_ASAP7_75t_SL g238 ( .A1(n_239), .A2(n_242), .B1(n_252), .B2(n_259), .C1(n_262), .C2(n_266), .Y(n_238) );
CKINVDCx16_ASAP7_75t_R g239 ( .A(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_L g242 ( .A(n_243), .B(n_251), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g363 ( .A(n_243), .B(n_312), .Y(n_363) );
AND2x4_ASAP7_75t_L g379 ( .A(n_243), .B(n_290), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_245), .B(n_249), .Y(n_244) );
INVx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
NAND2xp5_ASAP7_75t_SL g253 ( .A(n_254), .B(n_256), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g304 ( .A(n_255), .B(n_305), .Y(n_304) );
AOI222xp33_ASAP7_75t_L g269 ( .A1(n_256), .A2(n_270), .B1(n_275), .B2(n_280), .C1(n_288), .C2(n_832), .Y(n_269) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
OR2x2_ASAP7_75t_L g408 ( .A(n_257), .B(n_312), .Y(n_408) );
OR2x2_ASAP7_75t_L g451 ( .A(n_257), .B(n_357), .Y(n_451) );
AND2x2_ASAP7_75t_L g280 ( .A(n_258), .B(n_281), .Y(n_280) );
INVx2_ASAP7_75t_L g341 ( .A(n_258), .Y(n_341) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_258), .Y(n_356) );
O2A1O1Ixp33_ASAP7_75t_L g369 ( .A1(n_259), .A2(n_370), .B(n_375), .C(n_376), .Y(n_369) );
INVx1_ASAP7_75t_SL g259 ( .A(n_260), .Y(n_259) );
INVx1_ASAP7_75t_L g397 ( .A(n_261), .Y(n_397) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
HB1xp67_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
INVx2_ASAP7_75t_L g327 ( .A(n_266), .Y(n_327) );
AND2x2_ASAP7_75t_L g311 ( .A(n_267), .B(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g320 ( .A(n_267), .B(n_321), .Y(n_320) );
INVx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
OAI31xp33_ASAP7_75t_L g362 ( .A1(n_270), .A2(n_288), .A3(n_363), .B(n_364), .Y(n_362) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
A2O1A1Ixp33_ASAP7_75t_L g364 ( .A1(n_271), .A2(n_321), .B(n_365), .C(n_366), .Y(n_364) );
OR2x2_ASAP7_75t_L g271 ( .A(n_272), .B(n_274), .Y(n_271) );
OR2x2_ASAP7_75t_L g353 ( .A(n_272), .B(n_302), .Y(n_353) );
INVx2_ASAP7_75t_SL g275 ( .A(n_276), .Y(n_275) );
OR2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
BUFx2_ASAP7_75t_L g321 ( .A(n_281), .Y(n_321) );
AND2x2_ASAP7_75t_L g330 ( .A(n_281), .B(n_331), .Y(n_330) );
INVx2_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
BUFx6f_ASAP7_75t_L g312 ( .A(n_282), .Y(n_312) );
AOI21x1_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_284), .B(n_287), .Y(n_282) );
AO21x2_ASAP7_75t_L g514 ( .A1(n_283), .A2(n_515), .B(n_523), .Y(n_514) );
AO21x2_ASAP7_75t_L g574 ( .A1(n_283), .A2(n_515), .B(n_523), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_290), .B(n_347), .Y(n_439) );
OAI211xp5_ASAP7_75t_L g291 ( .A1(n_292), .A2(n_303), .B(n_306), .C(n_328), .Y(n_291) );
INVxp33_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_SL g293 ( .A(n_294), .B(n_299), .Y(n_293) );
OR2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_297), .Y(n_294) );
INVx1_ASAP7_75t_SL g295 ( .A(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g332 ( .A(n_296), .B(n_325), .Y(n_332) );
OR2x2_ASAP7_75t_L g308 ( .A(n_297), .B(n_309), .Y(n_308) );
OR2x2_ASAP7_75t_L g338 ( .A(n_297), .B(n_312), .Y(n_338) );
INVx2_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g414 ( .A(n_298), .B(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g437 ( .A(n_299), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_301), .B(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_301), .B(n_372), .Y(n_371) );
AND2x2_ASAP7_75t_L g449 ( .A(n_301), .B(n_325), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_301), .B(n_455), .Y(n_454) );
AND2x2_ASAP7_75t_L g392 ( .A(n_302), .B(n_374), .Y(n_392) );
INVx1_ASAP7_75t_SL g303 ( .A(n_304), .Y(n_303) );
AOI322xp5_ASAP7_75t_L g446 ( .A1(n_305), .A2(n_325), .A3(n_379), .B1(n_404), .B2(n_447), .C1(n_449), .C2(n_450), .Y(n_446) );
AOI211xp5_ASAP7_75t_SL g306 ( .A1(n_307), .A2(n_311), .B(n_313), .C(n_322), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_309), .B(n_337), .Y(n_359) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g324 ( .A(n_310), .B(n_325), .Y(n_324) );
NOR2x1p5_ASAP7_75t_L g390 ( .A(n_310), .B(n_391), .Y(n_390) );
HB1xp67_ASAP7_75t_L g423 ( .A(n_310), .Y(n_423) );
O2A1O1Ixp33_ASAP7_75t_L g328 ( .A1(n_311), .A2(n_329), .B(n_332), .C(n_333), .Y(n_328) );
AND2x4_ASAP7_75t_L g347 ( .A(n_312), .B(n_331), .Y(n_347) );
INVx2_ASAP7_75t_L g357 ( .A(n_312), .Y(n_357) );
NAND2xp5_ASAP7_75t_SL g377 ( .A(n_312), .B(n_346), .Y(n_377) );
AND2x2_ASAP7_75t_L g419 ( .A(n_312), .B(n_420), .Y(n_419) );
NOR2xp33_ASAP7_75t_L g457 ( .A(n_312), .B(n_436), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_312), .B(n_340), .Y(n_458) );
AOI21xp33_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_317), .B(n_319), .Y(n_313) );
AND2x2_ASAP7_75t_L g409 ( .A(n_315), .B(n_410), .Y(n_409) );
INVx1_ASAP7_75t_SL g315 ( .A(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g337 ( .A(n_318), .Y(n_337) );
INVx2_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_323), .B(n_327), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_330), .B(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g424 ( .A(n_330), .Y(n_424) );
O2A1O1Ixp33_ASAP7_75t_SL g333 ( .A1(n_334), .A2(n_336), .B(n_338), .C(n_339), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
HB1xp67_ASAP7_75t_L g421 ( .A(n_337), .Y(n_421) );
INVx3_ASAP7_75t_SL g436 ( .A(n_340), .Y(n_436) );
NAND5xp2_ASAP7_75t_L g342 ( .A(n_343), .B(n_362), .C(n_369), .D(n_382), .E(n_393), .Y(n_342) );
AOI222xp33_ASAP7_75t_L g343 ( .A1(n_344), .A2(n_348), .B1(n_352), .B2(n_354), .C1(n_358), .C2(n_360), .Y(n_343) );
NOR2xp33_ASAP7_75t_L g344 ( .A(n_345), .B(n_347), .Y(n_344) );
AOI22xp5_ASAP7_75t_L g425 ( .A1(n_345), .A2(n_426), .B1(n_430), .B2(n_431), .Y(n_425) );
INVx2_ASAP7_75t_SL g345 ( .A(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g375 ( .A(n_346), .B(n_347), .Y(n_375) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_SL g352 ( .A(n_353), .Y(n_352) );
NOR2xp33_ASAP7_75t_L g354 ( .A(n_355), .B(n_357), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
NAND2xp5_ASAP7_75t_SL g442 ( .A(n_356), .B(n_443), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_357), .B(n_379), .Y(n_378) );
AND2x2_ASAP7_75t_L g394 ( .A(n_357), .B(n_395), .Y(n_394) );
OR2x2_ASAP7_75t_L g405 ( .A(n_357), .B(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_SL g360 ( .A(n_361), .Y(n_360) );
OR2x2_ASAP7_75t_L g435 ( .A(n_361), .B(n_436), .Y(n_435) );
OR2x2_ASAP7_75t_L g366 ( .A(n_367), .B(n_368), .Y(n_366) );
INVx1_ASAP7_75t_L g383 ( .A(n_368), .Y(n_383) );
INVxp67_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVxp67_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
HB1xp67_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
AOI21xp33_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_378), .B(n_380), .Y(n_376) );
AOI22xp33_ASAP7_75t_L g382 ( .A1(n_379), .A2(n_383), .B1(n_384), .B2(n_388), .Y(n_382) );
HB1xp67_ASAP7_75t_L g430 ( .A(n_379), .Y(n_430) );
INVx2_ASAP7_75t_SL g380 ( .A(n_381), .Y(n_380) );
AND2x2_ASAP7_75t_L g396 ( .A(n_381), .B(n_397), .Y(n_396) );
AND2x2_ASAP7_75t_L g401 ( .A(n_383), .B(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_SL g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_390), .B(n_392), .Y(n_389) );
INVx1_ASAP7_75t_SL g429 ( .A(n_392), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_394), .B(n_396), .Y(n_393) );
NOR3xp33_ASAP7_75t_L g398 ( .A(n_399), .B(n_417), .C(n_440), .Y(n_398) );
NAND2xp5_ASAP7_75t_SL g399 ( .A(n_400), .B(n_416), .Y(n_399) );
AOI221xp5_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_404), .B1(n_407), .B2(n_409), .C(n_412), .Y(n_400) );
INVx1_ASAP7_75t_SL g402 ( .A(n_403), .Y(n_402) );
OR2x2_ASAP7_75t_L g441 ( .A(n_403), .B(n_429), .Y(n_441) );
INVx1_ASAP7_75t_SL g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_SL g407 ( .A(n_408), .Y(n_407) );
HB1xp67_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_SL g413 ( .A(n_414), .Y(n_413) );
OAI321xp33_ASAP7_75t_L g417 ( .A1(n_418), .A2(n_421), .A3(n_422), .B1(n_424), .B2(n_425), .C(n_433), .Y(n_417) );
INVx1_ASAP7_75t_SL g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_SL g426 ( .A(n_427), .Y(n_426) );
OR2x2_ASAP7_75t_L g427 ( .A(n_428), .B(n_429), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g452 ( .A1(n_431), .A2(n_453), .B1(n_457), .B2(n_458), .Y(n_452) );
INVx1_ASAP7_75t_SL g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
OAI211xp5_ASAP7_75t_SL g440 ( .A1(n_441), .A2(n_442), .B(n_446), .C(n_452), .Y(n_440) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_SL g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVxp67_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
NOR2x1_ASAP7_75t_L g459 ( .A(n_460), .B(n_780), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_461), .B(n_730), .Y(n_460) );
OAI21xp5_ASAP7_75t_L g461 ( .A1(n_462), .A2(n_670), .B(n_729), .Y(n_461) );
NOR3xp33_ASAP7_75t_L g780 ( .A(n_462), .B(n_731), .C(n_781), .Y(n_780) );
INVx1_ASAP7_75t_L g823 ( .A(n_462), .Y(n_823) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_463), .B(n_634), .Y(n_462) );
NOR3xp33_ASAP7_75t_L g463 ( .A(n_464), .B(n_575), .C(n_604), .Y(n_463) );
NAND2xp5_ASAP7_75t_SL g464 ( .A(n_465), .B(n_564), .Y(n_464) );
AOI22xp5_ASAP7_75t_L g465 ( .A1(n_466), .A2(n_485), .B1(n_524), .B2(n_536), .Y(n_465) );
NAND2x1_ASAP7_75t_L g766 ( .A(n_466), .B(n_565), .Y(n_766) );
INVx2_ASAP7_75t_SL g466 ( .A(n_467), .Y(n_466) );
OR2x2_ASAP7_75t_L g467 ( .A(n_468), .B(n_477), .Y(n_467) );
INVx2_ASAP7_75t_L g538 ( .A(n_468), .Y(n_538) );
INVx4_ASAP7_75t_L g580 ( .A(n_468), .Y(n_580) );
BUFx6f_ASAP7_75t_L g600 ( .A(n_468), .Y(n_600) );
AND2x4_ASAP7_75t_L g611 ( .A(n_468), .B(n_579), .Y(n_611) );
AND2x2_ASAP7_75t_L g617 ( .A(n_468), .B(n_541), .Y(n_617) );
NOR2x1_ASAP7_75t_SL g690 ( .A(n_468), .B(n_552), .Y(n_690) );
OR2x6_ASAP7_75t_L g468 ( .A(n_469), .B(n_470), .Y(n_468) );
INVxp67_ASAP7_75t_L g491 ( .A(n_474), .Y(n_491) );
INVx2_ASAP7_75t_L g551 ( .A(n_474), .Y(n_551) );
INVx2_ASAP7_75t_L g583 ( .A(n_477), .Y(n_583) );
HB1xp67_ASAP7_75t_L g597 ( .A(n_477), .Y(n_597) );
INVx1_ASAP7_75t_L g608 ( .A(n_477), .Y(n_608) );
HB1xp67_ASAP7_75t_L g620 ( .A(n_477), .Y(n_620) );
AND2x2_ASAP7_75t_L g652 ( .A(n_477), .B(n_552), .Y(n_652) );
INVx1_ASAP7_75t_L g678 ( .A(n_477), .Y(n_678) );
AND2x2_ASAP7_75t_L g740 ( .A(n_477), .B(n_568), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_479), .B(n_480), .Y(n_478) );
AND2x2_ASAP7_75t_L g485 ( .A(n_486), .B(n_504), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
AND2x2_ASAP7_75t_L g633 ( .A(n_487), .B(n_572), .Y(n_633) );
INVx2_ASAP7_75t_L g675 ( .A(n_487), .Y(n_675) );
AND2x2_ASAP7_75t_L g777 ( .A(n_487), .B(n_504), .Y(n_777) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_488), .B(n_527), .Y(n_571) );
INVx2_ASAP7_75t_L g592 ( .A(n_488), .Y(n_592) );
AND2x4_ASAP7_75t_L g614 ( .A(n_488), .B(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g649 ( .A(n_488), .Y(n_649) );
AND2x2_ASAP7_75t_L g773 ( .A(n_488), .B(n_530), .Y(n_773) );
OR2x2_ASAP7_75t_L g488 ( .A(n_489), .B(n_497), .Y(n_488) );
AO21x2_ASAP7_75t_L g505 ( .A1(n_496), .A2(n_506), .B(n_512), .Y(n_505) );
AO21x2_ASAP7_75t_L g527 ( .A1(n_496), .A2(n_506), .B(n_512), .Y(n_527) );
OAI22xp5_ASAP7_75t_L g497 ( .A1(n_498), .A2(n_501), .B1(n_502), .B2(n_503), .Y(n_497) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g747 ( .A(n_504), .Y(n_747) );
AND2x2_ASAP7_75t_L g504 ( .A(n_505), .B(n_513), .Y(n_504) );
NOR2xp67_ASAP7_75t_L g622 ( .A(n_505), .B(n_592), .Y(n_622) );
AND2x2_ASAP7_75t_L g627 ( .A(n_505), .B(n_592), .Y(n_627) );
INVx2_ASAP7_75t_L g640 ( .A(n_505), .Y(n_640) );
NOR2x1_ASAP7_75t_L g705 ( .A(n_505), .B(n_706), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_507), .B(n_508), .Y(n_506) );
AND2x4_ASAP7_75t_L g613 ( .A(n_513), .B(n_526), .Y(n_613) );
AND2x2_ASAP7_75t_L g628 ( .A(n_513), .B(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g683 ( .A(n_513), .Y(n_683) );
INVx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_514), .B(n_530), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_514), .B(n_527), .Y(n_681) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_516), .B(n_522), .Y(n_515) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVxp33_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
NAND2x1p5_ASAP7_75t_L g525 ( .A(n_526), .B(n_528), .Y(n_525) );
INVx3_ASAP7_75t_L g589 ( .A(n_526), .Y(n_589) );
INVx3_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
HB1xp67_ASAP7_75t_L g587 ( .A(n_527), .Y(n_587) );
AND2x2_ASAP7_75t_L g701 ( .A(n_527), .B(n_702), .Y(n_701) );
INVx3_ASAP7_75t_L g644 ( .A(n_528), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_528), .B(n_683), .Y(n_724) );
BUFx3_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
AND2x2_ASAP7_75t_L g591 ( .A(n_529), .B(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
AND2x4_ASAP7_75t_L g572 ( .A(n_530), .B(n_573), .Y(n_572) );
INVx2_ASAP7_75t_L g615 ( .A(n_530), .Y(n_615) );
INVxp67_ASAP7_75t_L g629 ( .A(n_530), .Y(n_629) );
HB1xp67_ASAP7_75t_L g702 ( .A(n_530), .Y(n_702) );
INVx1_ASAP7_75t_L g706 ( .A(n_530), .Y(n_706) );
INVx1_ASAP7_75t_L g684 ( .A(n_536), .Y(n_684) );
NOR2x1_ASAP7_75t_L g536 ( .A(n_537), .B(n_539), .Y(n_536) );
NOR2x1_ASAP7_75t_L g661 ( .A(n_537), .B(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
AND2x2_ASAP7_75t_L g726 ( .A(n_538), .B(n_567), .Y(n_726) );
OR2x2_ASAP7_75t_L g778 ( .A(n_539), .B(n_779), .Y(n_778) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g677 ( .A(n_540), .B(n_678), .Y(n_677) );
AND2x2_ASAP7_75t_L g713 ( .A(n_540), .B(n_600), .Y(n_713) );
AND2x2_ASAP7_75t_L g540 ( .A(n_541), .B(n_552), .Y(n_540) );
AND2x4_ASAP7_75t_L g567 ( .A(n_541), .B(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g579 ( .A(n_541), .Y(n_579) );
INVx2_ASAP7_75t_L g596 ( .A(n_541), .Y(n_596) );
HB1xp67_ASAP7_75t_L g722 ( .A(n_541), .Y(n_722) );
AND2x2_ASAP7_75t_L g541 ( .A(n_542), .B(n_547), .Y(n_541) );
NOR3xp33_ASAP7_75t_L g543 ( .A(n_544), .B(n_545), .C(n_546), .Y(n_543) );
INVx3_ASAP7_75t_L g568 ( .A(n_552), .Y(n_568) );
INVx2_ASAP7_75t_L g662 ( .A(n_552), .Y(n_662) );
AND2x4_ASAP7_75t_L g552 ( .A(n_553), .B(n_554), .Y(n_552) );
OAI21xp5_ASAP7_75t_L g554 ( .A1(n_555), .A2(n_558), .B(n_563), .Y(n_554) );
OAI22xp5_ASAP7_75t_L g558 ( .A1(n_559), .A2(n_560), .B1(n_561), .B2(n_562), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_565), .B(n_569), .Y(n_564) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
NOR2xp33_ASAP7_75t_L g659 ( .A(n_566), .B(n_642), .Y(n_659) );
NOR2x1_ASAP7_75t_L g751 ( .A(n_566), .B(n_580), .Y(n_751) );
INVx4_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_567), .B(n_642), .Y(n_728) );
AND2x2_ASAP7_75t_L g595 ( .A(n_568), .B(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g609 ( .A(n_568), .Y(n_609) );
AOI22xp5_ASAP7_75t_SL g657 ( .A1(n_569), .A2(n_658), .B1(n_659), .B2(n_660), .Y(n_657) );
AND2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_572), .Y(n_569) );
NAND2x1p5_ASAP7_75t_L g654 ( .A(n_570), .B(n_628), .Y(n_654) );
INVx2_ASAP7_75t_SL g570 ( .A(n_571), .Y(n_570) );
OR2x2_ASAP7_75t_L g762 ( .A(n_571), .B(n_603), .Y(n_762) );
AND2x2_ASAP7_75t_L g585 ( .A(n_572), .B(n_586), .Y(n_585) );
AND2x4_ASAP7_75t_L g621 ( .A(n_572), .B(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g764 ( .A(n_572), .B(n_675), .Y(n_764) );
INVx2_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
AND2x4_ASAP7_75t_L g639 ( .A(n_574), .B(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g665 ( .A(n_574), .Y(n_665) );
AND2x2_ASAP7_75t_L g700 ( .A(n_574), .B(n_592), .Y(n_700) );
OAI221xp5_ASAP7_75t_L g575 ( .A1(n_576), .A2(n_584), .B1(n_588), .B2(n_593), .C(n_598), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_581), .Y(n_577) );
INVx1_ASAP7_75t_L g656 ( .A(n_578), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_578), .B(n_652), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_578), .B(n_740), .Y(n_739) );
AND2x4_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .Y(n_578) );
NOR2xp67_ASAP7_75t_SL g624 ( .A(n_580), .B(n_625), .Y(n_624) );
HB1xp67_ASAP7_75t_L g637 ( .A(n_580), .Y(n_637) );
AND2x4_ASAP7_75t_SL g721 ( .A(n_580), .B(n_722), .Y(n_721) );
OR2x2_ASAP7_75t_L g768 ( .A(n_580), .B(n_769), .Y(n_768) );
HB1xp67_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx3_ASAP7_75t_L g642 ( .A(n_582), .Y(n_642) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
HB1xp67_ASAP7_75t_L g779 ( .A(n_583), .Y(n_779) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
AOI221x1_ASAP7_75t_L g732 ( .A1(n_585), .A2(n_733), .B1(n_735), .B2(n_736), .C(n_738), .Y(n_732) );
AND2x2_ASAP7_75t_L g658 ( .A(n_586), .B(n_614), .Y(n_658) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
OR2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
AND2x2_ASAP7_75t_L g601 ( .A(n_589), .B(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_589), .B(n_591), .Y(n_775) );
INVx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
INVx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_595), .B(n_597), .Y(n_594) );
AND2x2_ASAP7_75t_SL g599 ( .A(n_595), .B(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_595), .B(n_608), .Y(n_625) );
INVx2_ASAP7_75t_L g632 ( .A(n_595), .Y(n_632) );
INVx1_ASAP7_75t_L g694 ( .A(n_596), .Y(n_694) );
BUFx2_ASAP7_75t_L g714 ( .A(n_597), .Y(n_714) );
NAND2xp33_ASAP7_75t_SL g598 ( .A(n_599), .B(n_601), .Y(n_598) );
OR2x6_ASAP7_75t_L g631 ( .A(n_600), .B(n_632), .Y(n_631) );
AND2x2_ASAP7_75t_L g760 ( .A(n_600), .B(n_652), .Y(n_760) );
INVx2_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_605), .B(n_623), .Y(n_604) );
AOI22xp5_ASAP7_75t_L g605 ( .A1(n_606), .A2(n_612), .B1(n_616), .B2(n_621), .Y(n_605) );
NOR2xp33_ASAP7_75t_L g606 ( .A(n_607), .B(n_610), .Y(n_606) );
AND2x2_ASAP7_75t_SL g669 ( .A(n_607), .B(n_611), .Y(n_669) );
AND2x4_ASAP7_75t_L g735 ( .A(n_607), .B(n_693), .Y(n_735) );
AND2x4_ASAP7_75t_SL g607 ( .A(n_608), .B(n_609), .Y(n_607) );
HB1xp67_ASAP7_75t_L g750 ( .A(n_608), .Y(n_750) );
INVx2_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
NOR2xp33_ASAP7_75t_L g650 ( .A(n_611), .B(n_651), .Y(n_650) );
HB1xp67_ASAP7_75t_L g703 ( .A(n_611), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_611), .B(n_642), .Y(n_734) );
AND2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
AND2x2_ASAP7_75t_L g755 ( .A(n_613), .B(n_674), .Y(n_755) );
INVx3_ASAP7_75t_L g666 ( .A(n_614), .Y(n_666) );
AND2x2_ASAP7_75t_L g687 ( .A(n_614), .B(n_639), .Y(n_687) );
NAND2x1_ASAP7_75t_SL g758 ( .A(n_614), .B(n_665), .Y(n_758) );
AND2x2_ASAP7_75t_L g616 ( .A(n_617), .B(n_618), .Y(n_616) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
AOI22xp5_ASAP7_75t_L g623 ( .A1(n_624), .A2(n_626), .B1(n_630), .B2(n_633), .Y(n_623) );
BUFx2_ASAP7_75t_L g679 ( .A(n_625), .Y(n_679) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_626), .A2(n_717), .B1(n_726), .B2(n_727), .Y(n_725) );
AND2x2_ASAP7_75t_L g626 ( .A(n_627), .B(n_628), .Y(n_626) );
NAND2x1p5_ASAP7_75t_L g682 ( .A(n_627), .B(n_683), .Y(n_682) );
AND2x2_ASAP7_75t_L g647 ( .A(n_628), .B(n_648), .Y(n_647) );
INVx2_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
NAND3xp33_ASAP7_75t_L g711 ( .A(n_632), .B(n_712), .C(n_714), .Y(n_711) );
INVx1_ASAP7_75t_L g667 ( .A(n_633), .Y(n_667) );
AOI211x1_ASAP7_75t_L g634 ( .A1(n_635), .A2(n_643), .B(n_645), .C(n_663), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_637), .B(n_638), .Y(n_636) );
NAND2xp5_ASAP7_75t_SL g745 ( .A(n_638), .B(n_726), .Y(n_745) );
AND2x2_ASAP7_75t_L g638 ( .A(n_639), .B(n_641), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_639), .B(n_674), .Y(n_673) );
AND2x2_ASAP7_75t_L g717 ( .A(n_639), .B(n_675), .Y(n_717) );
AND2x2_ASAP7_75t_L g772 ( .A(n_639), .B(n_773), .Y(n_772) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g695 ( .A(n_642), .Y(n_695) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
OR2x2_ASAP7_75t_L g737 ( .A(n_644), .B(n_682), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_646), .B(n_657), .Y(n_645) );
AOI22xp5_ASAP7_75t_SL g646 ( .A1(n_647), .A2(n_650), .B1(n_653), .B2(n_655), .Y(n_646) );
BUFx2_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
AND2x2_ASAP7_75t_L g710 ( .A(n_649), .B(n_705), .Y(n_710) );
INVx1_ASAP7_75t_SL g752 ( .A(n_649), .Y(n_752) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
AND2x2_ASAP7_75t_SL g720 ( .A(n_652), .B(n_721), .Y(n_720) );
INVx3_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVxp67_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
HB1xp67_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
AND2x2_ASAP7_75t_L g756 ( .A(n_661), .B(n_678), .Y(n_756) );
AOI21xp5_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_667), .B(n_668), .Y(n_663) );
OR2x2_ASAP7_75t_L g664 ( .A(n_665), .B(n_666), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_665), .B(n_710), .Y(n_709) );
OR2x2_ASAP7_75t_L g680 ( .A(n_666), .B(n_681), .Y(n_680) );
INVx1_ASAP7_75t_SL g668 ( .A(n_669), .Y(n_668) );
INVxp67_ASAP7_75t_SL g825 ( .A(n_670), .Y(n_825) );
NAND3x1_ASAP7_75t_L g670 ( .A(n_671), .B(n_707), .C(n_715), .Y(n_670) );
NAND4xp25_ASAP7_75t_L g781 ( .A(n_671), .B(n_707), .C(n_715), .D(n_782), .Y(n_781) );
NOR2x1_ASAP7_75t_L g671 ( .A(n_672), .B(n_685), .Y(n_671) );
OAI222xp33_ASAP7_75t_L g672 ( .A1(n_673), .A2(n_676), .B1(n_679), .B2(n_680), .C1(n_682), .C2(n_684), .Y(n_672) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
OAI21xp5_ASAP7_75t_SL g759 ( .A1(n_677), .A2(n_760), .B(n_761), .Y(n_759) );
NAND2xp5_ASAP7_75t_SL g742 ( .A(n_678), .B(n_693), .Y(n_742) );
OAI22xp5_ASAP7_75t_L g738 ( .A1(n_681), .A2(n_739), .B1(n_741), .B2(n_742), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_686), .B(n_696), .Y(n_685) );
NAND2xp5_ASAP7_75t_SL g686 ( .A(n_687), .B(n_688), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_689), .B(n_691), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_689), .B(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_692), .B(n_695), .Y(n_691) );
INVx2_ASAP7_75t_SL g692 ( .A(n_693), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_693), .B(n_695), .Y(n_698) );
INVx2_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
AOI22xp5_ASAP7_75t_L g696 ( .A1(n_697), .A2(n_699), .B1(n_703), .B2(n_704), .Y(n_696) );
AND2x4_ASAP7_75t_L g699 ( .A(n_700), .B(n_701), .Y(n_699) );
AND2x2_ASAP7_75t_L g704 ( .A(n_700), .B(n_705), .Y(n_704) );
NAND2xp5_ASAP7_75t_SL g707 ( .A(n_708), .B(n_711), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g741 ( .A(n_710), .Y(n_741) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
AND2x2_ASAP7_75t_L g715 ( .A(n_716), .B(n_725), .Y(n_715) );
AOI22xp5_ASAP7_75t_SL g716 ( .A1(n_717), .A2(n_718), .B1(n_720), .B2(n_723), .Y(n_716) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVxp67_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
NAND2xp33_ASAP7_75t_L g730 ( .A(n_729), .B(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g824 ( .A(n_731), .Y(n_824) );
NAND3x1_ASAP7_75t_L g731 ( .A(n_732), .B(n_743), .C(n_763), .Y(n_731) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
AOI22xp5_ASAP7_75t_L g754 ( .A1(n_735), .A2(n_755), .B1(n_756), .B2(n_757), .Y(n_754) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_SL g769 ( .A(n_740), .Y(n_769) );
NOR2x1_ASAP7_75t_L g743 ( .A(n_744), .B(n_753), .Y(n_743) );
AOI21xp5_ASAP7_75t_SL g744 ( .A1(n_745), .A2(n_746), .B(n_752), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_747), .B(n_748), .Y(n_746) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_750), .B(n_751), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_754), .B(n_759), .Y(n_753) );
INVx2_ASAP7_75t_SL g757 ( .A(n_758), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_758), .B(n_771), .Y(n_770) );
INVx1_ASAP7_75t_SL g761 ( .A(n_762), .Y(n_761) );
AOI221xp5_ASAP7_75t_L g763 ( .A1(n_764), .A2(n_765), .B1(n_767), .B2(n_770), .C(n_774), .Y(n_763) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
INVxp67_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
INVx2_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
AOI21xp5_ASAP7_75t_L g774 ( .A1(n_775), .A2(n_776), .B(n_778), .Y(n_774) );
INVx1_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
NOR2xp33_ASAP7_75t_L g782 ( .A(n_783), .B(n_784), .Y(n_782) );
INVxp67_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
NOR3xp33_ASAP7_75t_L g826 ( .A(n_786), .B(n_827), .C(n_828), .Y(n_826) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_787), .B(n_794), .Y(n_786) );
INVxp33_ASAP7_75t_L g801 ( .A(n_787), .Y(n_801) );
NOR2xp33_ASAP7_75t_L g787 ( .A(n_788), .B(n_790), .Y(n_787) );
CKINVDCx8_ASAP7_75t_R g788 ( .A(n_789), .Y(n_788) );
NOR2xp33_ASAP7_75t_L g790 ( .A(n_791), .B(n_792), .Y(n_790) );
CKINVDCx5p33_ASAP7_75t_R g798 ( .A(n_793), .Y(n_798) );
OAI32xp33_ASAP7_75t_L g799 ( .A1(n_793), .A2(n_800), .A3(n_801), .B1(n_802), .B2(n_833), .Y(n_799) );
CKINVDCx20_ASAP7_75t_R g800 ( .A(n_794), .Y(n_800) );
INVx1_ASAP7_75t_SL g795 ( .A(n_796), .Y(n_795) );
BUFx2_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
NOR2x1_ASAP7_75t_R g803 ( .A(n_797), .B(n_804), .Y(n_803) );
NOR2xp33_ASAP7_75t_L g806 ( .A(n_800), .B(n_807), .Y(n_806) );
INVx1_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
HB1xp67_ASAP7_75t_L g811 ( .A(n_804), .Y(n_811) );
AOI21xp5_ASAP7_75t_L g805 ( .A1(n_806), .A2(n_812), .B(n_826), .Y(n_805) );
HB1xp67_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
CKINVDCx5p33_ASAP7_75t_R g808 ( .A(n_809), .Y(n_808) );
BUFx3_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
CKINVDCx20_ASAP7_75t_R g810 ( .A(n_811), .Y(n_810) );
AOI22xp33_ASAP7_75t_SL g813 ( .A1(n_814), .A2(n_815), .B1(n_821), .B2(n_822), .Y(n_813) );
INVx1_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
OAI22xp5_ASAP7_75t_L g815 ( .A1(n_816), .A2(n_817), .B1(n_819), .B2(n_820), .Y(n_815) );
INVx1_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
CKINVDCx5p33_ASAP7_75t_R g819 ( .A(n_820), .Y(n_819) );
INVx1_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
AND3x2_ASAP7_75t_L g822 ( .A(n_823), .B(n_824), .C(n_825), .Y(n_822) );
endmodule