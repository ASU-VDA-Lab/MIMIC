module fake_jpeg_111_n_110 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_110);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_110;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx16f_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_37),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_41),
.B(n_43),
.Y(n_45)
);

INVxp67_ASAP7_75t_SL g42 ( 
.A(n_37),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_44),
.Y(n_50)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

BUFx4f_ASAP7_75t_SL g44 ( 
.A(n_33),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_43),
.A2(n_34),
.B1(n_31),
.B2(n_28),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g54 ( 
.A1(n_46),
.A2(n_49),
.B(n_44),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_41),
.A2(n_36),
.B1(n_33),
.B2(n_29),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_47),
.A2(n_48),
.B1(n_38),
.B2(n_3),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_41),
.A2(n_34),
.B1(n_28),
.B2(n_35),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_39),
.A2(n_32),
.B1(n_36),
.B2(n_30),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_30),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_27),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_62),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_44),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_58),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_52),
.Y(n_56)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_57),
.B(n_59),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_0),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_1),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_60),
.B(n_61),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_45),
.B(n_1),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_26),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_23),
.Y(n_68)
);

AOI32xp33_ASAP7_75t_L g65 ( 
.A1(n_63),
.A2(n_47),
.A3(n_38),
.B1(n_5),
.B2(n_6),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_2),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_68),
.B(n_69),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_54),
.C(n_62),
.Y(n_69)
);

O2A1O1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_54),
.A2(n_53),
.B(n_3),
.C(n_5),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_70),
.B(n_7),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_53),
.C(n_22),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_74),
.C(n_66),
.Y(n_83)
);

AND2x4_ASAP7_75t_L g74 ( 
.A(n_54),
.B(n_20),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_74),
.Y(n_76)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_71),
.Y(n_75)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_75),
.Y(n_95)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_19),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_82),
.C(n_11),
.Y(n_94)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_74),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_79),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_66),
.A2(n_2),
.B1(n_6),
.B2(n_7),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_81),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_18),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_83),
.B(n_14),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_84),
.B(n_85),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_SL g86 ( 
.A(n_80),
.B(n_73),
.Y(n_86)
);

OA21x2_ASAP7_75t_SL g99 ( 
.A1(n_86),
.A2(n_89),
.B(n_91),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_8),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_92),
.B(n_94),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_10),
.Y(n_93)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_93),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_95),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_96),
.B(n_100),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_87),
.A2(n_76),
.B(n_79),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_97),
.A2(n_90),
.B1(n_92),
.B2(n_88),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_101),
.B(n_97),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_103),
.B(n_102),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_104),
.B(n_99),
.Y(n_105)
);

O2A1O1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_105),
.A2(n_86),
.B(n_98),
.C(n_100),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_106),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_94),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_13),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_109),
.B(n_11),
.Y(n_110)
);


endmodule