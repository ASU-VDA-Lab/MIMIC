module fake_jpeg_23660_n_183 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_183);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_183;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_31),
.A2(n_14),
.B1(n_18),
.B2(n_15),
.Y(n_55)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx3_ASAP7_75t_SL g40 ( 
.A(n_33),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_20),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_38),
.Y(n_41)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_25),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_43),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_31),
.A2(n_21),
.B1(n_17),
.B2(n_25),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_43),
.A2(n_50),
.B1(n_19),
.B2(n_16),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_26),
.Y(n_44)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_26),
.Y(n_45)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_20),
.Y(n_46)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_38),
.A2(n_17),
.B1(n_21),
.B2(n_25),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_37),
.A2(n_21),
.B1(n_17),
.B2(n_23),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_51),
.A2(n_50),
.B1(n_55),
.B2(n_14),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_32),
.B(n_18),
.Y(n_53)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_55),
.A2(n_28),
.B1(n_38),
.B2(n_19),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_41),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_58),
.B(n_63),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_59),
.A2(n_70),
.B1(n_40),
.B2(n_47),
.Y(n_83)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_61),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_32),
.Y(n_62)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_62),
.Y(n_87)
);

BUFx2_ASAP7_75t_SL g64 ( 
.A(n_54),
.Y(n_64)
);

INVxp33_ASAP7_75t_L g92 ( 
.A(n_64),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_65),
.B(n_68),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_51),
.A2(n_28),
.B1(n_16),
.B2(n_15),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_66),
.A2(n_47),
.B1(n_49),
.B2(n_52),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g68 ( 
.A(n_45),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_72),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_41),
.B(n_27),
.Y(n_73)
);

BUFx24_ASAP7_75t_SL g76 ( 
.A(n_73),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_58),
.A2(n_39),
.B(n_38),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_74),
.B(n_86),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_61),
.B(n_40),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_80),
.Y(n_95)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_63),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_84),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_83),
.A2(n_88),
.B1(n_89),
.B2(n_82),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_63),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_39),
.Y(n_86)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_83),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_57),
.A2(n_56),
.B(n_65),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_90),
.B(n_91),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_56),
.B(n_30),
.Y(n_91)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_92),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_107),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_96),
.A2(n_101),
.B1(n_104),
.B2(n_105),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_97),
.B(n_102),
.Y(n_113)
);

AOI21xp33_ASAP7_75t_L g99 ( 
.A1(n_81),
.A2(n_69),
.B(n_71),
.Y(n_99)
);

NAND3xp33_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_79),
.C(n_76),
.Y(n_112)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_80),
.B(n_69),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_103),
.B(n_106),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_84),
.A2(n_40),
.B1(n_71),
.B2(n_49),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_77),
.A2(n_40),
.B1(n_49),
.B2(n_52),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_48),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_85),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_81),
.A2(n_48),
.B1(n_27),
.B2(n_19),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_108),
.Y(n_116)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_109),
.B(n_79),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_102),
.B(n_91),
.Y(n_110)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_110),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_74),
.C(n_87),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_111),
.B(n_107),
.C(n_108),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_112),
.A2(n_117),
.B1(n_120),
.B2(n_105),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_98),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_114),
.B(n_93),
.Y(n_128)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_118),
.B(n_119),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_109),
.A2(n_88),
.B(n_27),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_96),
.A2(n_48),
.B1(n_67),
.B2(n_36),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_104),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_123),
.Y(n_130)
);

AOI322xp5_ASAP7_75t_L g124 ( 
.A1(n_98),
.A2(n_36),
.A3(n_33),
.B1(n_67),
.B2(n_27),
.C1(n_24),
.C2(n_75),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_124),
.B(n_125),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_94),
.B(n_75),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_126),
.B(n_128),
.C(n_134),
.Y(n_139)
);

XOR2x2_ASAP7_75t_L g127 ( 
.A(n_114),
.B(n_125),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_127),
.A2(n_0),
.B(n_1),
.Y(n_145)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_122),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_129),
.B(n_131),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_123),
.A2(n_97),
.B1(n_24),
.B2(n_27),
.Y(n_133)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_133),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_75),
.C(n_24),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_13),
.C(n_12),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_136),
.B(n_1),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_116),
.A2(n_118),
.B1(n_111),
.B2(n_119),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_137),
.A2(n_116),
.B1(n_120),
.B2(n_113),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_140),
.A2(n_142),
.B1(n_2),
.B2(n_3),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_130),
.A2(n_115),
.B(n_121),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_134),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_143),
.B(n_144),
.Y(n_150)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_132),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_145),
.B(n_127),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_136),
.B(n_13),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_146),
.B(n_148),
.Y(n_156)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_137),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_149),
.B(n_126),
.C(n_138),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_151),
.B(n_153),
.Y(n_163)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_152),
.Y(n_160)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_142),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_139),
.B(n_128),
.C(n_135),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_154),
.B(n_157),
.C(n_143),
.Y(n_159)
);

NOR3xp33_ASAP7_75t_SL g155 ( 
.A(n_145),
.B(n_141),
.C(n_144),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_155),
.B(n_5),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_139),
.B(n_135),
.C(n_3),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_158),
.A2(n_147),
.B1(n_149),
.B2(n_4),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_159),
.B(n_154),
.C(n_152),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_161),
.B(n_165),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_150),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_162),
.B(n_164),
.Y(n_169)
);

OAI22xp33_ASAP7_75t_L g165 ( 
.A1(n_155),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_166),
.B(n_171),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_159),
.B(n_156),
.C(n_7),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_167),
.B(n_168),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_163),
.B(n_6),
.C(n_9),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_162),
.B(n_6),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_169),
.B(n_164),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_174),
.B(n_175),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_170),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_172),
.B(n_160),
.C(n_165),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_176),
.B(n_177),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_173),
.B(n_10),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_178),
.B(n_11),
.Y(n_180)
);

INVxp33_ASAP7_75t_L g181 ( 
.A(n_180),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_181),
.B(n_179),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_182),
.B(n_11),
.Y(n_183)
);


endmodule