module fake_jpeg_8872_n_250 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_250);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_250;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

HB1xp67_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_16),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_16),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_37),
.B(n_41),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_20),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_44),
.B(n_37),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_28),
.A2(n_20),
.B1(n_13),
.B2(n_23),
.Y(n_45)
);

OAI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_45),
.A2(n_28),
.B1(n_15),
.B2(n_23),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_28),
.B(n_24),
.Y(n_47)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_52),
.Y(n_56)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_55),
.B(n_58),
.Y(n_76)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_38),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_51),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_59),
.B(n_60),
.Y(n_88)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_24),
.Y(n_61)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

INVx3_ASAP7_75t_SL g62 ( 
.A(n_39),
.Y(n_62)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

NOR2x1_ASAP7_75t_R g64 ( 
.A(n_41),
.B(n_36),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_67),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_65),
.A2(n_70),
.B1(n_34),
.B2(n_50),
.Y(n_71)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_69),
.Y(n_79)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_71),
.A2(n_73),
.B1(n_78),
.B2(n_84),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_66),
.A2(n_32),
.B1(n_34),
.B2(n_46),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_77),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_64),
.A2(n_32),
.B1(n_34),
.B2(n_13),
.Y(n_78)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_82),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_55),
.A2(n_52),
.B1(n_49),
.B2(n_42),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_63),
.A2(n_53),
.B1(n_30),
.B2(n_31),
.Y(n_85)
);

O2A1O1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_85),
.A2(n_48),
.B(n_57),
.C(n_53),
.Y(n_99)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_86),
.Y(n_96)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_63),
.A2(n_36),
.B(n_30),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_89),
.B(n_67),
.C(n_56),
.Y(n_92)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_90),
.B(n_98),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_92),
.A2(n_107),
.B(n_77),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_80),
.A2(n_60),
.B1(n_27),
.B2(n_30),
.Y(n_93)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_80),
.A2(n_31),
.B1(n_43),
.B2(n_70),
.Y(n_94)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_94),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_89),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_95),
.B(n_102),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_80),
.A2(n_31),
.B1(n_43),
.B2(n_68),
.Y(n_97)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_97),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_88),
.Y(n_98)
);

OAI32xp33_ASAP7_75t_L g125 ( 
.A1(n_99),
.A2(n_86),
.A3(n_33),
.B1(n_14),
.B2(n_18),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_79),
.A2(n_32),
.B1(n_15),
.B2(n_26),
.Y(n_101)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_101),
.Y(n_128)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_74),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_105),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_29),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_106),
.B(n_108),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_83),
.B(n_0),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_81),
.B(n_29),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_106),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_109),
.B(n_116),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_108),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_112),
.B(n_115),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_83),
.C(n_81),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_114),
.B(n_119),
.C(n_122),
.Y(n_142)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_104),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_90),
.B(n_21),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_118),
.B(n_21),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_92),
.B(n_82),
.C(n_74),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_120),
.B(n_97),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_74),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_121),
.B(n_127),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_94),
.B(n_29),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_125),
.A2(n_111),
.B1(n_126),
.B2(n_124),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_75),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_129),
.B(n_136),
.Y(n_150)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_123),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_131),
.A2(n_132),
.B1(n_139),
.B2(n_145),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_111),
.A2(n_102),
.B1(n_100),
.B2(n_93),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_123),
.Y(n_135)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_135),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_107),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_120),
.B(n_99),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_137),
.B(n_143),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_126),
.A2(n_103),
.B1(n_91),
.B2(n_75),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_138),
.A2(n_141),
.B(n_147),
.Y(n_167)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_113),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_110),
.A2(n_91),
.B1(n_103),
.B2(n_72),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_140),
.A2(n_122),
.B1(n_121),
.B2(n_117),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_110),
.A2(n_104),
.B(n_96),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_119),
.B(n_29),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_113),
.Y(n_144)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_144),
.Y(n_152)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_118),
.Y(n_146)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_146),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_127),
.A2(n_124),
.B(n_112),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_148),
.Y(n_157)
);

HB1xp67_ASAP7_75t_L g149 ( 
.A(n_115),
.Y(n_149)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_149),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_133),
.B(n_128),
.Y(n_154)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_154),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_133),
.B(n_128),
.Y(n_155)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_155),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_130),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_156),
.B(n_161),
.Y(n_179)
);

AO21x2_ASAP7_75t_L g159 ( 
.A1(n_141),
.A2(n_125),
.B(n_116),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_159),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_134),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_162),
.A2(n_166),
.B1(n_33),
.B2(n_25),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_147),
.B(n_117),
.Y(n_163)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_163),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_140),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_165),
.B(n_168),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_137),
.A2(n_72),
.B1(n_26),
.B2(n_54),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_145),
.Y(n_168)
);

HB1xp67_ASAP7_75t_L g169 ( 
.A(n_138),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_169),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_150),
.B(n_142),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_170),
.B(n_178),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_164),
.A2(n_142),
.B1(n_129),
.B2(n_136),
.Y(n_171)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_171),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_159),
.A2(n_143),
.B1(n_25),
.B2(n_19),
.Y(n_172)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_172),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_150),
.B(n_29),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_176),
.B(n_184),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_153),
.B(n_33),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_180),
.A2(n_151),
.B1(n_152),
.B2(n_159),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_159),
.A2(n_19),
.B1(n_18),
.B2(n_25),
.Y(n_181)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_181),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_153),
.B(n_19),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_163),
.B(n_18),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_185),
.B(n_162),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_159),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_186),
.B(n_167),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_170),
.B(n_167),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_187),
.B(n_184),
.Y(n_205)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_192),
.Y(n_214)
);

A2O1A1Ixp33_ASAP7_75t_L g193 ( 
.A1(n_175),
.A2(n_173),
.B(n_155),
.C(n_154),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_193),
.A2(n_157),
.B1(n_1),
.B2(n_2),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_194),
.B(n_199),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g195 ( 
.A(n_183),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_195),
.B(n_197),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_196),
.B(n_198),
.Y(n_210)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_179),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_185),
.B(n_160),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_178),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_182),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_200),
.A2(n_177),
.B1(n_174),
.B2(n_160),
.Y(n_203)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_203),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_190),
.A2(n_193),
.B1(n_183),
.B2(n_191),
.Y(n_204)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_204),
.Y(n_222)
);

MAJx2_ASAP7_75t_L g220 ( 
.A(n_205),
.B(n_2),
.C(n_3),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_188),
.A2(n_158),
.B(n_166),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_206),
.A2(n_209),
.B(n_3),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_187),
.B(n_158),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_208),
.B(n_12),
.C(n_5),
.Y(n_221)
);

OAI221xp5_ASAP7_75t_L g211 ( 
.A1(n_200),
.A2(n_201),
.B1(n_189),
.B2(n_195),
.C(n_4),
.Y(n_211)
);

OR2x2_ASAP7_75t_L g216 ( 
.A(n_211),
.B(n_212),
.Y(n_216)
);

NAND2x1p5_ASAP7_75t_L g212 ( 
.A(n_201),
.B(n_7),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_197),
.B(n_7),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_213),
.B(n_0),
.Y(n_215)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_215),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_202),
.B(n_2),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_218),
.B(n_224),
.Y(n_228)
);

INVx11_ASAP7_75t_L g219 ( 
.A(n_212),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_219),
.A2(n_203),
.B1(n_8),
.B2(n_9),
.Y(n_230)
);

NOR2x1_ASAP7_75t_SL g227 ( 
.A(n_220),
.B(n_6),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_221),
.B(n_223),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_205),
.B(n_3),
.C(n_5),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_207),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_225),
.B(n_210),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_225),
.B(n_208),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_226),
.B(n_219),
.Y(n_236)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_227),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_216),
.B(n_214),
.Y(n_229)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_229),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_230),
.A2(n_232),
.B(n_217),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_231),
.B(n_216),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_234),
.B(n_239),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_236),
.B(n_237),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_228),
.B(n_222),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_238),
.A2(n_229),
.B(n_233),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_242),
.A2(n_243),
.B(n_241),
.Y(n_244)
);

NOR2xp67_ASAP7_75t_L g243 ( 
.A(n_235),
.B(n_220),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_244),
.B(n_245),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_240),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_246),
.B(n_6),
.C(n_9),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_247),
.B(n_11),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_248),
.B(n_11),
.C(n_12),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_249),
.B(n_11),
.Y(n_250)
);


endmodule