module fake_jpeg_11503_n_176 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_176);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_176;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx6f_ASAP7_75t_SL g52 ( 
.A(n_18),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_11),
.Y(n_54)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_1),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_12),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_31),
.Y(n_59)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_24),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_6),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_16),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_37),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_16),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_14),
.B(n_22),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_43),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_47),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_11),
.B(n_1),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_73),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_0),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_80),
.B(n_83),
.Y(n_85)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_82),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_0),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_84),
.B(n_56),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_84),
.B(n_57),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_92),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_79),
.A2(n_53),
.B1(n_52),
.B2(n_50),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_87),
.A2(n_60),
.B1(n_68),
.B2(n_62),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_82),
.A2(n_78),
.B1(n_81),
.B2(n_66),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_89),
.A2(n_97),
.B1(n_60),
.B2(n_55),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_59),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_75),
.B(n_66),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_94),
.B(n_72),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_81),
.A2(n_49),
.B1(n_67),
.B2(n_50),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_56),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_99),
.B(n_2),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_100),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_86),
.A2(n_49),
.B1(n_67),
.B2(n_57),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_101),
.A2(n_103),
.B1(n_8),
.B2(n_9),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_99),
.B(n_71),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_102),
.B(n_105),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_90),
.A2(n_49),
.B1(n_67),
.B2(n_71),
.Y(n_103)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_106),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_107),
.A2(n_109),
.B1(n_6),
.B2(n_7),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_26),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_90),
.A2(n_51),
.B1(n_55),
.B2(n_65),
.Y(n_109)
);

A2O1A1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_88),
.A2(n_70),
.B(n_3),
.C(n_4),
.Y(n_110)
);

NOR2xp67_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_5),
.Y(n_125)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_111),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_91),
.A2(n_65),
.B1(n_3),
.B2(n_4),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_112),
.B(n_10),
.C(n_12),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_113),
.B(n_117),
.Y(n_123)
);

NOR2x1_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_85),
.Y(n_114)
);

NOR2x1_ASAP7_75t_L g128 ( 
.A(n_114),
.B(n_103),
.Y(n_128)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

INVx11_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_116),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_2),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_95),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_118),
.B(n_119),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_93),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_88),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_120),
.B(n_13),
.Y(n_141)
);

OAI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_109),
.A2(n_107),
.B1(n_101),
.B2(n_112),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_122),
.A2(n_126),
.B1(n_15),
.B2(n_20),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_104),
.B(n_5),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_124),
.B(n_128),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_125),
.B(n_127),
.Y(n_148)
);

NOR2x1_ASAP7_75t_L g129 ( 
.A(n_114),
.B(n_7),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_129),
.B(n_135),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_110),
.B(n_8),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_131),
.B(n_132),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_116),
.B(n_27),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_134),
.A2(n_14),
.B1(n_15),
.B2(n_17),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_115),
.B(n_9),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_106),
.B(n_10),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_136),
.B(n_137),
.Y(n_154)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_141),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_114),
.B(n_13),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_142),
.B(n_25),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_140),
.B(n_33),
.C(n_45),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_143),
.B(n_146),
.C(n_157),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_145),
.B(n_149),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_138),
.B(n_34),
.C(n_19),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_121),
.Y(n_149)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_139),
.Y(n_152)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_152),
.Y(n_159)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_139),
.Y(n_153)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_153),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_155),
.Y(n_164)
);

NAND3xp33_ASAP7_75t_L g163 ( 
.A(n_156),
.B(n_28),
.C(n_35),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_123),
.B(n_46),
.C(n_32),
.Y(n_157)
);

AOI322xp5_ASAP7_75t_L g158 ( 
.A1(n_147),
.A2(n_133),
.A3(n_122),
.B1(n_128),
.B2(n_137),
.C1(n_129),
.C2(n_130),
.Y(n_158)
);

AO221x1_ASAP7_75t_L g168 ( 
.A1(n_158),
.A2(n_163),
.B1(n_154),
.B2(n_148),
.C(n_150),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_159),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_165),
.B(n_166),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_164),
.A2(n_133),
.B1(n_134),
.B2(n_151),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_161),
.B(n_149),
.C(n_132),
.Y(n_167)
);

A2O1A1Ixp33_ASAP7_75t_L g170 ( 
.A1(n_167),
.A2(n_168),
.B(n_144),
.C(n_157),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_170),
.A2(n_167),
.B(n_160),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_171),
.B(n_169),
.C(n_143),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_162),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_173),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_174),
.A2(n_163),
.B(n_146),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_175),
.B(n_166),
.Y(n_176)
);


endmodule