module fake_jpeg_2349_n_381 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_381);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_381;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_292;
wire n_213;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_15),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_8),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

INVx11_ASAP7_75t_SL g39 ( 
.A(n_8),
.Y(n_39)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_1),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_44),
.Y(n_106)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_45),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_46),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g108 ( 
.A(n_49),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_29),
.B(n_13),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_50),
.B(n_52),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_51),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_24),
.B(n_13),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_53),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_54),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_55),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_59),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_27),
.B(n_23),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_60),
.B(n_71),
.Y(n_107)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_62),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_63),
.Y(n_105)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_64),
.B(n_65),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_29),
.B(n_11),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_66),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_67),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_17),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_68),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_69),
.Y(n_131)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_70),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_36),
.B(n_11),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_72),
.B(n_74),
.Y(n_102)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

INVx11_ASAP7_75t_L g118 ( 
.A(n_73),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_24),
.B(n_11),
.Y(n_74)
);

OA22x2_ASAP7_75t_L g75 ( 
.A1(n_27),
.A2(n_10),
.B1(n_1),
.B2(n_2),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_75),
.B(n_76),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_31),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_29),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_77),
.B(n_78),
.Y(n_101)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_34),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_38),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_79),
.Y(n_84)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_80),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_34),
.Y(n_81)
);

INVx11_ASAP7_75t_L g122 ( 
.A(n_81),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_34),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_26),
.Y(n_104)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_26),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_83),
.B(n_25),
.Y(n_110)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

INVx13_ASAP7_75t_L g176 ( 
.A(n_89),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_60),
.A2(n_41),
.B1(n_30),
.B2(n_20),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_91),
.A2(n_32),
.B1(n_37),
.B2(n_43),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_71),
.A2(n_25),
.B1(n_41),
.B2(n_42),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_93),
.A2(n_109),
.B1(n_132),
.B2(n_6),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_104),
.B(n_19),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_81),
.A2(n_25),
.B1(n_41),
.B2(n_42),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_110),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_75),
.B(n_28),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_111),
.B(n_119),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_82),
.B(n_31),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_112),
.B(n_116),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_46),
.A2(n_30),
.B1(n_20),
.B2(n_19),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_113),
.A2(n_32),
.B1(n_40),
.B2(n_2),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_67),
.B(n_35),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_59),
.B(n_43),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_69),
.B(n_35),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_123),
.B(n_125),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_79),
.B(n_30),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_63),
.B(n_16),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_28),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_47),
.B(n_20),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_128),
.B(n_129),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_66),
.B(n_37),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_51),
.A2(n_42),
.B1(n_19),
.B2(n_43),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_121),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_133),
.Y(n_213)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_121),
.Y(n_134)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_134),
.Y(n_211)
);

XNOR2x1_ASAP7_75t_SL g199 ( 
.A(n_135),
.B(n_177),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_136),
.A2(n_145),
.B1(n_153),
.B2(n_159),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_95),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_138),
.B(n_140),
.Y(n_198)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_106),
.Y(n_139)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_139),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_101),
.Y(n_140)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_106),
.Y(n_141)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_141),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_95),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_142),
.B(n_151),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_100),
.A2(n_58),
.B1(n_56),
.B2(n_55),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_114),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_146),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_111),
.A2(n_28),
.B(n_16),
.Y(n_147)
);

O2A1O1Ixp33_ASAP7_75t_L g212 ( 
.A1(n_147),
.A2(n_150),
.B(n_89),
.C(n_118),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_148),
.B(n_87),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_107),
.A2(n_102),
.B1(n_104),
.B2(n_128),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_149),
.Y(n_181)
);

OA22x2_ASAP7_75t_L g150 ( 
.A1(n_91),
.A2(n_54),
.B1(n_16),
.B2(n_40),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_95),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_114),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_154),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_122),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_155),
.A2(n_172),
.B1(n_175),
.B2(n_84),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_108),
.Y(n_156)
);

NAND3xp33_ASAP7_75t_L g192 ( 
.A(n_156),
.B(n_166),
.C(n_170),
.Y(n_192)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_119),
.Y(n_157)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_157),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_127),
.A2(n_10),
.B1(n_2),
.B2(n_3),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_130),
.Y(n_160)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_160),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_103),
.A2(n_1),
.B1(n_3),
.B2(n_5),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_161),
.A2(n_163),
.B1(n_94),
.B2(n_97),
.Y(n_197)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_130),
.Y(n_162)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_162),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_107),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_163)
);

NAND2xp33_ASAP7_75t_SL g164 ( 
.A(n_98),
.B(n_3),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_164),
.Y(n_216)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_92),
.Y(n_165)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_165),
.Y(n_195)
);

OR2x2_ASAP7_75t_L g166 ( 
.A(n_96),
.B(n_5),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_167),
.A2(n_87),
.B1(n_126),
.B2(n_99),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_86),
.B(n_6),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_168),
.B(n_117),
.Y(n_184)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_90),
.Y(n_169)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_169),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_108),
.Y(n_170)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_92),
.Y(n_171)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_171),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_122),
.A2(n_7),
.B1(n_9),
.B2(n_84),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_94),
.Y(n_173)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_173),
.Y(n_210)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_90),
.Y(n_174)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_174),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_103),
.A2(n_7),
.B1(n_9),
.B2(n_105),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_98),
.B(n_9),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_157),
.B(n_85),
.C(n_117),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_178),
.B(n_202),
.C(n_150),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_146),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_182),
.B(n_184),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_185),
.B(n_187),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_176),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_190),
.B(n_212),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_140),
.B(n_126),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_193),
.B(n_197),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_137),
.A2(n_108),
.B1(n_131),
.B2(n_85),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_194),
.A2(n_205),
.B1(n_175),
.B2(n_170),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_137),
.B(n_148),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_200),
.B(n_201),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_149),
.A2(n_120),
.B1(n_105),
.B2(n_97),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_135),
.B(n_120),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_135),
.B(n_158),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_204),
.B(n_136),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_145),
.A2(n_131),
.B1(n_115),
.B2(n_99),
.Y(n_205)
);

XNOR2x1_ASAP7_75t_L g241 ( 
.A(n_206),
.B(n_205),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_154),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_209),
.B(n_215),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_143),
.B(n_115),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_200),
.B(n_144),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_218),
.B(n_239),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_204),
.B(n_144),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_221),
.B(n_232),
.Y(n_266)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_203),
.Y(n_222)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_222),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_188),
.A2(n_147),
.B1(n_152),
.B2(n_150),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_223),
.A2(n_235),
.B1(n_245),
.B2(n_201),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_212),
.A2(n_164),
.B(n_176),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_225),
.A2(n_227),
.B(n_236),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_216),
.A2(n_166),
.B(n_177),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_226),
.A2(n_207),
.B(n_179),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_216),
.A2(n_177),
.B(n_151),
.Y(n_227)
);

CKINVDCx14_ASAP7_75t_R g228 ( 
.A(n_198),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_228),
.B(n_231),
.Y(n_260)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_196),
.Y(n_229)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_229),
.Y(n_254)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_196),
.Y(n_230)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_230),
.Y(n_255)
);

OAI221xp5_ASAP7_75t_L g232 ( 
.A1(n_199),
.A2(n_150),
.B1(n_159),
.B2(n_174),
.C(n_169),
.Y(n_232)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_214),
.Y(n_234)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_234),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_188),
.A2(n_181),
.B1(n_183),
.B2(n_190),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_192),
.A2(n_142),
.B(n_139),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_237),
.B(n_242),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_L g272 ( 
.A1(n_238),
.A2(n_191),
.B1(n_186),
.B2(n_210),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_199),
.B(n_162),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_214),
.Y(n_240)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_240),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_SL g263 ( 
.A(n_241),
.B(n_247),
.C(n_185),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_183),
.B(n_161),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_202),
.B(n_160),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_243),
.B(n_244),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_178),
.B(n_156),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_197),
.A2(n_88),
.B1(n_124),
.B2(n_134),
.Y(n_245)
);

AOI32xp33_ASAP7_75t_L g247 ( 
.A1(n_182),
.A2(n_173),
.A3(n_171),
.B1(n_165),
.B2(n_141),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_179),
.B(n_88),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_248),
.B(n_189),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_250),
.A2(n_265),
.B1(n_272),
.B2(n_274),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_228),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_251),
.B(n_263),
.Y(n_278)
);

INVx13_ASAP7_75t_L g253 ( 
.A(n_227),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_253),
.Y(n_282)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_258),
.Y(n_292)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_229),
.Y(n_259)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_259),
.Y(n_298)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_230),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_264),
.B(n_267),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_223),
.A2(n_211),
.B1(n_180),
.B2(n_189),
.Y(n_265)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_222),
.Y(n_267)
);

NOR2x1_ASAP7_75t_L g268 ( 
.A(n_237),
.B(n_226),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_268),
.B(n_271),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_224),
.A2(n_206),
.B1(n_211),
.B2(n_124),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_269),
.A2(n_232),
.B1(n_238),
.B2(n_220),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_270),
.B(n_246),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_246),
.Y(n_271)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_234),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_273),
.B(n_248),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_231),
.A2(n_133),
.B1(n_186),
.B2(n_191),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_250),
.A2(n_220),
.B1(n_224),
.B2(n_219),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_276),
.A2(n_285),
.B1(n_262),
.B2(n_274),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_249),
.A2(n_236),
.B(n_225),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_277),
.A2(n_249),
.B(n_253),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_260),
.B(n_239),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_279),
.B(n_280),
.C(n_288),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_260),
.B(n_244),
.C(n_218),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_254),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_281),
.B(n_284),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_283),
.Y(n_300)
);

NOR2xp67_ASAP7_75t_SL g284 ( 
.A(n_267),
.B(n_217),
.Y(n_284)
);

FAx1_ASAP7_75t_SL g286 ( 
.A(n_261),
.B(n_235),
.CI(n_268),
.CON(n_286),
.SN(n_286)
);

A2O1A1O1Ixp25_ASAP7_75t_L g304 ( 
.A1(n_286),
.A2(n_287),
.B(n_262),
.C(n_270),
.D(n_252),
.Y(n_304)
);

A2O1A1Ixp33_ASAP7_75t_L g287 ( 
.A1(n_266),
.A2(n_217),
.B(n_219),
.C(n_242),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_261),
.B(n_243),
.C(n_240),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_261),
.B(n_233),
.C(n_221),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_289),
.B(n_296),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_271),
.B(n_233),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_294),
.B(n_297),
.Y(n_308)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_295),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_275),
.B(n_207),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_275),
.B(n_247),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_290),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_301),
.B(n_310),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_290),
.B(n_251),
.Y(n_302)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_302),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_303),
.A2(n_304),
.B1(n_313),
.B2(n_314),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_306),
.B(n_309),
.Y(n_328)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_298),
.Y(n_307)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_307),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_295),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_292),
.B(n_252),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_291),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_311),
.Y(n_326)
);

OAI32xp33_ASAP7_75t_L g312 ( 
.A1(n_291),
.A2(n_263),
.A3(n_273),
.B1(n_255),
.B2(n_257),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_312),
.A2(n_318),
.B1(n_180),
.B2(n_241),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_293),
.A2(n_269),
.B1(n_265),
.B2(n_264),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_276),
.A2(n_285),
.B1(n_297),
.B2(n_287),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_282),
.A2(n_259),
.B1(n_257),
.B2(n_256),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_315),
.B(n_277),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_278),
.A2(n_256),
.B1(n_255),
.B2(n_254),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_316),
.B(n_279),
.C(n_280),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_322),
.B(n_329),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_323),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_316),
.B(n_283),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_324),
.B(n_333),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_311),
.A2(n_278),
.B1(n_282),
.B2(n_289),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_325),
.A2(n_331),
.B1(n_334),
.B2(n_305),
.Y(n_347)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_302),
.Y(n_327)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_327),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_317),
.B(n_288),
.C(n_296),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_317),
.B(n_300),
.C(n_308),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_330),
.B(n_335),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_303),
.A2(n_286),
.B1(n_298),
.B2(n_245),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_314),
.B(n_286),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_318),
.B(n_195),
.C(n_208),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_329),
.B(n_312),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_337),
.B(n_341),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_322),
.B(n_306),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_332),
.B(n_299),
.Y(n_342)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_342),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_321),
.A2(n_309),
.B1(n_305),
.B2(n_313),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_343),
.A2(n_331),
.B1(n_304),
.B2(n_333),
.Y(n_353)
);

CKINVDCx16_ASAP7_75t_R g344 ( 
.A(n_328),
.Y(n_344)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_344),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_326),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_345),
.A2(n_319),
.B1(n_320),
.B2(n_307),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_347),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_324),
.B(n_315),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_L g357 ( 
.A1(n_348),
.A2(n_330),
.B(n_195),
.Y(n_357)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_350),
.Y(n_360)
);

AOI22xp33_ASAP7_75t_SL g351 ( 
.A1(n_346),
.A2(n_335),
.B1(n_325),
.B2(n_323),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g363 ( 
.A(n_351),
.Y(n_363)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_353),
.Y(n_366)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_343),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_356),
.B(n_347),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_357),
.B(n_336),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_337),
.A2(n_213),
.B1(n_208),
.B2(n_133),
.Y(n_358)
);

OR2x2_ASAP7_75t_L g362 ( 
.A(n_358),
.B(n_348),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_355),
.B(n_338),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_359),
.B(n_361),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_362),
.B(n_364),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_355),
.B(n_341),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_365),
.B(n_340),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_360),
.B(n_352),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_368),
.Y(n_375)
);

AOI322xp5_ASAP7_75t_L g369 ( 
.A1(n_366),
.A2(n_354),
.A3(n_349),
.B1(n_339),
.B2(n_340),
.C1(n_351),
.C2(n_336),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_369),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_361),
.B(n_349),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_SL g374 ( 
.A1(n_370),
.A2(n_372),
.B(n_363),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_374),
.A2(n_367),
.B(n_363),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_L g376 ( 
.A1(n_373),
.A2(n_371),
.B(n_367),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g378 ( 
.A1(n_376),
.A2(n_377),
.B(n_375),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_378),
.B(n_213),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_379),
.B(n_210),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_380),
.B(n_118),
.Y(n_381)
);


endmodule