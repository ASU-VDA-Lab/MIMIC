module fake_jpeg_19007_n_300 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_300);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_300;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

BUFx16f_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx2_ASAP7_75t_SL g16 ( 
.A(n_13),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_4),
.B(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_35),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_24),
.Y(n_53)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_27),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_44),
.Y(n_57)
);

AND2x2_ASAP7_75t_SL g44 ( 
.A(n_39),
.B(n_23),
.Y(n_44)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_38),
.A2(n_16),
.B1(n_29),
.B2(n_30),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_47),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_32),
.A2(n_29),
.B1(n_16),
.B2(n_18),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_50),
.A2(n_16),
.B1(n_17),
.B2(n_30),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_27),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_52),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_33),
.B(n_23),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_53),
.B(n_24),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_49),
.A2(n_16),
.B1(n_29),
.B2(n_20),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_55),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_56),
.Y(n_104)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_58),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_33),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_60),
.B(n_66),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_49),
.A2(n_16),
.B1(n_20),
.B2(n_17),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_61),
.A2(n_42),
.B1(n_46),
.B2(n_49),
.Y(n_89)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_62),
.Y(n_111)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_64),
.A2(n_77),
.B1(n_80),
.B2(n_35),
.Y(n_85)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_65),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_37),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_67),
.B(n_70),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_68),
.B(n_31),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_37),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_69),
.A2(n_48),
.B1(n_15),
.B2(n_26),
.Y(n_110)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_71),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_72),
.Y(n_86)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_73),
.B(n_76),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_52),
.A2(n_18),
.B1(n_20),
.B2(n_24),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_74),
.A2(n_31),
.B1(n_22),
.B2(n_21),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_36),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_75),
.B(n_36),
.Y(n_102)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_44),
.A2(n_35),
.B1(n_30),
.B2(n_21),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_42),
.Y(n_101)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_79),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_44),
.A2(n_51),
.B1(n_47),
.B2(n_46),
.Y(n_80)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_82),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_85),
.A2(n_93),
.B1(n_96),
.B2(n_81),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_88),
.B(n_108),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_89),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_59),
.B(n_57),
.C(n_71),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_91),
.B(n_48),
.Y(n_114)
);

O2A1O1Ixp33_ASAP7_75t_L g93 ( 
.A1(n_82),
.A2(n_44),
.B(n_45),
.C(n_46),
.Y(n_93)
);

OA22x2_ASAP7_75t_L g94 ( 
.A1(n_76),
.A2(n_80),
.B1(n_83),
.B2(n_69),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_94),
.B(n_63),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_59),
.A2(n_57),
.B1(n_60),
.B2(n_66),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_69),
.A2(n_45),
.B(n_48),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_99),
.A2(n_110),
.B(n_67),
.Y(n_119)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_101),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_102),
.B(n_109),
.Y(n_127)
);

AND2x2_ASAP7_75t_SL g105 ( 
.A(n_75),
.B(n_34),
.Y(n_105)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_105),
.Y(n_131)
);

AOI32xp33_ASAP7_75t_L g106 ( 
.A1(n_79),
.A2(n_42),
.A3(n_34),
.B1(n_26),
.B2(n_21),
.Y(n_106)
);

AOI32xp33_ASAP7_75t_L g117 ( 
.A1(n_106),
.A2(n_81),
.A3(n_78),
.B1(n_58),
.B2(n_26),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_77),
.B(n_42),
.Y(n_109)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_112),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_103),
.A2(n_64),
.B1(n_62),
.B2(n_65),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_113),
.A2(n_133),
.B1(n_137),
.B2(n_93),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_114),
.B(n_123),
.C(n_105),
.Y(n_143)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_111),
.Y(n_115)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_115),
.Y(n_161)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_111),
.Y(n_116)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_116),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_117),
.A2(n_119),
.B(n_122),
.Y(n_149)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_95),
.Y(n_120)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_120),
.Y(n_166)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_101),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_121),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_91),
.B(n_25),
.Y(n_123)
);

BUFx2_ASAP7_75t_SL g124 ( 
.A(n_86),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_124),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_125),
.A2(n_93),
.B1(n_102),
.B2(n_107),
.Y(n_141)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_90),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_126),
.B(n_130),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_84),
.B(n_56),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_128),
.B(n_84),
.Y(n_140)
);

BUFx2_ASAP7_75t_L g130 ( 
.A(n_86),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_103),
.A2(n_31),
.B(n_22),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_132),
.A2(n_129),
.B(n_88),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_109),
.A2(n_22),
.B1(n_28),
.B2(n_23),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_104),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_135),
.B(n_136),
.Y(n_168)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_90),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_99),
.A2(n_28),
.B1(n_23),
.B2(n_19),
.Y(n_137)
);

INVx4_ASAP7_75t_SL g138 ( 
.A(n_87),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_138),
.A2(n_98),
.B1(n_87),
.B2(n_106),
.Y(n_142)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_104),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_139),
.B(n_97),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_140),
.B(n_147),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_141),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_196)
);

CKINVDCx14_ASAP7_75t_R g174 ( 
.A(n_142),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_143),
.B(n_160),
.Y(n_200)
);

FAx1_ASAP7_75t_SL g144 ( 
.A(n_123),
.B(n_96),
.CI(n_100),
.CON(n_144),
.SN(n_144)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_144),
.B(n_146),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_139),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_148),
.B(n_169),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_134),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_150),
.B(n_151),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_134),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_152),
.A2(n_153),
.B1(n_112),
.B2(n_28),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_118),
.A2(n_92),
.B1(n_98),
.B2(n_107),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_128),
.B(n_107),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_154),
.B(n_133),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_122),
.A2(n_94),
.B(n_105),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_155),
.B(n_159),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_114),
.B(n_94),
.C(n_105),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_156),
.B(n_158),
.C(n_120),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_125),
.B(n_94),
.C(n_85),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_127),
.B(n_100),
.Y(n_159)
);

MAJx2_ASAP7_75t_L g160 ( 
.A(n_119),
.B(n_94),
.C(n_110),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_122),
.A2(n_97),
.B1(n_108),
.B2(n_72),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_162),
.A2(n_165),
.B1(n_72),
.B2(n_28),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_113),
.A2(n_118),
.B1(n_127),
.B2(n_131),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_130),
.Y(n_169)
);

OR2x2_ASAP7_75t_L g170 ( 
.A(n_131),
.B(n_132),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_170),
.B(n_72),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_171),
.B(n_176),
.Y(n_206)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_168),
.Y(n_172)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_172),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_143),
.B(n_138),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_175),
.B(n_178),
.Y(n_208)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_164),
.Y(n_177)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_177),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_179),
.A2(n_170),
.B1(n_167),
.B2(n_154),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_182),
.A2(n_185),
.B1(n_186),
.B2(n_190),
.Y(n_204)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_170),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_183),
.B(n_184),
.Y(n_210)
);

OAI32xp33_ASAP7_75t_L g184 ( 
.A1(n_159),
.A2(n_19),
.A3(n_25),
.B1(n_15),
.B2(n_9),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_158),
.A2(n_19),
.B1(n_25),
.B2(n_15),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_165),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_186)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_169),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_187),
.B(n_188),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_161),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_144),
.B(n_14),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_189),
.B(n_9),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_148),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_161),
.Y(n_191)
);

OR2x2_ASAP7_75t_L g218 ( 
.A(n_191),
.B(n_166),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_156),
.B(n_14),
.C(n_13),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_192),
.B(n_152),
.C(n_149),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_144),
.B(n_140),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_194),
.B(n_145),
.Y(n_216)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_163),
.Y(n_195)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_195),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_196),
.A2(n_157),
.B1(n_5),
.B2(n_6),
.Y(n_221)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_163),
.Y(n_198)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_198),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_162),
.A2(n_0),
.B1(n_3),
.B2(n_5),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_199),
.A2(n_141),
.B1(n_151),
.B2(n_150),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_201),
.A2(n_189),
.B(n_173),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_175),
.B(n_149),
.C(n_155),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_202),
.B(n_214),
.C(n_178),
.Y(n_227)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_209),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_212),
.A2(n_215),
.B1(n_220),
.B2(n_221),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_200),
.B(n_160),
.C(n_147),
.Y(n_214)
);

OAI22x1_ASAP7_75t_L g215 ( 
.A1(n_174),
.A2(n_146),
.B1(n_167),
.B2(n_145),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_216),
.B(n_217),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_218),
.Y(n_226)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_181),
.Y(n_219)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_219),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_180),
.A2(n_166),
.B1(n_157),
.B2(n_6),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_197),
.B(n_3),
.Y(n_222)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_222),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_224),
.B(n_227),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_215),
.A2(n_213),
.B(n_218),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_229),
.B(n_231),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_210),
.A2(n_182),
.B1(n_190),
.B2(n_185),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_230),
.B(n_236),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_208),
.B(n_200),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_208),
.B(n_194),
.C(n_193),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_232),
.B(n_234),
.C(n_237),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_216),
.B(n_192),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_233),
.B(n_239),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_214),
.B(n_197),
.C(n_176),
.Y(n_234)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_205),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_202),
.B(n_176),
.C(n_179),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_201),
.B(n_184),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_206),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_240),
.B(n_220),
.Y(n_247)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_226),
.Y(n_242)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_242),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_235),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_243),
.B(n_248),
.Y(n_260)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_238),
.Y(n_244)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_244),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_223),
.A2(n_210),
.B1(n_186),
.B2(n_183),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_245),
.A2(n_252),
.B1(n_254),
.B2(n_196),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_231),
.B(n_206),
.C(n_209),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_246),
.B(n_241),
.C(n_250),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_247),
.Y(n_264)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_228),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_239),
.A2(n_221),
.B1(n_199),
.B2(n_204),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_240),
.B(n_203),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_253),
.B(n_187),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_233),
.A2(n_204),
.B1(n_211),
.B2(n_207),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_246),
.B(n_234),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_256),
.B(n_257),
.C(n_261),
.Y(n_271)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_258),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_259),
.A2(n_245),
.B1(n_225),
.B2(n_217),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_255),
.B(n_227),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_254),
.B(n_222),
.Y(n_263)
);

CKINVDCx14_ASAP7_75t_R g270 ( 
.A(n_263),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_255),
.B(n_237),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_265),
.B(n_267),
.C(n_261),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_241),
.B(n_232),
.Y(n_267)
);

OR2x2_ASAP7_75t_L g268 ( 
.A(n_260),
.B(n_250),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_268),
.A2(n_276),
.B1(n_266),
.B2(n_265),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_264),
.B(n_247),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_269),
.B(n_274),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_272),
.B(n_10),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_262),
.B(n_249),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_257),
.B(n_251),
.C(n_252),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_275),
.B(n_277),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_267),
.B(n_251),
.C(n_225),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_278),
.B(n_282),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_271),
.B(n_256),
.C(n_269),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_281),
.B(n_285),
.C(n_10),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_273),
.B(n_270),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_274),
.B(n_12),
.Y(n_283)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_283),
.Y(n_286)
);

FAx1_ASAP7_75t_L g284 ( 
.A(n_276),
.B(n_12),
.CI(n_11),
.CON(n_284),
.SN(n_284)
);

NOR2xp67_ASAP7_75t_SL g290 ( 
.A(n_284),
.B(n_3),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_288),
.B(n_289),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_281),
.B(n_11),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_290),
.B(n_286),
.Y(n_292)
);

AO21x1_ASAP7_75t_L g294 ( 
.A1(n_292),
.A2(n_293),
.B(n_279),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_287),
.B(n_280),
.Y(n_293)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_294),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_291),
.Y(n_295)
);

OAI321xp33_ASAP7_75t_L g297 ( 
.A1(n_296),
.A2(n_295),
.A3(n_284),
.B1(n_7),
.B2(n_8),
.C(n_6),
.Y(n_297)
);

A2O1A1Ixp33_ASAP7_75t_L g298 ( 
.A1(n_297),
.A2(n_284),
.B(n_7),
.C(n_8),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_298),
.B(n_5),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_299),
.B(n_5),
.Y(n_300)
);


endmodule