module fake_netlist_6_2374_n_464 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_464);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_464;

wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_209;
wire n_367;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_342;
wire n_358;
wire n_160;
wire n_449;
wire n_188;
wire n_310;
wire n_186;
wire n_245;
wire n_368;
wire n_396;
wire n_350;
wire n_392;
wire n_442;
wire n_382;
wire n_180;
wire n_349;
wire n_233;
wire n_255;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_443;
wire n_246;
wire n_289;
wire n_421;
wire n_424;
wire n_181;
wire n_182;
wire n_238;
wire n_202;
wire n_320;
wire n_327;
wire n_369;
wire n_280;
wire n_287;
wire n_353;
wire n_389;
wire n_415;
wire n_230;
wire n_461;
wire n_383;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_300;
wire n_179;
wire n_248;
wire n_222;
wire n_229;
wire n_305;
wire n_173;
wire n_250;
wire n_372;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_375;
wire n_338;
wire n_360;
wire n_235;
wire n_191;
wire n_340;
wire n_387;
wire n_452;
wire n_344;
wire n_428;
wire n_432;
wire n_167;
wire n_174;
wire n_371;
wire n_189;
wire n_405;
wire n_213;
wire n_294;
wire n_302;
wire n_380;
wire n_197;
wire n_343;
wire n_448;
wire n_397;
wire n_445;
wire n_425;
wire n_454;
wire n_218;
wire n_234;
wire n_381;
wire n_236;
wire n_172;
wire n_270;
wire n_239;
wire n_414;
wire n_290;
wire n_220;
wire n_224;
wire n_196;
wire n_402;
wire n_352;
wire n_460;
wire n_417;
wire n_446;
wire n_374;
wire n_366;
wire n_407;
wire n_450;
wire n_272;
wire n_185;
wire n_348;
wire n_376;
wire n_390;
wire n_293;
wire n_334;
wire n_370;
wire n_458;
wire n_232;
wire n_163;
wire n_330;
wire n_298;
wire n_281;
wire n_258;
wire n_456;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_279;
wire n_252;
wire n_228;
wire n_356;
wire n_166;
wire n_184;
wire n_216;
wire n_455;
wire n_363;
wire n_395;
wire n_323;
wire n_393;
wire n_411;
wire n_321;
wire n_331;
wire n_227;
wire n_406;
wire n_204;
wire n_261;
wire n_420;
wire n_312;
wire n_394;
wire n_164;
wire n_292;
wire n_307;
wire n_433;
wire n_291;
wire n_219;
wire n_357;
wire n_264;
wire n_263;
wire n_325;
wire n_329;
wire n_408;
wire n_237;
wire n_244;
wire n_399;
wire n_243;
wire n_282;
wire n_436;
wire n_211;
wire n_175;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_240;
wire n_319;
wire n_273;
wire n_311;
wire n_403;
wire n_253;
wire n_249;
wire n_201;
wire n_386;
wire n_162;
wire n_241;
wire n_275;
wire n_276;
wire n_441;
wire n_221;
wire n_444;
wire n_423;
wire n_318;
wire n_303;
wire n_306;
wire n_269;
wire n_193;
wire n_359;
wire n_346;
wire n_416;
wire n_277;
wire n_418;
wire n_199;
wire n_266;
wire n_296;
wire n_268;
wire n_271;
wire n_404;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_206;
wire n_453;
wire n_333;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_426;
wire n_317;
wire n_431;
wire n_347;
wire n_459;
wire n_328;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_257;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_401;
wire n_324;
wire n_335;
wire n_430;
wire n_463;
wire n_205;
wire n_251;
wire n_301;
wire n_274;
wire n_412;
wire n_267;
wire n_438;
wire n_339;
wire n_434;
wire n_315;
wire n_288;
wire n_427;
wire n_422;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_391;
wire n_457;
wire n_364;
wire n_295;
wire n_385;
wire n_388;
wire n_190;
wire n_262;
wire n_187;
wire n_361;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_194;
wire n_171;
wire n_192;
wire n_169;
wire n_283;

INVxp67_ASAP7_75t_L g160 ( 
.A(n_49),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_156),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_125),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_10),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_21),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_30),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_98),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_142),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_63),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_6),
.Y(n_169)
);

INVxp33_ASAP7_75t_SL g170 ( 
.A(n_83),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_24),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_1),
.Y(n_172)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_20),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_127),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_79),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_55),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_141),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_43),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_40),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_4),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_52),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_148),
.Y(n_182)
);

NOR2xp67_ASAP7_75t_L g183 ( 
.A(n_51),
.B(n_27),
.Y(n_183)
);

INVxp33_ASAP7_75t_L g184 ( 
.A(n_146),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_112),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_32),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_54),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_118),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_48),
.B(n_60),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_14),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_19),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_100),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_143),
.Y(n_193)
);

NOR2xp67_ASAP7_75t_L g194 ( 
.A(n_88),
.B(n_96),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_8),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_31),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_123),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_80),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_3),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_37),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_47),
.Y(n_201)
);

INVxp67_ASAP7_75t_SL g202 ( 
.A(n_101),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_107),
.Y(n_203)
);

INVxp67_ASAP7_75t_SL g204 ( 
.A(n_69),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_144),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_150),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_155),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_46),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_140),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_71),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_94),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_65),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_151),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_130),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_25),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_139),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_38),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_64),
.B(n_110),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_103),
.Y(n_219)
);

BUFx2_ASAP7_75t_L g220 ( 
.A(n_102),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_149),
.B(n_126),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_137),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_53),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_7),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_91),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_72),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_108),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_77),
.Y(n_228)
);

INVxp33_ASAP7_75t_SL g229 ( 
.A(n_17),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_104),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_75),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_5),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_34),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_92),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_28),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_74),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_154),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_158),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_95),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_87),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_73),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_128),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_1),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_44),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_134),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_111),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_2),
.Y(n_247)
);

INVxp67_ASAP7_75t_SL g248 ( 
.A(n_115),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_152),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_58),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_57),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_33),
.Y(n_252)
);

INVxp67_ASAP7_75t_SL g253 ( 
.A(n_67),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_159),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_22),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_132),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_81),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_109),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_78),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_45),
.Y(n_260)
);

INVxp67_ASAP7_75t_SL g261 ( 
.A(n_36),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_R g262 ( 
.A(n_136),
.B(n_70),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_89),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_121),
.B(n_84),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_23),
.Y(n_265)
);

INVxp67_ASAP7_75t_SL g266 ( 
.A(n_122),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_26),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_11),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_76),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_157),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_120),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_153),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_116),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_113),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_9),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_35),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_3),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_93),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_106),
.B(n_66),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_82),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_135),
.B(n_147),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_199),
.Y(n_282)
);

BUFx10_ASAP7_75t_L g283 ( 
.A(n_172),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_243),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_220),
.B(n_0),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_233),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_162),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_L g288 ( 
.A1(n_171),
.A2(n_0),
.B1(n_2),
.B2(n_12),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_164),
.Y(n_289)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_277),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_167),
.Y(n_291)
);

AND2x6_ASAP7_75t_L g292 ( 
.A(n_218),
.B(n_13),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_177),
.Y(n_293)
);

INVx4_ASAP7_75t_L g294 ( 
.A(n_165),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_168),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_197),
.Y(n_296)
);

OR2x2_ASAP7_75t_L g297 ( 
.A(n_173),
.B(n_15),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_179),
.A2(n_16),
.B1(n_18),
.B2(n_29),
.Y(n_298)
);

BUFx4f_ASAP7_75t_L g299 ( 
.A(n_178),
.Y(n_299)
);

BUFx2_ASAP7_75t_L g300 ( 
.A(n_247),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_182),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_161),
.A2(n_39),
.B1(n_41),
.B2(n_42),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_190),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_180),
.B(n_50),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_192),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_265),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_198),
.Y(n_307)
);

BUFx2_ASAP7_75t_L g308 ( 
.A(n_163),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_234),
.B(n_184),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_160),
.B(n_56),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_201),
.Y(n_311)
);

INVx1_ASAP7_75t_SL g312 ( 
.A(n_166),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_174),
.B(n_59),
.Y(n_313)
);

AND3x2_ASAP7_75t_L g314 ( 
.A(n_264),
.B(n_61),
.C(n_62),
.Y(n_314)
);

BUFx6f_ASAP7_75t_SL g315 ( 
.A(n_203),
.Y(n_315)
);

AND2x6_ASAP7_75t_L g316 ( 
.A(n_264),
.B(n_68),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_230),
.B(n_85),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_255),
.B(n_86),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_258),
.B(n_90),
.Y(n_319)
);

INVx5_ASAP7_75t_L g320 ( 
.A(n_183),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_207),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_267),
.B(n_97),
.Y(n_322)
);

AND2x4_ASAP7_75t_L g323 ( 
.A(n_208),
.B(n_99),
.Y(n_323)
);

BUFx3_ASAP7_75t_L g324 ( 
.A(n_169),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_268),
.B(n_105),
.Y(n_325)
);

OAI22xp33_ASAP7_75t_L g326 ( 
.A1(n_209),
.A2(n_114),
.B1(n_117),
.B2(n_119),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_210),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_170),
.B(n_229),
.Y(n_328)
);

INVxp67_ASAP7_75t_SL g329 ( 
.A(n_274),
.Y(n_329)
);

AND2x6_ASAP7_75t_L g330 ( 
.A(n_279),
.B(n_124),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_212),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_223),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_226),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_227),
.Y(n_334)
);

INVx4_ASAP7_75t_L g335 ( 
.A(n_175),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_275),
.B(n_129),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_289),
.B(n_228),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_295),
.B(n_324),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_290),
.B(n_232),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_309),
.A2(n_235),
.B1(n_280),
.B2(n_260),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_328),
.B(n_238),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_L g342 ( 
.A1(n_285),
.A2(n_225),
.B1(n_231),
.B2(n_242),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g343 ( 
.A(n_284),
.B(n_176),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g344 ( 
.A1(n_322),
.A2(n_279),
.B(n_204),
.Y(n_344)
);

BUFx8_ASAP7_75t_SL g345 ( 
.A(n_300),
.Y(n_345)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_329),
.B(n_224),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_299),
.A2(n_253),
.B(n_248),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_333),
.A2(n_286),
.B(n_325),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_310),
.A2(n_202),
.B(n_261),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_306),
.A2(n_222),
.B1(n_256),
.B2(n_276),
.Y(n_350)
);

A2O1A1Ixp33_ASAP7_75t_L g351 ( 
.A1(n_336),
.A2(n_194),
.B(n_189),
.C(n_221),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_335),
.B(n_241),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_296),
.Y(n_353)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_313),
.A2(n_266),
.B(n_278),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_294),
.B(n_244),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_304),
.B(n_205),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_317),
.A2(n_249),
.B(n_252),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_323),
.B(n_254),
.Y(n_358)
);

OAI21xp33_ASAP7_75t_L g359 ( 
.A1(n_297),
.A2(n_281),
.B(n_257),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_320),
.B(n_296),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_318),
.A2(n_270),
.B(n_271),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_L g362 ( 
.A1(n_319),
.A2(n_214),
.B(n_269),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_320),
.B(n_213),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_L g364 ( 
.A1(n_291),
.A2(n_211),
.B(n_263),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_301),
.A2(n_311),
.B(n_332),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_303),
.B(n_273),
.Y(n_366)
);

AOI22xp33_ASAP7_75t_L g367 ( 
.A1(n_316),
.A2(n_206),
.B1(n_251),
.B2(n_245),
.Y(n_367)
);

NAND2xp33_ASAP7_75t_L g368 ( 
.A(n_288),
.B(n_262),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_283),
.B(n_196),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_327),
.Y(n_370)
);

O2A1O1Ixp33_ASAP7_75t_L g371 ( 
.A1(n_282),
.A2(n_200),
.B(n_219),
.C(n_217),
.Y(n_371)
);

AOI21xp5_ASAP7_75t_L g372 ( 
.A1(n_305),
.A2(n_321),
.B(n_307),
.Y(n_372)
);

AOI21x1_ASAP7_75t_L g373 ( 
.A1(n_287),
.A2(n_193),
.B(n_195),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_SL g374 ( 
.A1(n_351),
.A2(n_298),
.B(n_292),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_368),
.A2(n_316),
.B1(n_330),
.B2(n_272),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_344),
.B(n_330),
.Y(n_376)
);

O2A1O1Ixp33_ASAP7_75t_SL g377 ( 
.A1(n_358),
.A2(n_326),
.B(n_331),
.C(n_293),
.Y(n_377)
);

AOI211xp5_ASAP7_75t_L g378 ( 
.A1(n_359),
.A2(n_312),
.B(n_308),
.C(n_334),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_353),
.Y(n_379)
);

INVx4_ASAP7_75t_L g380 ( 
.A(n_370),
.Y(n_380)
);

INVxp67_ASAP7_75t_SL g381 ( 
.A(n_370),
.Y(n_381)
);

AND2x4_ASAP7_75t_L g382 ( 
.A(n_338),
.B(n_215),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_370),
.Y(n_383)
);

AOI21xp33_ASAP7_75t_SL g384 ( 
.A1(n_350),
.A2(n_302),
.B(n_237),
.Y(n_384)
);

AOI221xp5_ASAP7_75t_L g385 ( 
.A1(n_342),
.A2(n_186),
.B1(n_191),
.B2(n_187),
.C(n_185),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_360),
.Y(n_386)
);

AO31x2_ASAP7_75t_L g387 ( 
.A1(n_357),
.A2(n_361),
.A3(n_341),
.B(n_354),
.Y(n_387)
);

BUFx2_ASAP7_75t_L g388 ( 
.A(n_345),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_367),
.B(n_181),
.Y(n_389)
);

INVx5_ASAP7_75t_L g390 ( 
.A(n_343),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_339),
.Y(n_391)
);

O2A1O1Ixp33_ASAP7_75t_L g392 ( 
.A1(n_337),
.A2(n_330),
.B(n_316),
.C(n_292),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_366),
.Y(n_393)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_373),
.Y(n_394)
);

INVx3_ASAP7_75t_SL g395 ( 
.A(n_369),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_346),
.B(n_239),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_348),
.B(n_292),
.Y(n_397)
);

OR2x6_ASAP7_75t_L g398 ( 
.A(n_371),
.B(n_327),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_379),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_391),
.B(n_340),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_386),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_383),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_395),
.B(n_363),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_387),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_387),
.Y(n_405)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_393),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_380),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_381),
.Y(n_408)
);

HB1xp67_ASAP7_75t_L g409 ( 
.A(n_398),
.Y(n_409)
);

HB1xp67_ASAP7_75t_L g410 ( 
.A(n_398),
.Y(n_410)
);

OR2x6_ASAP7_75t_L g411 ( 
.A(n_388),
.B(n_372),
.Y(n_411)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_394),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_397),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_376),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_390),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_382),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_377),
.Y(n_417)
);

NAND3xp33_ASAP7_75t_L g418 ( 
.A(n_414),
.B(n_384),
.C(n_385),
.Y(n_418)
);

NAND3xp33_ASAP7_75t_L g419 ( 
.A(n_400),
.B(n_378),
.C(n_389),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_413),
.A2(n_375),
.B1(n_374),
.B2(n_390),
.Y(n_420)
);

AOI21xp5_ASAP7_75t_L g421 ( 
.A1(n_412),
.A2(n_392),
.B(n_396),
.Y(n_421)
);

NAND3xp33_ASAP7_75t_L g422 ( 
.A(n_401),
.B(n_356),
.C(n_390),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_406),
.B(n_355),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_406),
.B(n_349),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_403),
.B(n_352),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_417),
.B(n_412),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_408),
.B(n_347),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_404),
.B(n_364),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_416),
.B(n_365),
.Y(n_429)
);

NAND3xp33_ASAP7_75t_L g430 ( 
.A(n_409),
.B(n_236),
.C(n_216),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g431 ( 
.A(n_410),
.B(n_240),
.Y(n_431)
);

AOI22xp33_ASAP7_75t_L g432 ( 
.A1(n_405),
.A2(n_399),
.B1(n_415),
.B2(n_402),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_425),
.B(n_411),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_423),
.B(n_407),
.Y(n_434)
);

OR2x2_ASAP7_75t_L g435 ( 
.A(n_419),
.B(n_418),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_431),
.Y(n_436)
);

AND2x4_ASAP7_75t_L g437 ( 
.A(n_429),
.B(n_411),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_426),
.Y(n_438)
);

OAI22xp33_ASAP7_75t_L g439 ( 
.A1(n_418),
.A2(n_246),
.B1(n_259),
.B2(n_250),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_432),
.B(n_188),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_420),
.B(n_314),
.Y(n_441)
);

NOR2x1p5_ASAP7_75t_L g442 ( 
.A(n_435),
.B(n_422),
.Y(n_442)
);

INVx1_ASAP7_75t_SL g443 ( 
.A(n_433),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_438),
.Y(n_444)
);

AOI22xp33_ASAP7_75t_L g445 ( 
.A1(n_437),
.A2(n_430),
.B1(n_428),
.B2(n_427),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_437),
.B(n_424),
.Y(n_446)
);

INVx1_ASAP7_75t_SL g447 ( 
.A(n_434),
.Y(n_447)
);

INVx2_ASAP7_75t_SL g448 ( 
.A(n_440),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_447),
.B(n_436),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_444),
.B(n_439),
.Y(n_450)
);

NOR2x1_ASAP7_75t_L g451 ( 
.A(n_442),
.B(n_441),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_443),
.B(n_262),
.Y(n_452)
);

NOR2x1_ASAP7_75t_L g453 ( 
.A(n_451),
.B(n_446),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_450),
.B(n_448),
.Y(n_454)
);

XNOR2x1_ASAP7_75t_L g455 ( 
.A(n_449),
.B(n_443),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_452),
.B(n_315),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_454),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_453),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_458),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_457),
.B(n_455),
.Y(n_460)
);

OR2x2_ASAP7_75t_L g461 ( 
.A(n_459),
.B(n_456),
.Y(n_461)
);

OAI21x1_ASAP7_75t_L g462 ( 
.A1(n_461),
.A2(n_460),
.B(n_421),
.Y(n_462)
);

OAI21xp5_ASAP7_75t_SL g463 ( 
.A1(n_462),
.A2(n_445),
.B(n_362),
.Y(n_463)
);

OAI221xp5_ASAP7_75t_R g464 ( 
.A1(n_463),
.A2(n_131),
.B1(n_133),
.B2(n_138),
.C(n_145),
.Y(n_464)
);


endmodule