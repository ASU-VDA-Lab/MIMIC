module real_aes_14945_n_8 (n_4, n_0, n_3, n_5, n_2, n_7, n_6, n_1, n_8);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_7;
input n_6;
input n_1;
output n_8;
wire n_28;
wire n_17;
wire n_22;
wire n_13;
wire n_24;
wire n_12;
wire n_19;
wire n_25;
wire n_32;
wire n_30;
wire n_14;
wire n_11;
wire n_16;
wire n_15;
wire n_27;
wire n_23;
wire n_9;
wire n_29;
wire n_20;
wire n_18;
wire n_26;
wire n_21;
wire n_31;
wire n_10;
wire n_33;
BUFx10_ASAP7_75t_L g20 ( .A(n_0), .Y(n_20) );
HB1xp67_ASAP7_75t_L g16 ( .A(n_1), .Y(n_16) );
INVx1_ASAP7_75t_L g23 ( .A(n_2), .Y(n_23) );
INVx1_ASAP7_75t_L g33 ( .A(n_3), .Y(n_33) );
HB1xp67_ASAP7_75t_L g27 ( .A(n_4), .Y(n_27) );
INVx1_ASAP7_75t_L g13 ( .A(n_5), .Y(n_13) );
HB1xp67_ASAP7_75t_L g18 ( .A(n_6), .Y(n_18) );
AND2x4_ASAP7_75t_L g22 ( .A(n_7), .B(n_23), .Y(n_22) );
INVx1_ASAP7_75t_L g30 ( .A(n_7), .Y(n_30) );
AOI31xp33_ASAP7_75t_L g8 ( .A1(n_9), .A2(n_14), .A3(n_27), .B(n_28), .Y(n_8) );
INVxp67_ASAP7_75t_L g9 ( .A(n_10), .Y(n_9) );
BUFx6f_ASAP7_75t_SL g10 ( .A(n_11), .Y(n_10) );
INVx1_ASAP7_75t_L g11 ( .A(n_12), .Y(n_11) );
BUFx2_ASAP7_75t_L g12 ( .A(n_13), .Y(n_12) );
OAI22xp33_ASAP7_75t_L g14 ( .A1(n_15), .A2(n_19), .B1(n_24), .B2(n_25), .Y(n_14) );
NAND2xp5_ASAP7_75t_L g15 ( .A(n_16), .B(n_17), .Y(n_15) );
NAND2xp5_ASAP7_75t_L g24 ( .A(n_16), .B(n_18), .Y(n_24) );
INVx1_ASAP7_75t_L g17 ( .A(n_18), .Y(n_17) );
OR2x6_ASAP7_75t_SL g19 ( .A(n_20), .B(n_21), .Y(n_19) );
NAND2xp5_ASAP7_75t_L g26 ( .A(n_20), .B(n_22), .Y(n_26) );
INVx1_ASAP7_75t_L g21 ( .A(n_22), .Y(n_21) );
HB1xp67_ASAP7_75t_L g31 ( .A(n_23), .Y(n_31) );
BUFx2_ASAP7_75t_L g25 ( .A(n_26), .Y(n_25) );
INVx1_ASAP7_75t_L g28 ( .A(n_29), .Y(n_28) );
NAND3xp33_ASAP7_75t_SL g29 ( .A(n_30), .B(n_31), .C(n_32), .Y(n_29) );
INVx1_ASAP7_75t_L g32 ( .A(n_33), .Y(n_32) );
endmodule