module real_jpeg_15086_n_16 (n_5, n_4, n_8, n_0, n_12, n_274, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_274;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_215;
wire n_176;
wire n_166;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_238;
wire n_76;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_137;
wire n_31;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_74;
wire n_70;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_225;
wire n_103;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_216;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_89;

BUFx2_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx4f_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_2),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_3),
.A2(n_43),
.B1(n_44),
.B2(n_46),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_3),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_3),
.A2(n_46),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_3),
.A2(n_29),
.B1(n_33),
.B2(n_46),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_4),
.A2(n_73),
.B1(n_74),
.B2(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_4),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_4),
.A2(n_61),
.B1(n_62),
.B2(n_134),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_4),
.A2(n_43),
.B1(n_44),
.B2(n_134),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_L g230 ( 
.A1(n_4),
.A2(n_29),
.B1(n_33),
.B2(n_134),
.Y(n_230)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_6),
.A2(n_73),
.B1(n_74),
.B2(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_6),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_6),
.A2(n_61),
.B1(n_62),
.B2(n_81),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_6),
.A2(n_43),
.B1(n_44),
.B2(n_81),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_6),
.A2(n_29),
.B1(n_33),
.B2(n_81),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_7),
.A2(n_73),
.B1(n_74),
.B2(n_159),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_7),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_7),
.A2(n_61),
.B1(n_62),
.B2(n_159),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_7),
.A2(n_43),
.B1(n_44),
.B2(n_159),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_7),
.A2(n_29),
.B1(n_33),
.B2(n_159),
.Y(n_238)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_8),
.Y(n_62)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_9),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_10),
.A2(n_43),
.B1(n_44),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_10),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_10),
.A2(n_55),
.B1(n_61),
.B2(n_62),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_10),
.A2(n_29),
.B1(n_33),
.B2(n_55),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_11),
.A2(n_29),
.B1(n_33),
.B2(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_11),
.A2(n_37),
.B1(n_61),
.B2(n_62),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_11),
.A2(n_37),
.B1(n_43),
.B2(n_44),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_11),
.A2(n_37),
.B1(n_73),
.B2(n_74),
.Y(n_113)
);

BUFx8_ASAP7_75t_L g72 ( 
.A(n_12),
.Y(n_72)
);

O2A1O1Ixp33_ASAP7_75t_L g148 ( 
.A1(n_13),
.A2(n_72),
.B(n_73),
.C(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_13),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_13),
.A2(n_73),
.B1(n_74),
.B2(n_150),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_13),
.B(n_83),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_13),
.A2(n_43),
.B1(n_44),
.B2(n_150),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_13),
.A2(n_101),
.B1(n_102),
.B2(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_13),
.B(n_89),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_14),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_14),
.A2(n_32),
.B1(n_73),
.B2(n_74),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_14),
.A2(n_32),
.B1(n_43),
.B2(n_44),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_14),
.A2(n_32),
.B1(n_61),
.B2(n_62),
.Y(n_130)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_137),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_135),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_115),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_19),
.B(n_115),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_85),
.B2(n_114),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_56),
.C(n_68),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_22),
.A2(n_23),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_39),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_24),
.A2(n_25),
.B1(n_39),
.B2(n_40),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_34),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_26),
.A2(n_101),
.B(n_232),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_28),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_33),
.Y(n_38)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_27),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_27),
.A2(n_38),
.B1(n_125),
.B2(n_146),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_27),
.A2(n_38),
.B1(n_229),
.B2(n_231),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_28),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_28),
.A2(n_38),
.B(n_127),
.Y(n_203)
);

CKINVDCx6p67_ASAP7_75t_R g33 ( 
.A(n_29),
.Y(n_33)
);

OA22x2_ASAP7_75t_L g52 ( 
.A1(n_29),
.A2(n_33),
.B1(n_49),
.B2(n_50),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_33),
.B(n_50),
.C(n_150),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_33),
.B(n_236),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_34),
.A2(n_102),
.B(n_147),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_38),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_36),
.B(n_102),
.Y(n_127)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_38),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_47),
.B1(n_53),
.B2(n_54),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_42),
.A2(n_52),
.B(n_94),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_43),
.A2(n_44),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

OA22x2_ASAP7_75t_SL g57 ( 
.A1(n_43),
.A2(n_44),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

O2A1O1Ixp33_ASAP7_75t_SL g199 ( 
.A1(n_43),
.A2(n_58),
.B(n_200),
.C(n_202),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_43),
.B(n_222),
.Y(n_221)
);

INVx6_ASAP7_75t_SL g43 ( 
.A(n_44),
.Y(n_43)
);

NOR3xp33_ASAP7_75t_L g202 ( 
.A(n_44),
.B(n_59),
.C(n_61),
.Y(n_202)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_47),
.B(n_95),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_47),
.A2(n_54),
.B(n_106),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_47),
.A2(n_93),
.B(n_106),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_47),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_47),
.A2(n_53),
.B1(n_207),
.B2(n_215),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_47),
.A2(n_53),
.B1(n_224),
.B2(n_225),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_47),
.A2(n_53),
.B1(n_215),
.B2(n_225),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_52),
.Y(n_47)
);

CKINVDCx14_ASAP7_75t_SL g49 ( 
.A(n_50),
.Y(n_49)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_52),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_52),
.B(n_96),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_52),
.B(n_150),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_53),
.B(n_93),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_56),
.B(n_68),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_60),
.B(n_63),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_57),
.B(n_67),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_57),
.A2(n_154),
.B1(n_187),
.B2(n_189),
.Y(n_186)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_58),
.A2(n_59),
.B1(n_61),
.B2(n_62),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_60),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_61),
.A2(n_62),
.B1(n_72),
.B2(n_77),
.Y(n_78)
);

OAI21xp33_ASAP7_75t_L g149 ( 
.A1(n_61),
.A2(n_77),
.B(n_150),
.Y(n_149)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

HAxp5_ASAP7_75t_SL g201 ( 
.A(n_62),
.B(n_150),
.CON(n_201),
.SN(n_201)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_64),
.B(n_66),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_64),
.A2(n_88),
.B1(n_89),
.B2(n_90),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_64),
.A2(n_130),
.B(n_131),
.Y(n_129)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_64),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_64),
.A2(n_89),
.B1(n_153),
.B2(n_172),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_64),
.A2(n_89),
.B1(n_188),
.B2(n_201),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_69),
.A2(n_79),
.B(n_82),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_69),
.A2(n_111),
.B(n_112),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_69),
.A2(n_78),
.B1(n_157),
.B2(n_160),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_70),
.A2(n_80),
.B1(n_83),
.B2(n_133),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_70),
.A2(n_83),
.B1(n_158),
.B2(n_174),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_78),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_73),
.B1(n_74),
.B2(n_77),
.Y(n_71)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_72),
.Y(n_77)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_84),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_83),
.B(n_113),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_84),
.Y(n_111)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_85),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_98),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_91),
.B(n_97),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_87),
.B(n_91),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_89),
.B(n_130),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_94),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_92),
.A2(n_205),
.B(n_206),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_107),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_104),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_100),
.A2(n_108),
.B1(n_109),
.B2(n_110),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_100),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_100),
.A2(n_104),
.B1(n_105),
.B2(n_108),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_102),
.B(n_103),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_101),
.A2(n_124),
.B(n_126),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_101),
.A2(n_102),
.B1(n_230),
.B2(n_238),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_102),
.B(n_150),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_120),
.C(n_121),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_116),
.A2(n_117),
.B1(n_120),
.B2(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_120),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_121),
.B(n_270),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_129),
.C(n_132),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_122),
.B(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_128),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_123),
.B(n_128),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_129),
.B(n_132),
.Y(n_164)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_133),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_267),
.B(n_272),
.Y(n_137)
);

AOI221xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_176),
.B1(n_192),
.B2(n_266),
.C(n_274),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_140),
.B(n_165),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_140),
.B(n_165),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_161),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_141),
.B(n_162),
.C(n_163),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_151),
.C(n_156),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_142),
.A2(n_143),
.B1(n_167),
.B2(n_168),
.Y(n_166)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_148),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_144),
.A2(n_145),
.B1(n_148),
.B2(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_148),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g168 ( 
.A(n_151),
.B(n_156),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_154),
.B(n_155),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_163),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_169),
.C(n_175),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_166),
.B(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_169),
.B(n_175),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.C(n_173),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_170),
.B(n_171),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_172),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_173),
.B(n_179),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_190),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_177),
.B(n_190),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_180),
.C(n_182),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_178),
.B(n_262),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_180),
.B(n_182),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.C(n_186),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_183),
.A2(n_184),
.B1(n_185),
.B2(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_183),
.Y(n_210)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_186),
.B(n_209),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_265),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_194),
.A2(n_260),
.B(n_264),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_216),
.B(n_259),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_196),
.B(n_211),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_196),
.B(n_211),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_208),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_204),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_198),
.B(n_204),
.C(n_208),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_203),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_199),
.B(n_203),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.C(n_214),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_212),
.B(n_256),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_213),
.B(n_214),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_217),
.A2(n_254),
.B(n_258),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_244),
.B(n_253),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_233),
.B(n_243),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_220),
.B(n_228),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_220),
.B(n_228),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_223),
.B1(n_226),
.B2(n_227),
.Y(n_220)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_221),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_223),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_223),
.B(n_226),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_239),
.B(n_242),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_237),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_240),
.B(n_241),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_245),
.B(n_246),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_247),
.B(n_249),
.C(n_252),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_250),
.B1(n_251),
.B2(n_252),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_251),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_255),
.B(n_257),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_255),
.B(n_257),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_261),
.B(n_263),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_261),
.B(n_263),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_268),
.B(n_269),
.Y(n_272)
);


endmodule