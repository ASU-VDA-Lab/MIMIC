module fake_jpeg_18418_n_157 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_157);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_157;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_93;
wire n_91;
wire n_54;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_1),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_18),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_19),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_7),
.Y(n_56)
);

INVx11_ASAP7_75t_SL g57 ( 
.A(n_1),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_39),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_11),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_12),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_15),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_0),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_45),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_10),
.Y(n_66)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

AOI21xp33_ASAP7_75t_L g69 ( 
.A1(n_37),
.A2(n_7),
.B(n_36),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_2),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_0),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_4),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_13),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_17),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_74),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_74),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_75),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_80),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

INVx3_ASAP7_75t_SL g86 ( 
.A(n_81),
.Y(n_86)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_83),
.Y(n_90)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_80),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_85),
.B(n_88),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_77),
.B(n_47),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_80),
.A2(n_56),
.B1(n_67),
.B2(n_59),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_92),
.A2(n_73),
.B1(n_65),
.B2(n_53),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_95),
.A2(n_48),
.B1(n_61),
.B2(n_62),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_86),
.A2(n_72),
.B1(n_70),
.B2(n_71),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_96),
.A2(n_98),
.B1(n_100),
.B2(n_106),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_87),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_97),
.B(n_93),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_86),
.A2(n_72),
.B1(n_70),
.B2(n_63),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

O2A1O1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_92),
.A2(n_94),
.B(n_91),
.C(n_89),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_101),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_90),
.A2(n_46),
.B1(n_58),
.B2(n_60),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_102),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_84),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_103),
.B(n_48),
.Y(n_110)
);

AOI21xp33_ASAP7_75t_L g104 ( 
.A1(n_84),
.A2(n_69),
.B(n_68),
.Y(n_104)
);

FAx1_ASAP7_75t_SL g122 ( 
.A(n_104),
.B(n_3),
.CI(n_4),
.CON(n_122),
.SN(n_122)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_93),
.A2(n_51),
.B1(n_52),
.B2(n_64),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_105),
.B(n_55),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_107),
.A2(n_120),
.B(n_122),
.Y(n_130)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_108),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_97),
.B(n_65),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_109),
.B(n_110),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_66),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_112),
.B(n_115),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_114),
.A2(n_119),
.B1(n_27),
.B2(n_42),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_101),
.B(n_54),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_50),
.Y(n_116)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_116),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_105),
.B(n_49),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_118),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_100),
.A2(n_24),
.B1(n_44),
.B2(n_43),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_105),
.B(n_2),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_101),
.Y(n_121)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_121),
.Y(n_126)
);

NAND2x1_ASAP7_75t_SL g127 ( 
.A(n_123),
.B(n_5),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g137 ( 
.A(n_127),
.Y(n_137)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_117),
.Y(n_128)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_128),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_113),
.Y(n_131)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_131),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_123),
.A2(n_5),
.B(n_6),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_134),
.A2(n_135),
.B1(n_8),
.B2(n_9),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_124),
.A2(n_111),
.B1(n_107),
.B2(n_114),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_138),
.A2(n_142),
.B1(n_133),
.B2(n_125),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_129),
.B(n_122),
.C(n_113),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_140),
.B(n_130),
.C(n_134),
.Y(n_145)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_126),
.Y(n_141)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_141),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_143),
.B(n_145),
.C(n_140),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_145),
.C(n_139),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_144),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_136),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_132),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_133),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_137),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_137),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_153),
.B(n_127),
.Y(n_154)
);

AOI322xp5_ASAP7_75t_L g155 ( 
.A1(n_154),
.A2(n_26),
.A3(n_40),
.B1(n_14),
.B2(n_16),
.C1(n_20),
.C2(n_21),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_155),
.A2(n_28),
.B(n_35),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_22),
.Y(n_157)
);


endmodule