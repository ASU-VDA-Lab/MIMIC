module fake_jpeg_24160_n_102 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_102);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_102;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_5),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_0),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx8_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_24),
.Y(n_25)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_24),
.B(n_0),
.C(n_2),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_20),
.C(n_16),
.Y(n_37)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_27),
.B(n_33),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_12),
.B(n_0),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_28),
.B(n_31),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_15),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_30),
.A2(n_23),
.B1(n_22),
.B2(n_21),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_12),
.B(n_4),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_32),
.B(n_34),
.Y(n_49)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_18),
.B(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_31),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_35),
.B(n_40),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g53 ( 
.A1(n_37),
.A2(n_24),
.B(n_23),
.Y(n_53)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_19),
.Y(n_42)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_43),
.A2(n_45),
.B(n_33),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_19),
.Y(n_44)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_26),
.B(n_22),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_48),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_25),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_47),
.Y(n_62)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_25),
.B(n_21),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_47),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_50),
.B(n_51),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_41),
.Y(n_51)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_53),
.B(n_65),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_54),
.B(n_57),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_55),
.A2(n_56),
.B1(n_39),
.B2(n_36),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_37),
.A2(n_39),
.B1(n_46),
.B2(n_36),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_40),
.A2(n_20),
.B1(n_16),
.B2(n_13),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_58),
.A2(n_38),
.B1(n_14),
.B2(n_17),
.Y(n_69)
);

AND2x2_ASAP7_75t_SL g59 ( 
.A(n_35),
.B(n_29),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_59),
.B(n_60),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_29),
.Y(n_60)
);

OAI32xp33_ASAP7_75t_L g65 ( 
.A1(n_49),
.A2(n_14),
.A3(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_66),
.B(n_67),
.Y(n_80)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_75),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_52),
.A2(n_39),
.B1(n_17),
.B2(n_9),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_71),
.A2(n_57),
.B1(n_56),
.B2(n_55),
.Y(n_82)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_74),
.Y(n_77)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_60),
.A2(n_6),
.B1(n_7),
.B2(n_10),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_76),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_72),
.B(n_52),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_59),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_82),
.B(n_84),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_72),
.A2(n_54),
.B(n_53),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_83),
.B(n_73),
.Y(n_87)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

INVxp67_ASAP7_75t_SL g85 ( 
.A(n_77),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_74),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_83),
.B(n_70),
.C(n_73),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_86),
.B(n_87),
.Y(n_93)
);

AOI322xp5_ASAP7_75t_L g88 ( 
.A1(n_80),
.A2(n_59),
.A3(n_69),
.B1(n_65),
.B2(n_76),
.C1(n_71),
.C2(n_64),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_88),
.A2(n_90),
.B(n_78),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_91),
.B(n_86),
.C(n_87),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_92),
.B(n_94),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_89),
.B(n_64),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_96),
.B(n_81),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_SL g97 ( 
.A(n_93),
.B(n_82),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_97),
.B(n_90),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_98),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_100),
.A2(n_81),
.B1(n_99),
.B2(n_95),
.Y(n_101)
);

AOI221xp5_ASAP7_75t_L g102 ( 
.A1(n_101),
.A2(n_79),
.B1(n_92),
.B2(n_63),
.C(n_6),
.Y(n_102)
);


endmodule