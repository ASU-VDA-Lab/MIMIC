module fake_jpeg_24362_n_257 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_257);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_257;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx6_ASAP7_75t_SL g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx6_ASAP7_75t_SL g27 ( 
.A(n_1),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_29),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_31),
.Y(n_42)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_17),
.B(n_0),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_17),
.Y(n_47)
);

BUFx8_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_34),
.B(n_28),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_6),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_35),
.B(n_19),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_39),
.A2(n_21),
.B1(n_29),
.B2(n_20),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_41),
.A2(n_50),
.B1(n_57),
.B2(n_14),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_33),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_45),
.B(n_47),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_52),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_35),
.B(n_19),
.Y(n_48)
);

OAI21xp33_ASAP7_75t_L g76 ( 
.A1(n_48),
.A2(n_54),
.B(n_56),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_39),
.A2(n_21),
.B1(n_29),
.B2(n_20),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_51),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_27),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_19),
.Y(n_54)
);

OAI21xp33_ASAP7_75t_SL g56 ( 
.A1(n_36),
.A2(n_26),
.B(n_14),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_30),
.A2(n_21),
.B1(n_29),
.B2(n_20),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_58),
.B(n_18),
.Y(n_64)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_59),
.B(n_62),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_45),
.A2(n_28),
.B1(n_31),
.B2(n_26),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_60),
.A2(n_71),
.B(n_73),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_61),
.A2(n_67),
.B1(n_68),
.B2(n_69),
.Y(n_81)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_64),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_65),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_L g67 ( 
.A1(n_41),
.A2(n_20),
.B1(n_27),
.B2(n_22),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_47),
.A2(n_17),
.B1(n_18),
.B2(n_16),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_44),
.A2(n_18),
.B1(n_15),
.B2(n_16),
.Y(n_69)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_56),
.A2(n_25),
.B1(n_15),
.B2(n_16),
.Y(n_71)
);

AND2x4_ASAP7_75t_L g73 ( 
.A(n_52),
.B(n_34),
.Y(n_73)
);

FAx1_ASAP7_75t_SL g74 ( 
.A(n_41),
.B(n_38),
.CI(n_32),
.CON(n_74),
.SN(n_74)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_74),
.B(n_79),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_75),
.Y(n_95)
);

A2O1A1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_52),
.A2(n_22),
.B(n_27),
.C(n_15),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_46),
.Y(n_83)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_49),
.C(n_42),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_84),
.B(n_76),
.C(n_77),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_54),
.Y(n_85)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_85),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_48),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_87),
.B(n_74),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_61),
.A2(n_51),
.B1(n_50),
.B2(n_57),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_88),
.A2(n_93),
.B1(n_100),
.B2(n_81),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_68),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_92),
.Y(n_104)
);

OA21x2_ASAP7_75t_L g90 ( 
.A1(n_73),
.A2(n_38),
.B(n_32),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_90),
.A2(n_79),
.B(n_74),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_64),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_73),
.A2(n_58),
.B1(n_40),
.B2(n_49),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_72),
.B(n_42),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_94),
.B(n_98),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_69),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_96),
.Y(n_105)
);

OA22x2_ASAP7_75t_L g97 ( 
.A1(n_73),
.A2(n_43),
.B1(n_53),
.B2(n_24),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_97),
.A2(n_70),
.B1(n_77),
.B2(n_43),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_23),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_23),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_101),
.B(n_86),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_80),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_103),
.B(n_107),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_80),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_82),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_108),
.B(n_115),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_109),
.A2(n_116),
.B1(n_117),
.B2(n_105),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_87),
.B(n_91),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_111),
.B(n_112),
.C(n_114),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_113),
.B(n_118),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_84),
.B(n_100),
.C(n_91),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_82),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_89),
.A2(n_96),
.B1(n_88),
.B2(n_81),
.Y(n_116)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_99),
.Y(n_119)
);

INVx11_ASAP7_75t_L g130 ( 
.A(n_119),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_94),
.B(n_65),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_120),
.B(n_123),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_121),
.A2(n_97),
.B1(n_22),
.B2(n_95),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_122),
.B(n_90),
.Y(n_129)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_101),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_111),
.B(n_85),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_124),
.B(n_143),
.C(n_137),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_116),
.A2(n_90),
.B1(n_97),
.B2(n_83),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_126),
.A2(n_131),
.B1(n_132),
.B2(n_108),
.Y(n_148)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_113),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_128),
.Y(n_150)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_120),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_129),
.B(n_16),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_105),
.A2(n_90),
.B1(n_97),
.B2(n_92),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_102),
.B(n_86),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_133),
.B(n_136),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_135),
.A2(n_24),
.B1(n_23),
.B2(n_7),
.Y(n_166)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_107),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_109),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_138),
.B(n_140),
.Y(n_167)
);

A2O1A1Ixp33_ASAP7_75t_SL g139 ( 
.A1(n_117),
.A2(n_97),
.B(n_104),
.C(n_115),
.Y(n_139)
);

OA22x2_ASAP7_75t_L g162 ( 
.A1(n_139),
.A2(n_75),
.B1(n_24),
.B2(n_25),
.Y(n_162)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_119),
.Y(n_140)
);

INVx13_ASAP7_75t_L g141 ( 
.A(n_118),
.Y(n_141)
);

INVx11_ASAP7_75t_L g163 ( 
.A(n_141),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_114),
.A2(n_25),
.B(n_99),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_112),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_122),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_146),
.B(n_152),
.C(n_158),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_142),
.B(n_110),
.Y(n_147)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_147),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_148),
.A2(n_161),
.B1(n_164),
.B2(n_130),
.Y(n_177)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_136),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_149),
.B(n_165),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_125),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_151),
.B(n_154),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_135),
.A2(n_102),
.B1(n_106),
.B2(n_123),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_153),
.A2(n_157),
.B1(n_166),
.B2(n_139),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_134),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_142),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_155),
.B(n_156),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_144),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_138),
.A2(n_106),
.B1(n_110),
.B2(n_99),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_144),
.B(n_65),
.Y(n_160)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_160),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_126),
.A2(n_63),
.B1(n_62),
.B2(n_59),
.Y(n_161)
);

AO22x1_ASAP7_75t_L g182 ( 
.A1(n_162),
.A2(n_139),
.B1(n_130),
.B2(n_143),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_132),
.A2(n_75),
.B1(n_24),
.B2(n_23),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_140),
.Y(n_165)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_160),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_172),
.B(n_174),
.Y(n_192)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_150),
.Y(n_174)
);

FAx1_ASAP7_75t_SL g175 ( 
.A(n_147),
.B(n_137),
.CI(n_129),
.CON(n_175),
.SN(n_175)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_175),
.B(n_177),
.Y(n_197)
);

AOI21x1_ASAP7_75t_L g176 ( 
.A1(n_157),
.A2(n_139),
.B(n_141),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_176),
.A2(n_182),
.B1(n_162),
.B2(n_1),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_152),
.B(n_124),
.C(n_145),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_179),
.B(n_180),
.C(n_148),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_146),
.B(n_158),
.C(n_156),
.Y(n_180)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_181),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_154),
.B(n_6),
.Y(n_183)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_183),
.Y(n_191)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_159),
.Y(n_184)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_184),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_163),
.B(n_7),
.Y(n_185)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_185),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_167),
.Y(n_186)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_186),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_153),
.B(n_5),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_187),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_188),
.B(n_173),
.C(n_172),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_179),
.B(n_149),
.C(n_161),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_189),
.B(n_193),
.C(n_199),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_169),
.B(n_180),
.C(n_171),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_182),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_198),
.B(n_162),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_169),
.B(n_165),
.C(n_164),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_171),
.B(n_166),
.C(n_163),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_200),
.B(n_184),
.C(n_173),
.Y(n_211)
);

NOR2xp67_ASAP7_75t_L g202 ( 
.A(n_182),
.B(n_162),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_202),
.B(n_170),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_203),
.B(n_181),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_192),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_205),
.B(n_212),
.Y(n_226)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_206),
.Y(n_222)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_207),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_199),
.B(n_189),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_208),
.B(n_191),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_209),
.B(n_210),
.C(n_211),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_193),
.B(n_188),
.C(n_197),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_196),
.B(n_174),
.Y(n_212)
);

FAx1_ASAP7_75t_SL g213 ( 
.A(n_200),
.B(n_176),
.CI(n_168),
.CON(n_213),
.SN(n_213)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_213),
.B(n_215),
.Y(n_225)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_214),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_201),
.B(n_178),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_190),
.B(n_168),
.C(n_175),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_216),
.B(n_8),
.C(n_12),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_203),
.B(n_175),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_217),
.B(n_5),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_211),
.A2(n_195),
.B(n_194),
.Y(n_218)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_218),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_220),
.B(n_223),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_221),
.B(n_224),
.C(n_8),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_204),
.B(n_0),
.C(n_2),
.Y(n_224)
);

NOR2xp67_ASAP7_75t_SL g229 ( 
.A(n_225),
.B(n_204),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_229),
.A2(n_234),
.B(n_236),
.Y(n_243)
);

AO21x1_ASAP7_75t_L g230 ( 
.A1(n_227),
.A2(n_207),
.B(n_213),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_230),
.B(n_232),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_222),
.A2(n_216),
.B1(n_217),
.B2(n_9),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_231),
.A2(n_4),
.B1(n_9),
.B2(n_10),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_226),
.B(n_4),
.Y(n_234)
);

NOR2xp67_ASAP7_75t_SL g236 ( 
.A(n_219),
.B(n_4),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_228),
.B(n_0),
.Y(n_237)
);

INVxp33_ASAP7_75t_L g239 ( 
.A(n_237),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_235),
.A2(n_219),
.B(n_221),
.Y(n_238)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_238),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_233),
.B(n_224),
.C(n_223),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_240),
.B(n_244),
.C(n_237),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_242),
.B(n_13),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_230),
.B(n_10),
.C(n_13),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_245),
.B(n_247),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_241),
.A2(n_10),
.B(n_13),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_246),
.A2(n_239),
.B(n_2),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_243),
.B(n_0),
.Y(n_247)
);

NOR3xp33_ASAP7_75t_L g251 ( 
.A(n_249),
.B(n_239),
.C(n_2),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_251),
.Y(n_254)
);

OAI21x1_ASAP7_75t_L g253 ( 
.A1(n_252),
.A2(n_247),
.B(n_245),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_253),
.B(n_250),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_255),
.A2(n_248),
.B1(n_254),
.B2(n_3),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_256),
.B(n_3),
.Y(n_257)
);


endmodule