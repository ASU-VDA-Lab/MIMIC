module real_aes_7955_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_349;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g107 ( .A(n_0), .B(n_86), .C(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g451 ( .A(n_0), .Y(n_451) );
A2O1A1Ixp33_ASAP7_75t_L g214 ( .A1(n_1), .A2(n_130), .B(n_134), .C(n_215), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_2), .A2(n_164), .B(n_242), .Y(n_241) );
INVx1_ASAP7_75t_L g509 ( .A(n_3), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_4), .B(n_231), .Y(n_250) );
AOI21xp33_ASAP7_75t_L g474 ( .A1(n_5), .A2(n_164), .B(n_475), .Y(n_474) );
AND2x6_ASAP7_75t_L g130 ( .A(n_6), .B(n_131), .Y(n_130) );
INVx1_ASAP7_75t_L g205 ( .A(n_7), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g105 ( .A(n_8), .B(n_42), .Y(n_105) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_9), .A2(n_163), .B(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_10), .B(n_142), .Y(n_217) );
INVx1_ASAP7_75t_L g479 ( .A(n_11), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_12), .B(n_245), .Y(n_534) );
INVx1_ASAP7_75t_L g150 ( .A(n_13), .Y(n_150) );
INVx1_ASAP7_75t_L g546 ( .A(n_14), .Y(n_546) );
A2O1A1Ixp33_ASAP7_75t_L g226 ( .A1(n_15), .A2(n_140), .B(n_227), .C(n_229), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_16), .B(n_231), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_17), .B(n_497), .Y(n_560) );
NAND2xp5_ASAP7_75t_SL g519 ( .A(n_18), .B(n_164), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_19), .B(n_176), .Y(n_175) );
A2O1A1Ixp33_ASAP7_75t_L g259 ( .A1(n_20), .A2(n_245), .B(n_260), .C(n_262), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_21), .B(n_231), .Y(n_500) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_22), .B(n_142), .Y(n_187) );
A2O1A1Ixp33_ASAP7_75t_L g544 ( .A1(n_23), .A2(n_172), .B(n_229), .C(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_SL g141 ( .A(n_24), .B(n_142), .Y(n_141) );
CKINVDCx16_ASAP7_75t_R g181 ( .A(n_25), .Y(n_181) );
INVx1_ASAP7_75t_L g138 ( .A(n_26), .Y(n_138) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_27), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g213 ( .A(n_28), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_29), .B(n_142), .Y(n_510) );
OAI22xp5_ASAP7_75t_SL g740 ( .A1(n_30), .A2(n_31), .B1(n_741), .B2(n_742), .Y(n_740) );
INVx1_ASAP7_75t_L g742 ( .A(n_30), .Y(n_742) );
CKINVDCx20_ASAP7_75t_R g741 ( .A(n_31), .Y(n_741) );
INVx1_ASAP7_75t_L g170 ( .A(n_32), .Y(n_170) );
INVx1_ASAP7_75t_L g488 ( .A(n_33), .Y(n_488) );
AOI222xp33_ASAP7_75t_L g457 ( .A1(n_34), .A2(n_458), .B1(n_740), .B2(n_743), .C1(n_746), .C2(n_747), .Y(n_457) );
INVx2_ASAP7_75t_L g128 ( .A(n_35), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g219 ( .A(n_36), .Y(n_219) );
A2O1A1Ixp33_ASAP7_75t_L g244 ( .A1(n_37), .A2(n_245), .B(n_246), .C(n_248), .Y(n_244) );
INVxp67_ASAP7_75t_L g171 ( .A(n_38), .Y(n_171) );
A2O1A1Ixp33_ASAP7_75t_L g133 ( .A1(n_39), .A2(n_134), .B(n_137), .C(n_145), .Y(n_133) );
CKINVDCx14_ASAP7_75t_R g243 ( .A(n_40), .Y(n_243) );
A2O1A1Ixp33_ASAP7_75t_L g520 ( .A1(n_41), .A2(n_130), .B(n_134), .C(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g487 ( .A(n_43), .Y(n_487) );
A2O1A1Ixp33_ASAP7_75t_L g202 ( .A1(n_44), .A2(n_189), .B(n_203), .C(n_204), .Y(n_202) );
NAND2xp5_ASAP7_75t_SL g559 ( .A(n_45), .B(n_142), .Y(n_559) );
CKINVDCx20_ASAP7_75t_R g152 ( .A(n_46), .Y(n_152) );
CKINVDCx20_ASAP7_75t_R g166 ( .A(n_47), .Y(n_166) );
NAND2xp5_ASAP7_75t_SL g452 ( .A(n_48), .B(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g258 ( .A(n_49), .Y(n_258) );
CKINVDCx16_ASAP7_75t_R g489 ( .A(n_50), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_51), .B(n_164), .Y(n_536) );
AOI22xp5_ASAP7_75t_L g101 ( .A1(n_52), .A2(n_102), .B1(n_111), .B2(n_752), .Y(n_101) );
AOI22xp5_ASAP7_75t_L g485 ( .A1(n_53), .A2(n_134), .B1(n_262), .B2(n_486), .Y(n_485) );
CKINVDCx20_ASAP7_75t_R g525 ( .A(n_54), .Y(n_525) );
CKINVDCx16_ASAP7_75t_R g506 ( .A(n_55), .Y(n_506) );
CKINVDCx14_ASAP7_75t_R g201 ( .A(n_56), .Y(n_201) );
A2O1A1Ixp33_ASAP7_75t_L g477 ( .A1(n_57), .A2(n_203), .B(n_248), .C(n_478), .Y(n_477) );
CKINVDCx20_ASAP7_75t_R g562 ( .A(n_58), .Y(n_562) );
INVx1_ASAP7_75t_L g476 ( .A(n_59), .Y(n_476) );
AOI22xp5_ASAP7_75t_L g443 ( .A1(n_60), .A2(n_88), .B1(n_444), .B2(n_445), .Y(n_443) );
CKINVDCx20_ASAP7_75t_R g445 ( .A(n_60), .Y(n_445) );
INVx1_ASAP7_75t_L g131 ( .A(n_61), .Y(n_131) );
INVx1_ASAP7_75t_L g149 ( .A(n_62), .Y(n_149) );
INVx1_ASAP7_75t_SL g247 ( .A(n_63), .Y(n_247) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_64), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_65), .B(n_231), .Y(n_264) );
INVx1_ASAP7_75t_L g184 ( .A(n_66), .Y(n_184) );
A2O1A1Ixp33_ASAP7_75t_SL g496 ( .A1(n_67), .A2(n_248), .B(n_497), .C(n_498), .Y(n_496) );
INVxp67_ASAP7_75t_L g499 ( .A(n_68), .Y(n_499) );
INVx1_ASAP7_75t_L g110 ( .A(n_69), .Y(n_110) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_70), .A2(n_164), .B(n_200), .Y(n_199) );
CKINVDCx20_ASAP7_75t_R g193 ( .A(n_71), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_72), .A2(n_164), .B(n_224), .Y(n_223) );
CKINVDCx20_ASAP7_75t_R g491 ( .A(n_73), .Y(n_491) );
INVx1_ASAP7_75t_L g556 ( .A(n_74), .Y(n_556) );
AOI21xp5_ASAP7_75t_L g162 ( .A1(n_75), .A2(n_163), .B(n_165), .Y(n_162) );
CKINVDCx16_ASAP7_75t_R g132 ( .A(n_76), .Y(n_132) );
INVx1_ASAP7_75t_L g225 ( .A(n_77), .Y(n_225) );
A2O1A1Ixp33_ASAP7_75t_L g557 ( .A1(n_78), .A2(n_130), .B(n_134), .C(n_558), .Y(n_557) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_79), .A2(n_164), .B(n_257), .Y(n_256) );
INVx1_ASAP7_75t_L g228 ( .A(n_80), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_81), .B(n_139), .Y(n_522) );
INVx2_ASAP7_75t_L g147 ( .A(n_82), .Y(n_147) );
INVx1_ASAP7_75t_L g216 ( .A(n_83), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_84), .B(n_497), .Y(n_523) );
A2O1A1Ixp33_ASAP7_75t_L g507 ( .A1(n_85), .A2(n_130), .B(n_134), .C(n_508), .Y(n_507) );
OR2x2_ASAP7_75t_L g448 ( .A(n_86), .B(n_449), .Y(n_448) );
OR2x2_ASAP7_75t_L g461 ( .A(n_86), .B(n_450), .Y(n_461) );
INVx2_ASAP7_75t_L g465 ( .A(n_86), .Y(n_465) );
A2O1A1Ixp33_ASAP7_75t_L g182 ( .A1(n_87), .A2(n_134), .B(n_183), .C(n_191), .Y(n_182) );
CKINVDCx20_ASAP7_75t_R g444 ( .A(n_88), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_89), .B(n_146), .Y(n_480) );
CKINVDCx20_ASAP7_75t_R g513 ( .A(n_90), .Y(n_513) );
A2O1A1Ixp33_ASAP7_75t_L g531 ( .A1(n_91), .A2(n_130), .B(n_134), .C(n_532), .Y(n_531) );
CKINVDCx20_ASAP7_75t_R g538 ( .A(n_92), .Y(n_538) );
INVx1_ASAP7_75t_L g495 ( .A(n_93), .Y(n_495) );
CKINVDCx16_ASAP7_75t_R g543 ( .A(n_94), .Y(n_543) );
NAND2xp5_ASAP7_75t_SL g533 ( .A(n_95), .B(n_139), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_96), .B(n_154), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_97), .B(n_154), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_98), .B(n_110), .Y(n_109) );
INVx2_ASAP7_75t_L g261 ( .A(n_99), .Y(n_261) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_100), .A2(n_164), .B(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
CKINVDCx12_ASAP7_75t_R g754 ( .A(n_104), .Y(n_754) );
AND2x2_ASAP7_75t_L g104 ( .A(n_105), .B(n_106), .Y(n_104) );
AND2x2_ASAP7_75t_L g450 ( .A(n_105), .B(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
AO21x2_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_116), .B(n_456), .Y(n_111) );
HB1xp67_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx2_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx1_ASAP7_75t_L g751 ( .A(n_115), .Y(n_751) );
OAI21xp5_ASAP7_75t_SL g116 ( .A1(n_117), .A2(n_446), .B(n_452), .Y(n_116) );
XOR2xp5_ASAP7_75t_L g117 ( .A(n_118), .B(n_443), .Y(n_117) );
OAI22xp5_ASAP7_75t_L g458 ( .A1(n_118), .A2(n_459), .B1(n_462), .B2(n_466), .Y(n_458) );
INVx1_ASAP7_75t_L g744 ( .A(n_118), .Y(n_744) );
OR4x2_ASAP7_75t_L g118 ( .A(n_119), .B(n_333), .C(n_380), .D(n_420), .Y(n_118) );
NAND3xp33_ASAP7_75t_SL g119 ( .A(n_120), .B(n_279), .C(n_308), .Y(n_119) );
AOI211xp5_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_194), .B(n_232), .C(n_272), .Y(n_120) );
O2A1O1Ixp33_ASAP7_75t_L g308 ( .A1(n_121), .A2(n_292), .B(n_309), .C(n_313), .Y(n_308) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g122 ( .A(n_123), .B(n_156), .Y(n_122) );
NAND2xp5_ASAP7_75t_SL g270 ( .A(n_123), .B(n_271), .Y(n_270) );
INVx3_ASAP7_75t_SL g275 ( .A(n_123), .Y(n_275) );
HB1xp67_ASAP7_75t_L g287 ( .A(n_123), .Y(n_287) );
AND2x4_ASAP7_75t_L g291 ( .A(n_123), .B(n_239), .Y(n_291) );
AND2x2_ASAP7_75t_L g302 ( .A(n_123), .B(n_179), .Y(n_302) );
OR2x2_ASAP7_75t_L g326 ( .A(n_123), .B(n_235), .Y(n_326) );
AND2x2_ASAP7_75t_L g339 ( .A(n_123), .B(n_240), .Y(n_339) );
AND2x2_ASAP7_75t_L g379 ( .A(n_123), .B(n_365), .Y(n_379) );
AND2x2_ASAP7_75t_L g386 ( .A(n_123), .B(n_349), .Y(n_386) );
AND2x2_ASAP7_75t_L g416 ( .A(n_123), .B(n_157), .Y(n_416) );
OR2x6_ASAP7_75t_L g123 ( .A(n_124), .B(n_151), .Y(n_123) );
O2A1O1Ixp33_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_132), .B(n_133), .C(n_146), .Y(n_124) );
OAI21xp5_ASAP7_75t_L g180 ( .A1(n_125), .A2(n_181), .B(n_182), .Y(n_180) );
OAI21xp5_ASAP7_75t_L g212 ( .A1(n_125), .A2(n_213), .B(n_214), .Y(n_212) );
OAI22xp33_ASAP7_75t_L g484 ( .A1(n_125), .A2(n_174), .B1(n_485), .B2(n_489), .Y(n_484) );
OAI21xp5_ASAP7_75t_L g505 ( .A1(n_125), .A2(n_506), .B(n_507), .Y(n_505) );
OAI21xp5_ASAP7_75t_L g555 ( .A1(n_125), .A2(n_556), .B(n_557), .Y(n_555) );
NAND2x1p5_ASAP7_75t_L g125 ( .A(n_126), .B(n_130), .Y(n_125) );
AND2x4_ASAP7_75t_L g164 ( .A(n_126), .B(n_130), .Y(n_164) );
AND2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_129), .Y(n_126) );
INVx1_ASAP7_75t_L g144 ( .A(n_127), .Y(n_144) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx2_ASAP7_75t_L g135 ( .A(n_128), .Y(n_135) );
INVx1_ASAP7_75t_L g263 ( .A(n_128), .Y(n_263) );
INVx1_ASAP7_75t_L g136 ( .A(n_129), .Y(n_136) );
INVx3_ASAP7_75t_L g140 ( .A(n_129), .Y(n_140) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_129), .Y(n_142) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_129), .Y(n_173) );
INVx1_ASAP7_75t_L g497 ( .A(n_129), .Y(n_497) );
BUFx3_ASAP7_75t_L g145 ( .A(n_130), .Y(n_145) );
INVx4_ASAP7_75t_SL g174 ( .A(n_130), .Y(n_174) );
INVx5_ASAP7_75t_L g167 ( .A(n_134), .Y(n_167) );
AND2x6_ASAP7_75t_L g134 ( .A(n_135), .B(n_136), .Y(n_134) );
BUFx3_ASAP7_75t_L g190 ( .A(n_135), .Y(n_190) );
BUFx6f_ASAP7_75t_L g249 ( .A(n_135), .Y(n_249) );
O2A1O1Ixp33_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_139), .B(n_141), .C(n_143), .Y(n_137) );
OAI22xp33_ASAP7_75t_L g169 ( .A1(n_139), .A2(n_170), .B1(n_171), .B2(n_172), .Y(n_169) );
O2A1O1Ixp33_ASAP7_75t_L g508 ( .A1(n_139), .A2(n_509), .B(n_510), .C(n_511), .Y(n_508) );
INVx5_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
NOR2xp33_ASAP7_75t_L g204 ( .A(n_140), .B(n_205), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g478 ( .A(n_140), .B(n_479), .Y(n_478) );
NOR2xp33_ASAP7_75t_L g498 ( .A(n_140), .B(n_499), .Y(n_498) );
INVx2_ASAP7_75t_L g203 ( .A(n_142), .Y(n_203) );
INVx4_ASAP7_75t_L g245 ( .A(n_142), .Y(n_245) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
NAND2xp5_ASAP7_75t_SL g168 ( .A(n_144), .B(n_169), .Y(n_168) );
INVx2_ASAP7_75t_L g177 ( .A(n_146), .Y(n_177) );
OA21x2_ASAP7_75t_L g198 ( .A1(n_146), .A2(n_199), .B(n_206), .Y(n_198) );
INVx1_ASAP7_75t_L g211 ( .A(n_146), .Y(n_211) );
OA21x2_ASAP7_75t_L g540 ( .A1(n_146), .A2(n_541), .B(n_547), .Y(n_540) );
AND2x2_ASAP7_75t_SL g146 ( .A(n_147), .B(n_148), .Y(n_146) );
AND2x2_ASAP7_75t_L g155 ( .A(n_147), .B(n_148), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_149), .B(n_150), .Y(n_148) );
NOR2xp33_ASAP7_75t_L g151 ( .A(n_152), .B(n_153), .Y(n_151) );
AO21x2_ASAP7_75t_L g179 ( .A1(n_153), .A2(n_180), .B(n_192), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_153), .B(n_219), .Y(n_218) );
INVx3_ASAP7_75t_L g231 ( .A(n_153), .Y(n_231) );
NOR2xp33_ASAP7_75t_SL g524 ( .A(n_153), .B(n_525), .Y(n_524) );
INVx4_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
HB1xp67_ASAP7_75t_L g222 ( .A(n_154), .Y(n_222) );
OA21x2_ASAP7_75t_L g492 ( .A1(n_154), .A2(n_493), .B(n_500), .Y(n_492) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx1_ASAP7_75t_L g161 ( .A(n_155), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_156), .B(n_343), .Y(n_355) );
AND2x2_ASAP7_75t_L g156 ( .A(n_157), .B(n_178), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_157), .B(n_286), .Y(n_285) );
OR2x2_ASAP7_75t_L g293 ( .A(n_157), .B(n_178), .Y(n_293) );
BUFx3_ASAP7_75t_L g301 ( .A(n_157), .Y(n_301) );
OR2x2_ASAP7_75t_L g322 ( .A(n_157), .B(n_197), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_157), .B(n_343), .Y(n_433) );
OA21x2_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_162), .B(n_175), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
AO21x2_ASAP7_75t_L g235 ( .A1(n_159), .A2(n_236), .B(n_237), .Y(n_235) );
AO21x2_ASAP7_75t_L g554 ( .A1(n_159), .A2(n_555), .B(n_561), .Y(n_554) );
INVx1_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
AOI21xp5_ASAP7_75t_SL g518 ( .A1(n_160), .A2(n_519), .B(n_520), .Y(n_518) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
AO21x2_ASAP7_75t_L g483 ( .A1(n_161), .A2(n_484), .B(n_490), .Y(n_483) );
NOR2xp33_ASAP7_75t_L g490 ( .A(n_161), .B(n_491), .Y(n_490) );
AO21x2_ASAP7_75t_L g504 ( .A1(n_161), .A2(n_505), .B(n_512), .Y(n_504) );
INVx1_ASAP7_75t_L g236 ( .A(n_162), .Y(n_236) );
BUFx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
O2A1O1Ixp33_ASAP7_75t_SL g165 ( .A1(n_166), .A2(n_167), .B(n_168), .C(n_174), .Y(n_165) );
O2A1O1Ixp33_ASAP7_75t_SL g200 ( .A1(n_167), .A2(n_174), .B(n_201), .C(n_202), .Y(n_200) );
O2A1O1Ixp33_ASAP7_75t_SL g224 ( .A1(n_167), .A2(n_174), .B(n_225), .C(n_226), .Y(n_224) );
O2A1O1Ixp33_ASAP7_75t_L g242 ( .A1(n_167), .A2(n_174), .B(n_243), .C(n_244), .Y(n_242) );
O2A1O1Ixp33_ASAP7_75t_SL g257 ( .A1(n_167), .A2(n_174), .B(n_258), .C(n_259), .Y(n_257) );
O2A1O1Ixp33_ASAP7_75t_L g475 ( .A1(n_167), .A2(n_174), .B(n_476), .C(n_477), .Y(n_475) );
O2A1O1Ixp33_ASAP7_75t_L g494 ( .A1(n_167), .A2(n_174), .B(n_495), .C(n_496), .Y(n_494) );
O2A1O1Ixp33_ASAP7_75t_L g542 ( .A1(n_167), .A2(n_174), .B(n_543), .C(n_544), .Y(n_542) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_172), .B(n_228), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g260 ( .A(n_172), .B(n_261), .Y(n_260) );
NOR2xp33_ASAP7_75t_L g545 ( .A(n_172), .B(n_546), .Y(n_545) );
INVx4_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx2_ASAP7_75t_L g186 ( .A(n_173), .Y(n_186) );
OAI22xp5_ASAP7_75t_SL g486 ( .A1(n_173), .A2(n_186), .B1(n_487), .B2(n_488), .Y(n_486) );
INVx1_ASAP7_75t_L g191 ( .A(n_174), .Y(n_191) );
INVx1_ASAP7_75t_L g237 ( .A(n_175), .Y(n_237) );
INVx1_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_177), .B(n_193), .Y(n_192) );
AO21x2_ASAP7_75t_L g529 ( .A1(n_177), .A2(n_530), .B(n_537), .Y(n_529) );
AND2x2_ASAP7_75t_L g238 ( .A(n_178), .B(n_239), .Y(n_238) );
INVx1_ASAP7_75t_L g286 ( .A(n_178), .Y(n_286) );
AND2x2_ASAP7_75t_L g349 ( .A(n_178), .B(n_240), .Y(n_349) );
AOI221xp5_ASAP7_75t_L g351 ( .A1(n_178), .A2(n_352), .B1(n_354), .B2(n_356), .C(n_357), .Y(n_351) );
AND2x2_ASAP7_75t_L g365 ( .A(n_178), .B(n_235), .Y(n_365) );
AND2x2_ASAP7_75t_L g391 ( .A(n_178), .B(n_275), .Y(n_391) );
INVx2_ASAP7_75t_SL g178 ( .A(n_179), .Y(n_178) );
AND2x2_ASAP7_75t_L g271 ( .A(n_179), .B(n_240), .Y(n_271) );
BUFx2_ASAP7_75t_L g405 ( .A(n_179), .Y(n_405) );
O2A1O1Ixp33_ASAP7_75t_L g183 ( .A1(n_184), .A2(n_185), .B(n_187), .C(n_188), .Y(n_183) );
O2A1O1Ixp5_ASAP7_75t_L g215 ( .A1(n_185), .A2(n_188), .B(n_216), .C(n_217), .Y(n_215) );
INVx2_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_188), .A2(n_522), .B(n_523), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g558 ( .A1(n_188), .A2(n_559), .B(n_560), .Y(n_558) );
INVx2_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVx1_ASAP7_75t_L g229 ( .A(n_190), .Y(n_229) );
INVx1_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
OAI32xp33_ASAP7_75t_L g371 ( .A1(n_195), .A2(n_332), .A3(n_346), .B1(n_372), .B2(n_373), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_196), .B(n_207), .Y(n_195) );
AND2x2_ASAP7_75t_L g312 ( .A(n_196), .B(n_254), .Y(n_312) );
INVx1_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
OR2x2_ASAP7_75t_L g294 ( .A(n_197), .B(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_197), .B(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g366 ( .A(n_197), .B(n_254), .Y(n_366) );
AND2x2_ASAP7_75t_L g377 ( .A(n_197), .B(n_269), .Y(n_377) );
BUFx3_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
OR2x2_ASAP7_75t_L g278 ( .A(n_198), .B(n_255), .Y(n_278) );
AND2x2_ASAP7_75t_L g282 ( .A(n_198), .B(n_255), .Y(n_282) );
AND2x2_ASAP7_75t_L g317 ( .A(n_198), .B(n_268), .Y(n_317) );
AND2x2_ASAP7_75t_L g324 ( .A(n_198), .B(n_220), .Y(n_324) );
OAI211xp5_ASAP7_75t_L g329 ( .A1(n_198), .A2(n_275), .B(n_286), .C(n_330), .Y(n_329) );
INVx2_ASAP7_75t_L g383 ( .A(n_198), .Y(n_383) );
NOR2xp33_ASAP7_75t_L g394 ( .A(n_198), .B(n_209), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_207), .B(n_266), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_207), .B(n_282), .Y(n_372) );
INVx1_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
OR2x2_ASAP7_75t_L g277 ( .A(n_208), .B(n_278), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_209), .B(n_220), .Y(n_208) );
AND2x2_ASAP7_75t_L g269 ( .A(n_209), .B(n_221), .Y(n_269) );
OR2x2_ASAP7_75t_L g284 ( .A(n_209), .B(n_221), .Y(n_284) );
AND2x2_ASAP7_75t_L g307 ( .A(n_209), .B(n_268), .Y(n_307) );
INVx1_ASAP7_75t_L g311 ( .A(n_209), .Y(n_311) );
AND2x2_ASAP7_75t_L g330 ( .A(n_209), .B(n_267), .Y(n_330) );
OAI22xp33_ASAP7_75t_L g340 ( .A1(n_209), .A2(n_295), .B1(n_341), .B2(n_342), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_209), .B(n_383), .Y(n_407) );
AND2x2_ASAP7_75t_L g422 ( .A(n_209), .B(n_282), .Y(n_422) );
INVx4_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
BUFx3_ASAP7_75t_L g252 ( .A(n_210), .Y(n_252) );
AND2x2_ASAP7_75t_L g296 ( .A(n_210), .B(n_221), .Y(n_296) );
AND2x2_ASAP7_75t_L g298 ( .A(n_210), .B(n_254), .Y(n_298) );
AND3x2_ASAP7_75t_L g360 ( .A(n_210), .B(n_324), .C(n_361), .Y(n_360) );
AO21x2_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_212), .B(n_218), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_211), .B(n_513), .Y(n_512) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_211), .B(n_538), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g561 ( .A(n_211), .B(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g395 ( .A(n_220), .B(n_267), .Y(n_395) );
INVx1_ASAP7_75t_SL g220 ( .A(n_221), .Y(n_220) );
AND2x2_ASAP7_75t_L g254 ( .A(n_221), .B(n_255), .Y(n_254) );
HB1xp67_ASAP7_75t_L g305 ( .A(n_221), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_221), .B(n_266), .Y(n_328) );
NAND3xp33_ASAP7_75t_L g435 ( .A(n_221), .B(n_307), .C(n_383), .Y(n_435) );
OA21x2_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_223), .B(n_230), .Y(n_221) );
OA21x2_ASAP7_75t_L g240 ( .A1(n_222), .A2(n_241), .B(n_250), .Y(n_240) );
OA21x2_ASAP7_75t_L g255 ( .A1(n_222), .A2(n_256), .B(n_264), .Y(n_255) );
OA21x2_ASAP7_75t_L g473 ( .A1(n_231), .A2(n_474), .B(n_480), .Y(n_473) );
OAI22xp5_ASAP7_75t_L g232 ( .A1(n_233), .A2(n_251), .B1(n_265), .B2(n_270), .Y(n_232) );
INVx1_ASAP7_75t_SL g233 ( .A(n_234), .Y(n_233) );
AND2x2_ASAP7_75t_L g234 ( .A(n_235), .B(n_238), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_235), .B(n_332), .Y(n_331) );
INVx1_ASAP7_75t_SL g347 ( .A(n_235), .Y(n_347) );
OAI31xp33_ASAP7_75t_L g363 ( .A1(n_238), .A2(n_364), .A3(n_365), .B(n_366), .Y(n_363) );
AND2x2_ASAP7_75t_L g388 ( .A(n_238), .B(n_275), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_238), .B(n_301), .Y(n_434) );
AND2x2_ASAP7_75t_L g343 ( .A(n_239), .B(n_275), .Y(n_343) );
AND2x2_ASAP7_75t_L g404 ( .A(n_239), .B(n_405), .Y(n_404) );
INVx2_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_L g274 ( .A(n_240), .B(n_275), .Y(n_274) );
INVx1_ASAP7_75t_L g332 ( .A(n_240), .Y(n_332) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_245), .B(n_247), .Y(n_246) );
INVx3_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
HB1xp67_ASAP7_75t_L g535 ( .A(n_249), .Y(n_535) );
OR2x2_ASAP7_75t_L g251 ( .A(n_252), .B(n_253), .Y(n_251) );
CKINVDCx16_ASAP7_75t_R g353 ( .A(n_252), .Y(n_353) );
NOR2xp33_ASAP7_75t_L g406 ( .A(n_253), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_SL g253 ( .A(n_254), .Y(n_253) );
AOI221x1_ASAP7_75t_SL g320 ( .A1(n_254), .A2(n_321), .B1(n_323), .B2(n_325), .C(n_327), .Y(n_320) );
INVx2_ASAP7_75t_L g268 ( .A(n_255), .Y(n_268) );
HB1xp67_ASAP7_75t_L g362 ( .A(n_255), .Y(n_362) );
INVx2_ASAP7_75t_L g511 ( .A(n_262), .Y(n_511) );
INVx3_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
INVx1_ASAP7_75t_L g350 ( .A(n_265), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_266), .B(n_269), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_266), .B(n_283), .Y(n_375) );
INVx1_ASAP7_75t_SL g438 ( .A(n_266), .Y(n_438) );
INVx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g356 ( .A(n_269), .B(n_282), .Y(n_356) );
INVx1_ASAP7_75t_L g424 ( .A(n_270), .Y(n_424) );
NOR2xp33_ASAP7_75t_L g437 ( .A(n_270), .B(n_353), .Y(n_437) );
INVx2_ASAP7_75t_SL g276 ( .A(n_271), .Y(n_276) );
AND2x2_ASAP7_75t_L g319 ( .A(n_271), .B(n_275), .Y(n_319) );
NOR2xp33_ASAP7_75t_L g325 ( .A(n_271), .B(n_326), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_271), .B(n_346), .Y(n_373) );
AOI21xp33_ASAP7_75t_SL g272 ( .A1(n_273), .A2(n_276), .B(n_277), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_274), .B(n_346), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_274), .B(n_301), .Y(n_442) );
OR2x2_ASAP7_75t_L g314 ( .A(n_275), .B(n_293), .Y(n_314) );
AND2x2_ASAP7_75t_L g413 ( .A(n_275), .B(n_404), .Y(n_413) );
OAI22xp5_ASAP7_75t_SL g288 ( .A1(n_276), .A2(n_289), .B1(n_294), .B2(n_297), .Y(n_288) );
NOR2xp33_ASAP7_75t_L g321 ( .A(n_276), .B(n_322), .Y(n_321) );
OR2x2_ASAP7_75t_L g336 ( .A(n_278), .B(n_284), .Y(n_336) );
INVx1_ASAP7_75t_L g400 ( .A(n_278), .Y(n_400) );
AOI311xp33_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_285), .A3(n_287), .B(n_288), .C(n_299), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
AOI221xp5_ASAP7_75t_L g426 ( .A1(n_283), .A2(n_415), .B1(n_427), .B2(n_430), .C(n_432), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_283), .B(n_438), .Y(n_440) );
INVx2_ASAP7_75t_SL g283 ( .A(n_284), .Y(n_283) );
INVx1_ASAP7_75t_L g337 ( .A(n_285), .Y(n_337) );
AOI211xp5_ASAP7_75t_L g327 ( .A1(n_286), .A2(n_328), .B(n_329), .C(n_331), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_290), .B(n_292), .Y(n_289) );
O2A1O1Ixp33_ASAP7_75t_SL g396 ( .A1(n_290), .A2(n_292), .B(n_397), .C(n_398), .Y(n_396) );
INVx3_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_291), .B(n_365), .Y(n_431) );
INVx1_ASAP7_75t_SL g292 ( .A(n_293), .Y(n_292) );
OAI221xp5_ASAP7_75t_L g313 ( .A1(n_294), .A2(n_314), .B1(n_315), .B2(n_318), .C(n_320), .Y(n_313) );
INVx1_ASAP7_75t_SL g295 ( .A(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g316 ( .A(n_296), .B(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g399 ( .A(n_296), .B(n_400), .Y(n_399) );
INVx1_ASAP7_75t_SL g297 ( .A(n_298), .Y(n_297) );
NOR2xp33_ASAP7_75t_L g299 ( .A(n_300), .B(n_303), .Y(n_299) );
A2O1A1Ixp33_ASAP7_75t_L g357 ( .A1(n_300), .A2(n_358), .B(n_359), .C(n_363), .Y(n_357) );
NAND2xp5_ASAP7_75t_SL g300 ( .A(n_301), .B(n_302), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_301), .B(n_391), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_301), .B(n_404), .Y(n_403) );
OR2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_306), .Y(n_303) );
INVxp67_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g323 ( .A(n_307), .B(n_324), .Y(n_323) );
INVx1_ASAP7_75t_SL g309 ( .A(n_310), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_311), .B(n_312), .Y(n_310) );
NOR2xp33_ASAP7_75t_L g382 ( .A(n_311), .B(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g425 ( .A(n_314), .Y(n_425) );
INVx1_ASAP7_75t_SL g315 ( .A(n_316), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_317), .B(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g352 ( .A(n_317), .B(n_353), .Y(n_352) );
INVx1_ASAP7_75t_SL g429 ( .A(n_317), .Y(n_429) );
INVx1_ASAP7_75t_SL g318 ( .A(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g370 ( .A(n_319), .B(n_346), .Y(n_370) );
INVx1_ASAP7_75t_SL g364 ( .A(n_326), .Y(n_364) );
INVx1_ASAP7_75t_L g341 ( .A(n_332), .Y(n_341) );
NAND3xp33_ASAP7_75t_SL g333 ( .A(n_334), .B(n_351), .C(n_367), .Y(n_333) );
AOI322xp5_ASAP7_75t_L g334 ( .A1(n_335), .A2(n_337), .A3(n_338), .B1(n_340), .B2(n_344), .C1(n_348), .C2(n_350), .Y(n_334) );
AOI211xp5_ASAP7_75t_L g387 ( .A1(n_335), .A2(n_388), .B(n_389), .C(n_396), .Y(n_387) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
OAI22xp5_ASAP7_75t_L g389 ( .A1(n_338), .A2(n_359), .B1(n_390), .B2(n_392), .Y(n_389) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g348 ( .A(n_346), .B(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g385 ( .A(n_346), .B(n_386), .Y(n_385) );
AOI32xp33_ASAP7_75t_L g436 ( .A1(n_346), .A2(n_437), .A3(n_438), .B1(n_439), .B2(n_441), .Y(n_436) );
INVx2_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g358 ( .A(n_349), .Y(n_358) );
AOI221xp5_ASAP7_75t_L g401 ( .A1(n_349), .A2(n_402), .B1(n_406), .B2(n_408), .C(n_411), .Y(n_401) );
AND2x2_ASAP7_75t_L g415 ( .A(n_349), .B(n_416), .Y(n_415) );
AND2x2_ASAP7_75t_L g418 ( .A(n_353), .B(n_419), .Y(n_418) );
OR2x2_ASAP7_75t_L g428 ( .A(n_353), .B(n_429), .Y(n_428) );
INVxp67_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx2_ASAP7_75t_SL g359 ( .A(n_360), .Y(n_359) );
INVxp67_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g419 ( .A(n_362), .B(n_383), .Y(n_419) );
AOI211xp5_ASAP7_75t_L g367 ( .A1(n_368), .A2(n_370), .B(n_371), .C(n_374), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
AOI21xp33_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_376), .B(n_378), .Y(n_374) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
OAI211xp5_ASAP7_75t_SL g380 ( .A1(n_381), .A2(n_384), .B(n_387), .C(n_401), .Y(n_380) );
INVxp67_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_394), .B(n_395), .Y(n_393) );
NAND2xp5_ASAP7_75t_SL g409 ( .A(n_395), .B(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g410 ( .A(n_407), .Y(n_410) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
AOI21xp33_ASAP7_75t_L g411 ( .A1(n_412), .A2(n_414), .B(n_417), .Y(n_411) );
INVx1_ASAP7_75t_SL g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
OAI211xp5_ASAP7_75t_SL g420 ( .A1(n_421), .A2(n_423), .B(n_426), .C(n_436), .Y(n_420) );
CKINVDCx20_ASAP7_75t_R g421 ( .A(n_422), .Y(n_421) );
NOR2xp33_ASAP7_75t_L g423 ( .A(n_424), .B(n_425), .Y(n_423) );
INVx1_ASAP7_75t_SL g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
AOI21xp33_ASAP7_75t_L g432 ( .A1(n_433), .A2(n_434), .B(n_435), .Y(n_432) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
HB1xp67_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
BUFx2_ASAP7_75t_L g455 ( .A(n_448), .Y(n_455) );
NOR2x2_ASAP7_75t_L g749 ( .A(n_449), .B(n_465), .Y(n_749) );
INVx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
OR2x2_ASAP7_75t_L g464 ( .A(n_450), .B(n_465), .Y(n_464) );
AOI21xp33_ASAP7_75t_L g456 ( .A1(n_452), .A2(n_457), .B(n_750), .Y(n_456) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
BUFx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
OAI22x1_ASAP7_75t_L g743 ( .A1(n_459), .A2(n_462), .B1(n_744), .B2(n_745), .Y(n_743) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVxp67_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
BUFx2_ASAP7_75t_L g745 ( .A(n_467), .Y(n_745) );
BUFx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
AND3x1_ASAP7_75t_L g468 ( .A(n_469), .B(n_662), .C(n_707), .Y(n_468) );
NOR4xp25_ASAP7_75t_L g469 ( .A(n_470), .B(n_585), .C(n_626), .D(n_643), .Y(n_469) );
A2O1A1Ixp33_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_501), .B(n_515), .C(n_548), .Y(n_470) );
OR2x2_ASAP7_75t_L g471 ( .A(n_472), .B(n_481), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_472), .B(n_502), .Y(n_501) );
NOR4xp25_ASAP7_75t_L g609 ( .A(n_472), .B(n_603), .C(n_610), .D(n_616), .Y(n_609) );
AND2x2_ASAP7_75t_L g682 ( .A(n_472), .B(n_571), .Y(n_682) );
AND2x2_ASAP7_75t_L g701 ( .A(n_472), .B(n_647), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_472), .B(n_696), .Y(n_710) );
AND2x2_ASAP7_75t_L g723 ( .A(n_472), .B(n_514), .Y(n_723) );
INVx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx1_ASAP7_75t_SL g568 ( .A(n_473), .Y(n_568) );
AND2x2_ASAP7_75t_L g575 ( .A(n_473), .B(n_576), .Y(n_575) );
OR2x2_ASAP7_75t_L g625 ( .A(n_473), .B(n_482), .Y(n_625) );
AND2x2_ASAP7_75t_SL g636 ( .A(n_473), .B(n_571), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_473), .B(n_482), .Y(n_640) );
AND2x2_ASAP7_75t_L g649 ( .A(n_473), .B(n_574), .Y(n_649) );
BUFx2_ASAP7_75t_L g672 ( .A(n_473), .Y(n_672) );
AND2x2_ASAP7_75t_L g676 ( .A(n_473), .B(n_492), .Y(n_676) );
OR2x2_ASAP7_75t_L g481 ( .A(n_482), .B(n_492), .Y(n_481) );
AND2x2_ASAP7_75t_L g514 ( .A(n_482), .B(n_492), .Y(n_514) );
BUFx2_ASAP7_75t_L g578 ( .A(n_482), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_482), .A2(n_611), .B1(n_613), .B2(n_614), .Y(n_610) );
OR2x2_ASAP7_75t_L g632 ( .A(n_482), .B(n_504), .Y(n_632) );
AND2x2_ASAP7_75t_L g696 ( .A(n_482), .B(n_574), .Y(n_696) );
INVx3_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
AND2x2_ASAP7_75t_L g564 ( .A(n_483), .B(n_504), .Y(n_564) );
AND2x2_ASAP7_75t_L g571 ( .A(n_483), .B(n_492), .Y(n_571) );
HB1xp67_ASAP7_75t_L g613 ( .A(n_483), .Y(n_613) );
OR2x2_ASAP7_75t_L g648 ( .A(n_483), .B(n_503), .Y(n_648) );
INVx1_ASAP7_75t_L g567 ( .A(n_492), .Y(n_567) );
INVx3_ASAP7_75t_L g576 ( .A(n_492), .Y(n_576) );
BUFx2_ASAP7_75t_L g600 ( .A(n_492), .Y(n_600) );
AND2x2_ASAP7_75t_L g633 ( .A(n_492), .B(n_568), .Y(n_633) );
OAI22xp5_ASAP7_75t_L g718 ( .A1(n_501), .A2(n_719), .B1(n_720), .B2(n_721), .Y(n_718) );
AND2x2_ASAP7_75t_L g502 ( .A(n_503), .B(n_514), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_503), .B(n_576), .Y(n_580) );
INVx1_ASAP7_75t_L g608 ( .A(n_503), .Y(n_608) );
INVx3_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx3_ASAP7_75t_L g574 ( .A(n_504), .Y(n_574) );
INVx1_ASAP7_75t_L g586 ( .A(n_514), .Y(n_586) );
NAND2x1_ASAP7_75t_SL g515 ( .A(n_516), .B(n_526), .Y(n_515) );
AND2x2_ASAP7_75t_L g584 ( .A(n_516), .B(n_539), .Y(n_584) );
HB1xp67_ASAP7_75t_L g658 ( .A(n_516), .Y(n_658) );
AND2x2_ASAP7_75t_L g685 ( .A(n_516), .B(n_605), .Y(n_685) );
AND2x2_ASAP7_75t_L g693 ( .A(n_516), .B(n_655), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_516), .B(n_551), .Y(n_720) );
INVx3_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
AND2x2_ASAP7_75t_L g552 ( .A(n_517), .B(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g569 ( .A(n_517), .B(n_570), .Y(n_569) );
INVx2_ASAP7_75t_L g590 ( .A(n_517), .Y(n_590) );
INVx1_ASAP7_75t_L g596 ( .A(n_517), .Y(n_596) );
NOR2xp33_ASAP7_75t_L g611 ( .A(n_517), .B(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g629 ( .A(n_517), .B(n_554), .Y(n_629) );
OR2x2_ASAP7_75t_L g667 ( .A(n_517), .B(n_622), .Y(n_667) );
AOI32xp33_ASAP7_75t_L g679 ( .A1(n_517), .A2(n_680), .A3(n_683), .B1(n_684), .B2(n_685), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_517), .B(n_655), .Y(n_719) );
NOR2xp33_ASAP7_75t_L g730 ( .A(n_517), .B(n_615), .Y(n_730) );
OR2x6_ASAP7_75t_L g517 ( .A(n_518), .B(n_524), .Y(n_517) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
OR2x2_ASAP7_75t_L g641 ( .A(n_527), .B(n_642), .Y(n_641) );
OR2x2_ASAP7_75t_L g527 ( .A(n_528), .B(n_539), .Y(n_527) );
INVx1_ASAP7_75t_L g603 ( .A(n_528), .Y(n_603) );
AND2x2_ASAP7_75t_L g605 ( .A(n_528), .B(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_528), .B(n_553), .Y(n_622) );
AND2x2_ASAP7_75t_L g655 ( .A(n_528), .B(n_631), .Y(n_655) );
AND2x2_ASAP7_75t_L g692 ( .A(n_528), .B(n_554), .Y(n_692) );
INVx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g551 ( .A(n_529), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_529), .B(n_553), .Y(n_582) );
AND2x2_ASAP7_75t_L g589 ( .A(n_529), .B(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g630 ( .A(n_529), .B(n_631), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_531), .B(n_536), .Y(n_530) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_533), .A2(n_534), .B(n_535), .Y(n_532) );
INVx2_ASAP7_75t_L g606 ( .A(n_539), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_539), .B(n_553), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_539), .B(n_597), .Y(n_678) );
INVx1_ASAP7_75t_L g700 ( .A(n_539), .Y(n_700) );
INVx1_ASAP7_75t_L g717 ( .A(n_539), .Y(n_717) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g570 ( .A(n_540), .B(n_553), .Y(n_570) );
AND2x2_ASAP7_75t_L g592 ( .A(n_540), .B(n_554), .Y(n_592) );
INVx1_ASAP7_75t_L g631 ( .A(n_540), .Y(n_631) );
AOI221x1_ASAP7_75t_SL g548 ( .A1(n_549), .A2(n_563), .B1(n_569), .B2(n_571), .C(n_572), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g702 ( .A1(n_549), .A2(n_636), .B1(n_703), .B2(n_704), .Y(n_702) );
AND2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_552), .Y(n_549) );
AND2x2_ASAP7_75t_L g594 ( .A(n_550), .B(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g689 ( .A(n_550), .B(n_569), .Y(n_689) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g645 ( .A(n_551), .B(n_570), .Y(n_645) );
INVx1_ASAP7_75t_L g657 ( .A(n_552), .Y(n_657) );
AND2x2_ASAP7_75t_L g668 ( .A(n_552), .B(n_655), .Y(n_668) );
AND2x2_ASAP7_75t_L g735 ( .A(n_552), .B(n_630), .Y(n_735) );
INVx2_ASAP7_75t_L g597 ( .A(n_553), .Y(n_597) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_564), .B(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g687 ( .A(n_564), .Y(n_687) );
NOR2xp33_ASAP7_75t_L g651 ( .A(n_565), .B(n_648), .Y(n_651) );
INVx3_ASAP7_75t_SL g565 ( .A(n_566), .Y(n_565) );
AOI21xp5_ASAP7_75t_L g731 ( .A1(n_566), .A2(n_687), .B(n_732), .Y(n_731) );
AND2x4_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
NOR2xp33_ASAP7_75t_SL g709 ( .A(n_569), .B(n_595), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_570), .B(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g661 ( .A(n_570), .B(n_589), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_570), .B(n_596), .Y(n_738) );
AND2x2_ASAP7_75t_L g607 ( .A(n_571), .B(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g674 ( .A(n_571), .Y(n_674) );
AOI21xp33_ASAP7_75t_L g572 ( .A1(n_573), .A2(n_577), .B(n_581), .Y(n_572) );
NAND2x1_ASAP7_75t_L g573 ( .A(n_574), .B(n_575), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_574), .B(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g623 ( .A(n_574), .B(n_624), .Y(n_623) );
INVx1_ASAP7_75t_SL g635 ( .A(n_574), .Y(n_635) );
NOR2xp33_ASAP7_75t_L g680 ( .A(n_574), .B(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g659 ( .A(n_575), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_575), .B(n_696), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_575), .B(n_578), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_578), .B(n_579), .Y(n_577) );
AOI211xp5_ASAP7_75t_L g646 ( .A1(n_578), .A2(n_617), .B(n_647), .C(n_649), .Y(n_646) );
AOI221xp5_ASAP7_75t_L g664 ( .A1(n_578), .A2(n_665), .B1(n_668), .B2(n_669), .C(n_673), .Y(n_664) );
AND2x2_ASAP7_75t_L g660 ( .A(n_579), .B(n_613), .Y(n_660) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
OR2x2_ASAP7_75t_L g581 ( .A(n_582), .B(n_583), .Y(n_581) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g620 ( .A(n_584), .B(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g691 ( .A(n_584), .B(n_692), .Y(n_691) );
OAI211xp5_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_587), .B(n_593), .C(n_618), .Y(n_585) );
NAND3xp33_ASAP7_75t_SL g704 ( .A(n_586), .B(n_705), .C(n_706), .Y(n_704) );
OR2x2_ASAP7_75t_L g587 ( .A(n_588), .B(n_591), .Y(n_587) );
OR2x2_ASAP7_75t_L g677 ( .A(n_588), .B(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AOI221xp5_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_598), .B1(n_601), .B2(n_607), .C(n_609), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_595), .B(n_605), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_595), .B(n_638), .Y(n_637) );
AND2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g617 ( .A(n_600), .Y(n_617) );
OAI22xp5_ASAP7_75t_L g656 ( .A1(n_600), .A2(n_657), .B1(n_658), .B2(n_659), .Y(n_656) );
OR2x2_ASAP7_75t_L g737 ( .A(n_600), .B(n_648), .Y(n_737) );
NAND2xp5_ASAP7_75t_SL g601 ( .A(n_602), .B(n_604), .Y(n_601) );
INVxp67_ASAP7_75t_L g711 ( .A(n_603), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_605), .B(n_726), .Y(n_725) );
INVxp67_ASAP7_75t_L g612 ( .A(n_606), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_608), .B(n_617), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_608), .B(n_655), .Y(n_654) );
NOR2xp33_ASAP7_75t_L g714 ( .A(n_608), .B(n_675), .Y(n_714) );
HB1xp67_ASAP7_75t_L g638 ( .A(n_612), .Y(n_638) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
OR2x2_ASAP7_75t_L g728 ( .A(n_617), .B(n_648), .Y(n_728) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g619 ( .A(n_620), .B(n_623), .Y(n_619) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx1_ASAP7_75t_SL g706 ( .A(n_623), .Y(n_706) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
OAI322xp33_ASAP7_75t_SL g626 ( .A1(n_627), .A2(n_632), .A3(n_633), .B1(n_634), .B2(n_637), .C1(n_639), .C2(n_641), .Y(n_626) );
OAI322xp33_ASAP7_75t_L g708 ( .A1(n_627), .A2(n_709), .A3(n_710), .B1(n_711), .B2(n_712), .C1(n_713), .C2(n_715), .Y(n_708) );
CKINVDCx16_ASAP7_75t_R g627 ( .A(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g628 ( .A(n_629), .B(n_630), .Y(n_628) );
INVx4_ASAP7_75t_L g642 ( .A(n_629), .Y(n_642) );
AND2x2_ASAP7_75t_L g703 ( .A(n_629), .B(n_655), .Y(n_703) );
AND2x2_ASAP7_75t_L g716 ( .A(n_629), .B(n_717), .Y(n_716) );
CKINVDCx16_ASAP7_75t_R g727 ( .A(n_632), .Y(n_727) );
INVx1_ASAP7_75t_L g705 ( .A(n_633), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_635), .B(n_636), .Y(n_634) );
OR2x2_ASAP7_75t_L g639 ( .A(n_635), .B(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_L g722 ( .A(n_635), .B(n_723), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_635), .B(n_676), .Y(n_733) );
OR2x2_ASAP7_75t_L g666 ( .A(n_638), .B(n_667), .Y(n_666) );
INVxp33_ASAP7_75t_L g683 ( .A(n_638), .Y(n_683) );
OAI221xp5_ASAP7_75t_SL g643 ( .A1(n_642), .A2(n_644), .B1(n_646), .B2(n_650), .C(n_652), .Y(n_643) );
NOR2xp67_ASAP7_75t_L g699 ( .A(n_642), .B(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g726 ( .A(n_642), .Y(n_726) );
INVx1_ASAP7_75t_SL g644 ( .A(n_645), .Y(n_644) );
INVx3_ASAP7_75t_SL g647 ( .A(n_648), .Y(n_647) );
AOI322xp5_ASAP7_75t_L g690 ( .A1(n_649), .A2(n_674), .A3(n_691), .B1(n_693), .B2(n_694), .C1(n_697), .C2(n_701), .Y(n_690) );
INVxp67_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
AOI22xp5_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_656), .B1(n_660), .B2(n_661), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
NOR2xp33_ASAP7_75t_L g662 ( .A(n_663), .B(n_686), .Y(n_662) );
NAND2xp5_ASAP7_75t_SL g663 ( .A(n_664), .B(n_679), .Y(n_663) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
NAND2xp5_ASAP7_75t_SL g697 ( .A(n_667), .B(n_698), .Y(n_697) );
INVx1_ASAP7_75t_SL g669 ( .A(n_670), .Y(n_669) );
NAND2xp33_ASAP7_75t_SL g684 ( .A(n_670), .B(n_681), .Y(n_684) );
INVx1_ASAP7_75t_SL g671 ( .A(n_672), .Y(n_671) );
OAI322xp33_ASAP7_75t_L g724 ( .A1(n_672), .A2(n_725), .A3(n_727), .B1(n_728), .B2(n_729), .C1(n_731), .C2(n_734), .Y(n_724) );
AOI21xp33_ASAP7_75t_SL g673 ( .A1(n_674), .A2(n_675), .B(n_677), .Y(n_673) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx2_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_682), .B(n_730), .Y(n_739) );
OAI211xp5_ASAP7_75t_SL g686 ( .A1(n_687), .A2(n_688), .B(n_690), .C(n_702), .Y(n_686) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
NOR4xp25_ASAP7_75t_L g707 ( .A(n_708), .B(n_718), .C(n_724), .D(n_736), .Y(n_707) );
INVxp67_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_SL g721 ( .A(n_722), .Y(n_721) );
INVxp67_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
CKINVDCx14_ASAP7_75t_R g734 ( .A(n_735), .Y(n_734) );
OAI21xp5_ASAP7_75t_SL g736 ( .A1(n_737), .A2(n_738), .B(n_739), .Y(n_736) );
INVx1_ASAP7_75t_L g746 ( .A(n_740), .Y(n_746) );
INVx1_ASAP7_75t_SL g747 ( .A(n_748), .Y(n_747) );
INVx2_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
endmodule