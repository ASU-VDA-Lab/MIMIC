module fake_jpeg_1242_n_577 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_577);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_577;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g19 ( 
.A(n_18),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_1),
.B(n_6),
.Y(n_37)
);

BUFx24_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_10),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_11),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_15),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_53),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_54),
.Y(n_115)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_55),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_56),
.Y(n_143)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_57),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_58),
.Y(n_144)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

INVx4_ASAP7_75t_SL g129 ( 
.A(n_59),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_35),
.B(n_16),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_60),
.B(n_74),
.Y(n_135)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_61),
.Y(n_114)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_62),
.Y(n_127)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_63),
.Y(n_156)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx11_ASAP7_75t_L g117 ( 
.A(n_64),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_65),
.Y(n_166)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_66),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_37),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_67),
.B(n_76),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_68),
.Y(n_169)
);

BUFx10_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx3_ASAP7_75t_SL g164 ( 
.A(n_69),
.Y(n_164)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_70),
.Y(n_120)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_71),
.Y(n_131)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_72),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_73),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_35),
.B(n_16),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_75),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_29),
.Y(n_76)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g133 ( 
.A(n_77),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_22),
.B(n_18),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_78),
.B(n_93),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_29),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_79),
.B(n_81),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_80),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_46),
.B(n_18),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g136 ( 
.A(n_82),
.Y(n_136)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_83),
.Y(n_141)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_38),
.Y(n_84)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_29),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_85),
.B(n_94),
.Y(n_121)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_36),
.Y(n_86)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_86),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_87),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_51),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g140 ( 
.A(n_88),
.Y(n_140)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_38),
.Y(n_89)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_89),
.Y(n_123)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_22),
.Y(n_90)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_90),
.Y(n_132)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_31),
.Y(n_91)
);

INVx6_ASAP7_75t_SL g150 ( 
.A(n_91),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g145 ( 
.A(n_92),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_50),
.B(n_14),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_19),
.B(n_15),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_32),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_95),
.B(n_41),
.Y(n_147)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_30),
.Y(n_96)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_96),
.Y(n_159)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_97),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_49),
.B(n_13),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_98),
.B(n_99),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_50),
.B(n_21),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_30),
.Y(n_100)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_100),
.Y(n_172)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_36),
.Y(n_101)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_20),
.Y(n_102)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_102),
.Y(n_152)
);

BUFx5_ASAP7_75t_L g103 ( 
.A(n_31),
.Y(n_103)
);

BUFx2_ASAP7_75t_R g162 ( 
.A(n_103),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_20),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_104),
.Y(n_111)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_20),
.Y(n_105)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_105),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_32),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g116 ( 
.A(n_106),
.Y(n_116)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_43),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_107),
.Y(n_160)
);

NAND2xp33_ASAP7_75t_SL g122 ( 
.A(n_100),
.B(n_43),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g211 ( 
.A(n_122),
.B(n_124),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_81),
.B(n_19),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_94),
.B(n_49),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_138),
.B(n_153),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_71),
.B(n_21),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_139),
.B(n_45),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_107),
.A2(n_41),
.B1(n_32),
.B2(n_45),
.Y(n_146)
);

OA22x2_ASAP7_75t_L g205 ( 
.A1(n_146),
.A2(n_69),
.B1(n_54),
.B2(n_87),
.Y(n_205)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_147),
.Y(n_178)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_72),
.Y(n_149)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_149),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_86),
.B(n_40),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_59),
.B(n_34),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_154),
.B(n_155),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_62),
.B(n_34),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_104),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_158),
.B(n_55),
.Y(n_174)
);

NAND2xp33_ASAP7_75t_SL g161 ( 
.A(n_101),
.B(n_56),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_161),
.B(n_103),
.Y(n_212)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_105),
.Y(n_163)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_163),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_106),
.A2(n_41),
.B1(n_25),
.B2(n_40),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_165),
.A2(n_64),
.B1(n_91),
.B2(n_92),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_65),
.B(n_39),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_168),
.B(n_170),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_80),
.B(n_39),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_80),
.B(n_25),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_171),
.B(n_2),
.Y(n_222)
);

BUFx12_ASAP7_75t_L g173 ( 
.A(n_150),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_173),
.Y(n_236)
);

CKINVDCx14_ASAP7_75t_R g274 ( 
.A(n_174),
.Y(n_274)
);

NAND2xp33_ASAP7_75t_SL g175 ( 
.A(n_162),
.B(n_77),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_175),
.Y(n_283)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_112),
.Y(n_176)
);

INVx3_ASAP7_75t_SL g258 ( 
.A(n_176),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_118),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_177),
.B(n_179),
.Y(n_268)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_112),
.Y(n_180)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_180),
.Y(n_244)
);

BUFx12f_ASAP7_75t_L g182 ( 
.A(n_142),
.Y(n_182)
);

INVx5_ASAP7_75t_L g254 ( 
.A(n_182),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_115),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_183),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_135),
.B(n_33),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_184),
.B(n_191),
.Y(n_237)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_134),
.Y(n_185)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_185),
.Y(n_240)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_126),
.Y(n_186)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_186),
.Y(n_249)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_142),
.Y(n_188)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_188),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_121),
.A2(n_63),
.B1(n_70),
.B2(n_73),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_189),
.A2(n_197),
.B1(n_157),
.B2(n_169),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_132),
.B(n_33),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_192),
.A2(n_207),
.B1(n_110),
.B2(n_164),
.Y(n_256)
);

BUFx2_ASAP7_75t_L g193 ( 
.A(n_126),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_193),
.Y(n_284)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_130),
.Y(n_194)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_194),
.Y(n_263)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_130),
.Y(n_195)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_195),
.Y(n_265)
);

NAND2x1_ASAP7_75t_L g196 ( 
.A(n_124),
.B(n_97),
.Y(n_196)
);

OR2x2_ASAP7_75t_L g286 ( 
.A(n_196),
.B(n_221),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_119),
.A2(n_75),
.B1(n_68),
.B2(n_88),
.Y(n_197)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_152),
.Y(n_198)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_198),
.Y(n_285)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_113),
.Y(n_200)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_200),
.Y(n_245)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_152),
.Y(n_201)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_201),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_115),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_202),
.Y(n_266)
);

INVx8_ASAP7_75t_L g203 ( 
.A(n_140),
.Y(n_203)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_203),
.Y(n_246)
);

INVx8_ASAP7_75t_L g204 ( 
.A(n_140),
.Y(n_204)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_204),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_205),
.A2(n_208),
.B1(n_166),
.B2(n_117),
.Y(n_262)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_143),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_206),
.Y(n_272)
);

OAI22xp33_ASAP7_75t_L g207 ( 
.A1(n_146),
.A2(n_82),
.B1(n_58),
.B2(n_102),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_161),
.A2(n_69),
.B1(n_89),
.B2(n_84),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_148),
.B(n_13),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_209),
.B(n_213),
.Y(n_239)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_114),
.Y(n_210)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_210),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_212),
.B(n_232),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_111),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_144),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_214),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_151),
.B(n_1),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_216),
.B(n_222),
.Y(n_241)
);

INVx8_ASAP7_75t_L g217 ( 
.A(n_140),
.Y(n_217)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_217),
.Y(n_260)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_127),
.Y(n_218)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_218),
.Y(n_264)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_127),
.Y(n_219)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_219),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_144),
.Y(n_220)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_220),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_122),
.B(n_1),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_109),
.B(n_2),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_223),
.B(n_227),
.Y(n_251)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_172),
.Y(n_224)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_224),
.Y(n_273)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_143),
.Y(n_225)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_225),
.Y(n_278)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_167),
.Y(n_226)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_226),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_125),
.B(n_2),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_160),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_228),
.B(n_229),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_116),
.Y(n_229)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_166),
.Y(n_230)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_230),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_141),
.B(n_3),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_231),
.B(n_234),
.Y(n_289)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_131),
.Y(n_232)
);

INVx6_ASAP7_75t_L g233 ( 
.A(n_169),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_233),
.Y(n_261)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_159),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_129),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_235),
.Y(n_276)
);

AOI32xp33_ASAP7_75t_L g238 ( 
.A1(n_190),
.A2(n_110),
.A3(n_123),
.B1(n_137),
.B2(n_162),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_238),
.B(n_287),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_L g242 ( 
.A1(n_207),
.A2(n_136),
.B1(n_129),
.B2(n_120),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_242),
.A2(n_247),
.B1(n_279),
.B2(n_208),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_L g247 ( 
.A1(n_211),
.A2(n_136),
.B1(n_120),
.B2(n_157),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_181),
.B(n_133),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_248),
.B(n_250),
.C(n_286),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_196),
.B(n_211),
.C(n_178),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_252),
.B(n_205),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_221),
.A2(n_164),
.B(n_123),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_253),
.A2(n_192),
.B(n_204),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_256),
.A2(n_283),
.B1(n_243),
.B2(n_261),
.Y(n_309)
);

OAI21xp33_ASAP7_75t_SL g302 ( 
.A1(n_262),
.A2(n_269),
.B(n_205),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_212),
.A2(n_175),
.B1(n_201),
.B2(n_198),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_L g279 ( 
.A1(n_187),
.A2(n_133),
.B1(n_156),
.B2(n_117),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_215),
.B(n_156),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_280),
.B(n_288),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_193),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_199),
.B(n_128),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_280),
.B(n_206),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_292),
.B(n_297),
.Y(n_341)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_288),
.Y(n_293)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_293),
.Y(n_343)
);

BUFx2_ASAP7_75t_L g380 ( 
.A(n_295),
.Y(n_380)
);

CKINVDCx14_ASAP7_75t_R g345 ( 
.A(n_296),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_274),
.B(n_186),
.Y(n_297)
);

BUFx2_ASAP7_75t_L g298 ( 
.A(n_258),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_298),
.Y(n_361)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_258),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_299),
.Y(n_368)
);

INVx11_ASAP7_75t_L g300 ( 
.A(n_258),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_300),
.Y(n_357)
);

CKINVDCx14_ASAP7_75t_R g301 ( 
.A(n_243),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_301),
.B(n_304),
.Y(n_344)
);

OR2x2_ASAP7_75t_L g365 ( 
.A(n_302),
.B(n_316),
.Y(n_365)
);

INVx13_ASAP7_75t_L g303 ( 
.A(n_236),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g359 ( 
.A(n_303),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_239),
.B(n_182),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_245),
.Y(n_305)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_305),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_248),
.B(n_182),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_306),
.B(n_310),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_307),
.B(n_337),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_250),
.B(n_230),
.C(n_225),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_308),
.B(n_335),
.C(n_246),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_309),
.A2(n_320),
.B1(n_329),
.B2(n_340),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_237),
.B(n_268),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_289),
.B(n_195),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_311),
.B(n_314),
.Y(n_352)
);

INVx2_ASAP7_75t_SL g312 ( 
.A(n_271),
.Y(n_312)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_312),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_276),
.B(n_176),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_313),
.B(n_318),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_251),
.B(n_194),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_286),
.B(n_180),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_315),
.B(n_325),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_275),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_317),
.B(n_328),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_245),
.B(n_233),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_259),
.B(n_217),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_319),
.B(n_321),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_283),
.A2(n_108),
.B1(n_214),
.B2(n_202),
.Y(n_320)
);

CKINVDCx16_ASAP7_75t_R g321 ( 
.A(n_253),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_252),
.A2(n_128),
.B1(n_108),
.B2(n_183),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_322),
.A2(n_257),
.B1(n_254),
.B2(n_27),
.Y(n_382)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_259),
.Y(n_323)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_323),
.Y(n_374)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_273),
.Y(n_324)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_324),
.Y(n_379)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_273),
.Y(n_325)
);

OA21x2_ASAP7_75t_L g326 ( 
.A1(n_243),
.A2(n_173),
.B(n_203),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_326),
.B(n_327),
.Y(n_360)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_281),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_284),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_L g329 ( 
.A1(n_285),
.A2(n_220),
.B1(n_27),
.B2(n_173),
.Y(n_329)
);

BUFx3_ASAP7_75t_L g330 ( 
.A(n_236),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_330),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_241),
.B(n_272),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_331),
.B(n_332),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_272),
.B(n_145),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_281),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_333),
.B(n_334),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_SL g334 ( 
.A(n_278),
.B(n_27),
.Y(n_334)
);

MAJx2_ASAP7_75t_L g335 ( 
.A(n_264),
.B(n_27),
.C(n_145),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_271),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_336),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_278),
.B(n_145),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_270),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_338),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_264),
.B(n_3),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_339),
.B(n_240),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_266),
.A2(n_277),
.B1(n_270),
.B2(n_244),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_321),
.A2(n_266),
.B1(n_277),
.B2(n_244),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_342),
.B(n_349),
.Y(n_394)
);

XNOR2x1_ASAP7_75t_L g397 ( 
.A(n_348),
.B(n_378),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_296),
.A2(n_290),
.B1(n_285),
.B2(n_282),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g351 ( 
.A1(n_294),
.A2(n_282),
.B(n_267),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_L g403 ( 
.A1(n_351),
.A2(n_328),
.B(n_339),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_296),
.A2(n_290),
.B1(n_265),
.B2(n_263),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_354),
.B(n_364),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_337),
.Y(n_362)
);

INVx13_ASAP7_75t_L g422 ( 
.A(n_362),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_293),
.A2(n_265),
.B1(n_263),
.B2(n_255),
.Y(n_364)
);

OA21x2_ASAP7_75t_L g366 ( 
.A1(n_316),
.A2(n_260),
.B(n_255),
.Y(n_366)
);

O2A1O1Ixp33_ASAP7_75t_L g399 ( 
.A1(n_366),
.A2(n_326),
.B(n_334),
.C(n_324),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_309),
.A2(n_267),
.B1(n_249),
.B2(n_260),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_369),
.B(n_372),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_317),
.A2(n_246),
.B1(n_249),
.B2(n_257),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_376),
.B(n_381),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_307),
.B(n_240),
.Y(n_378)
);

CKINVDCx16_ASAP7_75t_R g381 ( 
.A(n_297),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_382),
.A2(n_295),
.B1(n_320),
.B2(n_326),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_311),
.Y(n_383)
);

NOR3xp33_ASAP7_75t_L g405 ( 
.A(n_383),
.B(n_333),
.C(n_312),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_308),
.B(n_254),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_384),
.B(n_335),
.Y(n_391)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_350),
.Y(n_385)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_385),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_386),
.A2(n_393),
.B1(n_407),
.B2(n_413),
.Y(n_438)
);

OAI32xp33_ASAP7_75t_L g387 ( 
.A1(n_343),
.A2(n_291),
.A3(n_292),
.B1(n_314),
.B2(n_305),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_387),
.B(n_395),
.Y(n_425)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_350),
.Y(n_388)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_388),
.Y(n_437)
);

INVx3_ASAP7_75t_L g389 ( 
.A(n_363),
.Y(n_389)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_389),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_391),
.B(n_414),
.Y(n_441)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_374),
.Y(n_392)
);

INVx1_ASAP7_75t_SL g434 ( 
.A(n_392),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_380),
.A2(n_291),
.B1(n_315),
.B2(n_322),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_347),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_375),
.B(n_323),
.Y(n_396)
);

NAND3xp33_ASAP7_75t_L g445 ( 
.A(n_396),
.B(n_404),
.C(n_406),
.Y(n_445)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_342),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_398),
.B(n_400),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g444 ( 
.A1(n_399),
.A2(n_345),
.B(n_369),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_341),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_353),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_402),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_403),
.B(n_410),
.Y(n_431)
);

NAND3xp33_ASAP7_75t_L g404 ( 
.A(n_367),
.B(n_325),
.C(n_327),
.Y(n_404)
);

INVxp33_ASAP7_75t_L g442 ( 
.A(n_405),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_344),
.B(n_330),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_380),
.A2(n_312),
.B1(n_336),
.B2(n_338),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_351),
.B(n_352),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_SL g429 ( 
.A(n_408),
.B(n_409),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_352),
.B(n_299),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_374),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_365),
.A2(n_340),
.B(n_298),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_SL g430 ( 
.A1(n_412),
.A2(n_366),
.B(n_360),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_380),
.A2(n_338),
.B1(n_298),
.B2(n_300),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_378),
.B(n_303),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_SL g415 ( 
.A(n_383),
.B(n_303),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_SL g443 ( 
.A(n_415),
.B(n_417),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_343),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g455 ( 
.A1(n_416),
.A2(n_356),
.B1(n_358),
.B2(n_361),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_377),
.B(n_5),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_341),
.B(n_5),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_418),
.B(n_421),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_373),
.B(n_5),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_SL g453 ( 
.A(n_419),
.B(n_356),
.Y(n_453)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_363),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_420),
.Y(n_440)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_379),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_395),
.B(n_373),
.Y(n_424)
);

NAND3xp33_ASAP7_75t_L g462 ( 
.A(n_424),
.B(n_435),
.C(n_436),
.Y(n_462)
);

OA22x2_ASAP7_75t_L g426 ( 
.A1(n_398),
.A2(n_366),
.B1(n_382),
.B2(n_365),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_426),
.B(n_452),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_397),
.B(n_384),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_427),
.B(n_451),
.Y(n_467)
);

CKINVDCx16_ASAP7_75t_R g428 ( 
.A(n_403),
.Y(n_428)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_428),
.Y(n_474)
);

OAI21xp5_ASAP7_75t_SL g463 ( 
.A1(n_430),
.A2(n_444),
.B(n_446),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_402),
.B(n_362),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_SL g478 ( 
.A(n_432),
.B(n_433),
.Y(n_478)
);

AOI21xp33_ASAP7_75t_L g433 ( 
.A1(n_412),
.A2(n_360),
.B(n_355),
.Y(n_433)
);

NOR4xp25_ASAP7_75t_L g435 ( 
.A(n_400),
.B(n_355),
.C(n_348),
.D(n_371),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_415),
.B(n_359),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g446 ( 
.A1(n_399),
.A2(n_349),
.B(n_346),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_390),
.B(n_376),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_447),
.B(n_448),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_418),
.B(n_371),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_397),
.B(n_379),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_394),
.B(n_370),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_453),
.B(n_416),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_414),
.B(n_354),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_454),
.B(n_387),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_L g471 ( 
.A1(n_455),
.A2(n_438),
.B1(n_446),
.B2(n_386),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_449),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_457),
.B(n_479),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_451),
.B(n_391),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_458),
.B(n_468),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_459),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_443),
.B(n_389),
.Y(n_461)
);

NAND3xp33_ASAP7_75t_L g506 ( 
.A(n_461),
.B(n_472),
.C(n_483),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_425),
.A2(n_394),
.B1(n_411),
.B2(n_401),
.Y(n_464)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_464),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_427),
.B(n_421),
.C(n_385),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_466),
.B(n_469),
.C(n_470),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_441),
.B(n_393),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_441),
.B(n_454),
.C(n_428),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_L g508 ( 
.A1(n_471),
.A2(n_476),
.B1(n_481),
.B2(n_455),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_443),
.B(n_420),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_440),
.B(n_392),
.Y(n_473)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_473),
.Y(n_498)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_437),
.Y(n_475)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_475),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_423),
.A2(n_411),
.B1(n_407),
.B2(n_401),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_425),
.A2(n_422),
.B1(n_410),
.B2(n_388),
.Y(n_477)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_477),
.Y(n_496)
);

HB1xp67_ASAP7_75t_L g479 ( 
.A(n_453),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_423),
.B(n_370),
.C(n_422),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_480),
.B(n_485),
.C(n_466),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_L g481 ( 
.A1(n_445),
.A2(n_358),
.B1(n_413),
.B2(n_368),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_437),
.Y(n_482)
);

INVx2_ASAP7_75t_SL g495 ( 
.A(n_482),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_431),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_438),
.A2(n_368),
.B1(n_361),
.B2(n_357),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_484),
.B(n_426),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_431),
.B(n_6),
.C(n_7),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_477),
.Y(n_486)
);

NAND3xp33_ASAP7_75t_L g521 ( 
.A(n_486),
.B(n_499),
.C(n_456),
.Y(n_521)
);

OAI21xp5_ASAP7_75t_L g489 ( 
.A1(n_463),
.A2(n_449),
.B(n_444),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g527 ( 
.A(n_489),
.B(n_503),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_490),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_457),
.A2(n_452),
.B1(n_435),
.B2(n_442),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_493),
.A2(n_508),
.B1(n_484),
.B2(n_474),
.Y(n_514)
);

AOI21xp5_ASAP7_75t_L g497 ( 
.A1(n_463),
.A2(n_430),
.B(n_440),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_497),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_478),
.B(n_429),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_475),
.B(n_482),
.Y(n_500)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_500),
.Y(n_512)
);

BUFx24_ASAP7_75t_SL g502 ( 
.A(n_462),
.Y(n_502)
);

BUFx24_ASAP7_75t_SL g523 ( 
.A(n_502),
.Y(n_523)
);

XOR2xp5_ASAP7_75t_SL g503 ( 
.A(n_468),
.B(n_426),
.Y(n_503)
);

OAI21x1_ASAP7_75t_SL g504 ( 
.A1(n_460),
.A2(n_439),
.B(n_426),
.Y(n_504)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_504),
.Y(n_513)
);

BUFx24_ASAP7_75t_SL g505 ( 
.A(n_465),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_505),
.Y(n_525)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_507),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_L g509 ( 
.A1(n_476),
.A2(n_429),
.B1(n_439),
.B2(n_450),
.Y(n_509)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_509),
.Y(n_526)
);

AO22x1_ASAP7_75t_L g510 ( 
.A1(n_496),
.A2(n_464),
.B1(n_474),
.B2(n_460),
.Y(n_510)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_510),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_L g542 ( 
.A1(n_514),
.A2(n_518),
.B1(n_521),
.B2(n_495),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_488),
.B(n_470),
.C(n_469),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_516),
.B(n_517),
.C(n_507),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_488),
.B(n_480),
.C(n_467),
.Y(n_517)
);

AOI221xp5_ASAP7_75t_L g518 ( 
.A1(n_492),
.A2(n_473),
.B1(n_434),
.B2(n_450),
.C(n_485),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_506),
.B(n_500),
.Y(n_519)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_519),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_487),
.B(n_434),
.Y(n_520)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_520),
.Y(n_532)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_487),
.Y(n_522)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_522),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_SL g524 ( 
.A1(n_494),
.A2(n_456),
.B1(n_458),
.B2(n_467),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_524),
.B(n_503),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_529),
.B(n_530),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_515),
.B(n_491),
.C(n_496),
.Y(n_530)
);

CKINVDCx16_ASAP7_75t_R g533 ( 
.A(n_519),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_533),
.B(n_534),
.Y(n_556)
);

AOI21xp5_ASAP7_75t_L g535 ( 
.A1(n_511),
.A2(n_489),
.B(n_497),
.Y(n_535)
);

OAI21xp5_ASAP7_75t_L g552 ( 
.A1(n_535),
.A2(n_536),
.B(n_537),
.Y(n_552)
);

AOI21xp5_ASAP7_75t_L g536 ( 
.A1(n_526),
.A2(n_493),
.B(n_490),
.Y(n_536)
);

OAI21xp5_ASAP7_75t_SL g537 ( 
.A1(n_513),
.A2(n_494),
.B(n_498),
.Y(n_537)
);

XOR2xp5_ASAP7_75t_L g539 ( 
.A(n_527),
.B(n_491),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_539),
.B(n_543),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_517),
.B(n_495),
.C(n_501),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_541),
.B(n_544),
.C(n_524),
.Y(n_550)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_542),
.Y(n_549)
);

XOR2xp5_ASAP7_75t_L g543 ( 
.A(n_527),
.B(n_495),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_516),
.B(n_7),
.C(n_8),
.Y(n_544)
);

OAI22xp5_ASAP7_75t_SL g547 ( 
.A1(n_538),
.A2(n_536),
.B1(n_540),
.B2(n_514),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_547),
.B(n_551),
.Y(n_560)
);

OAI21x1_ASAP7_75t_L g548 ( 
.A1(n_535),
.A2(n_512),
.B(n_520),
.Y(n_548)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_548),
.Y(n_559)
);

XOR2xp5_ASAP7_75t_L g563 ( 
.A(n_550),
.B(n_553),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_541),
.B(n_528),
.C(n_510),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_L g553 ( 
.A1(n_531),
.A2(n_528),
.B1(n_510),
.B2(n_523),
.Y(n_553)
);

OAI21x1_ASAP7_75t_L g554 ( 
.A1(n_540),
.A2(n_525),
.B(n_9),
.Y(n_554)
);

OAI21xp33_ASAP7_75t_L g561 ( 
.A1(n_554),
.A2(n_8),
.B(n_9),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_SL g555 ( 
.A(n_529),
.B(n_8),
.Y(n_555)
);

OAI21xp5_ASAP7_75t_L g557 ( 
.A1(n_555),
.A2(n_532),
.B(n_544),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_557),
.B(n_558),
.Y(n_564)
);

AOI22xp5_ASAP7_75t_SL g558 ( 
.A1(n_556),
.A2(n_532),
.B1(n_531),
.B2(n_530),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_SL g567 ( 
.A(n_561),
.B(n_562),
.Y(n_567)
);

INVx6_ASAP7_75t_L g562 ( 
.A(n_545),
.Y(n_562)
);

NOR2xp67_ASAP7_75t_L g565 ( 
.A(n_559),
.B(n_552),
.Y(n_565)
);

AOI21x1_ASAP7_75t_L g570 ( 
.A1(n_565),
.A2(n_552),
.B(n_549),
.Y(n_570)
);

INVxp67_ASAP7_75t_L g566 ( 
.A(n_560),
.Y(n_566)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_566),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_564),
.B(n_562),
.Y(n_569)
);

AOI322xp5_ASAP7_75t_L g571 ( 
.A1(n_569),
.A2(n_570),
.A3(n_537),
.B1(n_546),
.B2(n_563),
.C1(n_567),
.C2(n_551),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_571),
.B(n_572),
.C(n_9),
.Y(n_573)
);

AOI322xp5_ASAP7_75t_L g572 ( 
.A1(n_568),
.A2(n_546),
.A3(n_550),
.B1(n_543),
.B2(n_539),
.C1(n_561),
.C2(n_12),
.Y(n_572)
);

BUFx24_ASAP7_75t_SL g574 ( 
.A(n_573),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_574),
.B(n_10),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_575),
.B(n_11),
.C(n_12),
.Y(n_576)
);

XOR2xp5_ASAP7_75t_L g577 ( 
.A(n_576),
.B(n_11),
.Y(n_577)
);


endmodule