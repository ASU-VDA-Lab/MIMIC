module fake_jpeg_3374_n_541 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_541);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_541;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx10_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx4f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_15),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_16),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx4f_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

INVx6_ASAP7_75t_SL g44 ( 
.A(n_7),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_10),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_3),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_14),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_16),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_32),
.B(n_17),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_52),
.B(n_53),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_54),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_55),
.Y(n_115)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_56),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_39),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_57),
.B(n_59),
.Y(n_106)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_58),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_39),
.Y(n_59)
);

AND2x2_ASAP7_75t_SL g60 ( 
.A(n_41),
.B(n_0),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_60),
.B(n_90),
.Y(n_119)
);

BUFx4f_ASAP7_75t_SL g61 ( 
.A(n_44),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_61),
.Y(n_132)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_62),
.Y(n_130)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_63),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_64),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_65),
.Y(n_139)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_66),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_32),
.B(n_17),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_67),
.B(n_77),
.Y(n_107)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_68),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_69),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_28),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_70),
.Y(n_169)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_71),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_28),
.Y(n_72)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_72),
.Y(n_110)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_21),
.Y(n_73)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_73),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_39),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_74),
.B(n_86),
.Y(n_116)
);

INVx6_ASAP7_75t_SL g75 ( 
.A(n_20),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_75),
.Y(n_118)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_21),
.Y(n_76)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_76),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_34),
.B(n_0),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_34),
.B(n_0),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_78),
.B(n_91),
.Y(n_127)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_21),
.Y(n_79)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_79),
.Y(n_134)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_41),
.Y(n_80)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_80),
.Y(n_153)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_21),
.Y(n_81)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_81),
.Y(n_149)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_31),
.Y(n_82)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_82),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_83),
.Y(n_164)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_41),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g108 ( 
.A(n_84),
.Y(n_108)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_28),
.Y(n_85)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_85),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_23),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_28),
.Y(n_87)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_87),
.Y(n_123)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_31),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_88),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_89),
.Y(n_158)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_36),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_36),
.Y(n_91)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_41),
.Y(n_92)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_92),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_37),
.B(n_1),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_93),
.B(n_101),
.Y(n_135)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_38),
.Y(n_94)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_94),
.Y(n_159)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_95),
.B(n_96),
.Y(n_131)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_24),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_97),
.B(n_99),
.Y(n_144)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_19),
.Y(n_98)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_98),
.Y(n_166)
);

INVx2_ASAP7_75t_SL g99 ( 
.A(n_42),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_23),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_104),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_51),
.B(n_1),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_42),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_102),
.B(n_103),
.Y(n_143)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_42),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_23),
.Y(n_104)
);

AOI21xp33_ASAP7_75t_SL g111 ( 
.A1(n_60),
.A2(n_42),
.B(n_50),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_111),
.B(n_89),
.C(n_83),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_96),
.A2(n_22),
.B1(n_51),
.B2(n_42),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_114),
.A2(n_121),
.B1(n_129),
.B2(n_54),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_62),
.A2(n_22),
.B1(n_51),
.B2(n_33),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_60),
.A2(n_45),
.B1(n_38),
.B2(n_50),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_128),
.A2(n_151),
.B1(n_152),
.B2(n_161),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_63),
.A2(n_22),
.B1(n_33),
.B2(n_19),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_55),
.A2(n_27),
.B1(n_47),
.B2(n_46),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_133),
.A2(n_142),
.B1(n_18),
.B2(n_24),
.Y(n_216)
);

OA22x2_ASAP7_75t_L g136 ( 
.A1(n_66),
.A2(n_38),
.B1(n_45),
.B2(n_18),
.Y(n_136)
);

OA22x2_ASAP7_75t_L g223 ( 
.A1(n_136),
.A2(n_154),
.B1(n_15),
.B2(n_9),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_75),
.B(n_49),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_138),
.B(n_140),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_61),
.B(n_49),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_65),
.A2(n_47),
.B1(n_46),
.B2(n_29),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_61),
.B(n_91),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_145),
.B(n_148),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_53),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_88),
.B(n_37),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_150),
.B(n_163),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_58),
.A2(n_45),
.B1(n_38),
.B2(n_19),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_69),
.A2(n_87),
.B1(n_72),
.B2(n_70),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_68),
.A2(n_45),
.B1(n_43),
.B2(n_40),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_95),
.A2(n_18),
.B(n_40),
.Y(n_156)
);

A2O1A1Ixp33_ASAP7_75t_L g221 ( 
.A1(n_156),
.A2(n_6),
.B(n_7),
.C(n_8),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_85),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_160),
.B(n_162),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_56),
.A2(n_43),
.B1(n_35),
.B2(n_29),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_90),
.B(n_35),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_73),
.B(n_27),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_64),
.B(n_1),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_165),
.B(n_2),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_76),
.B(n_2),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_168),
.B(n_99),
.Y(n_175)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_153),
.Y(n_170)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_170),
.Y(n_276)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_112),
.Y(n_171)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_171),
.Y(n_245)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_153),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g257 ( 
.A(n_173),
.Y(n_257)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_141),
.Y(n_174)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_174),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_175),
.B(n_185),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_178),
.B(n_183),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_119),
.B(n_103),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g263 ( 
.A(n_179),
.B(n_180),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_119),
.B(n_102),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_127),
.B(n_81),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_181),
.B(n_182),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_143),
.B(n_130),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_105),
.B(n_97),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_131),
.B(n_99),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_184),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_131),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_186),
.B(n_223),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_157),
.B(n_79),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_187),
.B(n_201),
.Y(n_236)
);

INVx11_ASAP7_75t_L g188 ( 
.A(n_108),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_188),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_107),
.B(n_92),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_189),
.B(n_195),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_190),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_151),
.A2(n_33),
.B1(n_98),
.B2(n_84),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_191),
.A2(n_194),
.B1(n_218),
.B2(n_110),
.Y(n_267)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_120),
.Y(n_192)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_192),
.Y(n_250)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_144),
.Y(n_193)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_193),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_128),
.A2(n_98),
.B1(n_71),
.B2(n_80),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_167),
.B(n_94),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_112),
.Y(n_196)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_196),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_118),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_197),
.B(n_200),
.Y(n_259)
);

AOI32xp33_ASAP7_75t_L g198 ( 
.A1(n_111),
.A2(n_18),
.A3(n_24),
.B1(n_4),
.B2(n_5),
.Y(n_198)
);

AOI32xp33_ASAP7_75t_L g255 ( 
.A1(n_198),
.A2(n_125),
.A3(n_164),
.B1(n_12),
.B2(n_13),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_135),
.B(n_2),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_199),
.B(n_210),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_132),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_126),
.B(n_156),
.Y(n_201)
);

OR2x2_ASAP7_75t_SL g202 ( 
.A(n_120),
.B(n_18),
.Y(n_202)
);

A2O1A1Ixp33_ASAP7_75t_L g251 ( 
.A1(n_202),
.A2(n_203),
.B(n_154),
.C(n_164),
.Y(n_251)
);

OR2x2_ASAP7_75t_SL g203 ( 
.A(n_109),
.B(n_18),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_113),
.Y(n_204)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_204),
.Y(n_258)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_113),
.Y(n_206)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_206),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_115),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_207),
.Y(n_285)
);

BUFx12f_ASAP7_75t_L g208 ( 
.A(n_158),
.Y(n_208)
);

INVx6_ASAP7_75t_L g280 ( 
.A(n_208),
.Y(n_280)
);

BUFx2_ASAP7_75t_L g209 ( 
.A(n_166),
.Y(n_209)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_209),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_106),
.B(n_2),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_116),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_211),
.B(n_213),
.Y(n_260)
);

INVx13_ASAP7_75t_L g212 ( 
.A(n_122),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_212),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_109),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_117),
.B(n_3),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_214),
.B(n_220),
.Y(n_281)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_117),
.Y(n_215)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_215),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_216),
.A2(n_184),
.B1(n_203),
.B2(n_202),
.Y(n_243)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_134),
.Y(n_217)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_217),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_158),
.A2(n_137),
.B1(n_136),
.B2(n_122),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_137),
.B(n_4),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_219),
.B(n_9),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_134),
.B(n_6),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_221),
.A2(n_166),
.B(n_146),
.Y(n_254)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_146),
.Y(n_222)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_222),
.Y(n_246)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_149),
.Y(n_224)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_224),
.Y(n_277)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_149),
.Y(n_225)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_225),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_136),
.B(n_8),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_226),
.B(n_229),
.Y(n_237)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_155),
.Y(n_227)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_227),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_136),
.B(n_9),
.Y(n_229)
);

INVx2_ASAP7_75t_SL g230 ( 
.A(n_159),
.Y(n_230)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_230),
.Y(n_284)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_155),
.Y(n_231)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_231),
.Y(n_247)
);

AO21x2_ASAP7_75t_L g233 ( 
.A1(n_226),
.A2(n_152),
.B(n_161),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_233),
.A2(n_287),
.B1(n_208),
.B2(n_12),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_184),
.B(n_125),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_239),
.Y(n_292)
);

AND2x4_ASAP7_75t_SL g240 ( 
.A(n_201),
.B(n_108),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_240),
.A2(n_254),
.B(n_214),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_243),
.B(n_251),
.Y(n_309)
);

OR2x2_ASAP7_75t_L g307 ( 
.A(n_255),
.B(n_223),
.Y(n_307)
);

A2O1A1Ixp33_ASAP7_75t_L g256 ( 
.A1(n_186),
.A2(n_108),
.B(n_159),
.C(n_123),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_256),
.B(n_221),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_261),
.B(n_209),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_179),
.B(n_123),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_266),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_SL g336 ( 
.A1(n_267),
.A2(n_268),
.B1(n_239),
.B2(n_242),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_229),
.A2(n_124),
.B1(n_110),
.B2(n_169),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_268),
.A2(n_272),
.B1(n_275),
.B2(n_230),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_181),
.B(n_124),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_269),
.B(n_193),
.C(n_175),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_177),
.A2(n_169),
.B1(n_147),
.B2(n_139),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_180),
.B(n_187),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_273),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_228),
.B(n_147),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_274),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_177),
.A2(n_115),
.B1(n_139),
.B2(n_12),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_205),
.B(n_9),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_279),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_176),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_286),
.B(n_172),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_182),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_288),
.B(n_287),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_259),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_289),
.B(n_290),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_260),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_234),
.A2(n_233),
.B1(n_236),
.B2(n_243),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_291),
.A2(n_310),
.B1(n_331),
.B2(n_333),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_237),
.B(n_220),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_294),
.B(n_300),
.Y(n_340)
);

OAI21xp33_ASAP7_75t_L g358 ( 
.A1(n_295),
.A2(n_307),
.B(n_325),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_296),
.B(n_317),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_280),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_297),
.B(n_301),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_298),
.Y(n_349)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_284),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_299),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_237),
.B(n_223),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_280),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_281),
.B(n_223),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_302),
.B(n_306),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_263),
.B(n_174),
.C(n_217),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_303),
.B(n_316),
.C(n_264),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_304),
.A2(n_315),
.B1(n_321),
.B2(n_324),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_244),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_305),
.B(n_314),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_281),
.B(n_196),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_232),
.B(n_269),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_308),
.B(n_311),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_234),
.A2(n_230),
.B1(n_222),
.B2(n_227),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_232),
.B(n_206),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_248),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_233),
.A2(n_272),
.B1(n_275),
.B2(n_234),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_263),
.B(n_204),
.C(n_225),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_262),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_284),
.Y(n_318)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_318),
.Y(n_347)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_249),
.Y(n_319)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_319),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_236),
.B(n_224),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_320),
.B(n_326),
.Y(n_364)
);

AOI22xp33_ASAP7_75t_L g321 ( 
.A1(n_271),
.A2(n_231),
.B1(n_173),
.B2(n_170),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_262),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_322),
.B(n_323),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_233),
.A2(n_215),
.B1(n_171),
.B2(n_207),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_238),
.B(n_213),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_239),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_SL g328 ( 
.A1(n_271),
.A2(n_192),
.B1(n_208),
.B2(n_188),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_328),
.Y(n_365)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_249),
.Y(n_329)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_329),
.Y(n_355)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_258),
.Y(n_330)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_330),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_233),
.A2(n_252),
.B1(n_235),
.B2(n_254),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_273),
.B(n_208),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_332),
.B(n_334),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_273),
.B(n_11),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_240),
.A2(n_212),
.B1(n_13),
.B2(n_14),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g356 ( 
.A1(n_335),
.A2(n_264),
.B(n_277),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_336),
.A2(n_276),
.B1(n_270),
.B2(n_278),
.Y(n_344)
);

A2O1A1O1Ixp25_ASAP7_75t_L g338 ( 
.A1(n_309),
.A2(n_256),
.B(n_251),
.C(n_240),
.D(n_242),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g386 ( 
.A(n_338),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_294),
.B(n_288),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_339),
.B(n_348),
.Y(n_408)
);

NAND2x1_ASAP7_75t_L g342 ( 
.A(n_309),
.B(n_266),
.Y(n_342)
);

INVx1_ASAP7_75t_SL g387 ( 
.A(n_342),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_344),
.A2(n_333),
.B1(n_326),
.B2(n_317),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_309),
.A2(n_276),
.B(n_266),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g379 ( 
.A1(n_345),
.A2(n_298),
.B(n_293),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_299),
.Y(n_346)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_346),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_315),
.A2(n_253),
.B1(n_278),
.B2(n_277),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_350),
.A2(n_370),
.B1(n_292),
.B2(n_310),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_314),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_354),
.B(n_359),
.Y(n_395)
);

INVx1_ASAP7_75t_SL g400 ( 
.A(n_356),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_325),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_L g361 ( 
.A1(n_309),
.A2(n_241),
.B(n_258),
.Y(n_361)
);

INVx1_ASAP7_75t_SL g401 ( 
.A(n_361),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_366),
.B(n_375),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_331),
.A2(n_270),
.B1(n_241),
.B2(n_246),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_367),
.A2(n_372),
.B1(n_330),
.B2(n_329),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_311),
.B(n_283),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_369),
.B(n_373),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_300),
.A2(n_307),
.B1(n_302),
.B2(n_336),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_332),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_371),
.B(n_378),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_291),
.A2(n_283),
.B1(n_265),
.B2(n_285),
.Y(n_372)
);

OAI32xp33_ASAP7_75t_L g373 ( 
.A1(n_312),
.A2(n_247),
.A3(n_245),
.B1(n_282),
.B2(n_250),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_308),
.B(n_245),
.Y(n_375)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_319),
.Y(n_377)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_377),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_316),
.B(n_282),
.C(n_250),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_379),
.Y(n_433)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_343),
.Y(n_381)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_381),
.Y(n_414)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_343),
.Y(n_382)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_382),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_376),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_383),
.B(n_392),
.Y(n_416)
);

OAI22x1_ASAP7_75t_SL g384 ( 
.A1(n_351),
.A2(n_324),
.B1(n_304),
.B2(n_335),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_384),
.A2(n_370),
.B1(n_358),
.B2(n_337),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_385),
.A2(n_398),
.B1(n_403),
.B2(n_367),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_389),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_351),
.A2(n_307),
.B1(n_320),
.B2(n_295),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_391),
.A2(n_363),
.B1(n_375),
.B2(n_348),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_352),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_355),
.Y(n_393)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_393),
.Y(n_431)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_355),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_394),
.B(n_397),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_349),
.A2(n_321),
.B(n_322),
.Y(n_397)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_362),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_399),
.B(n_404),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_350),
.A2(n_313),
.B1(n_306),
.B2(n_305),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_369),
.B(n_334),
.Y(n_404)
);

CKINVDCx14_ASAP7_75t_R g405 ( 
.A(n_341),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_405),
.B(n_406),
.Y(n_434)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_362),
.Y(n_406)
);

CKINVDCx14_ASAP7_75t_R g407 ( 
.A(n_353),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_407),
.B(n_409),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_374),
.B(n_289),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_364),
.B(n_357),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_410),
.B(n_411),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_364),
.B(n_297),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_377),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_412),
.B(n_413),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_SL g413 ( 
.A(n_360),
.B(n_296),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_408),
.B(n_366),
.C(n_339),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_417),
.B(n_430),
.C(n_395),
.Y(n_445)
);

AOI22xp33_ASAP7_75t_SL g449 ( 
.A1(n_418),
.A2(n_426),
.B1(n_400),
.B2(n_388),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_419),
.A2(n_428),
.B1(n_429),
.B2(n_432),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_408),
.B(n_340),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_420),
.B(n_421),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_390),
.B(n_340),
.Y(n_421)
);

XNOR2x2_ASAP7_75t_L g424 ( 
.A(n_403),
.B(n_360),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_424),
.B(n_439),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_425),
.B(n_398),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_409),
.A2(n_372),
.B1(n_290),
.B2(n_349),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_384),
.A2(n_361),
.B1(n_345),
.B2(n_356),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_400),
.A2(n_365),
.B1(n_338),
.B2(n_292),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_390),
.B(n_378),
.C(n_396),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_388),
.A2(n_363),
.B1(n_365),
.B2(n_347),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_396),
.B(n_342),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_437),
.B(n_438),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_391),
.B(n_342),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_410),
.B(n_303),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_386),
.B(n_387),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_440),
.B(n_441),
.C(n_428),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_387),
.B(n_368),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_413),
.B(n_368),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_442),
.B(n_401),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_445),
.B(n_456),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_417),
.B(n_430),
.C(n_420),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_446),
.B(n_462),
.C(n_467),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_447),
.B(n_452),
.Y(n_473)
);

OR2x2_ASAP7_75t_L g448 ( 
.A(n_435),
.B(n_395),
.Y(n_448)
);

CKINVDCx14_ASAP7_75t_R g474 ( 
.A(n_448),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_L g477 ( 
.A1(n_449),
.A2(n_440),
.B1(n_441),
.B2(n_431),
.Y(n_477)
);

BUFx24_ASAP7_75t_SL g451 ( 
.A(n_416),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_451),
.B(n_455),
.Y(n_478)
);

OAI221xp5_ASAP7_75t_L g452 ( 
.A1(n_443),
.A2(n_383),
.B1(n_404),
.B2(n_411),
.C(n_327),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_SL g453 ( 
.A(n_421),
.B(n_401),
.Y(n_453)
);

MAJx2_ASAP7_75t_L g488 ( 
.A(n_453),
.B(n_468),
.C(n_393),
.Y(n_488)
);

HB1xp67_ASAP7_75t_L g469 ( 
.A(n_454),
.Y(n_469)
);

CKINVDCx16_ASAP7_75t_R g455 ( 
.A(n_434),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_439),
.B(n_379),
.Y(n_456)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_436),
.Y(n_458)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_458),
.Y(n_470)
);

NAND3xp33_ASAP7_75t_L g459 ( 
.A(n_427),
.B(n_323),
.C(n_412),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_459),
.B(n_460),
.Y(n_483)
);

OAI21xp5_ASAP7_75t_SL g460 ( 
.A1(n_429),
.A2(n_397),
.B(n_385),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_442),
.B(n_432),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_461),
.B(n_463),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_437),
.B(n_392),
.C(n_352),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_424),
.B(n_381),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_414),
.Y(n_464)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_464),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_423),
.B(n_257),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_465),
.B(n_373),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_438),
.B(n_380),
.C(n_399),
.Y(n_467)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_471),
.Y(n_500)
);

BUFx12_ASAP7_75t_L g472 ( 
.A(n_467),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_472),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_SL g475 ( 
.A1(n_457),
.A2(n_433),
.B1(n_415),
.B2(n_422),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g505 ( 
.A1(n_475),
.A2(n_471),
.B1(n_483),
.B2(n_489),
.Y(n_505)
);

OAI21xp5_ASAP7_75t_SL g476 ( 
.A1(n_448),
.A2(n_433),
.B(n_419),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_SL g498 ( 
.A1(n_476),
.A2(n_489),
.B(n_265),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_477),
.A2(n_453),
.B1(n_444),
.B2(n_456),
.Y(n_491)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_454),
.Y(n_480)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_480),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_446),
.B(n_301),
.C(n_406),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_484),
.B(n_450),
.Y(n_490)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_462),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_485),
.B(n_257),
.Y(n_499)
);

OA21x2_ASAP7_75t_L g486 ( 
.A1(n_457),
.A2(n_389),
.B(n_394),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_486),
.A2(n_473),
.B1(n_470),
.B2(n_475),
.Y(n_506)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_488),
.B(n_285),
.Y(n_502)
);

AOI21xp5_ASAP7_75t_L g489 ( 
.A1(n_468),
.A2(n_382),
.B(n_380),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_490),
.B(n_492),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_491),
.B(n_498),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_484),
.B(n_445),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_481),
.B(n_450),
.C(n_466),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_493),
.B(n_494),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_481),
.B(n_466),
.C(n_444),
.Y(n_494)
);

AOI21xp5_ASAP7_75t_L g495 ( 
.A1(n_476),
.A2(n_318),
.B(n_402),
.Y(n_495)
);

OAI21xp5_ASAP7_75t_SL g507 ( 
.A1(n_495),
.A2(n_506),
.B(n_486),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_485),
.B(n_346),
.Y(n_496)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_496),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_474),
.B(n_402),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_497),
.B(n_479),
.Y(n_515)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_499),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_502),
.B(n_504),
.Y(n_509)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_488),
.B(n_477),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_SL g517 ( 
.A1(n_505),
.A2(n_486),
.B1(n_469),
.B2(n_479),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_507),
.B(n_515),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_SL g508 ( 
.A1(n_501),
.A2(n_487),
.B(n_480),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_508),
.B(n_513),
.Y(n_523)
);

OAI21xp5_ASAP7_75t_SL g513 ( 
.A1(n_501),
.A2(n_472),
.B(n_470),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_SL g522 ( 
.A1(n_517),
.A2(n_491),
.B1(n_500),
.B2(n_503),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_499),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_518),
.B(n_519),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_493),
.B(n_482),
.C(n_472),
.Y(n_519)
);

OAI21x1_ASAP7_75t_SL g521 ( 
.A1(n_514),
.A2(n_506),
.B(n_495),
.Y(n_521)
);

AOI21xp33_ASAP7_75t_L g531 ( 
.A1(n_521),
.A2(n_509),
.B(n_504),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_522),
.B(n_507),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_SL g525 ( 
.A(n_512),
.B(n_478),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_SL g528 ( 
.A(n_525),
.B(n_526),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_510),
.B(n_500),
.Y(n_526)
);

OAI21xp5_ASAP7_75t_SL g527 ( 
.A1(n_517),
.A2(n_503),
.B(n_505),
.Y(n_527)
);

OAI21xp5_ASAP7_75t_SL g530 ( 
.A1(n_527),
.A2(n_498),
.B(n_511),
.Y(n_530)
);

INVxp67_ASAP7_75t_L g535 ( 
.A(n_529),
.Y(n_535)
);

AOI21xp5_ASAP7_75t_L g533 ( 
.A1(n_530),
.A2(n_531),
.B(n_532),
.Y(n_533)
);

CKINVDCx14_ASAP7_75t_R g532 ( 
.A(n_524),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_528),
.B(n_523),
.C(n_519),
.Y(n_534)
);

OAI21xp5_ASAP7_75t_L g536 ( 
.A1(n_534),
.A2(n_520),
.B(n_527),
.Y(n_536)
);

AOI21xp5_ASAP7_75t_L g538 ( 
.A1(n_536),
.A2(n_537),
.B(n_533),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_535),
.B(n_522),
.C(n_494),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_538),
.B(n_516),
.Y(n_539)
);

AOI21xp5_ASAP7_75t_L g540 ( 
.A1(n_539),
.A2(n_516),
.B(n_482),
.Y(n_540)
);

AOI21xp5_ASAP7_75t_L g541 ( 
.A1(n_540),
.A2(n_502),
.B(n_509),
.Y(n_541)
);


endmodule