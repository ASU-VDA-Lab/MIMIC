module fake_jpeg_1627_n_83 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_83);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_83;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_19),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_21),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_36),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_28),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_34),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_0),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_25),
.Y(n_36)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_29),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_27),
.C(n_30),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_34),
.B(n_26),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_42),
.Y(n_47)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_40),
.A2(n_26),
.B1(n_30),
.B2(n_27),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g55 ( 
.A1(n_44),
.A2(n_48),
.B(n_43),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_41),
.A2(n_29),
.B(n_31),
.Y(n_48)
);

NAND3xp33_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_12),
.C(n_24),
.Y(n_58)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_50),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_42),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_52),
.B(n_53),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_48),
.B(n_40),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_49),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_54),
.A2(n_55),
.B1(n_46),
.B2(n_31),
.Y(n_60)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_56),
.B(n_50),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_0),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_58),
.Y(n_64)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_61),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_51),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_51),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_62),
.B(n_65),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_1),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_63),
.A2(n_46),
.B(n_31),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_66),
.B(n_1),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g67 ( 
.A(n_64),
.B(n_9),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_67),
.B(n_13),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_70),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_73),
.A2(n_75),
.B1(n_71),
.B2(n_69),
.Y(n_76)
);

A2O1A1Ixp33_ASAP7_75t_SL g77 ( 
.A1(n_74),
.A2(n_71),
.B(n_3),
.C(n_4),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

NOR2xp67_ASAP7_75t_SL g78 ( 
.A(n_76),
.B(n_77),
.Y(n_78)
);

AOI21xp33_ASAP7_75t_L g79 ( 
.A1(n_78),
.A2(n_72),
.B(n_15),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_79),
.A2(n_11),
.B(n_22),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_80),
.A2(n_8),
.B(n_20),
.Y(n_81)
);

OAI33xp33_ASAP7_75t_L g82 ( 
.A1(n_81),
.A2(n_17),
.A3(n_18),
.B1(n_23),
.B2(n_7),
.B3(n_2),
.Y(n_82)
);

AOI221xp5_ASAP7_75t_L g83 ( 
.A1(n_82),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.C(n_7),
.Y(n_83)
);


endmodule