module fake_jpeg_17393_n_127 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_127);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_127;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_49;
wire n_76;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx12_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_26),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

BUFx24_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_4),
.Y(n_56)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_1),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

BUFx10_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_3),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_42),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_68),
.B(n_69),
.Y(n_88)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_71),
.Y(n_74)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_73),
.Y(n_78)
);

CKINVDCx12_ASAP7_75t_R g79 ( 
.A(n_71),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_80),
.Y(n_94)
);

INVx13_ASAP7_75t_L g80 ( 
.A(n_73),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g97 ( 
.A(n_81),
.Y(n_97)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

INVx3_ASAP7_75t_SL g93 ( 
.A(n_83),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_66),
.A2(n_51),
.B1(n_63),
.B2(n_50),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_85),
.A2(n_86),
.B1(n_52),
.B2(n_53),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_66),
.A2(n_61),
.B1(n_64),
.B2(n_48),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_65),
.B(n_62),
.Y(n_87)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_90),
.B(n_92),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_91),
.Y(n_99)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_95),
.A2(n_81),
.B1(n_84),
.B2(n_74),
.Y(n_102)
);

O2A1O1Ixp33_ASAP7_75t_SL g96 ( 
.A1(n_88),
.A2(n_56),
.B(n_55),
.C(n_49),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_96),
.B(n_44),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_102),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_94),
.B(n_82),
.C(n_47),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_103),
.B(n_104),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_99),
.A2(n_89),
.B1(n_57),
.B2(n_98),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_107),
.A2(n_108),
.B1(n_0),
.B2(n_3),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_100),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_106),
.B(n_101),
.Y(n_109)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_109),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_105),
.A2(n_102),
.B1(n_93),
.B2(n_97),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_110),
.B(n_111),
.C(n_112),
.Y(n_114)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_105),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_113),
.B(n_110),
.C(n_52),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_115),
.B(n_116),
.Y(n_117)
);

XNOR2x1_ASAP7_75t_L g116 ( 
.A(n_114),
.B(n_44),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_22),
.C(n_5),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_118),
.A2(n_24),
.B1(n_6),
.B2(n_7),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_119),
.A2(n_29),
.B1(n_8),
.B2(n_9),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_31),
.C(n_10),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_121),
.B(n_32),
.Y(n_122)
);

OAI311xp33_ASAP7_75t_L g123 ( 
.A1(n_122),
.A2(n_33),
.A3(n_11),
.B1(n_12),
.C1(n_13),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_123),
.A2(n_36),
.B(n_14),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_37),
.C(n_16),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_125),
.A2(n_38),
.B(n_19),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_25),
.Y(n_127)
);


endmodule