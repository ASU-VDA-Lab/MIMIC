module fake_jpeg_7804_n_170 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_170);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_170;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_12),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx11_ASAP7_75t_SL g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_34),
.Y(n_45)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_22),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_37),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_15),
.B(n_0),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_39),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_31),
.A2(n_22),
.B1(n_27),
.B2(n_29),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_23),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_47),
.B(n_55),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_36),
.A2(n_27),
.B1(n_23),
.B2(n_16),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_50),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_L g53 ( 
.A1(n_39),
.A2(n_27),
.B1(n_35),
.B2(n_31),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_35),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_34),
.B(n_23),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_31),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_28),
.Y(n_57)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_61),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_60),
.A2(n_63),
.B1(n_62),
.B2(n_54),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_50),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_35),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_63),
.Y(n_81)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_28),
.Y(n_66)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_18),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_69),
.Y(n_82)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_52),
.B(n_29),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_71),
.B(n_17),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_17),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_72),
.A2(n_17),
.B(n_29),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_74),
.A2(n_78),
.B1(n_90),
.B2(n_25),
.Y(n_96)
);

AO22x1_ASAP7_75t_L g75 ( 
.A1(n_72),
.A2(n_54),
.B1(n_39),
.B2(n_32),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_80),
.Y(n_92)
);

NOR3xp33_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_71),
.C(n_67),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_60),
.A2(n_30),
.B1(n_34),
.B2(n_15),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_68),
.B(n_21),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_72),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_70),
.A2(n_30),
.B1(n_49),
.B2(n_44),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_84),
.A2(n_91),
.B1(n_14),
.B2(n_16),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_57),
.B(n_33),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_89),
.C(n_77),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_66),
.B(n_26),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_87),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_68),
.B(n_33),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_59),
.A2(n_30),
.B1(n_18),
.B2(n_26),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_58),
.A2(n_14),
.B1(n_25),
.B2(n_21),
.Y(n_91)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_93),
.B(n_96),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_107),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_97),
.B(n_99),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_98),
.A2(n_103),
.B1(n_65),
.B2(n_64),
.Y(n_122)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_69),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_102),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_101),
.B(n_105),
.C(n_88),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_61),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_74),
.A2(n_78),
.B1(n_90),
.B2(n_86),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_42),
.Y(n_104)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_104),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_76),
.B(n_33),
.C(n_50),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_91),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_106),
.B(n_80),
.Y(n_109)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_108),
.B(n_115),
.C(n_101),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_109),
.B(n_114),
.Y(n_126)
);

OA21x2_ASAP7_75t_L g112 ( 
.A1(n_93),
.A2(n_75),
.B(n_84),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_112),
.B(n_118),
.Y(n_132)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_104),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_102),
.B(n_75),
.C(n_49),
.Y(n_115)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_105),
.Y(n_119)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_119),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_94),
.B(n_64),
.Y(n_120)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_120),
.Y(n_127)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_103),
.Y(n_121)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_121),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_122),
.A2(n_107),
.B1(n_99),
.B2(n_65),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_123),
.B(n_134),
.C(n_110),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_125),
.B(n_128),
.Y(n_141)
);

NOR3xp33_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_92),
.C(n_97),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_115),
.A2(n_92),
.B(n_100),
.Y(n_129)
);

AO21x1_ASAP7_75t_L g144 ( 
.A1(n_129),
.A2(n_24),
.B(n_42),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g131 ( 
.A(n_112),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_131),
.B(n_133),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_113),
.A2(n_96),
.B1(n_94),
.B2(n_65),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_111),
.B(n_33),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_123),
.B(n_108),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_135),
.B(n_136),
.C(n_137),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_129),
.B(n_111),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_127),
.B(n_116),
.Y(n_138)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_138),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_126),
.B(n_114),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_139),
.B(n_140),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_124),
.B(n_110),
.C(n_122),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_134),
.B(n_112),
.Y(n_142)
);

AOI321xp33_ASAP7_75t_L g147 ( 
.A1(n_142),
.A2(n_144),
.A3(n_43),
.B1(n_1),
.B2(n_2),
.C(n_3),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_143),
.A2(n_130),
.B1(n_132),
.B2(n_131),
.Y(n_145)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_145),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_147),
.B(n_6),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_141),
.A2(n_8),
.B1(n_12),
.B2(n_11),
.Y(n_148)
);

CKINVDCx14_ASAP7_75t_R g158 ( 
.A(n_148),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_144),
.A2(n_8),
.B(n_11),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_151),
.B(n_152),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_137),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_150),
.B(n_136),
.C(n_6),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_154),
.B(n_156),
.Y(n_160)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_155),
.Y(n_162)
);

AOI21x1_ASAP7_75t_L g156 ( 
.A1(n_149),
.A2(n_146),
.B(n_152),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_153),
.A2(n_150),
.B1(n_10),
.B2(n_13),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_159),
.B(n_0),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_158),
.A2(n_13),
.B1(n_2),
.B2(n_4),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_161),
.B(n_0),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_157),
.B(n_155),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_154),
.Y(n_164)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_164),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_165),
.A2(n_166),
.B(n_163),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_160),
.C(n_162),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_169),
.B(n_167),
.Y(n_170)
);


endmodule