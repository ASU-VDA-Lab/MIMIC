module fake_jpeg_25417_n_304 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_304);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_304;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_14;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_273;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_303;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_294;
wire n_300;
wire n_211;
wire n_299;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx3_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx14_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_26),
.Y(n_27)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_17),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_29),
.B(n_30),
.Y(n_42)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_19),
.B(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_34),
.Y(n_44)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

OR2x2_ASAP7_75t_L g36 ( 
.A(n_35),
.B(n_20),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_36),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_27),
.A2(n_31),
.B1(n_30),
.B2(n_13),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_38),
.A2(n_47),
.B1(n_30),
.B2(n_34),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_27),
.A2(n_13),
.B1(n_18),
.B2(n_15),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_39),
.A2(n_27),
.B1(n_32),
.B2(n_28),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_20),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_45),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_27),
.A2(n_13),
.B1(n_26),
.B2(n_22),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_41),
.A2(n_30),
.B1(n_34),
.B2(n_32),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_20),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_27),
.A2(n_26),
.B1(n_22),
.B2(n_20),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_31),
.B(n_23),
.Y(n_48)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_50),
.A2(n_56),
.B1(n_41),
.B2(n_49),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_43),
.A2(n_17),
.B1(n_25),
.B2(n_15),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_49),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_43),
.A2(n_25),
.B1(n_18),
.B2(n_32),
.Y(n_56)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_29),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_62),
.B(n_70),
.Y(n_87)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_71),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_66),
.A2(n_68),
.B1(n_49),
.B2(n_30),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_32),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_67),
.A2(n_36),
.B(n_44),
.Y(n_76)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

BUFx24_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_45),
.B(n_28),
.C(n_32),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_76),
.A2(n_67),
.B(n_44),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_78),
.A2(n_95),
.B1(n_66),
.B2(n_67),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_29),
.Y(n_80)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_80),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_68),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_82),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_55),
.B(n_29),
.Y(n_84)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_84),
.Y(n_118)
);

INVx13_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_85),
.Y(n_108)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_53),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_90),
.B(n_91),
.Y(n_109)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_64),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_92),
.B(n_71),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_93),
.A2(n_57),
.B1(n_60),
.B2(n_39),
.Y(n_101)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_94),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_62),
.A2(n_45),
.B1(n_44),
.B2(n_38),
.Y(n_95)
);

BUFx8_ASAP7_75t_L g96 ( 
.A(n_63),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g121 ( 
.A(n_96),
.Y(n_121)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_72),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_97),
.B(n_103),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_95),
.B(n_59),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_117),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_101),
.A2(n_102),
.B1(n_89),
.B2(n_34),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_82),
.A2(n_70),
.B1(n_59),
.B2(n_57),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_78),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_52),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_SL g135 ( 
.A(n_104),
.B(n_115),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_105),
.A2(n_47),
.B1(n_49),
.B2(n_91),
.Y(n_128)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_106),
.B(n_112),
.Y(n_143)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_79),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_107),
.B(n_114),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_74),
.A2(n_87),
.B(n_76),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_110),
.A2(n_111),
.B(n_120),
.Y(n_144)
);

OR2x2_ASAP7_75t_SL g111 ( 
.A(n_81),
.B(n_52),
.Y(n_111)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_75),
.Y(n_112)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_93),
.Y(n_114)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_116),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_81),
.B(n_83),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_74),
.A2(n_49),
.B1(n_48),
.B2(n_58),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_119),
.A2(n_96),
.B1(n_73),
.B2(n_35),
.Y(n_147)
);

O2A1O1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_83),
.A2(n_46),
.B(n_48),
.C(n_28),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_86),
.B(n_36),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_122),
.B(n_36),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_117),
.B(n_86),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_123),
.B(n_152),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_104),
.B(n_36),
.C(n_92),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_124),
.B(n_136),
.C(n_137),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_126),
.B(n_130),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_128),
.A2(n_132),
.B1(n_134),
.B2(n_138),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_129),
.B(n_73),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_100),
.B(n_89),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_114),
.A2(n_90),
.B(n_96),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_131),
.A2(n_153),
.B(n_33),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_103),
.A2(n_99),
.B1(n_105),
.B2(n_110),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_102),
.A2(n_61),
.B1(n_69),
.B2(n_94),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_115),
.B(n_122),
.C(n_97),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_28),
.C(n_33),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_120),
.A2(n_75),
.B1(n_85),
.B2(n_88),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_77),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_139),
.B(n_146),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_119),
.B(n_28),
.C(n_35),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_141),
.B(n_77),
.C(n_35),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_109),
.A2(n_34),
.B1(n_47),
.B2(n_46),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_142),
.A2(n_145),
.B1(n_147),
.B2(n_151),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_111),
.A2(n_34),
.B1(n_46),
.B2(n_96),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_106),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_107),
.B(n_77),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_148),
.B(n_154),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_108),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_149),
.B(n_35),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_112),
.A2(n_24),
.B1(n_16),
.B2(n_14),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_150),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_98),
.A2(n_108),
.B1(n_14),
.B2(n_24),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_98),
.B(n_73),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_121),
.A2(n_23),
.B(n_16),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_121),
.A2(n_24),
.B1(n_16),
.B2(n_14),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_139),
.B(n_121),
.Y(n_155)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_155),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_135),
.B(n_33),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_156),
.B(n_159),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_148),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_157),
.B(n_161),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_134),
.B(n_121),
.Y(n_158)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_158),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_135),
.B(n_33),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_160),
.B(n_174),
.Y(n_210)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_143),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_133),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_162),
.B(n_168),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_166),
.B(n_33),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_151),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_138),
.Y(n_169)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_169),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_123),
.Y(n_170)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_170),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_137),
.Y(n_173)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_173),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_136),
.B(n_21),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_140),
.B(n_35),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_175),
.A2(n_181),
.B(n_185),
.Y(n_205)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_132),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_176),
.B(n_180),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_127),
.B(n_79),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_179),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_144),
.A2(n_0),
.B(n_1),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_130),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_182),
.B(n_186),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_124),
.B(n_35),
.C(n_33),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_183),
.B(n_184),
.C(n_147),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_129),
.B(n_126),
.C(n_125),
.Y(n_184)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_145),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_144),
.A2(n_0),
.B(n_1),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_187),
.A2(n_153),
.B1(n_154),
.B2(n_3),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_177),
.A2(n_125),
.B1(n_141),
.B2(n_131),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_188),
.A2(n_203),
.B1(n_209),
.B2(n_175),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_191),
.B(n_199),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_163),
.B(n_127),
.C(n_146),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_192),
.B(n_1),
.C(n_2),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_193),
.A2(n_12),
.B1(n_11),
.B2(n_3),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_186),
.A2(n_149),
.B1(n_142),
.B2(n_79),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_195),
.A2(n_204),
.B1(n_172),
.B2(n_166),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_163),
.B(n_79),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_201),
.B(n_183),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_177),
.A2(n_178),
.B1(n_165),
.B2(n_172),
.Y(n_202)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_202),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_178),
.A2(n_182),
.B1(n_184),
.B2(n_185),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_160),
.A2(n_22),
.B1(n_21),
.B2(n_3),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_161),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_206),
.B(n_171),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_167),
.B(n_22),
.Y(n_207)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_207),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_171),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_214),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_215),
.B(n_218),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_200),
.B(n_164),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_216),
.B(n_217),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_211),
.B(n_164),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_206),
.B(n_187),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_220),
.B(n_222),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_221),
.B(n_191),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_198),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_189),
.B(n_175),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_223),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_203),
.A2(n_159),
.B1(n_156),
.B2(n_174),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_226),
.A2(n_227),
.B(n_228),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_205),
.A2(n_181),
.B(n_2),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_198),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_196),
.B(n_21),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_229),
.B(n_231),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_230),
.Y(n_249)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_208),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_197),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_232),
.B(n_210),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_233),
.B(n_209),
.C(n_210),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_219),
.B(n_196),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_237),
.Y(n_253)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_239),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_219),
.B(n_192),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_240),
.B(n_229),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_216),
.Y(n_241)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_241),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_221),
.B(n_199),
.C(n_213),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_242),
.B(n_246),
.C(n_233),
.Y(n_255)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_245),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_226),
.B(n_201),
.C(n_188),
.Y(n_246)
);

NOR2xp67_ASAP7_75t_SL g250 ( 
.A(n_242),
.B(n_212),
.Y(n_250)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_250),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_243),
.B(n_234),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_252),
.B(n_258),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_254),
.B(n_255),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_247),
.A2(n_218),
.B1(n_224),
.B2(n_190),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_256),
.A2(n_259),
.B1(n_261),
.B2(n_263),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_244),
.A2(n_227),
.B(n_223),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_246),
.A2(n_194),
.B1(n_195),
.B2(n_217),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_249),
.A2(n_197),
.B1(n_215),
.B2(n_204),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_238),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_262),
.B(n_2),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_249),
.A2(n_225),
.B1(n_205),
.B2(n_207),
.Y(n_263)
);

OAI22xp33_ASAP7_75t_L g266 ( 
.A1(n_258),
.A2(n_248),
.B1(n_239),
.B2(n_237),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_266),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_282)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_257),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_267),
.B(n_271),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_259),
.A2(n_236),
.B1(n_235),
.B2(n_240),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_270),
.B(n_272),
.C(n_274),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_261),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_263),
.B(n_4),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_273),
.B(n_275),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_255),
.B(n_5),
.C(n_6),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_251),
.B(n_5),
.Y(n_275)
);

NOR2x1_ASAP7_75t_L g278 ( 
.A(n_268),
.B(n_260),
.Y(n_278)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_278),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_272),
.B(n_254),
.Y(n_279)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_279),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_269),
.B(n_253),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_280),
.B(n_282),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_264),
.B(n_253),
.Y(n_281)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_281),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_265),
.B(n_7),
.Y(n_283)
);

NAND2xp33_ASAP7_75t_SL g289 ( 
.A(n_283),
.B(n_285),
.Y(n_289)
);

OR2x2_ASAP7_75t_L g285 ( 
.A(n_274),
.B(n_7),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_281),
.A2(n_266),
.B(n_269),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_287),
.A2(n_276),
.B(n_277),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_284),
.B(n_270),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_290),
.B(n_293),
.Y(n_298)
);

NOR2x1_ASAP7_75t_L g293 ( 
.A(n_278),
.B(n_7),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_291),
.B(n_292),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_294),
.B(n_295),
.Y(n_299)
);

AOI21xp33_ASAP7_75t_L g296 ( 
.A1(n_288),
.A2(n_285),
.B(n_9),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_296),
.B(n_297),
.Y(n_300)
);

AO21x1_ASAP7_75t_L g297 ( 
.A1(n_286),
.A2(n_8),
.B(n_9),
.Y(n_297)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_300),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_301),
.B(n_298),
.C(n_299),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_302),
.B(n_289),
.C(n_293),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_303),
.A2(n_8),
.B1(n_10),
.B2(n_301),
.Y(n_304)
);


endmodule