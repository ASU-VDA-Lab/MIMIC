module fake_jpeg_22513_n_301 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_301);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_301;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_273;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_102;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx6_ASAP7_75t_SL g33 ( 
.A(n_15),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

CKINVDCx6p67_ASAP7_75t_R g46 ( 
.A(n_35),
.Y(n_46)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_18),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_26),
.Y(n_49)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

CKINVDCx6p67_ASAP7_75t_R g58 ( 
.A(n_40),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_20),
.B(n_6),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_42),
.Y(n_48)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_29),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_49),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_36),
.A2(n_21),
.B1(n_18),
.B2(n_26),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_47),
.A2(n_53),
.B1(n_17),
.B2(n_27),
.Y(n_76)
);

INVx2_ASAP7_75t_SL g50 ( 
.A(n_35),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_42),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_36),
.A2(n_21),
.B1(n_26),
.B2(n_20),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_51),
.A2(n_38),
.B1(n_42),
.B2(n_32),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_39),
.A2(n_21),
.B1(n_29),
.B2(n_20),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_59),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_56),
.Y(n_60)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_37),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_61),
.B(n_17),
.C(n_27),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_63),
.Y(n_102)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_65),
.B(n_73),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_48),
.Y(n_66)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_66),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_45),
.B(n_20),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_68),
.B(n_69),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_29),
.Y(n_69)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_70),
.A2(n_81),
.B1(n_87),
.B2(n_89),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_49),
.B(n_32),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_71),
.B(n_75),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_72),
.A2(n_92),
.B(n_25),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_58),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_58),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_74),
.B(n_78),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_32),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_76),
.A2(n_52),
.B1(n_55),
.B2(n_27),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_45),
.B(n_17),
.Y(n_77)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_77),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_58),
.Y(n_78)
);

A2O1A1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_47),
.A2(n_33),
.B(n_25),
.C(n_24),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_79),
.B(n_82),
.Y(n_113)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_80),
.Y(n_108)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_46),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_52),
.A2(n_34),
.B1(n_38),
.B2(n_40),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_83),
.A2(n_34),
.B1(n_54),
.B2(n_30),
.Y(n_107)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_46),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_85),
.B(n_88),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_43),
.B(n_23),
.Y(n_86)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_86),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_43),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_57),
.B(n_30),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_50),
.Y(n_112)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_91),
.A2(n_50),
.B1(n_57),
.B2(n_59),
.Y(n_101)
);

A2O1A1Ixp33_ASAP7_75t_L g92 ( 
.A1(n_55),
.A2(n_33),
.B(n_16),
.C(n_31),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_93),
.A2(n_60),
.B1(n_23),
.B2(n_9),
.Y(n_149)
);

NAND2xp33_ASAP7_75t_SL g95 ( 
.A(n_61),
.B(n_0),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_95),
.B(n_100),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_65),
.A2(n_76),
.B1(n_71),
.B2(n_69),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_96),
.A2(n_79),
.B1(n_90),
.B2(n_75),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_67),
.B(n_0),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_101),
.Y(n_139)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_66),
.B(n_33),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_68),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_111),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_67),
.B(n_0),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_105),
.A2(n_119),
.B(n_121),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_107),
.A2(n_115),
.B1(n_16),
.B2(n_19),
.Y(n_126)
);

XOR2x2_ASAP7_75t_SL g111 ( 
.A(n_67),
.B(n_33),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_112),
.B(n_63),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_92),
.A2(n_30),
.B1(n_31),
.B2(n_28),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_73),
.B(n_31),
.C(n_28),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_116),
.B(n_77),
.C(n_19),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_91),
.A2(n_28),
.B1(n_25),
.B2(n_24),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_118),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_91),
.A2(n_24),
.B1(n_22),
.B2(n_19),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_122),
.A2(n_135),
.B1(n_141),
.B2(n_109),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_114),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_123),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_124),
.A2(n_142),
.B(n_94),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g125 ( 
.A(n_119),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_125),
.B(n_0),
.Y(n_181)
);

OAI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_126),
.A2(n_149),
.B1(n_109),
.B2(n_60),
.Y(n_171)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_114),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_127),
.B(n_131),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_128),
.B(n_129),
.C(n_104),
.Y(n_155)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_106),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_113),
.A2(n_78),
.B1(n_74),
.B2(n_84),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_133),
.A2(n_137),
.B1(n_143),
.B2(n_147),
.Y(n_152)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_106),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_134),
.B(n_145),
.Y(n_167)
);

OA21x2_ASAP7_75t_L g135 ( 
.A1(n_113),
.A2(n_85),
.B(n_83),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_107),
.A2(n_80),
.B1(n_62),
.B2(n_82),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_108),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_138),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_108),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_140),
.Y(n_182)
);

OA21x2_ASAP7_75t_L g141 ( 
.A1(n_111),
.A2(n_16),
.B(n_22),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_97),
.A2(n_88),
.B(n_64),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_97),
.A2(n_64),
.B1(n_70),
.B2(n_81),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_112),
.B(n_70),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_144),
.B(n_150),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_120),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_96),
.A2(n_81),
.B1(n_60),
.B2(n_22),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_116),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_148),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_115),
.B(n_23),
.Y(n_150)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_143),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_153),
.B(n_158),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_154),
.A2(n_157),
.B(n_162),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_155),
.B(n_160),
.C(n_136),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_125),
.A2(n_98),
.B1(n_102),
.B2(n_110),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_156),
.A2(n_171),
.B1(n_173),
.B2(n_174),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_132),
.A2(n_99),
.B(n_94),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_142),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_137),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_159),
.B(n_163),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_144),
.B(n_99),
.C(n_117),
.Y(n_160)
);

XOR2x2_ASAP7_75t_L g162 ( 
.A(n_128),
.B(n_95),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_147),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_132),
.A2(n_103),
.B(n_102),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_164),
.A2(n_131),
.B(n_134),
.Y(n_191)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_138),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_165),
.B(n_169),
.Y(n_206)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_133),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_129),
.Y(n_170)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_170),
.Y(n_184)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_140),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_172),
.B(n_127),
.Y(n_186)
);

OAI22x1_ASAP7_75t_L g173 ( 
.A1(n_139),
.A2(n_103),
.B1(n_105),
.B2(n_100),
.Y(n_173)
);

XNOR2x1_ASAP7_75t_L g175 ( 
.A(n_136),
.B(n_105),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_175),
.B(n_130),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_126),
.Y(n_176)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_176),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_148),
.A2(n_110),
.B1(n_117),
.B2(n_100),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_177),
.A2(n_181),
.B1(n_146),
.B2(n_141),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_145),
.B(n_23),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_178),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_123),
.B(n_23),
.Y(n_179)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_179),
.Y(n_207)
);

A2O1A1Ixp33_ASAP7_75t_L g185 ( 
.A1(n_174),
.A2(n_162),
.B(n_173),
.C(n_166),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_185),
.A2(n_188),
.B(n_191),
.Y(n_226)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_186),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_156),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_187),
.B(n_190),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_166),
.B(n_124),
.Y(n_188)
);

OA21x2_ASAP7_75t_L g189 ( 
.A1(n_158),
.A2(n_135),
.B(n_141),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_189),
.A2(n_163),
.B(n_165),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_182),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_192),
.B(n_203),
.C(n_208),
.Y(n_211)
);

OAI32xp33_ASAP7_75t_L g193 ( 
.A1(n_151),
.A2(n_122),
.A3(n_135),
.B1(n_141),
.B2(n_150),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_193),
.B(n_194),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_161),
.B(n_130),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_195),
.B(n_164),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_168),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_200),
.B(n_202),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_154),
.B(n_180),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_201),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_157),
.B(n_130),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_180),
.A2(n_135),
.B1(n_2),
.B2(n_3),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_204),
.A2(n_152),
.B1(n_172),
.B2(n_11),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_160),
.B(n_1),
.C(n_2),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_167),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_209),
.A2(n_9),
.B1(n_4),
.B2(n_5),
.Y(n_224)
);

FAx1_ASAP7_75t_SL g210 ( 
.A(n_197),
.B(n_151),
.CI(n_175),
.CON(n_210),
.SN(n_210)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_210),
.B(n_220),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_212),
.B(n_219),
.C(n_203),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_187),
.A2(n_169),
.B1(n_159),
.B2(n_153),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_214),
.A2(n_199),
.B1(n_9),
.B2(n_11),
.Y(n_248)
);

OA21x2_ASAP7_75t_L g215 ( 
.A1(n_189),
.A2(n_182),
.B(n_168),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_215),
.A2(n_217),
.B(n_199),
.Y(n_241)
);

OAI21xp33_ASAP7_75t_L g216 ( 
.A1(n_194),
.A2(n_179),
.B(n_177),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_216),
.B(n_189),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_218),
.A2(n_224),
.B1(n_229),
.B2(n_209),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_192),
.B(n_155),
.C(n_152),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_206),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_205),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_221),
.A2(n_222),
.B1(n_185),
.B2(n_201),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_183),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_191),
.A2(n_3),
.B(n_5),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_204),
.B(n_7),
.Y(n_230)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_230),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_215),
.B(n_186),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_231),
.B(n_243),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_233),
.A2(n_237),
.B1(n_238),
.B2(n_239),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_219),
.B(n_197),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_234),
.B(n_240),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_215),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_235),
.B(n_241),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_227),
.A2(n_196),
.B1(n_198),
.B2(n_184),
.Y(n_238)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_213),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_242),
.B(n_244),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_221),
.B(n_207),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_225),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_211),
.B(n_207),
.C(n_208),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_245),
.B(n_211),
.C(n_223),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_227),
.A2(n_188),
.B1(n_193),
.B2(n_195),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_246),
.A2(n_248),
.B1(n_218),
.B2(n_222),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_223),
.B(n_188),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_247),
.B(n_228),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_249),
.B(n_258),
.C(n_262),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_247),
.B(n_214),
.Y(n_251)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_251),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_234),
.B(n_212),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_253),
.B(n_259),
.Y(n_264)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_255),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_245),
.B(n_240),
.C(n_228),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_236),
.B(n_226),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_246),
.B(n_226),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_238),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_261),
.B(n_237),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_241),
.A2(n_217),
.B(n_210),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_268),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_SL g267 ( 
.A(n_257),
.B(n_239),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_267),
.B(n_269),
.Y(n_278)
);

CKINVDCx14_ASAP7_75t_R g268 ( 
.A(n_250),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_256),
.B(n_232),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_270),
.B(n_272),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_254),
.B(n_248),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_259),
.B(n_210),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_273),
.B(n_260),
.C(n_258),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_252),
.B(n_229),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_274),
.B(n_251),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_271),
.B(n_249),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_275),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_276),
.B(n_264),
.C(n_267),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_277),
.A2(n_279),
.B(n_282),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_268),
.B(n_254),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_263),
.B(n_7),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_266),
.B(n_7),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_283),
.B(n_12),
.Y(n_287)
);

NOR2xp67_ASAP7_75t_L g285 ( 
.A(n_276),
.B(n_269),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_285),
.B(n_287),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_286),
.A2(n_290),
.B(n_14),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_SL g289 ( 
.A(n_278),
.B(n_273),
.Y(n_289)
);

INVx6_ASAP7_75t_L g292 ( 
.A(n_289),
.Y(n_292)
);

NOR3xp33_ASAP7_75t_L g290 ( 
.A(n_280),
.B(n_12),
.C(n_14),
.Y(n_290)
);

A2O1A1Ixp33_ASAP7_75t_SL g291 ( 
.A1(n_284),
.A2(n_278),
.B(n_281),
.C(n_14),
.Y(n_291)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_291),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_293),
.B(n_287),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_295),
.B(n_294),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_297),
.Y(n_298)
);

O2A1O1Ixp33_ASAP7_75t_L g299 ( 
.A1(n_298),
.A2(n_296),
.B(n_288),
.C(n_292),
.Y(n_299)
);

NAND2xp33_ASAP7_75t_SL g300 ( 
.A(n_299),
.B(n_15),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_300),
.B(n_15),
.Y(n_301)
);


endmodule