module real_aes_6773_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_726, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_726;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_666;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_310;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_417;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_713;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_717;
wire n_456;
wire n_712;
wire n_183;
wire n_312;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g468 ( .A1(n_0), .A2(n_206), .B(n_469), .C(n_472), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_1), .B(n_463), .Y(n_473) );
INVx1_ASAP7_75t_L g113 ( .A(n_2), .Y(n_113) );
INVx1_ASAP7_75t_L g241 ( .A(n_3), .Y(n_241) );
NAND2xp5_ASAP7_75t_SL g453 ( .A(n_4), .B(n_158), .Y(n_453) );
AOI21xp5_ASAP7_75t_L g545 ( .A1(n_5), .A2(n_458), .B(n_546), .Y(n_545) );
AO21x2_ASAP7_75t_L g507 ( .A1(n_6), .A2(n_181), .B(n_508), .Y(n_507) );
AOI22xp33_ASAP7_75t_L g205 ( .A1(n_7), .A2(n_38), .B1(n_151), .B2(n_175), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_8), .B(n_181), .Y(n_253) );
AND2x6_ASAP7_75t_L g166 ( .A(n_9), .B(n_167), .Y(n_166) );
A2O1A1Ixp33_ASAP7_75t_L g521 ( .A1(n_10), .A2(n_166), .B(n_449), .C(n_522), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_11), .B(n_39), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g128 ( .A(n_11), .B(n_39), .Y(n_128) );
INVx1_ASAP7_75t_L g147 ( .A(n_12), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_13), .B(n_156), .Y(n_189) );
INVx1_ASAP7_75t_L g233 ( .A(n_14), .Y(n_233) );
OAI22xp5_ASAP7_75t_SL g716 ( .A1(n_15), .A2(n_75), .B1(n_717), .B2(n_718), .Y(n_716) );
CKINVDCx20_ASAP7_75t_R g718 ( .A(n_15), .Y(n_718) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_16), .B(n_158), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_17), .B(n_182), .Y(n_220) );
AO32x2_ASAP7_75t_L g203 ( .A1(n_18), .A2(n_180), .A3(n_181), .B1(n_204), .B2(n_208), .Y(n_203) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_19), .B(n_151), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_20), .B(n_182), .Y(n_243) );
AOI22xp33_ASAP7_75t_L g207 ( .A1(n_21), .A2(n_55), .B1(n_151), .B2(n_175), .Y(n_207) );
AOI22xp33_ASAP7_75t_SL g178 ( .A1(n_22), .A2(n_83), .B1(n_151), .B2(n_156), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g162 ( .A(n_23), .B(n_151), .Y(n_162) );
A2O1A1Ixp33_ASAP7_75t_L g495 ( .A1(n_24), .A2(n_180), .B(n_449), .C(n_496), .Y(n_495) );
A2O1A1Ixp33_ASAP7_75t_L g510 ( .A1(n_25), .A2(n_180), .B(n_449), .C(n_511), .Y(n_510) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_26), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_27), .B(n_143), .Y(n_262) );
OAI22xp5_ASAP7_75t_SL g703 ( .A1(n_28), .A2(n_94), .B1(n_704), .B2(n_705), .Y(n_703) );
CKINVDCx20_ASAP7_75t_R g705 ( .A(n_28), .Y(n_705) );
AOI22xp5_ASAP7_75t_L g701 ( .A1(n_29), .A2(n_702), .B1(n_703), .B2(n_706), .Y(n_701) );
CKINVDCx20_ASAP7_75t_R g706 ( .A(n_29), .Y(n_706) );
AOI21xp5_ASAP7_75t_L g464 ( .A1(n_30), .A2(n_458), .B(n_465), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_31), .B(n_143), .Y(n_168) );
INVx2_ASAP7_75t_L g153 ( .A(n_32), .Y(n_153) );
A2O1A1Ixp33_ASAP7_75t_L g480 ( .A1(n_33), .A2(n_455), .B(n_481), .C(n_482), .Y(n_480) );
NAND2xp5_ASAP7_75t_SL g257 ( .A(n_34), .B(n_151), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_35), .B(n_143), .Y(n_196) );
OAI22xp5_ASAP7_75t_SL g721 ( .A1(n_36), .A2(n_43), .B1(n_439), .B2(n_722), .Y(n_721) );
CKINVDCx20_ASAP7_75t_R g722 ( .A(n_36), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_37), .B(n_191), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_40), .B(n_494), .Y(n_493) );
CKINVDCx20_ASAP7_75t_R g526 ( .A(n_41), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_42), .B(n_158), .Y(n_534) );
OAI22xp5_ASAP7_75t_SL g133 ( .A1(n_43), .A2(n_134), .B1(n_439), .B2(n_440), .Y(n_133) );
INVx1_ASAP7_75t_L g439 ( .A(n_43), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_44), .B(n_458), .Y(n_509) );
A2O1A1Ixp33_ASAP7_75t_L g531 ( .A1(n_45), .A2(n_455), .B(n_481), .C(n_532), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g248 ( .A(n_46), .B(n_151), .Y(n_248) );
INVx1_ASAP7_75t_L g470 ( .A(n_47), .Y(n_470) );
AOI22xp5_ASAP7_75t_SL g130 ( .A1(n_48), .A2(n_126), .B1(n_131), .B2(n_709), .Y(n_130) );
AOI22xp33_ASAP7_75t_L g174 ( .A1(n_49), .A2(n_92), .B1(n_175), .B2(n_176), .Y(n_174) );
INVx1_ASAP7_75t_L g533 ( .A(n_50), .Y(n_533) );
NAND2xp5_ASAP7_75t_SL g251 ( .A(n_51), .B(n_151), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_52), .B(n_151), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_53), .B(n_458), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_54), .B(n_239), .Y(n_252) );
AOI22xp33_ASAP7_75t_SL g224 ( .A1(n_56), .A2(n_60), .B1(n_151), .B2(n_156), .Y(n_224) );
CKINVDCx20_ASAP7_75t_R g501 ( .A(n_57), .Y(n_501) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_58), .B(n_151), .Y(n_188) );
NAND2xp5_ASAP7_75t_SL g261 ( .A(n_59), .B(n_151), .Y(n_261) );
INVx1_ASAP7_75t_L g167 ( .A(n_61), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_62), .B(n_458), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_63), .B(n_463), .Y(n_551) );
A2O1A1Ixp33_ASAP7_75t_L g548 ( .A1(n_64), .A2(n_236), .B(n_239), .C(n_549), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_65), .B(n_151), .Y(n_242) );
INVx1_ASAP7_75t_L g146 ( .A(n_66), .Y(n_146) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_67), .Y(n_122) );
NAND2xp5_ASAP7_75t_SL g486 ( .A(n_68), .B(n_158), .Y(n_486) );
AO32x2_ASAP7_75t_L g172 ( .A1(n_69), .A2(n_173), .A3(n_179), .B1(n_180), .B2(n_181), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_70), .B(n_159), .Y(n_523) );
INVx1_ASAP7_75t_L g260 ( .A(n_71), .Y(n_260) );
INVx1_ASAP7_75t_L g154 ( .A(n_72), .Y(n_154) );
CKINVDCx16_ASAP7_75t_R g466 ( .A(n_73), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_74), .B(n_485), .Y(n_497) );
CKINVDCx20_ASAP7_75t_R g717 ( .A(n_75), .Y(n_717) );
A2O1A1Ixp33_ASAP7_75t_L g448 ( .A1(n_76), .A2(n_449), .B(n_451), .C(n_455), .Y(n_448) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_77), .Y(n_129) );
NAND2xp5_ASAP7_75t_SL g155 ( .A(n_78), .B(n_156), .Y(n_155) );
CKINVDCx16_ASAP7_75t_R g547 ( .A(n_79), .Y(n_547) );
INVx1_ASAP7_75t_L g117 ( .A(n_80), .Y(n_117) );
NAND2xp5_ASAP7_75t_SL g498 ( .A(n_81), .B(n_484), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_82), .A2(n_105), .B1(n_118), .B2(n_724), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_84), .B(n_175), .Y(n_194) );
CKINVDCx20_ASAP7_75t_R g489 ( .A(n_85), .Y(n_489) );
NAND2xp5_ASAP7_75t_SL g163 ( .A(n_86), .B(n_156), .Y(n_163) );
INVx2_ASAP7_75t_L g144 ( .A(n_87), .Y(n_144) );
CKINVDCx20_ASAP7_75t_R g461 ( .A(n_88), .Y(n_461) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_89), .B(n_177), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_90), .B(n_156), .Y(n_249) );
INVx2_ASAP7_75t_L g114 ( .A(n_91), .Y(n_114) );
OR2x2_ASAP7_75t_L g125 ( .A(n_91), .B(n_126), .Y(n_125) );
AOI22xp33_ASAP7_75t_L g223 ( .A1(n_93), .A2(n_103), .B1(n_156), .B2(n_157), .Y(n_223) );
CKINVDCx20_ASAP7_75t_R g704 ( .A(n_94), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_95), .B(n_458), .Y(n_479) );
INVx1_ASAP7_75t_L g483 ( .A(n_96), .Y(n_483) );
INVxp67_ASAP7_75t_L g550 ( .A(n_97), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_98), .B(n_156), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_99), .B(n_117), .Y(n_116) );
INVx1_ASAP7_75t_L g452 ( .A(n_100), .Y(n_452) );
INVx1_ASAP7_75t_L g519 ( .A(n_101), .Y(n_519) );
AND2x2_ASAP7_75t_L g535 ( .A(n_102), .B(n_143), .Y(n_535) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_SL g724 ( .A(n_107), .Y(n_724) );
CKINVDCx9p33_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_109), .B(n_111), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_110), .Y(n_109) );
CKINVDCx14_ASAP7_75t_R g111 ( .A(n_112), .Y(n_111) );
NAND3xp33_ASAP7_75t_SL g112 ( .A(n_113), .B(n_114), .C(n_115), .Y(n_112) );
AND2x2_ASAP7_75t_L g127 ( .A(n_113), .B(n_128), .Y(n_127) );
AO22x2_ASAP7_75t_SL g132 ( .A1(n_114), .A2(n_133), .B1(n_441), .B2(n_700), .Y(n_132) );
INVx1_ASAP7_75t_L g700 ( .A(n_114), .Y(n_700) );
NOR2x2_ASAP7_75t_L g711 ( .A(n_114), .B(n_126), .Y(n_711) );
INVx1_ASAP7_75t_SL g115 ( .A(n_116), .Y(n_115) );
AOI22x1_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_130), .B1(n_712), .B2(n_713), .Y(n_118) );
NOR2xp33_ASAP7_75t_L g119 ( .A(n_120), .B(n_123), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx2_ASAP7_75t_SL g712 ( .A(n_121), .Y(n_712) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
AOI21xp5_ASAP7_75t_L g713 ( .A1(n_123), .A2(n_714), .B(n_723), .Y(n_713) );
NOR2xp33_ASAP7_75t_SL g123 ( .A(n_124), .B(n_129), .Y(n_123) );
HB1xp67_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
BUFx2_ASAP7_75t_L g723 ( .A(n_125), .Y(n_723) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
OAI22xp33_ASAP7_75t_SL g131 ( .A1(n_132), .A2(n_701), .B1(n_707), .B2(n_708), .Y(n_131) );
INVx1_ASAP7_75t_L g707 ( .A(n_132), .Y(n_707) );
INVx1_ASAP7_75t_L g440 ( .A(n_134), .Y(n_440) );
OAI22xp5_ASAP7_75t_SL g719 ( .A1(n_134), .A2(n_440), .B1(n_720), .B2(n_721), .Y(n_719) );
OR2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_360), .Y(n_134) );
NAND3xp33_ASAP7_75t_L g135 ( .A(n_136), .B(n_309), .C(n_351), .Y(n_135) );
AOI211xp5_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_214), .B(n_263), .C(n_285), .Y(n_136) );
OAI211xp5_ASAP7_75t_SL g137 ( .A1(n_138), .A2(n_169), .B(n_197), .C(n_209), .Y(n_137) );
INVxp67_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_139), .B(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g372 ( .A(n_139), .B(n_289), .Y(n_372) );
BUFx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
AND2x2_ASAP7_75t_L g274 ( .A(n_140), .B(n_200), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_140), .B(n_185), .Y(n_391) );
INVx1_ASAP7_75t_L g409 ( .A(n_140), .Y(n_409) );
AND2x2_ASAP7_75t_L g418 ( .A(n_140), .B(n_306), .Y(n_418) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
OR2x2_ASAP7_75t_L g301 ( .A(n_141), .B(n_185), .Y(n_301) );
AND2x2_ASAP7_75t_L g359 ( .A(n_141), .B(n_306), .Y(n_359) );
INVx1_ASAP7_75t_L g403 ( .A(n_141), .Y(n_403) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
OR2x2_ASAP7_75t_L g280 ( .A(n_142), .B(n_281), .Y(n_280) );
INVx2_ASAP7_75t_L g288 ( .A(n_142), .Y(n_288) );
HB1xp67_ASAP7_75t_L g328 ( .A(n_142), .Y(n_328) );
OA21x2_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_148), .B(n_168), .Y(n_142) );
INVx2_ASAP7_75t_L g179 ( .A(n_143), .Y(n_179) );
OA21x2_ASAP7_75t_L g185 ( .A1(n_143), .A2(n_186), .B(n_196), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_143), .A2(n_479), .B(n_480), .Y(n_478) );
INVx1_ASAP7_75t_L g502 ( .A(n_143), .Y(n_502) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_143), .A2(n_530), .B(n_531), .Y(n_529) );
AND2x2_ASAP7_75t_SL g143 ( .A(n_144), .B(n_145), .Y(n_143) );
AND2x2_ASAP7_75t_L g182 ( .A(n_144), .B(n_145), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_146), .B(n_147), .Y(n_145) );
OAI21xp5_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_161), .B(n_166), .Y(n_148) );
O2A1O1Ixp5_ASAP7_75t_SL g149 ( .A1(n_150), .A2(n_154), .B(n_155), .C(n_158), .Y(n_149) );
INVx3_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
HB1xp67_ASAP7_75t_L g454 ( .A(n_151), .Y(n_454) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g175 ( .A(n_152), .Y(n_175) );
BUFx3_ASAP7_75t_L g176 ( .A(n_152), .Y(n_176) );
AND2x6_ASAP7_75t_L g449 ( .A(n_152), .B(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx1_ASAP7_75t_L g157 ( .A(n_153), .Y(n_157) );
INVx1_ASAP7_75t_L g240 ( .A(n_153), .Y(n_240) );
INVx2_ASAP7_75t_L g234 ( .A(n_156), .Y(n_234) );
INVx3_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx2_ASAP7_75t_L g206 ( .A(n_158), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_158), .A2(n_248), .B(n_249), .Y(n_247) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_158), .A2(n_257), .B(n_258), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g549 ( .A(n_158), .B(n_550), .Y(n_549) );
INVx5_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
OAI22xp5_ASAP7_75t_SL g173 ( .A1(n_159), .A2(n_174), .B1(n_177), .B2(n_178), .Y(n_173) );
INVx3_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_160), .Y(n_165) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_160), .Y(n_177) );
INVx1_ASAP7_75t_L g191 ( .A(n_160), .Y(n_191) );
INVx1_ASAP7_75t_L g450 ( .A(n_160), .Y(n_450) );
AND2x2_ASAP7_75t_L g459 ( .A(n_160), .B(n_240), .Y(n_459) );
AOI21xp5_ASAP7_75t_L g161 ( .A1(n_162), .A2(n_163), .B(n_164), .Y(n_161) );
INVx1_ASAP7_75t_L g236 ( .A(n_164), .Y(n_236) );
INVx4_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx2_ASAP7_75t_L g485 ( .A(n_165), .Y(n_485) );
BUFx3_ASAP7_75t_L g180 ( .A(n_166), .Y(n_180) );
OAI21xp5_ASAP7_75t_L g186 ( .A1(n_166), .A2(n_187), .B(n_192), .Y(n_186) );
OAI21xp5_ASAP7_75t_L g231 ( .A1(n_166), .A2(n_232), .B(n_237), .Y(n_231) );
OAI21xp5_ASAP7_75t_L g246 ( .A1(n_166), .A2(n_247), .B(n_250), .Y(n_246) );
INVx4_ASAP7_75t_SL g456 ( .A(n_166), .Y(n_456) );
AND2x4_ASAP7_75t_L g458 ( .A(n_166), .B(n_459), .Y(n_458) );
NAND2x1p5_ASAP7_75t_L g520 ( .A(n_166), .B(n_459), .Y(n_520) );
INVxp67_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_171), .B(n_183), .Y(n_170) );
AND2x2_ASAP7_75t_L g267 ( .A(n_171), .B(n_268), .Y(n_267) );
INVx2_ASAP7_75t_L g300 ( .A(n_171), .Y(n_300) );
OR2x2_ASAP7_75t_L g426 ( .A(n_171), .B(n_427), .Y(n_426) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_171), .B(n_185), .Y(n_430) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx1_ASAP7_75t_L g200 ( .A(n_172), .Y(n_200) );
INVx1_ASAP7_75t_L g212 ( .A(n_172), .Y(n_212) );
AND2x2_ASAP7_75t_L g289 ( .A(n_172), .B(n_202), .Y(n_289) );
AND2x2_ASAP7_75t_L g329 ( .A(n_172), .B(n_203), .Y(n_329) );
INVx2_ASAP7_75t_L g472 ( .A(n_176), .Y(n_472) );
HB1xp67_ASAP7_75t_L g487 ( .A(n_176), .Y(n_487) );
INVx2_ASAP7_75t_L g195 ( .A(n_177), .Y(n_195) );
OAI22xp5_ASAP7_75t_L g204 ( .A1(n_177), .A2(n_205), .B1(n_206), .B2(n_207), .Y(n_204) );
OAI22xp5_ASAP7_75t_L g222 ( .A1(n_177), .A2(n_206), .B1(n_223), .B2(n_224), .Y(n_222) );
INVx4_ASAP7_75t_L g471 ( .A(n_177), .Y(n_471) );
INVx1_ASAP7_75t_L g499 ( .A(n_179), .Y(n_499) );
NAND3xp33_ASAP7_75t_L g221 ( .A(n_180), .B(n_222), .C(n_225), .Y(n_221) );
OAI21xp5_ASAP7_75t_L g255 ( .A1(n_180), .A2(n_256), .B(n_259), .Y(n_255) );
INVx4_ASAP7_75t_L g225 ( .A(n_181), .Y(n_225) );
OA21x2_ASAP7_75t_L g245 ( .A1(n_181), .A2(n_246), .B(n_253), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_181), .A2(n_509), .B(n_510), .Y(n_508) );
HB1xp67_ASAP7_75t_L g544 ( .A(n_181), .Y(n_544) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
INVx1_ASAP7_75t_L g208 ( .A(n_182), .Y(n_208) );
INVxp67_ASAP7_75t_L g371 ( .A(n_183), .Y(n_371) );
AND2x4_ASAP7_75t_L g396 ( .A(n_183), .B(n_289), .Y(n_396) );
BUFx3_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
AND2x2_ASAP7_75t_SL g287 ( .A(n_184), .B(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
AND2x2_ASAP7_75t_L g201 ( .A(n_185), .B(n_202), .Y(n_201) );
AND2x2_ASAP7_75t_L g275 ( .A(n_185), .B(n_203), .Y(n_275) );
INVx1_ASAP7_75t_L g281 ( .A(n_185), .Y(n_281) );
INVx2_ASAP7_75t_L g307 ( .A(n_185), .Y(n_307) );
AND2x2_ASAP7_75t_L g323 ( .A(n_185), .B(n_324), .Y(n_323) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_189), .B(n_190), .Y(n_187) );
INVx1_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_194), .B(n_195), .Y(n_192) );
O2A1O1Ixp5_ASAP7_75t_L g259 ( .A1(n_195), .A2(n_238), .B(n_260), .C(n_261), .Y(n_259) );
INVx1_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_198), .B(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g198 ( .A(n_199), .B(n_201), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
BUFx2_ASAP7_75t_L g278 ( .A(n_200), .Y(n_278) );
AND2x2_ASAP7_75t_L g386 ( .A(n_200), .B(n_202), .Y(n_386) );
AND2x2_ASAP7_75t_L g303 ( .A(n_201), .B(n_288), .Y(n_303) );
AND2x2_ASAP7_75t_L g402 ( .A(n_201), .B(n_403), .Y(n_402) );
NOR2xp67_ASAP7_75t_L g324 ( .A(n_202), .B(n_325), .Y(n_324) );
OR2x2_ASAP7_75t_L g427 ( .A(n_202), .B(n_288), .Y(n_427) );
INVx2_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
BUFx2_ASAP7_75t_L g213 ( .A(n_203), .Y(n_213) );
AND2x2_ASAP7_75t_L g306 ( .A(n_203), .B(n_307), .Y(n_306) );
O2A1O1Ixp33_ASAP7_75t_L g237 ( .A1(n_206), .A2(n_238), .B(n_241), .C(n_242), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_206), .A2(n_251), .B(n_252), .Y(n_250) );
INVx2_ASAP7_75t_L g230 ( .A(n_208), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_208), .B(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
AND2x2_ASAP7_75t_L g210 ( .A(n_211), .B(n_213), .Y(n_210) );
AND2x2_ASAP7_75t_L g352 ( .A(n_211), .B(n_287), .Y(n_352) );
HB1xp67_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_212), .B(n_288), .Y(n_337) );
INVx2_ASAP7_75t_L g336 ( .A(n_213), .Y(n_336) );
OAI222xp33_ASAP7_75t_L g340 ( .A1(n_213), .A2(n_280), .B1(n_341), .B2(n_343), .C1(n_344), .C2(n_347), .Y(n_340) );
INVx1_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_216), .B(n_226), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVx2_ASAP7_75t_L g265 ( .A(n_218), .Y(n_265) );
OR2x2_ASAP7_75t_L g376 ( .A(n_218), .B(n_377), .Y(n_376) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
INVx3_ASAP7_75t_L g298 ( .A(n_219), .Y(n_298) );
NOR2x1_ASAP7_75t_L g349 ( .A(n_219), .B(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g355 ( .A(n_219), .B(n_269), .Y(n_355) );
AND2x4_ASAP7_75t_L g219 ( .A(n_220), .B(n_221), .Y(n_219) );
INVx1_ASAP7_75t_L g316 ( .A(n_220), .Y(n_316) );
AO21x1_ASAP7_75t_L g315 ( .A1(n_222), .A2(n_225), .B(n_316), .Y(n_315) );
AO21x2_ASAP7_75t_L g446 ( .A1(n_225), .A2(n_447), .B(n_460), .Y(n_446) );
NOR2xp33_ASAP7_75t_L g460 ( .A(n_225), .B(n_461), .Y(n_460) );
INVx3_ASAP7_75t_L g463 ( .A(n_225), .Y(n_463) );
NOR2xp33_ASAP7_75t_L g488 ( .A(n_225), .B(n_489), .Y(n_488) );
AO21x2_ASAP7_75t_L g517 ( .A1(n_225), .A2(n_518), .B(n_525), .Y(n_517) );
AOI22xp5_ASAP7_75t_L g357 ( .A1(n_226), .A2(n_319), .B1(n_358), .B2(n_359), .Y(n_357) );
AND2x2_ASAP7_75t_L g226 ( .A(n_227), .B(n_244), .Y(n_226) );
INVx3_ASAP7_75t_L g291 ( .A(n_227), .Y(n_291) );
OR2x2_ASAP7_75t_L g424 ( .A(n_227), .B(n_300), .Y(n_424) );
INVx2_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
AND2x2_ASAP7_75t_L g297 ( .A(n_228), .B(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g313 ( .A(n_228), .B(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g321 ( .A(n_228), .B(n_269), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_228), .B(n_245), .Y(n_377) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
AND2x2_ASAP7_75t_L g268 ( .A(n_229), .B(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g272 ( .A(n_229), .B(n_245), .Y(n_272) );
AND2x2_ASAP7_75t_L g348 ( .A(n_229), .B(n_295), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_229), .B(n_254), .Y(n_388) );
OA21x2_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_231), .B(n_243), .Y(n_229) );
OA21x2_ASAP7_75t_L g254 ( .A1(n_230), .A2(n_255), .B(n_262), .Y(n_254) );
O2A1O1Ixp33_ASAP7_75t_L g232 ( .A1(n_233), .A2(n_234), .B(n_235), .C(n_236), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_234), .A2(n_512), .B(n_513), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_234), .A2(n_523), .B(n_524), .Y(n_522) );
O2A1O1Ixp33_ASAP7_75t_L g451 ( .A1(n_236), .A2(n_452), .B(n_453), .C(n_454), .Y(n_451) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_238), .A2(n_497), .B(n_498), .Y(n_496) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_244), .B(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g304 ( .A(n_244), .B(n_265), .Y(n_304) );
AND2x2_ASAP7_75t_L g308 ( .A(n_244), .B(n_298), .Y(n_308) );
AND2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_254), .Y(n_244) );
INVx3_ASAP7_75t_L g269 ( .A(n_245), .Y(n_269) );
AND2x2_ASAP7_75t_L g294 ( .A(n_245), .B(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g429 ( .A(n_245), .B(n_412), .Y(n_429) );
HB1xp67_ASAP7_75t_L g283 ( .A(n_254), .Y(n_283) );
INVx2_ASAP7_75t_L g295 ( .A(n_254), .Y(n_295) );
AND2x2_ASAP7_75t_L g339 ( .A(n_254), .B(n_315), .Y(n_339) );
INVx1_ASAP7_75t_L g382 ( .A(n_254), .Y(n_382) );
OR2x2_ASAP7_75t_L g413 ( .A(n_254), .B(n_315), .Y(n_413) );
AND2x2_ASAP7_75t_L g433 ( .A(n_254), .B(n_269), .Y(n_433) );
OAI21xp5_ASAP7_75t_L g263 ( .A1(n_264), .A2(n_266), .B(n_270), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
AND2x2_ASAP7_75t_L g271 ( .A(n_265), .B(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_265), .B(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g390 ( .A(n_267), .Y(n_390) );
INVx2_ASAP7_75t_SL g284 ( .A(n_268), .Y(n_284) );
AND2x2_ASAP7_75t_L g404 ( .A(n_268), .B(n_298), .Y(n_404) );
INVx2_ASAP7_75t_L g350 ( .A(n_269), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_269), .B(n_382), .Y(n_381) );
AOI22xp5_ASAP7_75t_L g270 ( .A1(n_271), .A2(n_273), .B1(n_276), .B2(n_282), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_272), .B(n_417), .Y(n_416) );
INVx1_ASAP7_75t_SL g438 ( .A(n_272), .Y(n_438) );
AND2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
INVx1_ASAP7_75t_L g363 ( .A(n_274), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_274), .B(n_306), .Y(n_375) );
NOR2xp33_ASAP7_75t_L g362 ( .A(n_275), .B(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g379 ( .A(n_275), .B(n_328), .Y(n_379) );
INVx2_ASAP7_75t_L g435 ( .A(n_275), .Y(n_435) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
AND2x2_ASAP7_75t_L g305 ( .A(n_278), .B(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_278), .B(n_323), .Y(n_356) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
NOR2xp33_ASAP7_75t_L g358 ( .A(n_280), .B(n_300), .Y(n_358) );
NOR2xp33_ASAP7_75t_L g282 ( .A(n_283), .B(n_284), .Y(n_282) );
INVx1_ASAP7_75t_L g417 ( .A(n_283), .Y(n_417) );
O2A1O1Ixp33_ASAP7_75t_SL g367 ( .A1(n_284), .A2(n_368), .B(n_370), .C(n_373), .Y(n_367) );
OR2x2_ASAP7_75t_L g394 ( .A(n_284), .B(n_298), .Y(n_394) );
OAI221xp5_ASAP7_75t_SL g285 ( .A1(n_286), .A2(n_290), .B1(n_292), .B2(n_299), .C(n_302), .Y(n_285) );
NAND2xp5_ASAP7_75t_SL g286 ( .A(n_287), .B(n_289), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_287), .B(n_336), .Y(n_343) );
AND2x2_ASAP7_75t_L g385 ( .A(n_287), .B(n_386), .Y(n_385) );
INVx2_ASAP7_75t_L g421 ( .A(n_287), .Y(n_421) );
HB1xp67_ASAP7_75t_L g312 ( .A(n_288), .Y(n_312) );
INVx1_ASAP7_75t_L g325 ( .A(n_288), .Y(n_325) );
NOR2xp67_ASAP7_75t_L g345 ( .A(n_291), .B(n_346), .Y(n_345) );
INVxp67_ASAP7_75t_L g399 ( .A(n_291), .Y(n_399) );
NAND2xp5_ASAP7_75t_SL g415 ( .A(n_291), .B(n_339), .Y(n_415) );
INVx2_ASAP7_75t_L g401 ( .A(n_292), .Y(n_401) );
OR2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_296), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g342 ( .A(n_294), .B(n_313), .Y(n_342) );
O2A1O1Ixp33_ASAP7_75t_L g351 ( .A1(n_294), .A2(n_310), .B(n_352), .C(n_353), .Y(n_351) );
AND2x2_ASAP7_75t_L g320 ( .A(n_295), .B(n_315), .Y(n_320) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
NOR2xp33_ASAP7_75t_L g397 ( .A(n_299), .B(n_398), .Y(n_397) );
OR2x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
OR2x2_ASAP7_75t_L g368 ( .A(n_300), .B(n_369), .Y(n_368) );
AOI22xp5_ASAP7_75t_L g302 ( .A1(n_303), .A2(n_304), .B1(n_305), .B2(n_308), .Y(n_302) );
INVx1_ASAP7_75t_L g422 ( .A(n_304), .Y(n_422) );
INVx1_ASAP7_75t_L g369 ( .A(n_306), .Y(n_369) );
INVx1_ASAP7_75t_L g420 ( .A(n_308), .Y(n_420) );
AOI211xp5_ASAP7_75t_SL g309 ( .A1(n_310), .A2(n_313), .B(n_317), .C(n_340), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
OR2x2_ASAP7_75t_L g332 ( .A(n_312), .B(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g383 ( .A(n_313), .Y(n_383) );
AND2x2_ASAP7_75t_L g432 ( .A(n_313), .B(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
OAI21xp33_ASAP7_75t_L g317 ( .A1(n_318), .A2(n_322), .B(n_330), .Y(n_317) );
INVx1_ASAP7_75t_SL g318 ( .A(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
INVx2_ASAP7_75t_L g346 ( .A(n_320), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_320), .B(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g338 ( .A(n_321), .B(n_339), .Y(n_338) );
INVx2_ASAP7_75t_L g414 ( .A(n_321), .Y(n_414) );
OAI32xp33_ASAP7_75t_L g425 ( .A1(n_321), .A2(n_373), .A3(n_380), .B1(n_421), .B2(n_426), .Y(n_425) );
NOR2xp33_ASAP7_75t_SL g322 ( .A(n_323), .B(n_326), .Y(n_322) );
INVx1_ASAP7_75t_SL g393 ( .A(n_323), .Y(n_393) );
AND2x2_ASAP7_75t_L g326 ( .A(n_327), .B(n_329), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx1_ASAP7_75t_SL g333 ( .A(n_329), .Y(n_333) );
OAI21xp33_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_334), .B(n_338), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
OAI22xp33_ASAP7_75t_L g405 ( .A1(n_332), .A2(n_380), .B1(n_406), .B2(n_408), .Y(n_405) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
OR2x2_ASAP7_75t_L g335 ( .A(n_336), .B(n_337), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_336), .B(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g373 ( .A(n_339), .Y(n_373) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
NAND2x1p5_ASAP7_75t_L g347 ( .A(n_348), .B(n_349), .Y(n_347) );
INVx1_ASAP7_75t_L g366 ( .A(n_350), .Y(n_366) );
OAI21xp5_ASAP7_75t_L g353 ( .A1(n_354), .A2(n_356), .B(n_357), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
AOI221xp5_ASAP7_75t_L g400 ( .A1(n_359), .A2(n_401), .B1(n_402), .B2(n_404), .C(n_405), .Y(n_400) );
NAND5xp2_ASAP7_75t_L g360 ( .A(n_361), .B(n_384), .C(n_400), .D(n_410), .E(n_428), .Y(n_360) );
AOI211xp5_ASAP7_75t_SL g361 ( .A1(n_362), .A2(n_364), .B(n_367), .C(n_374), .Y(n_361) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g431 ( .A(n_368), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_371), .B(n_372), .Y(n_370) );
OAI22xp33_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_376), .B1(n_378), .B2(n_380), .Y(n_374) );
INVx1_ASAP7_75t_SL g407 ( .A(n_377), .Y(n_407) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
OAI322xp33_ASAP7_75t_L g389 ( .A1(n_380), .A2(n_390), .A3(n_391), .B1(n_392), .B2(n_393), .C1(n_394), .C2(n_395), .Y(n_389) );
OR2x2_ASAP7_75t_L g380 ( .A(n_381), .B(n_383), .Y(n_380) );
INVx1_ASAP7_75t_L g392 ( .A(n_382), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_382), .B(n_407), .Y(n_406) );
AOI211xp5_ASAP7_75t_SL g384 ( .A1(n_385), .A2(n_387), .B(n_389), .C(n_397), .Y(n_384) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
OAI22xp33_ASAP7_75t_L g419 ( .A1(n_393), .A2(n_420), .B1(n_421), .B2(n_422), .Y(n_419) );
INVx1_ASAP7_75t_SL g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g436 ( .A(n_403), .Y(n_436) );
AOI221xp5_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_418), .B1(n_419), .B2(n_423), .C(n_425), .Y(n_410) );
OAI211xp5_ASAP7_75t_SL g411 ( .A1(n_412), .A2(n_414), .B(n_415), .C(n_416), .Y(n_411) );
INVx1_ASAP7_75t_SL g412 ( .A(n_413), .Y(n_412) );
OR2x2_ASAP7_75t_L g437 ( .A(n_413), .B(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
AOI221xp5_ASAP7_75t_L g428 ( .A1(n_429), .A2(n_430), .B1(n_431), .B2(n_432), .C(n_434), .Y(n_428) );
AOI21xp33_ASAP7_75t_SL g434 ( .A1(n_435), .A2(n_436), .B(n_437), .Y(n_434) );
NAND2x1p5_ASAP7_75t_L g441 ( .A(n_442), .B(n_643), .Y(n_441) );
AND4x1_ASAP7_75t_L g442 ( .A(n_443), .B(n_583), .C(n_598), .D(n_623), .Y(n_442) );
NOR2xp33_ASAP7_75t_SL g443 ( .A(n_444), .B(n_556), .Y(n_443) );
OAI21xp33_ASAP7_75t_L g444 ( .A1(n_445), .A2(n_474), .B(n_536), .Y(n_444) );
AND2x2_ASAP7_75t_L g586 ( .A(n_445), .B(n_491), .Y(n_586) );
AND2x2_ASAP7_75t_L g599 ( .A(n_445), .B(n_490), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_445), .B(n_475), .Y(n_649) );
INVx1_ASAP7_75t_L g653 ( .A(n_445), .Y(n_653) );
AND2x2_ASAP7_75t_L g445 ( .A(n_446), .B(n_462), .Y(n_445) );
INVx2_ASAP7_75t_L g570 ( .A(n_446), .Y(n_570) );
BUFx2_ASAP7_75t_L g597 ( .A(n_446), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_448), .B(n_457), .Y(n_447) );
INVx5_ASAP7_75t_L g467 ( .A(n_449), .Y(n_467) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
O2A1O1Ixp33_ASAP7_75t_SL g465 ( .A1(n_456), .A2(n_466), .B(n_467), .C(n_468), .Y(n_465) );
O2A1O1Ixp33_ASAP7_75t_L g546 ( .A1(n_456), .A2(n_467), .B(n_547), .C(n_548), .Y(n_546) );
BUFx2_ASAP7_75t_L g494 ( .A(n_458), .Y(n_494) );
AND2x2_ASAP7_75t_L g537 ( .A(n_462), .B(n_491), .Y(n_537) );
INVx2_ASAP7_75t_L g553 ( .A(n_462), .Y(n_553) );
AND2x2_ASAP7_75t_L g562 ( .A(n_462), .B(n_490), .Y(n_562) );
AND2x2_ASAP7_75t_L g641 ( .A(n_462), .B(n_570), .Y(n_641) );
OA21x2_ASAP7_75t_L g462 ( .A1(n_463), .A2(n_464), .B(n_473), .Y(n_462) );
INVx2_ASAP7_75t_L g481 ( .A(n_467), .Y(n_481) );
NOR2xp33_ASAP7_75t_L g469 ( .A(n_470), .B(n_471), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_475), .B(n_503), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_475), .B(n_568), .Y(n_606) );
INVx1_ASAP7_75t_L g694 ( .A(n_475), .Y(n_694) );
AND2x2_ASAP7_75t_L g475 ( .A(n_476), .B(n_490), .Y(n_475) );
AND2x2_ASAP7_75t_L g552 ( .A(n_476), .B(n_553), .Y(n_552) );
OR2x2_ASAP7_75t_L g566 ( .A(n_476), .B(n_567), .Y(n_566) );
HB1xp67_ASAP7_75t_L g595 ( .A(n_476), .Y(n_595) );
OR2x2_ASAP7_75t_L g627 ( .A(n_476), .B(n_569), .Y(n_627) );
AND2x2_ASAP7_75t_L g635 ( .A(n_476), .B(n_636), .Y(n_635) );
AND2x2_ASAP7_75t_L g668 ( .A(n_476), .B(n_637), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_476), .B(n_537), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_476), .B(n_597), .Y(n_693) );
AND2x2_ASAP7_75t_L g699 ( .A(n_476), .B(n_586), .Y(n_699) );
INVx5_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
BUFx2_ASAP7_75t_L g559 ( .A(n_477), .Y(n_559) );
AND2x2_ASAP7_75t_L g589 ( .A(n_477), .B(n_569), .Y(n_589) );
AND2x2_ASAP7_75t_L g622 ( .A(n_477), .B(n_582), .Y(n_622) );
AND2x2_ASAP7_75t_L g642 ( .A(n_477), .B(n_491), .Y(n_642) );
AND2x2_ASAP7_75t_L g676 ( .A(n_477), .B(n_542), .Y(n_676) );
OR2x6_ASAP7_75t_L g477 ( .A(n_478), .B(n_488), .Y(n_477) );
O2A1O1Ixp33_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_484), .B(n_486), .C(n_487), .Y(n_482) );
O2A1O1Ixp33_ASAP7_75t_L g532 ( .A1(n_484), .A2(n_487), .B(n_533), .C(n_534), .Y(n_532) );
INVx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
AND2x4_ASAP7_75t_L g582 ( .A(n_490), .B(n_553), .Y(n_582) );
AND2x2_ASAP7_75t_L g593 ( .A(n_490), .B(n_589), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_490), .B(n_569), .Y(n_632) );
INVx2_ASAP7_75t_L g647 ( .A(n_490), .Y(n_647) );
NOR2xp33_ASAP7_75t_L g670 ( .A(n_490), .B(n_581), .Y(n_670) );
AND2x2_ASAP7_75t_L g689 ( .A(n_490), .B(n_641), .Y(n_689) );
INVx5_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
HB1xp67_ASAP7_75t_L g588 ( .A(n_491), .Y(n_588) );
AND2x2_ASAP7_75t_L g596 ( .A(n_491), .B(n_597), .Y(n_596) );
AND2x4_ASAP7_75t_L g637 ( .A(n_491), .B(n_553), .Y(n_637) );
OR2x6_ASAP7_75t_L g491 ( .A(n_492), .B(n_500), .Y(n_491) );
AOI21xp5_ASAP7_75t_SL g492 ( .A1(n_493), .A2(n_495), .B(n_499), .Y(n_492) );
NOR2xp33_ASAP7_75t_L g500 ( .A(n_501), .B(n_502), .Y(n_500) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_505), .B(n_514), .Y(n_504) );
AND2x2_ASAP7_75t_L g560 ( .A(n_505), .B(n_543), .Y(n_560) );
INVx1_ASAP7_75t_SL g505 ( .A(n_506), .Y(n_505) );
NAND2xp5_ASAP7_75t_SL g540 ( .A(n_506), .B(n_517), .Y(n_540) );
OR2x2_ASAP7_75t_L g573 ( .A(n_506), .B(n_543), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_506), .B(n_543), .Y(n_578) );
AND2x2_ASAP7_75t_L g605 ( .A(n_506), .B(n_542), .Y(n_605) );
AND2x2_ASAP7_75t_L g657 ( .A(n_506), .B(n_516), .Y(n_657) );
INVx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_507), .B(n_527), .Y(n_565) );
AND2x2_ASAP7_75t_L g601 ( .A(n_507), .B(n_517), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_514), .B(n_665), .Y(n_664) );
INVx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
OR2x2_ASAP7_75t_L g591 ( .A(n_515), .B(n_573), .Y(n_591) );
OR2x2_ASAP7_75t_L g515 ( .A(n_516), .B(n_527), .Y(n_515) );
OAI322xp33_ASAP7_75t_L g556 ( .A1(n_516), .A2(n_557), .A3(n_561), .B1(n_563), .B2(n_566), .C1(n_571), .C2(n_579), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_516), .B(n_542), .Y(n_564) );
OR2x2_ASAP7_75t_L g574 ( .A(n_516), .B(n_528), .Y(n_574) );
AND2x2_ASAP7_75t_L g576 ( .A(n_516), .B(n_528), .Y(n_576) );
NOR2xp33_ASAP7_75t_L g577 ( .A(n_516), .B(n_578), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_516), .B(n_543), .Y(n_638) );
NOR2xp33_ASAP7_75t_L g671 ( .A(n_516), .B(n_672), .Y(n_671) );
INVx5_ASAP7_75t_SL g516 ( .A(n_517), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_517), .B(n_560), .Y(n_686) );
OAI21xp5_ASAP7_75t_L g518 ( .A1(n_519), .A2(n_520), .B(n_521), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_527), .B(n_542), .Y(n_541) );
AND2x2_ASAP7_75t_L g554 ( .A(n_527), .B(n_555), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_527), .B(n_605), .Y(n_604) );
OR2x2_ASAP7_75t_L g616 ( .A(n_527), .B(n_543), .Y(n_616) );
AOI211xp5_ASAP7_75t_SL g644 ( .A1(n_527), .A2(n_645), .B(n_648), .C(n_660), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_527), .B(n_651), .Y(n_650) );
AND2x2_ASAP7_75t_L g682 ( .A(n_527), .B(n_657), .Y(n_682) );
INVx5_ASAP7_75t_SL g527 ( .A(n_528), .Y(n_527) );
AND2x2_ASAP7_75t_L g610 ( .A(n_528), .B(n_543), .Y(n_610) );
HB1xp67_ASAP7_75t_L g619 ( .A(n_528), .Y(n_619) );
AND2x2_ASAP7_75t_L g659 ( .A(n_528), .B(n_657), .Y(n_659) );
AND2x2_ASAP7_75t_SL g690 ( .A(n_528), .B(n_560), .Y(n_690) );
AND2x2_ASAP7_75t_L g697 ( .A(n_528), .B(n_656), .Y(n_697) );
OR2x6_ASAP7_75t_L g528 ( .A(n_529), .B(n_535), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_537), .A2(n_538), .B1(n_552), .B2(n_554), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_537), .B(n_559), .Y(n_607) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
OR2x2_ASAP7_75t_L g539 ( .A(n_540), .B(n_541), .Y(n_539) );
INVx1_ASAP7_75t_L g555 ( .A(n_540), .Y(n_555) );
OR2x2_ASAP7_75t_L g615 ( .A(n_540), .B(n_616), .Y(n_615) );
OAI221xp5_ASAP7_75t_SL g663 ( .A1(n_540), .A2(n_664), .B1(n_666), .B2(n_667), .C(n_669), .Y(n_663) );
INVx2_ASAP7_75t_L g602 ( .A(n_541), .Y(n_602) );
AND2x2_ASAP7_75t_L g575 ( .A(n_542), .B(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g665 ( .A(n_542), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_542), .B(n_657), .Y(n_678) );
INVx3_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVxp67_ASAP7_75t_L g620 ( .A(n_543), .Y(n_620) );
AND2x2_ASAP7_75t_L g656 ( .A(n_543), .B(n_657), .Y(n_656) );
OA21x2_ASAP7_75t_L g543 ( .A1(n_544), .A2(n_545), .B(n_551), .Y(n_543) );
AND2x2_ASAP7_75t_L g658 ( .A(n_552), .B(n_597), .Y(n_658) );
AND2x2_ASAP7_75t_L g568 ( .A(n_553), .B(n_569), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_553), .B(n_626), .Y(n_625) );
NOR2xp33_ASAP7_75t_SL g639 ( .A(n_555), .B(n_602), .Y(n_639) );
INVx1_ASAP7_75t_SL g557 ( .A(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_L g645 ( .A(n_558), .B(n_646), .Y(n_645) );
AND2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_560), .Y(n_558) );
OR2x2_ASAP7_75t_L g631 ( .A(n_559), .B(n_632), .Y(n_631) );
AND2x2_ASAP7_75t_L g696 ( .A(n_559), .B(n_641), .Y(n_696) );
INVx2_ASAP7_75t_L g629 ( .A(n_560), .Y(n_629) );
NAND4xp25_ASAP7_75t_SL g692 ( .A(n_561), .B(n_693), .C(n_694), .D(n_695), .Y(n_692) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_562), .B(n_626), .Y(n_661) );
OR2x2_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
INVx1_ASAP7_75t_SL g698 ( .A(n_565), .Y(n_698) );
O2A1O1Ixp33_ASAP7_75t_SL g660 ( .A1(n_566), .A2(n_629), .B(n_633), .C(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g655 ( .A(n_568), .B(n_647), .Y(n_655) );
HB1xp67_ASAP7_75t_L g581 ( .A(n_569), .Y(n_581) );
INVx1_ASAP7_75t_L g636 ( .A(n_569), .Y(n_636) );
INVx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
HB1xp67_ASAP7_75t_L g613 ( .A(n_570), .Y(n_613) );
AOI211xp5_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_574), .B(n_575), .C(n_577), .Y(n_571) );
AND2x2_ASAP7_75t_L g592 ( .A(n_572), .B(n_576), .Y(n_592) );
OAI322xp33_ASAP7_75t_SL g630 ( .A1(n_572), .A2(n_631), .A3(n_633), .B1(n_634), .B2(n_638), .C1(n_639), .C2(n_640), .Y(n_630) );
INVx1_ASAP7_75t_SL g572 ( .A(n_573), .Y(n_572) );
OR2x2_ASAP7_75t_L g652 ( .A(n_574), .B(n_578), .Y(n_652) );
INVx1_ASAP7_75t_L g633 ( .A(n_576), .Y(n_633) );
INVx1_ASAP7_75t_SL g651 ( .A(n_578), .Y(n_651) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_581), .B(n_582), .Y(n_580) );
AOI222xp33_ASAP7_75t_L g583 ( .A1(n_584), .A2(n_590), .B1(n_592), .B2(n_593), .C1(n_594), .C2(n_726), .Y(n_583) );
NAND2xp5_ASAP7_75t_SL g584 ( .A(n_585), .B(n_587), .Y(n_584) );
OAI322xp33_ASAP7_75t_L g673 ( .A1(n_585), .A2(n_647), .A3(n_652), .B1(n_674), .B2(n_675), .C1(n_677), .C2(n_678), .Y(n_673) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
AOI221xp5_ASAP7_75t_L g623 ( .A1(n_586), .A2(n_600), .B1(n_624), .B2(n_628), .C(n_630), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_588), .B(n_589), .Y(n_587) );
INVx1_ASAP7_75t_SL g590 ( .A(n_591), .Y(n_590) );
OAI222xp33_ASAP7_75t_L g603 ( .A1(n_591), .A2(n_604), .B1(n_606), .B2(n_607), .C1(n_608), .C2(n_611), .Y(n_603) );
AOI22xp5_ASAP7_75t_L g669 ( .A1(n_593), .A2(n_600), .B1(n_670), .B2(n_671), .Y(n_669) );
AND2x2_ASAP7_75t_L g594 ( .A(n_595), .B(n_596), .Y(n_594) );
AOI211xp5_ASAP7_75t_L g598 ( .A1(n_599), .A2(n_600), .B(n_603), .C(n_614), .Y(n_598) );
O2A1O1Ixp33_ASAP7_75t_L g679 ( .A1(n_600), .A2(n_637), .B(n_680), .C(n_683), .Y(n_679) );
AND2x4_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
AND2x2_ASAP7_75t_L g609 ( .A(n_601), .B(n_610), .Y(n_609) );
INVx1_ASAP7_75t_SL g672 ( .A(n_605), .Y(n_672) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_612), .B(n_637), .Y(n_666) );
BUFx2_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
AOI21xp33_ASAP7_75t_L g614 ( .A1(n_615), .A2(n_617), .B(n_621), .Y(n_614) );
OAI221xp5_ASAP7_75t_SL g683 ( .A1(n_615), .A2(n_684), .B1(n_685), .B2(n_686), .C(n_687), .Y(n_683) );
INVxp33_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
NOR2xp33_ASAP7_75t_L g618 ( .A(n_619), .B(n_620), .Y(n_618) );
NOR2xp33_ASAP7_75t_L g628 ( .A(n_619), .B(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_626), .B(n_637), .Y(n_677) );
INVx2_ASAP7_75t_SL g626 ( .A(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_635), .B(n_637), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_641), .B(n_642), .Y(n_640) );
AND2x2_ASAP7_75t_L g688 ( .A(n_641), .B(n_647), .Y(n_688) );
AND4x1_ASAP7_75t_L g643 ( .A(n_644), .B(n_662), .C(n_679), .D(n_691), .Y(n_643) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
OAI221xp5_ASAP7_75t_SL g648 ( .A1(n_649), .A2(n_650), .B1(n_652), .B2(n_653), .C(n_654), .Y(n_648) );
AOI22xp5_ASAP7_75t_L g654 ( .A1(n_655), .A2(n_656), .B1(n_658), .B2(n_659), .Y(n_654) );
INVx1_ASAP7_75t_L g684 ( .A(n_655), .Y(n_684) );
INVx1_ASAP7_75t_SL g674 ( .A(n_659), .Y(n_674) );
NOR2xp33_ASAP7_75t_SL g662 ( .A(n_663), .B(n_673), .Y(n_662) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
NOR2xp33_ASAP7_75t_L g680 ( .A(n_675), .B(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_682), .A2(n_688), .B1(n_689), .B2(n_690), .Y(n_687) );
AOI22xp5_ASAP7_75t_L g691 ( .A1(n_692), .A2(n_697), .B1(n_698), .B2(n_699), .Y(n_691) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g708 ( .A(n_701), .Y(n_708) );
CKINVDCx20_ASAP7_75t_R g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_SL g709 ( .A(n_710), .Y(n_709) );
INVx3_ASAP7_75t_SL g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
XNOR2xp5_ASAP7_75t_SL g715 ( .A(n_716), .B(n_719), .Y(n_715) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
endmodule