module real_aes_3257_n_234 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_913, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_38, n_155, n_118, n_143, n_139, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_234);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_913;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_234;
wire n_480;
wire n_476;
wire n_758;
wire n_887;
wire n_436;
wire n_599;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_285;
wire n_624;
wire n_618;
wire n_800;
wire n_778;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_852;
wire n_766;
wire n_857;
wire n_461;
wire n_242;
wire n_908;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_767;
wire n_889;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_763;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_415;
wire n_572;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_356;
wire n_478;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_352;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_746;
wire n_284;
wire n_656;
wire n_316;
wire n_532;
wire n_755;
wire n_409;
wire n_781;
wire n_748;
wire n_909;
wire n_298;
wire n_523;
wire n_860;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_874;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_671;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_903;
wire n_454;
wire n_812;
wire n_817;
wire n_565;
wire n_443;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_879;
wire n_331;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_807;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_632;
wire n_246;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_898;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_756;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_907;
wire n_847;
wire n_779;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_831;
wire n_290;
wire n_653;
wire n_899;
wire n_526;
wire n_365;
wire n_637;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_472;
wire n_866;
wire n_452;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_623;
wire n_249;
wire n_446;
wire n_721;
wire n_681;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_266;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_686;
wire n_279;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_911;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_668;
wire n_237;
wire n_797;
wire n_862;
AOI22xp5_ASAP7_75t_L g570 ( .A1(n_0), .A2(n_198), .B1(n_571), .B2(n_573), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_1), .A2(n_96), .B1(n_528), .B2(n_530), .Y(n_527) );
HB1xp67_ASAP7_75t_L g246 ( .A(n_2), .Y(n_246) );
AND2x4_ASAP7_75t_L g671 ( .A(n_2), .B(n_227), .Y(n_671) );
AND2x4_ASAP7_75t_L g676 ( .A(n_2), .B(n_677), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_3), .A2(n_194), .B1(n_485), .B2(n_522), .Y(n_521) );
AO22x1_ASAP7_75t_L g709 ( .A1(n_4), .A2(n_5), .B1(n_672), .B2(n_682), .Y(n_709) );
AOI22xp33_ASAP7_75t_L g674 ( .A1(n_6), .A2(n_176), .B1(n_675), .B2(n_678), .Y(n_674) );
INVx1_ASAP7_75t_L g341 ( .A(n_7), .Y(n_341) );
AOI22xp33_ASAP7_75t_L g539 ( .A1(n_8), .A2(n_57), .B1(n_321), .B2(n_507), .Y(n_539) );
AOI22xp5_ASAP7_75t_L g642 ( .A1(n_9), .A2(n_35), .B1(n_562), .B2(n_643), .Y(n_642) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_10), .A2(n_206), .B1(n_324), .B2(n_502), .Y(n_501) );
AOI22xp33_ASAP7_75t_L g492 ( .A1(n_11), .A2(n_56), .B1(n_493), .B2(n_494), .Y(n_492) );
AOI21xp33_ASAP7_75t_L g433 ( .A1(n_12), .A2(n_434), .B(n_435), .Y(n_433) );
AOI22xp33_ASAP7_75t_L g441 ( .A1(n_13), .A2(n_164), .B1(n_384), .B2(n_390), .Y(n_441) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_14), .A2(n_108), .B1(n_260), .B2(n_526), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_15), .A2(n_20), .B1(n_612), .B2(n_613), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_16), .A2(n_209), .B1(n_453), .B2(n_454), .Y(n_647) );
AOI22xp33_ASAP7_75t_L g410 ( .A1(n_17), .A2(n_231), .B1(n_386), .B2(n_387), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_18), .A2(n_139), .B1(n_392), .B2(n_393), .Y(n_584) );
AOI22xp33_ASAP7_75t_L g645 ( .A1(n_19), .A2(n_128), .B1(n_331), .B2(n_646), .Y(n_645) );
AOI22xp33_ASAP7_75t_L g484 ( .A1(n_21), .A2(n_49), .B1(n_300), .B2(n_485), .Y(n_484) );
AOI22xp5_ASAP7_75t_L g706 ( .A1(n_22), .A2(n_107), .B1(n_699), .B2(n_707), .Y(n_706) );
XNOR2x1_ASAP7_75t_L g543 ( .A(n_23), .B(n_544), .Y(n_543) );
AOI22xp33_ASAP7_75t_SL g568 ( .A1(n_24), .A2(n_186), .B1(n_304), .B2(n_569), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_25), .B(n_505), .Y(n_504) );
AOI22xp5_ASAP7_75t_L g888 ( .A1(n_26), .A2(n_123), .B1(n_260), .B2(n_889), .Y(n_888) );
AOI22xp33_ASAP7_75t_L g388 ( .A1(n_27), .A2(n_70), .B1(n_389), .B2(n_390), .Y(n_388) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_28), .A2(n_230), .B1(n_498), .B2(n_500), .Y(n_497) );
INVx1_ASAP7_75t_L g553 ( .A(n_29), .Y(n_553) );
AOI221xp5_ASAP7_75t_L g532 ( .A1(n_30), .A2(n_47), .B1(n_451), .B2(n_533), .C(n_535), .Y(n_532) );
AOI22xp5_ASAP7_75t_L g875 ( .A1(n_31), .A2(n_66), .B1(n_457), .B2(n_876), .Y(n_875) );
INVx1_ASAP7_75t_L g422 ( .A(n_32), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g487 ( .A1(n_33), .A2(n_177), .B1(n_311), .B2(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g536 ( .A(n_34), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_36), .B(n_183), .Y(n_244) );
INVx1_ASAP7_75t_L g282 ( .A(n_36), .Y(n_282) );
INVxp67_ASAP7_75t_L g352 ( .A(n_36), .Y(n_352) );
OA22x2_ASAP7_75t_L g580 ( .A1(n_37), .A2(n_581), .B1(n_592), .B2(n_593), .Y(n_580) );
INVx1_ASAP7_75t_L g593 ( .A(n_37), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g881 ( .A1(n_38), .A2(n_117), .B1(n_507), .B2(n_549), .Y(n_881) );
AOI22xp33_ASAP7_75t_L g421 ( .A1(n_39), .A2(n_126), .B1(n_371), .B2(n_376), .Y(n_421) );
AOI22xp33_ASAP7_75t_L g439 ( .A1(n_40), .A2(n_51), .B1(n_392), .B2(n_393), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_41), .B(n_555), .Y(n_644) );
INVx1_ASAP7_75t_L g378 ( .A(n_42), .Y(n_378) );
NAND2xp5_ASAP7_75t_SL g277 ( .A(n_43), .B(n_266), .Y(n_277) );
INVx1_ASAP7_75t_L g560 ( .A(n_44), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g303 ( .A1(n_45), .A2(n_146), .B1(n_304), .B2(n_307), .Y(n_303) );
AOI22xp33_ASAP7_75t_L g295 ( .A1(n_46), .A2(n_69), .B1(n_296), .B2(n_300), .Y(n_295) );
AOI22xp33_ASAP7_75t_L g452 ( .A1(n_48), .A2(n_226), .B1(n_453), .B2(n_454), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_50), .A2(n_199), .B1(n_260), .B2(n_485), .Y(n_650) );
AOI22xp33_ASAP7_75t_SL g372 ( .A1(n_52), .A2(n_187), .B1(n_373), .B2(n_374), .Y(n_372) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_53), .A2(n_191), .B1(n_606), .B2(n_607), .Y(n_605) );
AOI22xp5_ASAP7_75t_L g692 ( .A1(n_54), .A2(n_154), .B1(n_668), .B2(n_672), .Y(n_692) );
AOI21xp33_ASAP7_75t_L g375 ( .A1(n_55), .A2(n_376), .B(n_377), .Y(n_375) );
AOI22xp33_ASAP7_75t_SL g575 ( .A1(n_58), .A2(n_219), .B1(n_493), .B2(n_576), .Y(n_575) );
INVx2_ASAP7_75t_L g241 ( .A(n_59), .Y(n_241) );
AOI22xp33_ASAP7_75t_L g369 ( .A1(n_60), .A2(n_150), .B1(n_370), .B2(n_371), .Y(n_369) );
INVx1_ASAP7_75t_L g670 ( .A(n_61), .Y(n_670) );
AND2x4_ASAP7_75t_L g673 ( .A(n_61), .B(n_241), .Y(n_673) );
INVx1_ASAP7_75t_SL g705 ( .A(n_61), .Y(n_705) );
AOI22xp33_ASAP7_75t_SL g626 ( .A1(n_62), .A2(n_233), .B1(n_627), .B2(n_628), .Y(n_626) );
AOI22xp33_ASAP7_75t_L g766 ( .A1(n_63), .A2(n_166), .B1(n_682), .B2(n_689), .Y(n_766) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_64), .A2(n_87), .B1(n_370), .B2(n_374), .Y(n_416) );
INVx1_ASAP7_75t_L g460 ( .A(n_65), .Y(n_460) );
INVx1_ASAP7_75t_L g639 ( .A(n_67), .Y(n_639) );
BUFx6f_ASAP7_75t_L g266 ( .A(n_68), .Y(n_266) );
AOI22xp33_ASAP7_75t_L g651 ( .A1(n_71), .A2(n_171), .B1(n_528), .B2(n_530), .Y(n_651) );
AOI22xp5_ASAP7_75t_L g463 ( .A1(n_72), .A2(n_229), .B1(n_464), .B2(n_466), .Y(n_463) );
AOI22xp5_ASAP7_75t_L g696 ( .A1(n_73), .A2(n_147), .B1(n_675), .B2(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g547 ( .A(n_74), .Y(n_547) );
AOI21x1_ASAP7_75t_SL g334 ( .A1(n_75), .A2(n_335), .B(n_340), .Y(n_334) );
AOI22xp33_ASAP7_75t_L g320 ( .A1(n_76), .A2(n_143), .B1(n_321), .B2(n_324), .Y(n_320) );
AOI22xp5_ASAP7_75t_L g649 ( .A1(n_77), .A2(n_148), .B1(n_307), .B2(n_522), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_78), .A2(n_175), .B1(n_668), .B2(n_672), .Y(n_667) );
AOI22xp33_ASAP7_75t_L g681 ( .A1(n_79), .A2(n_157), .B1(n_672), .B2(n_682), .Y(n_681) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_80), .A2(n_202), .B1(n_383), .B2(n_389), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g327 ( .A1(n_81), .A2(n_105), .B1(n_328), .B2(n_331), .Y(n_327) );
INVx1_ASAP7_75t_L g267 ( .A(n_82), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_82), .B(n_181), .Y(n_349) );
AOI22xp33_ASAP7_75t_L g411 ( .A1(n_83), .A2(n_100), .B1(n_389), .B2(n_390), .Y(n_411) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_84), .A2(n_127), .B1(n_355), .B2(n_507), .Y(n_506) );
AOI22xp33_ASAP7_75t_L g310 ( .A1(n_85), .A2(n_155), .B1(n_311), .B2(n_315), .Y(n_310) );
AOI22xp33_ASAP7_75t_L g258 ( .A1(n_86), .A2(n_178), .B1(n_259), .B2(n_285), .Y(n_258) );
XNOR2x1_ASAP7_75t_L g426 ( .A(n_88), .B(n_427), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_89), .B(n_451), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g685 ( .A1(n_90), .A2(n_151), .B1(n_675), .B2(n_686), .Y(n_685) );
AOI22xp5_ASAP7_75t_L g583 ( .A1(n_91), .A2(n_228), .B1(n_386), .B2(n_387), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g683 ( .A1(n_92), .A2(n_103), .B1(n_675), .B2(n_678), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_93), .B(n_415), .Y(n_414) );
AOI22xp33_ASAP7_75t_L g455 ( .A1(n_94), .A2(n_119), .B1(n_456), .B2(n_457), .Y(n_455) );
AOI221xp5_ASAP7_75t_SL g587 ( .A1(n_95), .A2(n_210), .B1(n_373), .B2(n_432), .C(n_588), .Y(n_587) );
CKINVDCx5p33_ASAP7_75t_R g589 ( .A(n_97), .Y(n_589) );
AOI221xp5_ASAP7_75t_L g590 ( .A1(n_98), .A2(n_161), .B1(n_370), .B2(n_374), .C(n_591), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g440 ( .A1(n_99), .A2(n_204), .B1(n_387), .B2(n_389), .Y(n_440) );
AOI21xp33_ASAP7_75t_L g458 ( .A1(n_101), .A2(n_415), .B(n_459), .Y(n_458) );
AOI22xp33_ASAP7_75t_L g486 ( .A1(n_102), .A2(n_201), .B1(n_304), .B2(n_307), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_104), .A2(n_159), .B1(n_609), .B2(n_610), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g763 ( .A1(n_106), .A2(n_184), .B1(n_686), .B2(n_764), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_109), .B(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g619 ( .A(n_110), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_111), .B(n_432), .Y(n_431) );
AOI22xp5_ASAP7_75t_L g693 ( .A1(n_112), .A2(n_218), .B1(n_675), .B2(n_678), .Y(n_693) );
AOI22xp5_ASAP7_75t_L g882 ( .A1(n_113), .A2(n_162), .B1(n_368), .B2(n_883), .Y(n_882) );
AOI22xp5_ASAP7_75t_L g586 ( .A1(n_114), .A2(n_140), .B1(n_384), .B2(n_390), .Y(n_586) );
NAND2xp33_ASAP7_75t_L g871 ( .A(n_115), .B(n_464), .Y(n_871) );
AOI22xp33_ASAP7_75t_L g391 ( .A1(n_116), .A2(n_167), .B1(n_392), .B2(n_393), .Y(n_391) );
INVx1_ASAP7_75t_L g436 ( .A(n_118), .Y(n_436) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_120), .A2(n_179), .B1(n_564), .B2(n_565), .Y(n_563) );
AOI21xp33_ASAP7_75t_SL g615 ( .A1(n_121), .A2(n_616), .B(n_618), .Y(n_615) );
AOI22xp5_ASAP7_75t_L g540 ( .A1(n_122), .A2(n_174), .B1(n_331), .B2(n_541), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g438 ( .A1(n_124), .A2(n_217), .B1(n_373), .B2(n_386), .Y(n_438) );
AOI22xp5_ASAP7_75t_L g467 ( .A1(n_125), .A2(n_156), .B1(n_468), .B2(n_469), .Y(n_467) );
AOI22xp33_ASAP7_75t_SL g577 ( .A1(n_129), .A2(n_205), .B1(n_296), .B2(n_300), .Y(n_577) );
INVx1_ASAP7_75t_L g353 ( .A(n_130), .Y(n_353) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_131), .A2(n_189), .B1(n_370), .B2(n_371), .Y(n_430) );
AOI22xp5_ASAP7_75t_L g600 ( .A1(n_132), .A2(n_153), .B1(n_601), .B2(n_604), .Y(n_600) );
OAI22xp5_ASAP7_75t_L g901 ( .A1(n_133), .A2(n_902), .B1(n_907), .B2(n_908), .Y(n_901) );
CKINVDCx5p33_ASAP7_75t_R g907 ( .A(n_133), .Y(n_907) );
AOI22xp33_ASAP7_75t_L g385 ( .A1(n_134), .A2(n_182), .B1(n_386), .B2(n_387), .Y(n_385) );
AOI22xp33_ASAP7_75t_SL g474 ( .A1(n_135), .A2(n_224), .B1(n_475), .B2(n_476), .Y(n_474) );
AOI22xp5_ASAP7_75t_L g703 ( .A1(n_136), .A2(n_214), .B1(n_678), .B2(n_704), .Y(n_703) );
AO22x1_ASAP7_75t_L g591 ( .A1(n_137), .A2(n_197), .B1(n_371), .B2(n_434), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g382 ( .A1(n_138), .A2(n_203), .B1(n_383), .B2(n_384), .Y(n_382) );
AOI22x1_ASAP7_75t_L g596 ( .A1(n_141), .A2(n_597), .B1(n_598), .B2(n_631), .Y(n_596) );
INVx1_ASAP7_75t_L g631 ( .A(n_141), .Y(n_631) );
OAI22x1_ASAP7_75t_L g654 ( .A1(n_141), .A2(n_597), .B1(n_598), .B2(n_631), .Y(n_654) );
AOI22xp33_ASAP7_75t_L g409 ( .A1(n_142), .A2(n_208), .B1(n_383), .B2(n_384), .Y(n_409) );
INVx1_ASAP7_75t_L g550 ( .A(n_144), .Y(n_550) );
AOI22xp5_ASAP7_75t_L g471 ( .A1(n_145), .A2(n_225), .B1(n_472), .B2(n_473), .Y(n_471) );
XNOR2x1_ASAP7_75t_L g447 ( .A(n_147), .B(n_448), .Y(n_447) );
AOI22xp5_ASAP7_75t_L g698 ( .A1(n_149), .A2(n_188), .B1(n_668), .B2(n_699), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_152), .B(n_565), .Y(n_621) );
AO221x2_ASAP7_75t_L g708 ( .A1(n_158), .A2(n_195), .B1(n_675), .B2(n_697), .C(n_709), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g429 ( .A1(n_160), .A2(n_190), .B1(n_374), .B2(n_383), .Y(n_429) );
OA22x2_ASAP7_75t_L g272 ( .A1(n_163), .A2(n_183), .B1(n_266), .B2(n_270), .Y(n_272) );
INVx1_ASAP7_75t_L g292 ( .A(n_163), .Y(n_292) );
AOI22xp5_ASAP7_75t_L g886 ( .A1(n_165), .A2(n_180), .B1(n_475), .B2(n_887), .Y(n_886) );
XNOR2x1_ASAP7_75t_L g255 ( .A(n_168), .B(n_256), .Y(n_255) );
INVx1_ASAP7_75t_L g419 ( .A(n_169), .Y(n_419) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_170), .A2(n_212), .B1(n_307), .B2(n_524), .Y(n_523) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_172), .A2(n_222), .B1(n_668), .B2(n_689), .Y(n_688) );
AOI221x1_ASAP7_75t_L g872 ( .A1(n_173), .A2(n_211), .B1(n_472), .B2(n_476), .C(n_873), .Y(n_872) );
INVx1_ASAP7_75t_L g284 ( .A(n_181), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_181), .B(n_290), .Y(n_360) );
OAI21xp33_ASAP7_75t_L g293 ( .A1(n_183), .A2(n_192), .B(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g873 ( .A(n_185), .B(n_470), .Y(n_873) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_192), .B(n_220), .Y(n_245) );
INVx1_ASAP7_75t_L g269 ( .A(n_192), .Y(n_269) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_193), .A2(n_216), .B1(n_392), .B2(n_393), .Y(n_412) );
INVx1_ASAP7_75t_L g364 ( .A(n_195), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g877 ( .A(n_196), .B(n_878), .Y(n_877) );
AOI22xp33_ASAP7_75t_L g622 ( .A1(n_200), .A2(n_207), .B1(n_623), .B2(n_625), .Y(n_622) );
AOI22xp5_ASAP7_75t_L g652 ( .A1(n_213), .A2(n_223), .B1(n_524), .B2(n_653), .Y(n_652) );
NOR3xp33_ASAP7_75t_L g869 ( .A(n_214), .B(n_870), .C(n_874), .Y(n_869) );
AOI22xp5_ASAP7_75t_L g891 ( .A1(n_214), .A2(n_874), .B1(n_880), .B2(n_913), .Y(n_891) );
OAI21xp5_ASAP7_75t_L g892 ( .A1(n_214), .A2(n_870), .B(n_885), .Y(n_892) );
AOI22xp33_ASAP7_75t_L g898 ( .A1(n_214), .A2(n_899), .B1(n_901), .B2(n_909), .Y(n_898) );
INVx1_ASAP7_75t_L g556 ( .A(n_215), .Y(n_556) );
INVx1_ASAP7_75t_L g480 ( .A(n_218), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_220), .B(n_276), .Y(n_275) );
AOI21xp33_ASAP7_75t_L g417 ( .A1(n_221), .A2(n_373), .B(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g677 ( .A(n_227), .Y(n_677) );
XNOR2x1_ASAP7_75t_L g518 ( .A(n_232), .B(n_519), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_247), .B(n_656), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
BUFx3_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
HB1xp67_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
NAND3xp33_ASAP7_75t_L g238 ( .A(n_239), .B(n_242), .C(n_246), .Y(n_238) );
AND2x2_ASAP7_75t_L g895 ( .A(n_239), .B(n_896), .Y(n_895) );
AND2x2_ASAP7_75t_L g900 ( .A(n_239), .B(n_897), .Y(n_900) );
INVx1_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
OA21x2_ASAP7_75t_L g910 ( .A1(n_240), .A2(n_705), .B(n_911), .Y(n_910) );
HB1xp67_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
AND2x2_ASAP7_75t_L g669 ( .A(n_241), .B(n_670), .Y(n_669) );
AND3x4_ASAP7_75t_L g704 ( .A(n_241), .B(n_676), .C(n_705), .Y(n_704) );
NOR2xp33_ASAP7_75t_L g896 ( .A(n_242), .B(n_897), .Y(n_896) );
HB1xp67_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
AO21x2_ASAP7_75t_L g357 ( .A1(n_243), .A2(n_358), .B(n_359), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_244), .B(n_245), .Y(n_243) );
INVx1_ASAP7_75t_L g897 ( .A(n_246), .Y(n_897) );
OAI22xp5_ASAP7_75t_L g247 ( .A1(n_248), .A2(n_249), .B1(n_512), .B2(n_513), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
XNOR2xp5_ASAP7_75t_L g249 ( .A(n_250), .B(n_400), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
OAI22xp5_ASAP7_75t_L g251 ( .A1(n_252), .A2(n_361), .B1(n_395), .B2(n_399), .Y(n_251) );
INVxp67_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
HB1xp67_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
BUFx3_ASAP7_75t_L g398 ( .A(n_255), .Y(n_398) );
NAND4xp75_ASAP7_75t_SL g256 ( .A(n_257), .B(n_302), .C(n_319), .D(n_334), .Y(n_256) );
AND2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_295), .Y(n_257) );
BUFx12f_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
BUFx6f_ASAP7_75t_L g612 ( .A(n_260), .Y(n_612) );
BUFx12f_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
BUFx6f_ASAP7_75t_L g473 ( .A(n_261), .Y(n_473) );
BUFx6f_ASAP7_75t_L g493 ( .A(n_261), .Y(n_493) );
AND2x4_ASAP7_75t_L g261 ( .A(n_262), .B(n_273), .Y(n_261) );
AND2x4_ASAP7_75t_L g297 ( .A(n_262), .B(n_298), .Y(n_297) );
AND2x4_ASAP7_75t_L g312 ( .A(n_262), .B(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g316 ( .A(n_262), .B(n_317), .Y(n_316) );
AND2x4_ASAP7_75t_L g383 ( .A(n_262), .B(n_309), .Y(n_383) );
AND2x4_ASAP7_75t_L g389 ( .A(n_262), .B(n_273), .Y(n_389) );
AND2x4_ASAP7_75t_L g392 ( .A(n_262), .B(n_313), .Y(n_392) );
AND2x4_ASAP7_75t_L g393 ( .A(n_262), .B(n_317), .Y(n_393) );
AND2x4_ASAP7_75t_L g262 ( .A(n_263), .B(n_271), .Y(n_262) );
AND2x2_ASAP7_75t_L g323 ( .A(n_263), .B(n_272), .Y(n_323) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g306 ( .A(n_264), .B(n_272), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_265), .B(n_268), .Y(n_264) );
NAND2xp33_ASAP7_75t_L g265 ( .A(n_266), .B(n_267), .Y(n_265) );
INVx2_ASAP7_75t_L g270 ( .A(n_266), .Y(n_270) );
INVx3_ASAP7_75t_L g276 ( .A(n_266), .Y(n_276) );
NAND2xp33_ASAP7_75t_L g283 ( .A(n_266), .B(n_284), .Y(n_283) );
INVx1_ASAP7_75t_L g294 ( .A(n_266), .Y(n_294) );
HB1xp67_ASAP7_75t_L g348 ( .A(n_266), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_267), .B(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
OAI21xp5_ASAP7_75t_L g351 ( .A1(n_269), .A2(n_294), .B(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g350 ( .A(n_272), .B(n_351), .Y(n_350) );
AND2x4_ASAP7_75t_L g287 ( .A(n_273), .B(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g305 ( .A(n_273), .B(n_306), .Y(n_305) );
AND2x4_ASAP7_75t_L g386 ( .A(n_273), .B(n_306), .Y(n_386) );
AND2x4_ASAP7_75t_L g390 ( .A(n_273), .B(n_288), .Y(n_390) );
AND2x2_ASAP7_75t_L g470 ( .A(n_273), .B(n_306), .Y(n_470) );
AND2x4_ASAP7_75t_L g273 ( .A(n_274), .B(n_278), .Y(n_273) );
OR2x2_ASAP7_75t_L g299 ( .A(n_274), .B(n_279), .Y(n_299) );
AND2x4_ASAP7_75t_L g313 ( .A(n_274), .B(n_314), .Y(n_313) );
INVx2_ASAP7_75t_L g318 ( .A(n_274), .Y(n_318) );
AND2x2_ASAP7_75t_L g346 ( .A(n_274), .B(n_347), .Y(n_346) );
AND2x4_ASAP7_75t_L g274 ( .A(n_275), .B(n_277), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_276), .B(n_282), .Y(n_281) );
INVxp67_ASAP7_75t_L g290 ( .A(n_276), .Y(n_290) );
NAND3xp33_ASAP7_75t_L g359 ( .A(n_277), .B(n_289), .C(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
INVx1_ASAP7_75t_L g314 ( .A(n_280), .Y(n_314) );
AND2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_283), .Y(n_280) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx2_ASAP7_75t_L g468 ( .A(n_286), .Y(n_468) );
INVx4_ASAP7_75t_L g494 ( .A(n_286), .Y(n_494) );
INVx2_ASAP7_75t_SL g526 ( .A(n_286), .Y(n_526) );
INVx4_ASAP7_75t_L g576 ( .A(n_286), .Y(n_576) );
INVx2_ASAP7_75t_L g653 ( .A(n_286), .Y(n_653) );
INVx4_ASAP7_75t_L g887 ( .A(n_286), .Y(n_887) );
INVx8_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
AND2x4_ASAP7_75t_L g301 ( .A(n_288), .B(n_298), .Y(n_301) );
AND2x4_ASAP7_75t_L g333 ( .A(n_288), .B(n_317), .Y(n_333) );
AND2x4_ASAP7_75t_L g371 ( .A(n_288), .B(n_317), .Y(n_371) );
AND2x4_ASAP7_75t_L g384 ( .A(n_288), .B(n_298), .Y(n_384) );
AND2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_293), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
BUFx6f_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
BUFx6f_ASAP7_75t_L g472 ( .A(n_297), .Y(n_472) );
BUFx6f_ASAP7_75t_L g485 ( .A(n_297), .Y(n_485) );
BUFx6f_ASAP7_75t_L g603 ( .A(n_297), .Y(n_603) );
AND2x4_ASAP7_75t_L g387 ( .A(n_298), .B(n_306), .Y(n_387) );
INVx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx2_ASAP7_75t_L g309 ( .A(n_299), .Y(n_309) );
BUFx3_ASAP7_75t_L g604 ( .A(n_300), .Y(n_604) );
BUFx12f_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx6_ASAP7_75t_L g465 ( .A(n_301), .Y(n_465) );
AND2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_310), .Y(n_302) );
BUFx8_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
BUFx6f_ASAP7_75t_L g524 ( .A(n_305), .Y(n_524) );
AND2x4_ASAP7_75t_L g308 ( .A(n_306), .B(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g326 ( .A(n_306), .B(n_313), .Y(n_326) );
AND2x2_ASAP7_75t_L g339 ( .A(n_306), .B(n_317), .Y(n_339) );
AND2x4_ASAP7_75t_L g370 ( .A(n_306), .B(n_313), .Y(n_370) );
AND2x2_ASAP7_75t_L g434 ( .A(n_306), .B(n_317), .Y(n_434) );
BUFx6f_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
BUFx12f_ASAP7_75t_L g466 ( .A(n_308), .Y(n_466) );
BUFx3_ASAP7_75t_L g569 ( .A(n_308), .Y(n_569) );
BUFx6f_ASAP7_75t_L g889 ( .A(n_308), .Y(n_889) );
BUFx6f_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
BUFx12f_ASAP7_75t_L g476 ( .A(n_312), .Y(n_476) );
INVx3_ASAP7_75t_L g529 ( .A(n_312), .Y(n_529) );
AND2x4_ASAP7_75t_L g322 ( .A(n_313), .B(n_323), .Y(n_322) );
AND2x4_ASAP7_75t_L g373 ( .A(n_313), .B(n_323), .Y(n_373) );
AND2x4_ASAP7_75t_L g317 ( .A(n_314), .B(n_318), .Y(n_317) );
BUFx5_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
BUFx3_ASAP7_75t_L g475 ( .A(n_316), .Y(n_475) );
INVx1_ASAP7_75t_L g491 ( .A(n_316), .Y(n_491) );
BUFx6f_ASAP7_75t_L g530 ( .A(n_316), .Y(n_530) );
AND2x4_ASAP7_75t_L g330 ( .A(n_317), .B(n_323), .Y(n_330) );
AND2x2_ASAP7_75t_L g376 ( .A(n_317), .B(n_323), .Y(n_376) );
AND2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_327), .Y(n_319) );
BUFx6f_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
BUFx3_ASAP7_75t_L g456 ( .A(n_322), .Y(n_456) );
INVx1_ASAP7_75t_L g503 ( .A(n_322), .Y(n_503) );
BUFx3_ASAP7_75t_L g549 ( .A(n_322), .Y(n_549) );
INVx2_ASAP7_75t_L g551 ( .A(n_324), .Y(n_551) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
BUFx6f_ASAP7_75t_L g542 ( .A(n_325), .Y(n_542) );
INVx2_ASAP7_75t_L g876 ( .A(n_325), .Y(n_876) );
INVx2_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
BUFx6f_ASAP7_75t_L g453 ( .A(n_326), .Y(n_453) );
BUFx3_ASAP7_75t_L g630 ( .A(n_326), .Y(n_630) );
INVx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx3_ASAP7_75t_L g555 ( .A(n_329), .Y(n_555) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
BUFx6f_ASAP7_75t_L g432 ( .A(n_330), .Y(n_432) );
BUFx8_ASAP7_75t_SL g451 ( .A(n_330), .Y(n_451) );
INVx2_ASAP7_75t_L g499 ( .A(n_330), .Y(n_499) );
BUFx6f_ASAP7_75t_L g624 ( .A(n_330), .Y(n_624) );
BUFx3_ASAP7_75t_L g878 ( .A(n_330), .Y(n_878) );
INVx3_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx2_ASAP7_75t_L g558 ( .A(n_332), .Y(n_558) );
INVx3_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
BUFx6f_ASAP7_75t_L g457 ( .A(n_333), .Y(n_457) );
BUFx6f_ASAP7_75t_L g500 ( .A(n_333), .Y(n_500) );
HB1xp67_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
BUFx6f_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx2_ASAP7_75t_L g368 ( .A(n_338), .Y(n_368) );
INVx2_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
BUFx3_ASAP7_75t_L g415 ( .A(n_339), .Y(n_415) );
INVx3_ASAP7_75t_L g534 ( .A(n_339), .Y(n_534) );
OAI22xp5_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_342), .B1(n_353), .B2(n_354), .Y(n_340) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx4_ASAP7_75t_L g507 ( .A(n_344), .Y(n_507) );
INVx5_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
BUFx2_ASAP7_75t_L g454 ( .A(n_345), .Y(n_454) );
BUFx4f_ASAP7_75t_L g564 ( .A(n_345), .Y(n_564) );
AND2x4_ASAP7_75t_L g345 ( .A(n_346), .B(n_350), .Y(n_345) );
AND2x2_ASAP7_75t_L g374 ( .A(n_346), .B(n_350), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_348), .B(n_349), .Y(n_347) );
INVx1_ASAP7_75t_L g358 ( .A(n_348), .Y(n_358) );
INVx2_ASAP7_75t_SL g354 ( .A(n_355), .Y(n_354) );
INVx2_ASAP7_75t_SL g355 ( .A(n_356), .Y(n_355) );
BUFx6f_ASAP7_75t_L g461 ( .A(n_356), .Y(n_461) );
INVx2_ASAP7_75t_L g538 ( .A(n_356), .Y(n_538) );
NOR2xp33_ASAP7_75t_L g588 ( .A(n_356), .B(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g643 ( .A(n_356), .Y(n_643) );
BUFx6f_ASAP7_75t_L g884 ( .A(n_356), .Y(n_884) );
BUFx6f_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx3_ASAP7_75t_L g380 ( .A(n_357), .Y(n_380) );
INVx1_ASAP7_75t_SL g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g399 ( .A(n_363), .Y(n_399) );
AO21x2_ASAP7_75t_L g363 ( .A1(n_364), .A2(n_365), .B(n_394), .Y(n_363) );
NOR3xp33_ASAP7_75t_SL g394 ( .A(n_364), .B(n_366), .C(n_381), .Y(n_394) );
OR2x2_ASAP7_75t_L g365 ( .A(n_366), .B(n_381), .Y(n_365) );
NAND4xp75_ASAP7_75t_L g366 ( .A(n_367), .B(n_369), .C(n_372), .D(n_375), .Y(n_366) );
BUFx3_ASAP7_75t_L g505 ( .A(n_368), .Y(n_505) );
NOR2xp33_ASAP7_75t_L g377 ( .A(n_378), .B(n_379), .Y(n_377) );
NOR2xp33_ASAP7_75t_L g435 ( .A(n_379), .B(n_436), .Y(n_435) );
INVx4_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx3_ASAP7_75t_L g420 ( .A(n_380), .Y(n_420) );
NAND4xp25_ASAP7_75t_L g381 ( .A(n_382), .B(n_385), .C(n_388), .D(n_391), .Y(n_381) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
AOI22xp5_ASAP7_75t_SL g400 ( .A1(n_401), .A2(n_402), .B1(n_443), .B2(n_511), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
OAI22xp5_ASAP7_75t_L g402 ( .A1(n_403), .A2(n_423), .B1(n_424), .B2(n_442), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVxp33_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
HB1xp67_ASAP7_75t_L g442 ( .A(n_406), .Y(n_442) );
XOR2x2_ASAP7_75t_L g406 ( .A(n_407), .B(n_422), .Y(n_406) );
NOR2xp67_ASAP7_75t_L g407 ( .A(n_408), .B(n_413), .Y(n_407) );
NAND4xp25_ASAP7_75t_L g408 ( .A(n_409), .B(n_410), .C(n_411), .D(n_412), .Y(n_408) );
NAND4xp25_ASAP7_75t_L g413 ( .A(n_414), .B(n_416), .C(n_417), .D(n_421), .Y(n_413) );
BUFx3_ASAP7_75t_L g617 ( .A(n_415), .Y(n_617) );
NOR2xp33_ASAP7_75t_L g418 ( .A(n_419), .B(n_420), .Y(n_418) );
INVx4_ASAP7_75t_L g565 ( .A(n_420), .Y(n_565) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
NOR2x1_ASAP7_75t_L g427 ( .A(n_428), .B(n_437), .Y(n_427) );
NAND4xp25_ASAP7_75t_L g428 ( .A(n_429), .B(n_430), .C(n_431), .D(n_433), .Y(n_428) );
NAND4xp25_ASAP7_75t_L g437 ( .A(n_438), .B(n_439), .C(n_440), .D(n_441), .Y(n_437) );
INVx1_ASAP7_75t_L g511 ( .A(n_443), .Y(n_511) );
AOI22x1_ASAP7_75t_L g443 ( .A1(n_444), .A2(n_445), .B1(n_477), .B2(n_509), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_SL g446 ( .A(n_447), .Y(n_446) );
NOR2x1_ASAP7_75t_L g448 ( .A(n_449), .B(n_462), .Y(n_448) );
NAND4xp25_ASAP7_75t_L g449 ( .A(n_450), .B(n_452), .C(n_455), .D(n_458), .Y(n_449) );
BUFx2_ASAP7_75t_L g627 ( .A(n_456), .Y(n_627) );
NOR2xp33_ASAP7_75t_L g459 ( .A(n_460), .B(n_461), .Y(n_459) );
NAND4xp25_ASAP7_75t_L g462 ( .A(n_463), .B(n_467), .C(n_471), .D(n_474), .Y(n_462) );
INVx5_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx3_ASAP7_75t_L g522 ( .A(n_465), .Y(n_522) );
BUFx3_ASAP7_75t_L g607 ( .A(n_466), .Y(n_607) );
BUFx2_ASAP7_75t_SL g613 ( .A(n_468), .Y(n_613) );
BUFx4f_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
BUFx6f_ASAP7_75t_L g606 ( .A(n_470), .Y(n_606) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
BUFx2_ASAP7_75t_L g510 ( .A(n_479), .Y(n_510) );
AO21x2_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_481), .B(n_508), .Y(n_479) );
NOR3xp33_ASAP7_75t_SL g508 ( .A(n_480), .B(n_483), .C(n_496), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_482), .B(n_495), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
NAND4xp25_ASAP7_75t_SL g483 ( .A(n_484), .B(n_486), .C(n_487), .D(n_492), .Y(n_483) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
BUFx6f_ASAP7_75t_L g573 ( .A(n_490), .Y(n_573) );
INVx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
NAND4xp25_ASAP7_75t_L g496 ( .A(n_497), .B(n_501), .C(n_504), .D(n_506), .Y(n_496) );
INVx2_ASAP7_75t_SL g498 ( .A(n_499), .Y(n_498) );
BUFx3_ASAP7_75t_L g625 ( .A(n_500), .Y(n_625) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx2_ASAP7_75t_L g646 ( .A(n_503), .Y(n_646) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
XOR2xp5_ASAP7_75t_L g513 ( .A(n_514), .B(n_595), .Y(n_513) );
OAI22xp5_ASAP7_75t_L g514 ( .A1(n_515), .A2(n_516), .B1(n_578), .B2(n_594), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
XNOR2xp5_ASAP7_75t_L g516 ( .A(n_517), .B(n_543), .Y(n_516) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
NOR2x1_ASAP7_75t_L g519 ( .A(n_520), .B(n_531), .Y(n_519) );
NAND4xp25_ASAP7_75t_L g520 ( .A(n_521), .B(n_523), .C(n_525), .D(n_527), .Y(n_520) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx2_ASAP7_75t_L g572 ( .A(n_529), .Y(n_572) );
INVx1_ASAP7_75t_L g609 ( .A(n_529), .Y(n_609) );
BUFx2_ASAP7_75t_SL g610 ( .A(n_530), .Y(n_610) );
NAND3xp33_ASAP7_75t_L g531 ( .A(n_532), .B(n_539), .C(n_540), .Y(n_531) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx2_ASAP7_75t_L g562 ( .A(n_534), .Y(n_562) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_536), .B(n_537), .Y(n_535) );
INVx3_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
AND2x2_ASAP7_75t_L g544 ( .A(n_545), .B(n_566), .Y(n_544) );
NOR3xp33_ASAP7_75t_L g545 ( .A(n_546), .B(n_552), .C(n_559), .Y(n_545) );
OAI22xp5_ASAP7_75t_L g546 ( .A1(n_547), .A2(n_548), .B1(n_550), .B2(n_551), .Y(n_546) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
OAI22xp5_ASAP7_75t_L g552 ( .A1(n_553), .A2(n_554), .B1(n_556), .B2(n_557), .Y(n_552) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
OAI21xp33_ASAP7_75t_L g559 ( .A1(n_560), .A2(n_561), .B(n_563), .Y(n_559) );
INVx2_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx2_ASAP7_75t_SL g620 ( .A(n_564), .Y(n_620) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_567), .B(n_574), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_568), .B(n_570), .Y(n_567) );
BUFx4f_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_575), .B(n_577), .Y(n_574) );
INVx1_ASAP7_75t_SL g594 ( .A(n_578), .Y(n_594) );
BUFx4_ASAP7_75t_R g578 ( .A(n_579), .Y(n_578) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g592 ( .A(n_581), .Y(n_592) );
NAND3xp33_ASAP7_75t_L g581 ( .A(n_582), .B(n_587), .C(n_590), .Y(n_581) );
AND4x1_ASAP7_75t_L g582 ( .A(n_583), .B(n_584), .C(n_585), .D(n_586), .Y(n_582) );
OAI22xp5_ASAP7_75t_L g595 ( .A1(n_596), .A2(n_632), .B1(n_654), .B2(n_655), .Y(n_595) );
INVx2_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
OR2x2_ASAP7_75t_L g598 ( .A(n_599), .B(n_614), .Y(n_598) );
NAND4xp25_ASAP7_75t_SL g599 ( .A(n_600), .B(n_605), .C(n_608), .D(n_611), .Y(n_599) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
NAND3xp33_ASAP7_75t_L g614 ( .A(n_615), .B(n_622), .C(n_626), .Y(n_614) );
HB1xp67_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
OAI21xp33_ASAP7_75t_L g618 ( .A1(n_619), .A2(n_620), .B(n_621), .Y(n_618) );
BUFx3_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx2_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx2_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
HB1xp67_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
HB1xp67_ASAP7_75t_L g655 ( .A(n_634), .Y(n_655) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
XNOR2xp5_ASAP7_75t_L g637 ( .A(n_638), .B(n_640), .Y(n_637) );
CKINVDCx5p33_ASAP7_75t_R g638 ( .A(n_639), .Y(n_638) );
NOR2x1_ASAP7_75t_L g640 ( .A(n_641), .B(n_648), .Y(n_640) );
NAND4xp25_ASAP7_75t_L g641 ( .A(n_642), .B(n_644), .C(n_645), .D(n_647), .Y(n_641) );
NAND4xp25_ASAP7_75t_L g648 ( .A(n_649), .B(n_650), .C(n_651), .D(n_652), .Y(n_648) );
OAI221xp5_ASAP7_75t_L g656 ( .A1(n_657), .A2(n_863), .B1(n_865), .B2(n_893), .C(n_898), .Y(n_656) );
AND5x1_ASAP7_75t_L g657 ( .A(n_658), .B(n_800), .C(n_851), .D(n_856), .E(n_861), .Y(n_657) );
AOI21xp5_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_761), .B(n_767), .Y(n_658) );
NAND3xp33_ASAP7_75t_SL g659 ( .A(n_660), .B(n_721), .C(n_732), .Y(n_659) );
O2A1O1Ixp33_ASAP7_75t_L g660 ( .A1(n_661), .A2(n_690), .B(n_694), .C(n_710), .Y(n_660) );
AND2x2_ASAP7_75t_L g661 ( .A(n_662), .B(n_679), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g853 ( .A(n_662), .B(n_854), .Y(n_853) );
HB1xp67_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g725 ( .A(n_663), .Y(n_725) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g781 ( .A(n_664), .Y(n_781) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
OR2x2_ASAP7_75t_L g745 ( .A(n_665), .B(n_746), .Y(n_745) );
INVx2_ASAP7_75t_L g829 ( .A(n_665), .Y(n_829) );
INVx4_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
NOR2xp33_ASAP7_75t_L g690 ( .A(n_666), .B(n_691), .Y(n_690) );
OR2x2_ASAP7_75t_L g747 ( .A(n_666), .B(n_680), .Y(n_747) );
AND2x2_ASAP7_75t_L g757 ( .A(n_666), .B(n_746), .Y(n_757) );
OR2x2_ASAP7_75t_L g791 ( .A(n_666), .B(n_746), .Y(n_791) );
NOR2xp33_ASAP7_75t_L g840 ( .A(n_666), .B(n_770), .Y(n_840) );
AND2x2_ASAP7_75t_L g666 ( .A(n_667), .B(n_674), .Y(n_666) );
AND2x2_ASAP7_75t_L g668 ( .A(n_669), .B(n_671), .Y(n_668) );
AND2x4_ASAP7_75t_L g675 ( .A(n_669), .B(n_676), .Y(n_675) );
AND2x4_ASAP7_75t_L g682 ( .A(n_669), .B(n_671), .Y(n_682) );
AND2x2_ASAP7_75t_L g707 ( .A(n_669), .B(n_671), .Y(n_707) );
AND2x2_ASAP7_75t_L g672 ( .A(n_671), .B(n_673), .Y(n_672) );
AND2x4_ASAP7_75t_L g689 ( .A(n_671), .B(n_673), .Y(n_689) );
AND2x2_ASAP7_75t_L g699 ( .A(n_671), .B(n_673), .Y(n_699) );
AND2x4_ASAP7_75t_L g678 ( .A(n_673), .B(n_676), .Y(n_678) );
AND2x4_ASAP7_75t_L g697 ( .A(n_673), .B(n_676), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g864 ( .A(n_673), .B(n_676), .Y(n_864) );
INVx3_ASAP7_75t_L g765 ( .A(n_675), .Y(n_765) );
CKINVDCx5p33_ASAP7_75t_R g911 ( .A(n_676), .Y(n_911) );
INVx2_ASAP7_75t_SL g687 ( .A(n_678), .Y(n_687) );
INVx1_ASAP7_75t_L g720 ( .A(n_679), .Y(n_720) );
AND2x2_ASAP7_75t_L g679 ( .A(n_680), .B(n_684), .Y(n_679) );
INVx2_ASAP7_75t_L g746 ( .A(n_680), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_681), .B(n_683), .Y(n_680) );
INVx4_ASAP7_75t_L g759 ( .A(n_684), .Y(n_759) );
AND2x2_ASAP7_75t_L g771 ( .A(n_684), .B(n_744), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_684), .B(n_781), .Y(n_780) );
INVx1_ASAP7_75t_L g803 ( .A(n_684), .Y(n_803) );
AND2x2_ASAP7_75t_L g828 ( .A(n_684), .B(n_829), .Y(n_828) );
AND2x2_ASAP7_75t_L g684 ( .A(n_685), .B(n_688), .Y(n_684) );
INVx2_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g820 ( .A(n_690), .Y(n_820) );
NOR2xp33_ASAP7_75t_L g712 ( .A(n_691), .B(n_713), .Y(n_712) );
INVx3_ASAP7_75t_L g730 ( .A(n_691), .Y(n_730) );
INVx2_ASAP7_75t_L g743 ( .A(n_691), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_691), .B(n_757), .Y(n_756) );
INVx2_ASAP7_75t_L g770 ( .A(n_691), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_691), .B(n_759), .Y(n_799) );
AND2x2_ASAP7_75t_L g813 ( .A(n_691), .B(n_717), .Y(n_813) );
AND2x2_ASAP7_75t_L g691 ( .A(n_692), .B(n_693), .Y(n_691) );
AND2x2_ASAP7_75t_L g848 ( .A(n_694), .B(n_743), .Y(n_848) );
AND2x2_ASAP7_75t_L g694 ( .A(n_695), .B(n_700), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_695), .B(n_708), .Y(n_713) );
CKINVDCx6p67_ASAP7_75t_R g717 ( .A(n_695), .Y(n_717) );
AND2x2_ASAP7_75t_L g735 ( .A(n_695), .B(n_729), .Y(n_735) );
AND2x2_ASAP7_75t_L g738 ( .A(n_695), .B(n_739), .Y(n_738) );
AND2x2_ASAP7_75t_L g786 ( .A(n_695), .B(n_718), .Y(n_786) );
AND2x2_ASAP7_75t_L g787 ( .A(n_695), .B(n_702), .Y(n_787) );
NOR2xp33_ASAP7_75t_L g818 ( .A(n_695), .B(n_701), .Y(n_818) );
AND2x2_ASAP7_75t_L g695 ( .A(n_696), .B(n_698), .Y(n_695) );
INVx1_ASAP7_75t_L g755 ( .A(n_700), .Y(n_755) );
AND2x2_ASAP7_75t_L g805 ( .A(n_700), .B(n_717), .Y(n_805) );
AND2x2_ASAP7_75t_L g812 ( .A(n_700), .B(n_813), .Y(n_812) );
AND2x2_ASAP7_75t_L g700 ( .A(n_701), .B(n_708), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_701), .B(n_717), .Y(n_798) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
AND2x2_ASAP7_75t_L g718 ( .A(n_702), .B(n_719), .Y(n_718) );
OR2x2_ASAP7_75t_L g731 ( .A(n_702), .B(n_708), .Y(n_731) );
AND2x2_ASAP7_75t_L g736 ( .A(n_702), .B(n_708), .Y(n_736) );
OAI22xp33_ASAP7_75t_L g748 ( .A1(n_702), .A2(n_749), .B1(n_752), .B2(n_756), .Y(n_748) );
AND2x2_ASAP7_75t_L g702 ( .A(n_703), .B(n_706), .Y(n_702) );
INVx1_ASAP7_75t_L g719 ( .A(n_708), .Y(n_719) );
AND2x2_ASAP7_75t_L g774 ( .A(n_708), .B(n_717), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g832 ( .A(n_708), .B(n_735), .Y(n_832) );
AOI21xp5_ASAP7_75t_L g710 ( .A1(n_711), .A2(n_714), .B(n_720), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
O2A1O1Ixp33_ASAP7_75t_L g794 ( .A1(n_712), .A2(n_786), .B(n_790), .C(n_795), .Y(n_794) );
OAI322xp33_ASAP7_75t_L g801 ( .A1(n_714), .A2(n_717), .A3(n_744), .B1(n_745), .B2(n_789), .C1(n_802), .C2(n_804), .Y(n_801) );
INVx2_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
NOR2xp33_ASAP7_75t_L g760 ( .A(n_716), .B(n_741), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_717), .B(n_718), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_717), .B(n_728), .Y(n_727) );
AND2x2_ASAP7_75t_L g825 ( .A(n_717), .B(n_736), .Y(n_825) );
NAND2xp5_ASAP7_75t_L g846 ( .A(n_717), .B(n_847), .Y(n_846) );
INVx1_ASAP7_75t_L g754 ( .A(n_718), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g835 ( .A(n_718), .B(n_729), .Y(n_835) );
OAI211xp5_ASAP7_75t_SL g814 ( .A1(n_719), .A2(n_815), .B(n_817), .C(n_830), .Y(n_814) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_722), .B(n_726), .Y(n_721) );
HB1xp67_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
NOR2xp33_ASAP7_75t_L g821 ( .A(n_723), .B(n_822), .Y(n_821) );
HB1xp67_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g811 ( .A(n_725), .Y(n_811) );
NAND2xp5_ASAP7_75t_L g792 ( .A(n_726), .B(n_793), .Y(n_792) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g826 ( .A(n_728), .Y(n_826) );
O2A1O1Ixp33_ASAP7_75t_L g856 ( .A1(n_728), .A2(n_771), .B(n_857), .C(n_859), .Y(n_856) );
NOR2x1_ASAP7_75t_L g728 ( .A(n_729), .B(n_731), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_729), .B(n_750), .Y(n_749) );
AOI22xp5_ASAP7_75t_L g815 ( .A1(n_729), .A2(n_744), .B1(n_758), .B2(n_816), .Y(n_815) );
INVx3_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
AND2x2_ASAP7_75t_L g847 ( .A(n_730), .B(n_736), .Y(n_847) );
INVx1_ASAP7_75t_L g739 ( .A(n_731), .Y(n_739) );
AOI211xp5_ASAP7_75t_SL g795 ( .A1(n_731), .A2(n_745), .B(n_796), .C(n_799), .Y(n_795) );
AOI221xp5_ASAP7_75t_L g732 ( .A1(n_733), .A2(n_740), .B1(n_748), .B2(n_758), .C(n_760), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_734), .B(n_737), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_735), .B(n_736), .Y(n_734) );
AND2x2_ASAP7_75t_L g854 ( .A(n_735), .B(n_739), .Y(n_854) );
NAND2xp5_ASAP7_75t_L g822 ( .A(n_736), .B(n_813), .Y(n_822) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
AND2x2_ASAP7_75t_L g769 ( .A(n_738), .B(n_770), .Y(n_769) );
NAND3xp33_ASAP7_75t_L g839 ( .A(n_739), .B(n_777), .C(n_840), .Y(n_839) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_741), .B(n_747), .Y(n_740) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
AND2x2_ASAP7_75t_L g742 ( .A(n_743), .B(n_744), .Y(n_742) );
NOR2xp33_ASAP7_75t_L g772 ( .A(n_743), .B(n_773), .Y(n_772) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_743), .B(n_786), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_743), .B(n_787), .Y(n_809) );
NOR2xp33_ASAP7_75t_L g816 ( .A(n_743), .B(n_747), .Y(n_816) );
NOR2xp33_ASAP7_75t_L g849 ( .A(n_743), .B(n_850), .Y(n_849) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx2_ASAP7_75t_L g751 ( .A(n_746), .Y(n_751) );
INVxp67_ASAP7_75t_L g777 ( .A(n_746), .Y(n_777) );
AND2x2_ASAP7_75t_L g843 ( .A(n_746), .B(n_759), .Y(n_843) );
INVx1_ASAP7_75t_L g793 ( .A(n_747), .Y(n_793) );
NOR2xp33_ASAP7_75t_L g808 ( .A(n_747), .B(n_759), .Y(n_808) );
OAI22xp33_ASAP7_75t_L g859 ( .A1(n_747), .A2(n_809), .B1(n_837), .B2(n_860), .Y(n_859) );
OAI221xp5_ASAP7_75t_L g806 ( .A1(n_750), .A2(n_773), .B1(n_807), .B2(n_809), .C(n_810), .Y(n_806) );
INVx3_ASAP7_75t_SL g750 ( .A(n_751), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g837 ( .A(n_751), .B(n_759), .Y(n_837) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
AND2x2_ASAP7_75t_L g753 ( .A(n_754), .B(n_755), .Y(n_753) );
INVx1_ASAP7_75t_L g782 ( .A(n_757), .Y(n_782) );
NOR2xp33_ASAP7_75t_L g819 ( .A(n_758), .B(n_820), .Y(n_819) );
OAI21xp33_ASAP7_75t_L g851 ( .A1(n_758), .A2(n_852), .B(n_855), .Y(n_851) );
INVx2_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
OR2x2_ASAP7_75t_L g776 ( .A(n_759), .B(n_777), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_759), .B(n_790), .Y(n_789) );
AND2x2_ASAP7_75t_L g833 ( .A(n_759), .B(n_829), .Y(n_833) );
INVx2_ASAP7_75t_L g783 ( .A(n_761), .Y(n_783) );
OAI21xp5_ASAP7_75t_L g841 ( .A1(n_761), .A2(n_842), .B(n_844), .Y(n_841) );
CKINVDCx5p33_ASAP7_75t_R g761 ( .A(n_762), .Y(n_761) );
OAI211xp5_ASAP7_75t_L g836 ( .A1(n_762), .A2(n_837), .B(n_838), .C(n_839), .Y(n_836) );
AND2x2_ASAP7_75t_L g762 ( .A(n_763), .B(n_766), .Y(n_762) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
NAND4xp25_ASAP7_75t_SL g767 ( .A(n_768), .B(n_778), .C(n_792), .D(n_794), .Y(n_767) );
OAI31xp33_ASAP7_75t_L g768 ( .A1(n_769), .A2(n_771), .A3(n_772), .B(n_775), .Y(n_768) );
NOR2xp33_ASAP7_75t_L g857 ( .A(n_770), .B(n_858), .Y(n_857) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
INVx1_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
AOI22xp5_ASAP7_75t_L g778 ( .A1(n_779), .A2(n_784), .B1(n_787), .B2(n_788), .Y(n_778) );
AOI21xp33_ASAP7_75t_L g779 ( .A1(n_780), .A2(n_782), .B(n_783), .Y(n_779) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
INVx1_ASAP7_75t_L g850 ( .A(n_786), .Y(n_850) );
INVx1_ASAP7_75t_L g838 ( .A(n_787), .Y(n_838) );
INVx1_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
INVx1_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
AOI221xp5_ASAP7_75t_L g830 ( .A1(n_793), .A2(n_831), .B1(n_833), .B2(n_834), .C(n_836), .Y(n_830) );
INVx1_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
OAI31xp33_ASAP7_75t_SL g800 ( .A1(n_801), .A2(n_806), .A3(n_814), .B(n_841), .Y(n_800) );
INVx1_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
INVx1_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
NOR2xp33_ASAP7_75t_L g862 ( .A(n_807), .B(n_824), .Y(n_862) );
INVx1_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_811), .B(n_812), .Y(n_810) );
AOI211xp5_ASAP7_75t_L g817 ( .A1(n_818), .A2(n_819), .B(n_821), .C(n_823), .Y(n_817) );
INVx1_ASAP7_75t_L g858 ( .A(n_818), .Y(n_858) );
INVx1_ASAP7_75t_L g855 ( .A(n_822), .Y(n_855) );
AOI21xp33_ASAP7_75t_L g823 ( .A1(n_824), .A2(n_826), .B(n_827), .Y(n_823) );
INVx1_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
INVx1_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
AOI211xp5_ASAP7_75t_L g844 ( .A1(n_829), .A2(n_845), .B(n_848), .C(n_849), .Y(n_844) );
INVx1_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
INVx1_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
INVx1_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
INVx1_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
INVxp33_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
INVx1_ASAP7_75t_L g860 ( .A(n_854), .Y(n_860) );
INVxp67_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
BUFx2_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
HB1xp67_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
INVx1_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
INVx1_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
AO21x2_ASAP7_75t_L g868 ( .A1(n_869), .A2(n_879), .B(n_890), .Y(n_868) );
INVxp33_ASAP7_75t_SL g904 ( .A(n_870), .Y(n_904) );
NAND2xp5_ASAP7_75t_L g870 ( .A(n_871), .B(n_872), .Y(n_870) );
INVxp67_ASAP7_75t_L g905 ( .A(n_874), .Y(n_905) );
NAND2xp5_ASAP7_75t_SL g874 ( .A(n_875), .B(n_877), .Y(n_874) );
NOR2xp33_ASAP7_75t_L g879 ( .A(n_880), .B(n_885), .Y(n_879) );
INVxp33_ASAP7_75t_L g906 ( .A(n_880), .Y(n_906) );
NAND2xp5_ASAP7_75t_L g880 ( .A(n_881), .B(n_882), .Y(n_880) );
INVx2_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
INVxp67_ASAP7_75t_L g903 ( .A(n_885), .Y(n_903) );
NAND2x1_ASAP7_75t_SL g885 ( .A(n_886), .B(n_888), .Y(n_885) );
NAND2xp5_ASAP7_75t_L g890 ( .A(n_891), .B(n_892), .Y(n_890) );
INVx1_ASAP7_75t_L g893 ( .A(n_894), .Y(n_893) );
HB1xp67_ASAP7_75t_L g894 ( .A(n_895), .Y(n_894) );
BUFx3_ASAP7_75t_L g899 ( .A(n_900), .Y(n_899) );
INVx1_ASAP7_75t_L g908 ( .A(n_902), .Y(n_908) );
NAND4xp25_ASAP7_75t_L g902 ( .A(n_903), .B(n_904), .C(n_905), .D(n_906), .Y(n_902) );
HB1xp67_ASAP7_75t_L g909 ( .A(n_910), .Y(n_909) );
endmodule