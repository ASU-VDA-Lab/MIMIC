module real_jpeg_16384_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_202;
wire n_128;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx1_ASAP7_75t_SL g73 ( 
.A(n_0),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_1),
.A2(n_19),
.B(n_470),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_1),
.B(n_471),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_2),
.B(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_2),
.B(n_234),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_2),
.B(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_2),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_2),
.B(n_402),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_2),
.B(n_406),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_2),
.B(n_410),
.Y(n_409)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_3),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_3),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g356 ( 
.A(n_3),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_4),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_4),
.Y(n_78)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_4),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_4),
.Y(n_205)
);

BUFx5_ASAP7_75t_L g360 ( 
.A(n_4),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_4),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_5),
.B(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_5),
.B(n_95),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_5),
.B(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_5),
.B(n_311),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_6),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_6),
.B(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_6),
.B(n_134),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_6),
.B(n_105),
.Y(n_142)
);

AND2x2_ASAP7_75t_SL g197 ( 
.A(n_6),
.B(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_6),
.B(n_338),
.Y(n_337)
);

AND2x2_ASAP7_75t_SL g376 ( 
.A(n_6),
.B(n_377),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_7),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_7),
.B(n_75),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_7),
.B(n_36),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_7),
.B(n_120),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_7),
.B(n_138),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_7),
.B(n_91),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_7),
.B(n_118),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_7),
.B(n_456),
.Y(n_455)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_8),
.Y(n_194)
);

BUFx5_ASAP7_75t_L g379 ( 
.A(n_8),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_9),
.B(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_9),
.B(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_9),
.B(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_9),
.B(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_9),
.B(n_190),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_9),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_9),
.B(n_442),
.Y(n_441)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_10),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_10),
.Y(n_121)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_10),
.Y(n_131)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_10),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_11),
.Y(n_471)
);

AND2x2_ASAP7_75t_SL g46 ( 
.A(n_12),
.B(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_12),
.B(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_12),
.B(n_116),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_12),
.B(n_125),
.Y(n_196)
);

AND2x2_ASAP7_75t_SL g265 ( 
.A(n_12),
.B(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_12),
.B(n_358),
.Y(n_357)
);

AND2x2_ASAP7_75t_SL g374 ( 
.A(n_12),
.B(n_375),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_12),
.B(n_392),
.Y(n_391)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_13),
.Y(n_60)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_13),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_13),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_14),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx4f_ASAP7_75t_L g64 ( 
.A(n_15),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_15),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_16),
.B(n_31),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_16),
.B(n_58),
.Y(n_57)
);

AND2x2_ASAP7_75t_SL g229 ( 
.A(n_16),
.B(n_230),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_16),
.B(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_16),
.B(n_362),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_16),
.B(n_389),
.Y(n_388)
);

AND2x2_ASAP7_75t_SL g397 ( 
.A(n_16),
.B(n_398),
.Y(n_397)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_17),
.Y(n_69)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_17),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g294 ( 
.A(n_17),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_432),
.Y(n_19)
);

HB1xp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_315),
.Y(n_21)
);

A2O1A1O1Ixp25_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_216),
.B(n_274),
.C(n_275),
.D(n_314),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_24),
.B(n_276),
.Y(n_317)
);

AND2x2_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_177),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_25),
.B(n_177),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_99),
.Y(n_25)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_26),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_65),
.C(n_84),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_28),
.B(n_180),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_41),
.C(n_51),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_29),
.B(n_239),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_32),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_30),
.B(n_33),
.C(n_37),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_37),
.Y(n_32)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_36),
.Y(n_375)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_36),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_37),
.B(n_156),
.Y(n_330)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_38),
.B(n_90),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_38),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_41),
.A2(n_42),
.B1(n_51),
.B2(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_42),
.A2(n_43),
.B(n_46),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_46),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_44),
.B(n_45),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_45),
.B(n_461),
.Y(n_460)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_49),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_51),
.Y(n_240)
);

MAJx3_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_57),
.C(n_61),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_SL g184 ( 
.A(n_52),
.B(n_185),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_56),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_54),
.Y(n_312)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_55),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_56),
.B(n_332),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_57),
.B(n_61),
.Y(n_185)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_59),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_60),
.Y(n_118)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_64),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_65),
.A2(n_85),
.B1(n_86),
.B2(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_65),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_77),
.C(n_79),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_66),
.B(n_207),
.Y(n_206)
);

MAJx2_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_70),
.C(n_74),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_67),
.B(n_223),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_70),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_70),
.A2(n_202),
.B1(n_225),
.B2(n_258),
.Y(n_443)
);

OR2x2_ASAP7_75t_SL g70 ( 
.A(n_71),
.B(n_73),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_73),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_74),
.B(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_74),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_77),
.B(n_79),
.Y(n_207)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_83),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_83),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_88),
.Y(n_86)
);

MAJx2_ASAP7_75t_L g149 ( 
.A(n_87),
.B(n_89),
.C(n_94),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_93),
.B1(n_94),
.B2(n_98),
.Y(n_88)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_89),
.Y(n_98)
);

NAND2x1_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_91),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_90),
.B(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_90),
.B(n_154),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_90),
.B(n_157),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_90),
.B(n_203),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_90),
.B(n_292),
.Y(n_291)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_97),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_151),
.B1(n_175),
.B2(n_176),
.Y(n_99)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_100),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_139),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_101),
.B(n_148),
.C(n_281),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_113),
.C(n_127),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_102),
.B(n_113),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_108),
.Y(n_102)
);

OAI21xp33_ASAP7_75t_L g161 ( 
.A1(n_103),
.A2(n_110),
.B(n_111),
.Y(n_161)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_107),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_110),
.B1(n_111),
.B2(n_112),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_109),
.A2(n_110),
.B1(n_188),
.B2(n_189),
.Y(n_259)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_110),
.B(n_111),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_110),
.B(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_111),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_111),
.A2(n_112),
.B1(n_156),
.B2(n_158),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_111),
.B(n_153),
.C(n_158),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_111),
.B(n_337),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_112),
.B(n_337),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_119),
.C(n_122),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_114),
.A2(n_115),
.B1(n_122),
.B2(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_119),
.A2(n_209),
.B1(n_210),
.B2(n_212),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_119),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_119),
.A2(n_212),
.B1(n_310),
.B2(n_313),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_119),
.B(n_313),
.C(n_448),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx6_ASAP7_75t_L g201 ( 
.A(n_121),
.Y(n_201)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_122),
.Y(n_211)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g138 ( 
.A(n_126),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_126),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_127),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_132),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_128),
.B(n_133),
.C(n_147),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_131),
.Y(n_172)
);

INVxp67_ASAP7_75t_SL g402 ( 
.A(n_131),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_137),
.Y(n_132)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_137),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_148),
.B1(n_149),
.B2(n_150),
.Y(n_139)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_140),
.Y(n_150)
);

HB1xp67_ASAP7_75t_L g282 ( 
.A(n_140),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_146),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_143),
.B1(n_144),
.B2(n_145),
.Y(n_141)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_142),
.Y(n_145)
);

MAJx2_ASAP7_75t_L g287 ( 
.A(n_143),
.B(n_145),
.C(n_146),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_143),
.A2(n_144),
.B1(n_291),
.B2(n_295),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_143),
.B(n_291),
.C(n_464),
.Y(n_463)
);

INVx3_ASAP7_75t_SL g143 ( 
.A(n_144),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_147),
.B(n_460),
.Y(n_459)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_151),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_151),
.B(n_175),
.C(n_278),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_159),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_152),
.B(n_160),
.C(n_163),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_155),
.Y(n_152)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_156),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g298 ( 
.A1(n_156),
.A2(n_158),
.B1(n_202),
.B2(n_258),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_SL g445 ( 
.A(n_158),
.B(n_299),
.C(n_446),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_163),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_162),
.Y(n_160)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_162),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_162),
.A2(n_228),
.B1(n_325),
.B2(n_326),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_170),
.B1(n_173),
.B2(n_174),
.Y(n_164)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_165),
.Y(n_173)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_170),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_170),
.B(n_173),
.C(n_224),
.Y(n_306)
);

INVx6_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_182),
.C(n_213),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_179),
.B(n_213),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_182),
.B(n_242),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_206),
.C(n_208),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_183),
.B(n_220),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_186),
.C(n_195),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_184),
.B(n_252),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_186),
.A2(n_187),
.B1(n_195),
.B2(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx5_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx5_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx4_ASAP7_75t_L g412 ( 
.A(n_193),
.Y(n_412)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_195),
.Y(n_253)
);

MAJx2_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.C(n_202),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_196),
.A2(n_202),
.B1(n_257),
.B2(n_258),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_196),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_197),
.B(n_256),
.Y(n_255)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_201),
.Y(n_364)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_202),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g446 ( 
.A(n_202),
.Y(n_446)
);

BUFx2_ASAP7_75t_L g406 ( 
.A(n_203),
.Y(n_406)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx8_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_206),
.B(n_208),
.Y(n_220)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

AOI21x1_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_243),
.B(n_273),
.Y(n_216)
);

OR2x2_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_241),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_218),
.B(n_241),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_221),
.C(n_237),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_219),
.B(n_245),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_221),
.B(n_238),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_226),
.C(n_227),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_222),
.B(n_226),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_227),
.B(n_249),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.C(n_232),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_229),
.A2(n_232),
.B1(n_233),
.B2(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_SL g327 ( 
.A(n_229),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_236),
.Y(n_442)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_244),
.B(n_246),
.Y(n_243)
);

OR2x2_ASAP7_75t_L g316 ( 
.A(n_244),
.B(n_246),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_250),
.C(n_254),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_247),
.A2(n_248),
.B1(n_425),
.B2(n_426),
.Y(n_424)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_250),
.A2(n_251),
.B1(n_427),
.B2(n_428),
.Y(n_426)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_259),
.C(n_260),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_255),
.B(n_343),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_255),
.B(n_259),
.C(n_260),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_259),
.B(n_260),
.Y(n_343)
);

MAJx2_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_265),
.C(n_271),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_261),
.A2(n_262),
.B1(n_271),
.B2(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_264),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_265),
.B(n_366),
.Y(n_365)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g367 ( 
.A(n_271),
.Y(n_367)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_273),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_279),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_277),
.B(n_279),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_283),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_280),
.B(n_296),
.C(n_467),
.Y(n_466)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

XNOR2x1_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_296),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g467 ( 
.A(n_284),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_285),
.B(n_287),
.C(n_288),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_289),
.Y(n_464)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_291),
.Y(n_295)
);

INVx3_ASAP7_75t_SL g292 ( 
.A(n_293),
.Y(n_292)
);

INVx8_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

XNOR2x2_ASAP7_75t_SL g296 ( 
.A(n_297),
.B(n_305),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_297),
.B(n_306),
.C(n_307),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_304),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_309),
.Y(n_307)
);

INVxp33_ASAP7_75t_SL g448 ( 
.A(n_308),
.Y(n_448)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_310),
.Y(n_313)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

NAND4xp25_ASAP7_75t_SL g315 ( 
.A(n_316),
.B(n_317),
.C(n_318),
.D(n_319),
.Y(n_315)
);

OAI21x1_ASAP7_75t_SL g319 ( 
.A1(n_320),
.A2(n_423),
.B(n_431),
.Y(n_319)
);

AOI21x1_ASAP7_75t_SL g320 ( 
.A1(n_321),
.A2(n_368),
.B(n_422),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_322),
.B(n_344),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_322),
.B(n_344),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_342),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_328),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_324),
.B(n_328),
.C(n_430),
.Y(n_429)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_331),
.C(n_336),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_329),
.A2(n_330),
.B1(n_331),
.B2(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_331),
.Y(n_347)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_336),
.B(n_346),
.Y(n_345)
);

BUFx2_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx5_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g430 ( 
.A(n_342),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_348),
.C(n_365),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_345),
.B(n_383),
.Y(n_382)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_349),
.B(n_365),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_357),
.C(n_361),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_351),
.B(n_357),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_353),
.Y(n_351)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_361),
.B(n_372),
.Y(n_371)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

HB1xp67_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_SL g368 ( 
.A1(n_369),
.A2(n_384),
.B(n_421),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_382),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_370),
.B(n_382),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_373),
.C(n_380),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_371),
.B(n_418),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_373),
.A2(n_380),
.B1(n_381),
.B2(n_419),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_373),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_376),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_374),
.B(n_376),
.Y(n_394)
);

INVx3_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_385),
.A2(n_415),
.B(n_420),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_SL g385 ( 
.A1(n_386),
.A2(n_403),
.B(n_414),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_393),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_387),
.B(n_393),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_391),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_388),
.B(n_391),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_388),
.B(n_409),
.Y(n_408)
);

INVx3_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_395),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_394),
.B(n_397),
.C(n_400),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_396),
.A2(n_397),
.B1(n_400),
.B2(n_401),
.Y(n_395)
);

CKINVDCx16_ASAP7_75t_R g396 ( 
.A(n_397),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_404),
.A2(n_408),
.B(n_413),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_407),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_405),
.B(n_407),
.Y(n_413)
);

INVx2_ASAP7_75t_SL g410 ( 
.A(n_411),
.Y(n_410)
);

INVx5_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_417),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_416),
.B(n_417),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_429),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_424),
.B(n_429),
.Y(n_431)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_433),
.B(n_468),
.Y(n_432)
);

INVxp33_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_435),
.B(n_466),
.Y(n_434)
);

OR2x2_ASAP7_75t_L g469 ( 
.A(n_435),
.B(n_466),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_436),
.B(n_437),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_438),
.A2(n_439),
.B1(n_449),
.B2(n_450),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

XNOR2x2_ASAP7_75t_SL g439 ( 
.A(n_440),
.B(n_444),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_SL g440 ( 
.A(n_441),
.B(n_443),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_447),
.Y(n_444)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_451),
.B(n_465),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_452),
.A2(n_453),
.B1(n_462),
.B2(n_463),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_454),
.A2(n_455),
.B1(n_458),
.B2(n_459),
.Y(n_453)
);

CKINVDCx16_ASAP7_75t_R g454 ( 
.A(n_455),
.Y(n_454)
);

INVx4_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

INVxp33_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);


endmodule