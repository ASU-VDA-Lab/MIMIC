module fake_jpeg_23825_n_78 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_78);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_78;

wire n_10;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

BUFx16f_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_2),
.Y(n_11)
);

OR2x2_ASAP7_75t_L g12 ( 
.A(n_3),
.B(n_8),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_6),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_0),
.B(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_8),
.B(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_15),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_21),
.B(n_24),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_15),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_27),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_12),
.B(n_1),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_26),
.B(n_14),
.Y(n_34)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_12),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_33),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_21),
.B(n_14),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_35),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_33),
.A2(n_21),
.B1(n_24),
.B2(n_18),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_36),
.A2(n_39),
.B1(n_44),
.B2(n_17),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_30),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_37),
.B(n_38),
.Y(n_50)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

OAI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_29),
.A2(n_27),
.B1(n_23),
.B2(n_25),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_10),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_45),
.Y(n_46)
);

A2O1A1O1Ixp25_ASAP7_75t_L g42 ( 
.A1(n_31),
.A2(n_18),
.B(n_16),
.C(n_19),
.D(n_22),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_34),
.C(n_13),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_32),
.A2(n_17),
.B1(n_11),
.B2(n_13),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVxp67_ASAP7_75t_SL g47 ( 
.A(n_45),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

NOR2xp67_ASAP7_75t_R g57 ( 
.A(n_48),
.B(n_51),
.Y(n_57)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_53),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_37),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_52),
.B(n_43),
.Y(n_56)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_56),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_52),
.B(n_38),
.Y(n_59)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_59),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_48),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g64 ( 
.A(n_60),
.B(n_36),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_58),
.B(n_46),
.C(n_28),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_63),
.B(n_64),
.C(n_28),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_57),
.A2(n_42),
.B1(n_32),
.B2(n_23),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_SL g67 ( 
.A1(n_65),
.A2(n_28),
.B(n_27),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_66),
.B(n_68),
.C(n_69),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_67),
.A2(n_25),
.B(n_35),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_61),
.B(n_60),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_62),
.B(n_63),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_70),
.A2(n_55),
.B1(n_11),
.B2(n_22),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_66),
.B(n_64),
.C(n_35),
.Y(n_72)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_72),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_73),
.A2(n_20),
.B1(n_55),
.B2(n_4),
.Y(n_75)
);

AOI221xp5_ASAP7_75t_L g77 ( 
.A1(n_75),
.A2(n_76),
.B1(n_7),
.B2(n_20),
.C(n_5),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_74),
.A2(n_71),
.B1(n_7),
.B2(n_20),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_5),
.Y(n_78)
);


endmodule