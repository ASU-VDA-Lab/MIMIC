module fake_ariane_2604_n_1996 (n_295, n_356, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_516, n_332, n_294, n_197, n_463, n_176, n_34, n_404, n_172, n_347, n_423, n_183, n_469, n_479, n_373, n_299, n_499, n_12, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_522, n_319, n_49, n_20, n_416, n_283, n_50, n_187, n_525, n_367, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_443, n_57, n_424, n_528, n_387, n_406, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_466, n_346, n_214, n_348, n_2, n_462, n_32, n_410, n_379, n_445, n_515, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_441, n_385, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_23, n_399, n_520, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_473, n_186, n_202, n_145, n_193, n_500, n_59, n_336, n_315, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_339, n_487, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_446, n_143, n_152, n_405, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_401, n_485, n_267, n_495, n_504, n_483, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_481, n_398, n_62, n_210, n_200, n_529, n_502, n_166, n_253, n_218, n_79, n_3, n_271, n_465, n_486, n_507, n_247, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_420, n_518, n_439, n_222, n_478, n_510, n_256, n_326, n_227, n_48, n_188, n_323, n_330, n_400, n_11, n_129, n_126, n_282, n_328, n_368, n_277, n_248, n_301, n_467, n_432, n_293, n_228, n_325, n_276, n_93, n_427, n_108, n_497, n_303, n_442, n_168, n_81, n_1, n_206, n_352, n_511, n_238, n_365, n_429, n_455, n_136, n_334, n_192, n_488, n_300, n_505, n_14, n_163, n_88, n_141, n_390, n_498, n_104, n_501, n_438, n_314, n_16, n_440, n_273, n_305, n_312, n_233, n_56, n_60, n_388, n_333, n_449, n_413, n_392, n_376, n_512, n_459, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_237, n_175, n_453, n_74, n_491, n_19, n_40, n_181, n_53, n_260, n_362, n_310, n_236, n_281, n_24, n_7, n_461, n_209, n_262, n_490, n_17, n_225, n_235, n_464, n_297, n_503, n_290, n_527, n_46, n_84, n_371, n_199, n_107, n_217, n_452, n_178, n_42, n_308, n_417, n_201, n_70, n_343, n_10, n_414, n_287, n_302, n_380, n_6, n_94, n_284, n_4, n_448, n_249, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_278, n_255, n_450, n_257, n_148, n_451, n_475, n_135, n_409, n_171, n_519, n_384, n_468, n_61, n_526, n_102, n_182, n_482, n_316, n_196, n_125, n_43, n_407, n_13, n_27, n_254, n_476, n_460, n_219, n_55, n_231, n_366, n_234, n_492, n_280, n_215, n_252, n_161, n_454, n_298, n_68, n_415, n_78, n_63, n_99, n_216, n_5, n_514, n_418, n_223, n_403, n_25, n_83, n_389, n_513, n_288, n_179, n_395, n_195, n_213, n_110, n_304, n_67, n_509, n_306, n_313, n_92, n_430, n_493, n_203, n_378, n_436, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_337, n_437, n_111, n_21, n_274, n_472, n_296, n_265, n_208, n_456, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_521, n_51, n_496, n_76, n_342, n_26, n_246, n_517, n_0, n_428, n_159, n_358, n_105, n_30, n_494, n_131, n_263, n_434, n_360, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_523, n_268, n_266, n_470, n_457, n_164, n_157, n_184, n_177, n_477, n_364, n_258, n_425, n_431, n_508, n_118, n_121, n_411, n_484, n_353, n_22, n_241, n_29, n_357, n_412, n_447, n_191, n_382, n_489, n_80, n_480, n_211, n_97, n_408, n_322, n_251, n_506, n_116, n_397, n_471, n_351, n_39, n_393, n_474, n_359, n_155, n_127, n_1996);

input n_295;
input n_356;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_332;
input n_294;
input n_197;
input n_463;
input n_176;
input n_34;
input n_404;
input n_172;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_373;
input n_299;
input n_499;
input n_12;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_522;
input n_319;
input n_49;
input n_20;
input n_416;
input n_283;
input n_50;
input n_187;
input n_525;
input n_367;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_443;
input n_57;
input n_424;
input n_528;
input n_387;
input n_406;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_466;
input n_346;
input n_214;
input n_348;
input n_2;
input n_462;
input n_32;
input n_410;
input n_379;
input n_445;
input n_515;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_385;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_23;
input n_399;
input n_520;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_202;
input n_145;
input n_193;
input n_500;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_487;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_446;
input n_143;
input n_152;
input n_405;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_481;
input n_398;
input n_62;
input n_210;
input n_200;
input n_529;
input n_502;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_247;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_420;
input n_518;
input n_439;
input n_222;
input n_478;
input n_510;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_330;
input n_400;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_427;
input n_108;
input n_497;
input n_303;
input n_442;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_511;
input n_238;
input n_365;
input n_429;
input n_455;
input n_136;
input n_334;
input n_192;
input n_488;
input n_300;
input n_505;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_16;
input n_440;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_449;
input n_413;
input n_392;
input n_376;
input n_512;
input n_459;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_237;
input n_175;
input n_453;
input n_74;
input n_491;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_362;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_461;
input n_209;
input n_262;
input n_490;
input n_17;
input n_225;
input n_235;
input n_464;
input n_297;
input n_503;
input n_290;
input n_527;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_452;
input n_178;
input n_42;
input n_308;
input n_417;
input n_201;
input n_70;
input n_343;
input n_10;
input n_414;
input n_287;
input n_302;
input n_380;
input n_6;
input n_94;
input n_284;
input n_4;
input n_448;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_278;
input n_255;
input n_450;
input n_257;
input n_148;
input n_451;
input n_475;
input n_135;
input n_409;
input n_171;
input n_519;
input n_384;
input n_468;
input n_61;
input n_526;
input n_102;
input n_182;
input n_482;
input n_316;
input n_196;
input n_125;
input n_43;
input n_407;
input n_13;
input n_27;
input n_254;
input n_476;
input n_460;
input n_219;
input n_55;
input n_231;
input n_366;
input n_234;
input n_492;
input n_280;
input n_215;
input n_252;
input n_161;
input n_454;
input n_298;
input n_68;
input n_415;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_514;
input n_418;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_513;
input n_288;
input n_179;
input n_395;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_509;
input n_306;
input n_313;
input n_92;
input n_430;
input n_493;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_472;
input n_296;
input n_265;
input n_208;
input n_456;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_521;
input n_51;
input n_496;
input n_76;
input n_342;
input n_26;
input n_246;
input n_517;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_30;
input n_494;
input n_131;
input n_263;
input n_434;
input n_360;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_523;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_425;
input n_431;
input n_508;
input n_118;
input n_121;
input n_411;
input n_484;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_447;
input n_191;
input n_382;
input n_489;
input n_80;
input n_480;
input n_211;
input n_97;
input n_408;
input n_322;
input n_251;
input n_506;
input n_116;
input n_397;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_359;
input n_155;
input n_127;

output n_1996;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_1383;
wire n_603;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_1713;
wire n_1436;
wire n_690;
wire n_1109;
wire n_1430;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_1853;
wire n_764;
wire n_1503;
wire n_1196;
wire n_1181;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_1682;
wire n_1836;
wire n_870;
wire n_1453;
wire n_958;
wire n_945;
wire n_813;
wire n_1985;
wire n_995;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_1979;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_1944;
wire n_559;
wire n_1988;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_1636;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_1254;
wire n_929;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_661;
wire n_1751;
wire n_533;
wire n_1917;
wire n_1924;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_1396;
wire n_1230;
wire n_612;
wire n_1840;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_942;
wire n_1437;
wire n_1378;
wire n_1121;
wire n_1416;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_1716;
wire n_1872;
wire n_1585;
wire n_1432;
wire n_1108;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_652;
wire n_1819;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_696;
wire n_1442;
wire n_798;
wire n_577;
wire n_1833;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_1555;
wire n_1842;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_1376;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_815;
wire n_542;
wire n_1340;
wire n_1240;
wire n_1087;
wire n_632;
wire n_650;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_974;
wire n_1731;
wire n_799;
wire n_1147;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_698;
wire n_1674;
wire n_1992;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_1913;
wire n_1058;
wire n_1042;
wire n_1234;
wire n_1578;
wire n_1455;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_1237;
wire n_927;
wire n_1095;
wire n_1728;
wire n_706;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_1263;
wire n_1817;
wire n_552;
wire n_670;
wire n_1826;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_1611;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_1423;
wire n_600;
wire n_1609;
wire n_1053;
wire n_1939;
wire n_1906;
wire n_1899;
wire n_1467;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_677;
wire n_604;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_681;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_699;
wire n_590;
wire n_727;
wire n_1726;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_1098;
wire n_1490;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_1156;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_957;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_1859;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_1005;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_1708;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_1741;
wire n_745;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_1854;
wire n_666;
wire n_1747;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_1950;
wire n_805;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_1596;
wire n_1281;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_1476;
wire n_1733;
wire n_1856;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_1133;
wire n_883;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1288;
wire n_1201;
wire n_858;
wire n_1185;
wire n_1035;
wire n_1143;
wire n_1090;
wire n_1367;
wire n_928;
wire n_1153;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_1291;
wire n_562;
wire n_748;
wire n_1045;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_914;
wire n_689;
wire n_1116;
wire n_1958;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_728;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_673;
wire n_1038;
wire n_1978;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_1166;
wire n_1056;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_1986;
wire n_540;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_621;
wire n_1587;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_975;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_581;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1926;
wire n_1458;
wire n_679;
wire n_1630;
wire n_663;
wire n_1720;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_1358;
wire n_1200;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_1268;
wire n_917;
wire n_1271;
wire n_1530;
wire n_631;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_1813;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_784;
wire n_648;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_1344;
wire n_1390;
wire n_1792;
wire n_1141;
wire n_1629;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_1152;
wire n_1845;
wire n_1934;
wire n_921;
wire n_1615;
wire n_1236;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_904;
wire n_1696;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_1136;
wire n_1782;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_1964;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_1982;
wire n_662;
wire n_641;
wire n_910;
wire n_741;
wire n_939;
wire n_1410;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_1223;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_1347;
wire n_860;
wire n_1043;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_656;
wire n_574;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_1967;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_626;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_937;
wire n_1474;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_1827;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_1102;
wire n_1129;
wire n_1252;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_718;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_548;
wire n_1662;
wire n_1299;
wire n_1870;
wire n_1925;
wire n_782;
wire n_1861;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_849;
wire n_1820;
wire n_1251;
wire n_1989;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g530 ( 
.A(n_386),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g531 ( 
.A(n_126),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_274),
.Y(n_532)
);

CKINVDCx16_ASAP7_75t_R g533 ( 
.A(n_508),
.Y(n_533)
);

HB1xp67_ASAP7_75t_L g534 ( 
.A(n_252),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_26),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_400),
.Y(n_536)
);

CKINVDCx14_ASAP7_75t_R g537 ( 
.A(n_116),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_418),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_115),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_507),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_43),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_505),
.Y(n_542)
);

CKINVDCx16_ASAP7_75t_R g543 ( 
.A(n_61),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_266),
.Y(n_544)
);

INVx3_ASAP7_75t_L g545 ( 
.A(n_411),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_24),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_36),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_529),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_122),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_221),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_213),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_2),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g553 ( 
.A(n_216),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_181),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_443),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_430),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_425),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_256),
.Y(n_558)
);

BUFx3_ASAP7_75t_L g559 ( 
.A(n_217),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_414),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_506),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_427),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_376),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_52),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_390),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_218),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_150),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_52),
.Y(n_568)
);

INVx2_ASAP7_75t_SL g569 ( 
.A(n_304),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_4),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_367),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_204),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_59),
.Y(n_573)
);

BUFx2_ASAP7_75t_L g574 ( 
.A(n_120),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_500),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_463),
.Y(n_576)
);

INVx1_ASAP7_75t_SL g577 ( 
.A(n_306),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_51),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_488),
.Y(n_579)
);

CKINVDCx20_ASAP7_75t_R g580 ( 
.A(n_118),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_114),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_155),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_421),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_358),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_75),
.Y(n_585)
);

INVx1_ASAP7_75t_SL g586 ( 
.A(n_496),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_17),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_146),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_334),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_3),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_422),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_167),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_32),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_54),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_33),
.Y(n_595)
);

CKINVDCx16_ASAP7_75t_R g596 ( 
.A(n_272),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_244),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_242),
.Y(n_598)
);

CKINVDCx20_ASAP7_75t_R g599 ( 
.A(n_499),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_471),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_325),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_113),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_497),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_373),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_392),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_313),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_490),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_523),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_383),
.Y(n_609)
);

INVx2_ASAP7_75t_SL g610 ( 
.A(n_145),
.Y(n_610)
);

INVx1_ASAP7_75t_SL g611 ( 
.A(n_175),
.Y(n_611)
);

CKINVDCx20_ASAP7_75t_R g612 ( 
.A(n_72),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_176),
.Y(n_613)
);

HB1xp67_ASAP7_75t_L g614 ( 
.A(n_128),
.Y(n_614)
);

BUFx3_ASAP7_75t_L g615 ( 
.A(n_245),
.Y(n_615)
);

BUFx2_ASAP7_75t_SL g616 ( 
.A(n_270),
.Y(n_616)
);

BUFx2_ASAP7_75t_L g617 ( 
.A(n_30),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_501),
.Y(n_618)
);

BUFx3_ASAP7_75t_L g619 ( 
.A(n_492),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_290),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_479),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_407),
.Y(n_622)
);

INVx2_ASAP7_75t_SL g623 ( 
.A(n_103),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_83),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_101),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_89),
.Y(n_626)
);

INVxp33_ASAP7_75t_SL g627 ( 
.A(n_76),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_509),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_447),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_189),
.Y(n_630)
);

INVx1_ASAP7_75t_SL g631 ( 
.A(n_108),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_341),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_444),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_377),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_472),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_184),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_161),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_3),
.Y(n_638)
);

INVx1_ASAP7_75t_SL g639 ( 
.A(n_45),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_97),
.Y(n_640)
);

CKINVDCx16_ASAP7_75t_R g641 ( 
.A(n_279),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_322),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_516),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_434),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_435),
.Y(n_645)
);

CKINVDCx20_ASAP7_75t_R g646 ( 
.A(n_210),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_95),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_140),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_185),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_247),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_303),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_267),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_502),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_503),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_522),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_504),
.Y(n_656)
);

BUFx10_ASAP7_75t_L g657 ( 
.A(n_261),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_259),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_23),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_10),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_283),
.Y(n_661)
);

HB1xp67_ASAP7_75t_L g662 ( 
.A(n_498),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_450),
.Y(n_663)
);

CKINVDCx20_ASAP7_75t_R g664 ( 
.A(n_342),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_65),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_483),
.Y(n_666)
);

CKINVDCx20_ASAP7_75t_R g667 ( 
.A(n_149),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_375),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_520),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_188),
.Y(n_670)
);

BUFx3_ASAP7_75t_L g671 ( 
.A(n_125),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_310),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_81),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_494),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_200),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_475),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_405),
.Y(n_677)
);

BUFx10_ASAP7_75t_L g678 ( 
.A(n_453),
.Y(n_678)
);

CKINVDCx20_ASAP7_75t_R g679 ( 
.A(n_464),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_289),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_307),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_37),
.Y(n_682)
);

INVx1_ASAP7_75t_SL g683 ( 
.A(n_339),
.Y(n_683)
);

CKINVDCx20_ASAP7_75t_R g684 ( 
.A(n_456),
.Y(n_684)
);

HB1xp67_ASAP7_75t_L g685 ( 
.A(n_461),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_297),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_59),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_321),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_315),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_495),
.Y(n_690)
);

INVx1_ASAP7_75t_SL g691 ( 
.A(n_198),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_402),
.Y(n_692)
);

CKINVDCx20_ASAP7_75t_R g693 ( 
.A(n_351),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_282),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_203),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_38),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_243),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_513),
.Y(n_698)
);

CKINVDCx20_ASAP7_75t_R g699 ( 
.A(n_246),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_378),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_417),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_333),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_151),
.Y(n_703)
);

CKINVDCx20_ASAP7_75t_R g704 ( 
.A(n_44),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_546),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_578),
.Y(n_706)
);

HB1xp67_ASAP7_75t_L g707 ( 
.A(n_617),
.Y(n_707)
);

HB1xp67_ASAP7_75t_L g708 ( 
.A(n_543),
.Y(n_708)
);

CKINVDCx16_ASAP7_75t_R g709 ( 
.A(n_533),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_587),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_595),
.Y(n_711)
);

INVxp33_ASAP7_75t_SL g712 ( 
.A(n_535),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_624),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_660),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_665),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_531),
.Y(n_716)
);

INVxp67_ASAP7_75t_SL g717 ( 
.A(n_696),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_570),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_534),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_614),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_559),
.Y(n_721)
);

CKINVDCx16_ASAP7_75t_R g722 ( 
.A(n_596),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_662),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_685),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_574),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_657),
.Y(n_726)
);

INVxp67_ASAP7_75t_L g727 ( 
.A(n_547),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_657),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_678),
.Y(n_729)
);

BUFx3_ASAP7_75t_L g730 ( 
.A(n_678),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_530),
.Y(n_731)
);

INVxp67_ASAP7_75t_SL g732 ( 
.A(n_627),
.Y(n_732)
);

OR2x2_ASAP7_75t_L g733 ( 
.A(n_639),
.B(n_0),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_536),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_559),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_538),
.Y(n_736)
);

INVxp33_ASAP7_75t_SL g737 ( 
.A(n_552),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_540),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_544),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_548),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_549),
.Y(n_741)
);

HB1xp67_ASAP7_75t_L g742 ( 
.A(n_564),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_554),
.Y(n_743)
);

CKINVDCx20_ASAP7_75t_R g744 ( 
.A(n_553),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_615),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_615),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_556),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_558),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_580),
.Y(n_749)
);

CKINVDCx20_ASAP7_75t_R g750 ( 
.A(n_599),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_575),
.Y(n_751)
);

HB1xp67_ASAP7_75t_L g752 ( 
.A(n_568),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_646),
.Y(n_753)
);

BUFx3_ASAP7_75t_L g754 ( 
.A(n_619),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_664),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_576),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_589),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_606),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_608),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_613),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_667),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_618),
.Y(n_762)
);

CKINVDCx20_ASAP7_75t_R g763 ( 
.A(n_679),
.Y(n_763)
);

CKINVDCx20_ASAP7_75t_R g764 ( 
.A(n_684),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_635),
.Y(n_765)
);

CKINVDCx16_ASAP7_75t_R g766 ( 
.A(n_641),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_654),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_693),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_661),
.Y(n_769)
);

BUFx3_ASAP7_75t_L g770 ( 
.A(n_619),
.Y(n_770)
);

CKINVDCx14_ASAP7_75t_R g771 ( 
.A(n_537),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_669),
.Y(n_772)
);

BUFx2_ASAP7_75t_SL g773 ( 
.A(n_699),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_670),
.Y(n_774)
);

INVxp33_ASAP7_75t_SL g775 ( 
.A(n_573),
.Y(n_775)
);

INVxp33_ASAP7_75t_L g776 ( 
.A(n_598),
.Y(n_776)
);

INVxp67_ASAP7_75t_SL g777 ( 
.A(n_545),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_545),
.B(n_0),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_674),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_585),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_675),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_677),
.Y(n_782)
);

HB1xp67_ASAP7_75t_L g783 ( 
.A(n_590),
.Y(n_783)
);

CKINVDCx16_ASAP7_75t_R g784 ( 
.A(n_541),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_680),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_689),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_593),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_697),
.Y(n_788)
);

CKINVDCx20_ASAP7_75t_R g789 ( 
.A(n_612),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_594),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_700),
.B(n_701),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_671),
.Y(n_792)
);

BUFx3_ASAP7_75t_L g793 ( 
.A(n_671),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_626),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_638),
.Y(n_795)
);

BUFx2_ASAP7_75t_L g796 ( 
.A(n_659),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_673),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_682),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_687),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_598),
.Y(n_800)
);

CKINVDCx16_ASAP7_75t_R g801 ( 
.A(n_704),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_605),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_605),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_625),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_625),
.Y(n_805)
);

BUFx6f_ASAP7_75t_L g806 ( 
.A(n_754),
.Y(n_806)
);

BUFx2_ASAP7_75t_L g807 ( 
.A(n_708),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_705),
.Y(n_808)
);

BUFx6f_ASAP7_75t_L g809 ( 
.A(n_770),
.Y(n_809)
);

BUFx6f_ASAP7_75t_L g810 ( 
.A(n_793),
.Y(n_810)
);

INVx4_ASAP7_75t_L g811 ( 
.A(n_730),
.Y(n_811)
);

BUFx6f_ASAP7_75t_L g812 ( 
.A(n_718),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_800),
.Y(n_813)
);

AND2x4_ASAP7_75t_L g814 ( 
.A(n_726),
.B(n_569),
.Y(n_814)
);

AND2x4_ASAP7_75t_L g815 ( 
.A(n_728),
.B(n_610),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_721),
.Y(n_816)
);

INVx4_ASAP7_75t_L g817 ( 
.A(n_780),
.Y(n_817)
);

BUFx6f_ASAP7_75t_L g818 ( 
.A(n_735),
.Y(n_818)
);

BUFx6f_ASAP7_75t_L g819 ( 
.A(n_745),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_802),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_803),
.Y(n_821)
);

OAI21x1_ASAP7_75t_L g822 ( 
.A1(n_791),
.A2(n_734),
.B(n_731),
.Y(n_822)
);

OAI21x1_ASAP7_75t_L g823 ( 
.A1(n_736),
.A2(n_663),
.B(n_607),
.Y(n_823)
);

BUFx6f_ASAP7_75t_L g824 ( 
.A(n_746),
.Y(n_824)
);

INVx5_ASAP7_75t_L g825 ( 
.A(n_792),
.Y(n_825)
);

AOI22xp5_ASAP7_75t_L g826 ( 
.A1(n_732),
.A2(n_586),
.B1(n_611),
.B2(n_577),
.Y(n_826)
);

BUFx3_ASAP7_75t_L g827 ( 
.A(n_738),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_771),
.B(n_631),
.Y(n_828)
);

XNOR2x2_ASAP7_75t_L g829 ( 
.A(n_789),
.B(n_683),
.Y(n_829)
);

BUFx6f_ASAP7_75t_L g830 ( 
.A(n_706),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_804),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_710),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_771),
.B(n_691),
.Y(n_833)
);

BUFx6f_ASAP7_75t_L g834 ( 
.A(n_711),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_713),
.Y(n_835)
);

BUFx6f_ASAP7_75t_L g836 ( 
.A(n_714),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_776),
.B(n_616),
.Y(n_837)
);

OA21x2_ASAP7_75t_L g838 ( 
.A1(n_805),
.A2(n_778),
.B(n_740),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_715),
.Y(n_839)
);

AND2x4_ASAP7_75t_L g840 ( 
.A(n_729),
.B(n_623),
.Y(n_840)
);

HB1xp67_ASAP7_75t_L g841 ( 
.A(n_708),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_739),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_741),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_743),
.Y(n_844)
);

BUFx12f_ASAP7_75t_L g845 ( 
.A(n_716),
.Y(n_845)
);

INVx4_ASAP7_75t_L g846 ( 
.A(n_787),
.Y(n_846)
);

AND2x6_ASAP7_75t_L g847 ( 
.A(n_778),
.B(n_663),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_747),
.Y(n_848)
);

BUFx6f_ASAP7_75t_L g849 ( 
.A(n_748),
.Y(n_849)
);

CKINVDCx20_ASAP7_75t_R g850 ( 
.A(n_744),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_751),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_756),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_SL g853 ( 
.A(n_709),
.B(n_532),
.Y(n_853)
);

AND2x2_ASAP7_75t_L g854 ( 
.A(n_776),
.B(n_539),
.Y(n_854)
);

AOI22xp5_ASAP7_75t_L g855 ( 
.A1(n_732),
.A2(n_550),
.B1(n_551),
.B2(n_542),
.Y(n_855)
);

OAI22x1_ASAP7_75t_R g856 ( 
.A1(n_784),
.A2(n_560),
.B1(n_561),
.B2(n_555),
.Y(n_856)
);

CKINVDCx11_ASAP7_75t_R g857 ( 
.A(n_750),
.Y(n_857)
);

INVx2_ASAP7_75t_SL g858 ( 
.A(n_790),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_757),
.Y(n_859)
);

BUFx6f_ASAP7_75t_L g860 ( 
.A(n_758),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_759),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_760),
.Y(n_862)
);

NOR2x1_ASAP7_75t_L g863 ( 
.A(n_794),
.B(n_557),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_762),
.Y(n_864)
);

OAI22xp5_ASAP7_75t_L g865 ( 
.A1(n_707),
.A2(n_562),
.B1(n_565),
.B2(n_563),
.Y(n_865)
);

BUFx8_ASAP7_75t_L g866 ( 
.A(n_796),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_765),
.Y(n_867)
);

INVx4_ASAP7_75t_L g868 ( 
.A(n_799),
.Y(n_868)
);

BUFx2_ASAP7_75t_L g869 ( 
.A(n_742),
.Y(n_869)
);

INVx6_ASAP7_75t_L g870 ( 
.A(n_722),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_767),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_769),
.Y(n_872)
);

OAI22xp5_ASAP7_75t_L g873 ( 
.A1(n_707),
.A2(n_566),
.B1(n_571),
.B2(n_567),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_772),
.Y(n_874)
);

AND2x4_ASAP7_75t_L g875 ( 
.A(n_725),
.B(n_557),
.Y(n_875)
);

BUFx3_ASAP7_75t_L g876 ( 
.A(n_774),
.Y(n_876)
);

AND2x4_ASAP7_75t_L g877 ( 
.A(n_727),
.B(n_557),
.Y(n_877)
);

HB1xp67_ASAP7_75t_L g878 ( 
.A(n_742),
.Y(n_878)
);

AND2x4_ASAP7_75t_L g879 ( 
.A(n_727),
.B(n_557),
.Y(n_879)
);

AND2x4_ASAP7_75t_L g880 ( 
.A(n_719),
.B(n_572),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_779),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_781),
.Y(n_882)
);

BUFx6f_ASAP7_75t_L g883 ( 
.A(n_782),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_785),
.Y(n_884)
);

OA21x2_ASAP7_75t_L g885 ( 
.A1(n_786),
.A2(n_581),
.B(n_579),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_777),
.B(n_582),
.Y(n_886)
);

OAI22x1_ASAP7_75t_SL g887 ( 
.A1(n_763),
.A2(n_584),
.B1(n_588),
.B2(n_583),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_788),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_777),
.B(n_591),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_717),
.Y(n_890)
);

AND2x4_ASAP7_75t_L g891 ( 
.A(n_720),
.B(n_592),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_818),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_818),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_822),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_855),
.B(n_766),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_839),
.Y(n_896)
);

INVx3_ASAP7_75t_L g897 ( 
.A(n_849),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_837),
.B(n_795),
.Y(n_898)
);

INVx3_ASAP7_75t_L g899 ( 
.A(n_849),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_819),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_816),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_852),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_852),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_819),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_859),
.Y(n_905)
);

AND2x4_ASAP7_75t_L g906 ( 
.A(n_877),
.B(n_723),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_859),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_824),
.Y(n_908)
);

BUFx3_ASAP7_75t_L g909 ( 
.A(n_806),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_861),
.Y(n_910)
);

INVxp67_ASAP7_75t_L g911 ( 
.A(n_869),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_854),
.B(n_797),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_824),
.Y(n_913)
);

BUFx6f_ASAP7_75t_L g914 ( 
.A(n_812),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_861),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_812),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_862),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_862),
.Y(n_918)
);

CKINVDCx16_ASAP7_75t_R g919 ( 
.A(n_845),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_857),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_864),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_813),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_813),
.Y(n_923)
);

AND2x6_ASAP7_75t_L g924 ( 
.A(n_828),
.B(n_724),
.Y(n_924)
);

NAND2xp33_ASAP7_75t_SL g925 ( 
.A(n_858),
.B(n_733),
.Y(n_925)
);

BUFx6f_ASAP7_75t_L g926 ( 
.A(n_830),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_847),
.B(n_798),
.Y(n_927)
);

BUFx6f_ASAP7_75t_L g928 ( 
.A(n_830),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_864),
.Y(n_929)
);

OAI22xp5_ASAP7_75t_SL g930 ( 
.A1(n_850),
.A2(n_764),
.B1(n_801),
.B2(n_753),
.Y(n_930)
);

BUFx6f_ASAP7_75t_L g931 ( 
.A(n_834),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_820),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_881),
.Y(n_933)
);

HB1xp67_ASAP7_75t_L g934 ( 
.A(n_807),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_881),
.Y(n_935)
);

INVx3_ASAP7_75t_L g936 ( 
.A(n_860),
.Y(n_936)
);

BUFx6f_ASAP7_75t_L g937 ( 
.A(n_834),
.Y(n_937)
);

INVx3_ASAP7_75t_L g938 ( 
.A(n_860),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_838),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_847),
.B(n_712),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_847),
.B(n_737),
.Y(n_941)
);

HB1xp67_ASAP7_75t_L g942 ( 
.A(n_807),
.Y(n_942)
);

CKINVDCx20_ASAP7_75t_R g943 ( 
.A(n_870),
.Y(n_943)
);

INVx3_ASAP7_75t_L g944 ( 
.A(n_883),
.Y(n_944)
);

INVx3_ASAP7_75t_L g945 ( 
.A(n_883),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_808),
.Y(n_946)
);

HB1xp67_ASAP7_75t_L g947 ( 
.A(n_869),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_886),
.B(n_775),
.Y(n_948)
);

BUFx6f_ASAP7_75t_L g949 ( 
.A(n_836),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_832),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_820),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_889),
.B(n_783),
.Y(n_952)
);

BUFx6f_ASAP7_75t_L g953 ( 
.A(n_836),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_835),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_821),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_878),
.B(n_752),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_879),
.B(n_783),
.Y(n_957)
);

BUFx2_ASAP7_75t_L g958 ( 
.A(n_866),
.Y(n_958)
);

INVx1_ASAP7_75t_SL g959 ( 
.A(n_870),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_821),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_871),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_817),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_838),
.Y(n_963)
);

BUFx6f_ASAP7_75t_L g964 ( 
.A(n_823),
.Y(n_964)
);

HB1xp67_ASAP7_75t_L g965 ( 
.A(n_841),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_872),
.Y(n_966)
);

NAND2xp33_ASAP7_75t_SL g967 ( 
.A(n_846),
.B(n_752),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_831),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_842),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_831),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_843),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_844),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_848),
.Y(n_973)
);

BUFx6f_ASAP7_75t_L g974 ( 
.A(n_806),
.Y(n_974)
);

OA21x2_ASAP7_75t_L g975 ( 
.A1(n_851),
.A2(n_717),
.B(n_600),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_867),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_874),
.Y(n_977)
);

INVx3_ASAP7_75t_L g978 ( 
.A(n_882),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_884),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_888),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_827),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_890),
.B(n_597),
.Y(n_982)
);

INVx3_ASAP7_75t_L g983 ( 
.A(n_876),
.Y(n_983)
);

BUFx6f_ASAP7_75t_L g984 ( 
.A(n_809),
.Y(n_984)
);

AND2x4_ASAP7_75t_L g985 ( 
.A(n_959),
.B(n_868),
.Y(n_985)
);

AOI22xp33_ASAP7_75t_L g986 ( 
.A1(n_924),
.A2(n_885),
.B1(n_826),
.B2(n_773),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_948),
.B(n_833),
.Y(n_987)
);

BUFx6f_ASAP7_75t_L g988 ( 
.A(n_974),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_940),
.B(n_749),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_978),
.Y(n_990)
);

INVx5_ASAP7_75t_L g991 ( 
.A(n_926),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_L g992 ( 
.A(n_941),
.B(n_755),
.Y(n_992)
);

BUFx3_ASAP7_75t_L g993 ( 
.A(n_943),
.Y(n_993)
);

AND2x4_ASAP7_75t_L g994 ( 
.A(n_983),
.B(n_809),
.Y(n_994)
);

INVx3_ASAP7_75t_L g995 ( 
.A(n_974),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_978),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_902),
.Y(n_997)
);

AND2x2_ASAP7_75t_L g998 ( 
.A(n_911),
.B(n_761),
.Y(n_998)
);

AOI22xp33_ASAP7_75t_L g999 ( 
.A1(n_924),
.A2(n_885),
.B1(n_875),
.B2(n_880),
.Y(n_999)
);

INVx3_ASAP7_75t_L g1000 ( 
.A(n_974),
.Y(n_1000)
);

INVx3_ASAP7_75t_L g1001 ( 
.A(n_984),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_898),
.B(n_891),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_903),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_SL g1004 ( 
.A(n_962),
.B(n_853),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_983),
.B(n_865),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_976),
.Y(n_1006)
);

AOI22xp33_ASAP7_75t_L g1007 ( 
.A1(n_924),
.A2(n_814),
.B1(n_840),
.B2(n_815),
.Y(n_1007)
);

BUFx6f_ASAP7_75t_L g1008 ( 
.A(n_984),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_912),
.B(n_863),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_905),
.Y(n_1010)
);

NOR2xp33_ASAP7_75t_L g1011 ( 
.A(n_952),
.B(n_768),
.Y(n_1011)
);

BUFx3_ASAP7_75t_L g1012 ( 
.A(n_909),
.Y(n_1012)
);

OR2x6_ASAP7_75t_L g1013 ( 
.A(n_958),
.B(n_810),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_920),
.Y(n_1014)
);

OR2x6_ASAP7_75t_L g1015 ( 
.A(n_930),
.B(n_810),
.Y(n_1015)
);

INVx4_ASAP7_75t_L g1016 ( 
.A(n_984),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_956),
.B(n_811),
.Y(n_1017)
);

AND2x4_ASAP7_75t_L g1018 ( 
.A(n_897),
.B(n_899),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_919),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_934),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_907),
.B(n_873),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_910),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_915),
.Y(n_1023)
);

HB1xp67_ASAP7_75t_L g1024 ( 
.A(n_942),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_977),
.Y(n_1025)
);

INVx2_ASAP7_75t_SL g1026 ( 
.A(n_947),
.Y(n_1026)
);

AOI22xp33_ASAP7_75t_L g1027 ( 
.A1(n_924),
.A2(n_829),
.B1(n_825),
.B2(n_602),
.Y(n_1027)
);

INVx2_ASAP7_75t_SL g1028 ( 
.A(n_965),
.Y(n_1028)
);

AOI22xp5_ASAP7_75t_L g1029 ( 
.A1(n_927),
.A2(n_887),
.B1(n_603),
.B2(n_604),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_925),
.B(n_825),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_917),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_918),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_922),
.Y(n_1033)
);

BUFx10_ASAP7_75t_L g1034 ( 
.A(n_906),
.Y(n_1034)
);

INVx4_ASAP7_75t_L g1035 ( 
.A(n_926),
.Y(n_1035)
);

INVx3_ASAP7_75t_L g1036 ( 
.A(n_914),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_921),
.Y(n_1037)
);

INVx4_ASAP7_75t_SL g1038 ( 
.A(n_906),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_923),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_SL g1040 ( 
.A(n_926),
.B(n_825),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_929),
.Y(n_1041)
);

BUFx10_ASAP7_75t_L g1042 ( 
.A(n_946),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_L g1043 ( 
.A(n_895),
.B(n_601),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_932),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_951),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_955),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_933),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_935),
.Y(n_1048)
);

INVx4_ASAP7_75t_L g1049 ( 
.A(n_928),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_950),
.B(n_609),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_954),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_SL g1052 ( 
.A(n_928),
.B(n_620),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_961),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_966),
.B(n_621),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_960),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_968),
.Y(n_1056)
);

AOI22xp33_ASAP7_75t_L g1057 ( 
.A1(n_939),
.A2(n_628),
.B1(n_629),
.B2(n_622),
.Y(n_1057)
);

INVx3_ASAP7_75t_R g1058 ( 
.A(n_892),
.Y(n_1058)
);

AND2x2_ASAP7_75t_L g1059 ( 
.A(n_957),
.B(n_856),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_970),
.Y(n_1060)
);

OR2x2_ASAP7_75t_L g1061 ( 
.A(n_981),
.B(n_1),
.Y(n_1061)
);

AND2x4_ASAP7_75t_L g1062 ( 
.A(n_897),
.B(n_1),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_SL g1063 ( 
.A(n_928),
.B(n_931),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_899),
.B(n_2),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_901),
.Y(n_1065)
);

AND2x6_ASAP7_75t_L g1066 ( 
.A(n_939),
.B(n_90),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_896),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_969),
.Y(n_1068)
);

INVxp67_ASAP7_75t_SL g1069 ( 
.A(n_963),
.Y(n_1069)
);

NAND2xp33_ASAP7_75t_R g1070 ( 
.A(n_975),
.B(n_630),
.Y(n_1070)
);

BUFx8_ASAP7_75t_SL g1071 ( 
.A(n_893),
.Y(n_1071)
);

AND2x4_ASAP7_75t_L g1072 ( 
.A(n_936),
.B(n_938),
.Y(n_1072)
);

BUFx6f_ASAP7_75t_L g1073 ( 
.A(n_931),
.Y(n_1073)
);

AOI22xp5_ASAP7_75t_L g1074 ( 
.A1(n_975),
.A2(n_633),
.B1(n_634),
.B2(n_632),
.Y(n_1074)
);

AND2x6_ASAP7_75t_L g1075 ( 
.A(n_963),
.B(n_91),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_971),
.Y(n_1076)
);

INVx5_ASAP7_75t_L g1077 ( 
.A(n_931),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_972),
.Y(n_1078)
);

INVx1_ASAP7_75t_SL g1079 ( 
.A(n_937),
.Y(n_1079)
);

BUFx3_ASAP7_75t_L g1080 ( 
.A(n_937),
.Y(n_1080)
);

NAND2xp33_ASAP7_75t_SL g1081 ( 
.A(n_982),
.B(n_636),
.Y(n_1081)
);

INVx5_ASAP7_75t_L g1082 ( 
.A(n_937),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_973),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_987),
.B(n_979),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_1011),
.B(n_980),
.Y(n_1085)
);

NOR2xp67_ASAP7_75t_L g1086 ( 
.A(n_1014),
.B(n_936),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_SL g1087 ( 
.A(n_985),
.B(n_967),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_SL g1088 ( 
.A(n_985),
.B(n_949),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_1002),
.B(n_938),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_1069),
.A2(n_894),
.B(n_964),
.Y(n_1090)
);

INVx3_ASAP7_75t_L g1091 ( 
.A(n_993),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_SL g1092 ( 
.A(n_1028),
.B(n_998),
.Y(n_1092)
);

INVxp67_ASAP7_75t_L g1093 ( 
.A(n_1024),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_1021),
.B(n_944),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_1051),
.Y(n_1095)
);

NOR2xp33_ASAP7_75t_L g1096 ( 
.A(n_1020),
.B(n_944),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_1006),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_1025),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_989),
.B(n_945),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_992),
.B(n_945),
.Y(n_1100)
);

NAND3xp33_ASAP7_75t_L g1101 ( 
.A(n_1026),
.B(n_953),
.C(n_949),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_997),
.B(n_1003),
.Y(n_1102)
);

AO22x2_ASAP7_75t_L g1103 ( 
.A1(n_1059),
.A2(n_894),
.B1(n_916),
.B2(n_904),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_1010),
.B(n_949),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_1022),
.B(n_953),
.Y(n_1105)
);

A2O1A1Ixp33_ASAP7_75t_L g1106 ( 
.A1(n_1023),
.A2(n_964),
.B(n_908),
.C(n_913),
.Y(n_1106)
);

NOR2xp33_ASAP7_75t_L g1107 ( 
.A(n_1005),
.B(n_953),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1053),
.Y(n_1108)
);

AND2x4_ASAP7_75t_L g1109 ( 
.A(n_1038),
.B(n_900),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_1065),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_1031),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_1032),
.B(n_914),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_1067),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_1037),
.B(n_914),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_1033),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_1041),
.B(n_964),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_L g1117 ( 
.A(n_1004),
.B(n_637),
.Y(n_1117)
);

INVxp67_ASAP7_75t_L g1118 ( 
.A(n_1017),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_1039),
.Y(n_1119)
);

NOR2xp33_ASAP7_75t_L g1120 ( 
.A(n_1009),
.B(n_703),
.Y(n_1120)
);

NOR2xp67_ASAP7_75t_L g1121 ( 
.A(n_1019),
.B(n_640),
.Y(n_1121)
);

NOR2xp33_ASAP7_75t_L g1122 ( 
.A(n_1079),
.B(n_702),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_1047),
.B(n_642),
.Y(n_1123)
);

OAI22xp33_ASAP7_75t_L g1124 ( 
.A1(n_1061),
.A2(n_644),
.B1(n_645),
.B2(n_643),
.Y(n_1124)
);

INVx3_ASAP7_75t_L g1125 ( 
.A(n_1073),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1048),
.Y(n_1126)
);

BUFx3_ASAP7_75t_L g1127 ( 
.A(n_1012),
.Y(n_1127)
);

BUFx10_ASAP7_75t_L g1128 ( 
.A(n_994),
.Y(n_1128)
);

NAND3xp33_ASAP7_75t_L g1129 ( 
.A(n_1057),
.B(n_648),
.C(n_647),
.Y(n_1129)
);

NAND2xp33_ASAP7_75t_L g1130 ( 
.A(n_1066),
.B(n_1075),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_1044),
.Y(n_1131)
);

NAND2xp33_ASAP7_75t_L g1132 ( 
.A(n_1066),
.B(n_649),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_SL g1133 ( 
.A(n_1042),
.B(n_991),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_1055),
.B(n_650),
.Y(n_1134)
);

NOR2xp33_ASAP7_75t_L g1135 ( 
.A(n_1043),
.B(n_651),
.Y(n_1135)
);

NOR3xp33_ASAP7_75t_L g1136 ( 
.A(n_1050),
.B(n_653),
.C(n_652),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1045),
.B(n_655),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1054),
.A2(n_658),
.B(n_656),
.Y(n_1138)
);

OAI22xp5_ASAP7_75t_L g1139 ( 
.A1(n_999),
.A2(n_668),
.B1(n_672),
.B2(n_666),
.Y(n_1139)
);

INVx4_ASAP7_75t_L g1140 ( 
.A(n_991),
.Y(n_1140)
);

INVxp67_ASAP7_75t_L g1141 ( 
.A(n_994),
.Y(n_1141)
);

AOI22xp5_ASAP7_75t_L g1142 ( 
.A1(n_1074),
.A2(n_698),
.B1(n_681),
.B2(n_686),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_1046),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1056),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1060),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1068),
.B(n_1076),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1078),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_SL g1148 ( 
.A(n_991),
.B(n_676),
.Y(n_1148)
);

NOR2xp33_ASAP7_75t_L g1149 ( 
.A(n_1034),
.B(n_695),
.Y(n_1149)
);

AOI22xp33_ASAP7_75t_SL g1150 ( 
.A1(n_1015),
.A2(n_690),
.B1(n_692),
.B2(n_688),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1083),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_1013),
.Y(n_1152)
);

BUFx6f_ASAP7_75t_L g1153 ( 
.A(n_1073),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_990),
.Y(n_1154)
);

INVx3_ASAP7_75t_L g1155 ( 
.A(n_1013),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_SL g1156 ( 
.A(n_1077),
.B(n_694),
.Y(n_1156)
);

AOI22xp5_ASAP7_75t_L g1157 ( 
.A1(n_1062),
.A2(n_6),
.B1(n_4),
.B2(n_5),
.Y(n_1157)
);

BUFx6f_ASAP7_75t_SL g1158 ( 
.A(n_1015),
.Y(n_1158)
);

AOI22xp5_ASAP7_75t_L g1159 ( 
.A1(n_1062),
.A2(n_7),
.B1(n_5),
.B2(n_6),
.Y(n_1159)
);

AOI22xp33_ASAP7_75t_L g1160 ( 
.A1(n_1027),
.A2(n_9),
.B1(n_7),
.B2(n_8),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_986),
.B(n_996),
.Y(n_1161)
);

AOI22xp5_ASAP7_75t_L g1162 ( 
.A1(n_1070),
.A2(n_10),
.B1(n_8),
.B2(n_9),
.Y(n_1162)
);

NAND3xp33_ASAP7_75t_SL g1163 ( 
.A(n_1135),
.B(n_1029),
.C(n_1007),
.Y(n_1163)
);

INVx5_ASAP7_75t_L g1164 ( 
.A(n_1155),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1100),
.B(n_1038),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1146),
.Y(n_1166)
);

BUFx2_ASAP7_75t_L g1167 ( 
.A(n_1152),
.Y(n_1167)
);

AND2x4_ASAP7_75t_L g1168 ( 
.A(n_1127),
.B(n_1018),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_1110),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1095),
.Y(n_1170)
);

AND3x1_ASAP7_75t_SL g1171 ( 
.A(n_1108),
.B(n_11),
.C(n_12),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1085),
.B(n_1018),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_SL g1173 ( 
.A(n_1150),
.B(n_1077),
.Y(n_1173)
);

BUFx8_ASAP7_75t_L g1174 ( 
.A(n_1158),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1084),
.B(n_1072),
.Y(n_1175)
);

INVx5_ASAP7_75t_L g1176 ( 
.A(n_1128),
.Y(n_1176)
);

BUFx6f_ASAP7_75t_L g1177 ( 
.A(n_1153),
.Y(n_1177)
);

OAI22xp5_ASAP7_75t_SL g1178 ( 
.A1(n_1162),
.A2(n_1058),
.B1(n_1072),
.B2(n_1016),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_1113),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1118),
.B(n_988),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1111),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1102),
.B(n_988),
.Y(n_1182)
);

AND2x2_ASAP7_75t_L g1183 ( 
.A(n_1093),
.B(n_1080),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1089),
.B(n_1008),
.Y(n_1184)
);

OAI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1116),
.A2(n_1064),
.B(n_1081),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1126),
.Y(n_1186)
);

AND3x2_ASAP7_75t_SL g1187 ( 
.A(n_1115),
.B(n_1071),
.C(n_1058),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1147),
.Y(n_1188)
);

AND2x2_ASAP7_75t_L g1189 ( 
.A(n_1096),
.B(n_995),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1094),
.B(n_1008),
.Y(n_1190)
);

AND2x4_ASAP7_75t_L g1191 ( 
.A(n_1109),
.B(n_1077),
.Y(n_1191)
);

INVx3_ASAP7_75t_L g1192 ( 
.A(n_1128),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1151),
.Y(n_1193)
);

NOR2xp67_ASAP7_75t_L g1194 ( 
.A(n_1091),
.B(n_1082),
.Y(n_1194)
);

BUFx3_ASAP7_75t_L g1195 ( 
.A(n_1153),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1120),
.B(n_1036),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_SL g1197 ( 
.A(n_1099),
.B(n_1082),
.Y(n_1197)
);

AOI22x1_ASAP7_75t_L g1198 ( 
.A1(n_1090),
.A2(n_1049),
.B1(n_1035),
.B2(n_1001),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_1119),
.Y(n_1199)
);

AOI22xp33_ASAP7_75t_L g1200 ( 
.A1(n_1131),
.A2(n_1075),
.B1(n_1066),
.B2(n_1052),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1141),
.B(n_1000),
.Y(n_1201)
);

NOR2xp67_ASAP7_75t_L g1202 ( 
.A(n_1101),
.B(n_1082),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_SL g1203 ( 
.A(n_1153),
.B(n_1030),
.Y(n_1203)
);

INVx4_ASAP7_75t_L g1204 ( 
.A(n_1140),
.Y(n_1204)
);

O2A1O1Ixp5_ASAP7_75t_L g1205 ( 
.A1(n_1148),
.A2(n_1063),
.B(n_1040),
.C(n_1075),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_1143),
.Y(n_1206)
);

INVx3_ASAP7_75t_L g1207 ( 
.A(n_1140),
.Y(n_1207)
);

AND2x4_ASAP7_75t_SL g1208 ( 
.A(n_1109),
.B(n_11),
.Y(n_1208)
);

INVx3_ASAP7_75t_L g1209 ( 
.A(n_1125),
.Y(n_1209)
);

HB1xp67_ASAP7_75t_L g1210 ( 
.A(n_1092),
.Y(n_1210)
);

BUFx3_ASAP7_75t_L g1211 ( 
.A(n_1125),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1122),
.B(n_12),
.Y(n_1212)
);

NOR2xp33_ASAP7_75t_L g1213 ( 
.A(n_1087),
.B(n_13),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_1097),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1088),
.B(n_13),
.Y(n_1215)
);

BUFx12f_ASAP7_75t_L g1216 ( 
.A(n_1086),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_1117),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1144),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1145),
.Y(n_1219)
);

INVx5_ASAP7_75t_L g1220 ( 
.A(n_1154),
.Y(n_1220)
);

AOI22xp33_ASAP7_75t_L g1221 ( 
.A1(n_1160),
.A2(n_16),
.B1(n_14),
.B2(n_15),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1098),
.Y(n_1222)
);

BUFx3_ASAP7_75t_L g1223 ( 
.A(n_1149),
.Y(n_1223)
);

AOI22xp33_ASAP7_75t_L g1224 ( 
.A1(n_1161),
.A2(n_16),
.B1(n_14),
.B2(n_15),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1104),
.Y(n_1225)
);

INVx2_ASAP7_75t_SL g1226 ( 
.A(n_1133),
.Y(n_1226)
);

BUFx6f_ASAP7_75t_L g1227 ( 
.A(n_1105),
.Y(n_1227)
);

NOR2xp33_ASAP7_75t_R g1228 ( 
.A(n_1132),
.B(n_92),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_SL g1229 ( 
.A(n_1124),
.B(n_17),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_SL g1230 ( 
.A(n_1121),
.B(n_18),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1107),
.B(n_18),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_SL g1232 ( 
.A(n_1136),
.B(n_19),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1112),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1114),
.B(n_1103),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1103),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_SL g1236 ( 
.A(n_1142),
.B(n_19),
.Y(n_1236)
);

NOR2xp33_ASAP7_75t_L g1237 ( 
.A(n_1123),
.B(n_20),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1134),
.B(n_20),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1137),
.Y(n_1239)
);

INVx6_ASAP7_75t_L g1240 ( 
.A(n_1156),
.Y(n_1240)
);

NOR2xp33_ASAP7_75t_L g1241 ( 
.A(n_1129),
.B(n_21),
.Y(n_1241)
);

NOR2xp33_ASAP7_75t_L g1242 ( 
.A(n_1217),
.B(n_1157),
.Y(n_1242)
);

HB1xp67_ASAP7_75t_L g1243 ( 
.A(n_1183),
.Y(n_1243)
);

O2A1O1Ixp33_ASAP7_75t_L g1244 ( 
.A1(n_1212),
.A2(n_1130),
.B(n_1139),
.C(n_1106),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1166),
.B(n_1159),
.Y(n_1245)
);

AOI22xp33_ASAP7_75t_L g1246 ( 
.A1(n_1163),
.A2(n_1138),
.B1(n_23),
.B2(n_21),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1170),
.Y(n_1247)
);

INVx4_ASAP7_75t_L g1248 ( 
.A(n_1177),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_1169),
.Y(n_1249)
);

AND2x2_ASAP7_75t_L g1250 ( 
.A(n_1168),
.B(n_22),
.Y(n_1250)
);

INVx3_ASAP7_75t_L g1251 ( 
.A(n_1191),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1181),
.Y(n_1252)
);

INVxp67_ASAP7_75t_L g1253 ( 
.A(n_1210),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_1179),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_1199),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1168),
.B(n_22),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1186),
.Y(n_1257)
);

AND2x4_ASAP7_75t_L g1258 ( 
.A(n_1191),
.B(n_528),
.Y(n_1258)
);

INVx2_ASAP7_75t_L g1259 ( 
.A(n_1206),
.Y(n_1259)
);

HB1xp67_ASAP7_75t_L g1260 ( 
.A(n_1167),
.Y(n_1260)
);

INVx1_ASAP7_75t_SL g1261 ( 
.A(n_1223),
.Y(n_1261)
);

NOR2xp33_ASAP7_75t_L g1262 ( 
.A(n_1239),
.B(n_24),
.Y(n_1262)
);

INVx3_ASAP7_75t_L g1263 ( 
.A(n_1177),
.Y(n_1263)
);

BUFx3_ASAP7_75t_L g1264 ( 
.A(n_1174),
.Y(n_1264)
);

NOR2x1p5_ASAP7_75t_L g1265 ( 
.A(n_1216),
.B(n_25),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_1174),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1175),
.B(n_1172),
.Y(n_1267)
);

INVx2_ASAP7_75t_SL g1268 ( 
.A(n_1164),
.Y(n_1268)
);

AND2x4_ASAP7_75t_L g1269 ( 
.A(n_1195),
.B(n_527),
.Y(n_1269)
);

CKINVDCx5p33_ASAP7_75t_R g1270 ( 
.A(n_1211),
.Y(n_1270)
);

CKINVDCx10_ASAP7_75t_R g1271 ( 
.A(n_1187),
.Y(n_1271)
);

INVx3_ASAP7_75t_L g1272 ( 
.A(n_1227),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1189),
.B(n_25),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_SL g1274 ( 
.A(n_1165),
.B(n_26),
.Y(n_1274)
);

OR2x6_ASAP7_75t_L g1275 ( 
.A(n_1178),
.B(n_1194),
.Y(n_1275)
);

INVx2_ASAP7_75t_L g1276 ( 
.A(n_1214),
.Y(n_1276)
);

AND2x4_ASAP7_75t_L g1277 ( 
.A(n_1176),
.B(n_93),
.Y(n_1277)
);

BUFx3_ASAP7_75t_L g1278 ( 
.A(n_1164),
.Y(n_1278)
);

BUFx3_ASAP7_75t_L g1279 ( 
.A(n_1164),
.Y(n_1279)
);

BUFx12f_ASAP7_75t_SL g1280 ( 
.A(n_1204),
.Y(n_1280)
);

BUFx3_ASAP7_75t_L g1281 ( 
.A(n_1176),
.Y(n_1281)
);

BUFx3_ASAP7_75t_L g1282 ( 
.A(n_1176),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1218),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1188),
.Y(n_1284)
);

OR2x6_ASAP7_75t_L g1285 ( 
.A(n_1240),
.B(n_27),
.Y(n_1285)
);

BUFx3_ASAP7_75t_L g1286 ( 
.A(n_1240),
.Y(n_1286)
);

A2O1A1Ixp33_ASAP7_75t_L g1287 ( 
.A1(n_1237),
.A2(n_29),
.B(n_27),
.C(n_28),
.Y(n_1287)
);

INVx2_ASAP7_75t_L g1288 ( 
.A(n_1219),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1225),
.B(n_28),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1233),
.B(n_29),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1185),
.A2(n_96),
.B(n_94),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1182),
.B(n_30),
.Y(n_1292)
);

INVx3_ASAP7_75t_L g1293 ( 
.A(n_1227),
.Y(n_1293)
);

BUFx8_ASAP7_75t_L g1294 ( 
.A(n_1226),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1193),
.B(n_31),
.Y(n_1295)
);

HB1xp67_ASAP7_75t_L g1296 ( 
.A(n_1180),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_1222),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1196),
.B(n_31),
.Y(n_1298)
);

BUFx2_ASAP7_75t_L g1299 ( 
.A(n_1192),
.Y(n_1299)
);

AOI22xp5_ASAP7_75t_L g1300 ( 
.A1(n_1213),
.A2(n_34),
.B1(n_32),
.B2(n_33),
.Y(n_1300)
);

AO22x1_ASAP7_75t_L g1301 ( 
.A1(n_1241),
.A2(n_36),
.B1(n_34),
.B2(n_35),
.Y(n_1301)
);

BUFx6f_ASAP7_75t_L g1302 ( 
.A(n_1227),
.Y(n_1302)
);

BUFx2_ASAP7_75t_L g1303 ( 
.A(n_1209),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1184),
.B(n_35),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1190),
.B(n_37),
.Y(n_1305)
);

BUFx3_ASAP7_75t_L g1306 ( 
.A(n_1220),
.Y(n_1306)
);

NOR2xp33_ASAP7_75t_L g1307 ( 
.A(n_1173),
.B(n_38),
.Y(n_1307)
);

INVx3_ASAP7_75t_L g1308 ( 
.A(n_1207),
.Y(n_1308)
);

AND2x4_ASAP7_75t_L g1309 ( 
.A(n_1220),
.B(n_526),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1215),
.Y(n_1310)
);

INVx1_ASAP7_75t_SL g1311 ( 
.A(n_1208),
.Y(n_1311)
);

BUFx3_ASAP7_75t_L g1312 ( 
.A(n_1220),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1201),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1231),
.B(n_1238),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_1228),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1235),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1234),
.Y(n_1317)
);

OAI22xp5_ASAP7_75t_SL g1318 ( 
.A1(n_1224),
.A2(n_41),
.B1(n_39),
.B2(n_40),
.Y(n_1318)
);

INVx5_ASAP7_75t_L g1319 ( 
.A(n_1171),
.Y(n_1319)
);

NOR2xp33_ASAP7_75t_SL g1320 ( 
.A(n_1202),
.B(n_98),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1267),
.B(n_1230),
.Y(n_1321)
);

AOI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1291),
.A2(n_1197),
.B(n_1205),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1250),
.B(n_1229),
.Y(n_1323)
);

OAI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1314),
.A2(n_1236),
.B(n_1221),
.Y(n_1324)
);

OAI21x1_ASAP7_75t_L g1325 ( 
.A1(n_1244),
.A2(n_1198),
.B(n_1200),
.Y(n_1325)
);

OAI21x1_ASAP7_75t_L g1326 ( 
.A1(n_1272),
.A2(n_1203),
.B(n_1232),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1283),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1313),
.B(n_39),
.Y(n_1328)
);

AOI21xp5_ASAP7_75t_L g1329 ( 
.A1(n_1245),
.A2(n_40),
.B(n_41),
.Y(n_1329)
);

OAI21x1_ASAP7_75t_L g1330 ( 
.A1(n_1272),
.A2(n_100),
.B(n_99),
.Y(n_1330)
);

AOI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1320),
.A2(n_42),
.B(n_43),
.Y(n_1331)
);

OAI21xp33_ASAP7_75t_L g1332 ( 
.A1(n_1300),
.A2(n_42),
.B(n_44),
.Y(n_1332)
);

OAI21x1_ASAP7_75t_L g1333 ( 
.A1(n_1293),
.A2(n_104),
.B(n_102),
.Y(n_1333)
);

OAI21x1_ASAP7_75t_SL g1334 ( 
.A1(n_1298),
.A2(n_45),
.B(n_46),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1288),
.Y(n_1335)
);

OAI21x1_ASAP7_75t_L g1336 ( 
.A1(n_1293),
.A2(n_106),
.B(n_105),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1296),
.B(n_46),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1247),
.Y(n_1338)
);

BUFx2_ASAP7_75t_L g1339 ( 
.A(n_1243),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1262),
.B(n_47),
.Y(n_1340)
);

BUFx6f_ASAP7_75t_L g1341 ( 
.A(n_1286),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1252),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1256),
.B(n_47),
.Y(n_1343)
);

O2A1O1Ixp5_ASAP7_75t_L g1344 ( 
.A1(n_1301),
.A2(n_50),
.B(n_48),
.C(n_49),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1261),
.B(n_48),
.Y(n_1345)
);

AND2x2_ASAP7_75t_SL g1346 ( 
.A(n_1309),
.B(n_49),
.Y(n_1346)
);

OAI21x1_ASAP7_75t_L g1347 ( 
.A1(n_1257),
.A2(n_1284),
.B(n_1310),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1242),
.B(n_50),
.Y(n_1348)
);

AO31x2_ASAP7_75t_L g1349 ( 
.A1(n_1316),
.A2(n_109),
.A3(n_110),
.B(n_107),
.Y(n_1349)
);

OAI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1304),
.A2(n_112),
.B(n_111),
.Y(n_1350)
);

AO22x2_ASAP7_75t_L g1351 ( 
.A1(n_1317),
.A2(n_54),
.B1(n_51),
.B2(n_53),
.Y(n_1351)
);

AOI21xp5_ASAP7_75t_L g1352 ( 
.A1(n_1301),
.A2(n_53),
.B(n_55),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1251),
.B(n_55),
.Y(n_1353)
);

AOI21x1_ASAP7_75t_L g1354 ( 
.A1(n_1305),
.A2(n_119),
.B(n_117),
.Y(n_1354)
);

AND2x4_ASAP7_75t_L g1355 ( 
.A(n_1251),
.B(n_56),
.Y(n_1355)
);

NAND2x1p5_ASAP7_75t_L g1356 ( 
.A(n_1278),
.B(n_121),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1315),
.B(n_56),
.Y(n_1357)
);

NOR4xp25_ASAP7_75t_L g1358 ( 
.A(n_1287),
.B(n_1307),
.C(n_1246),
.D(n_1273),
.Y(n_1358)
);

OAI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1292),
.A2(n_124),
.B(n_123),
.Y(n_1359)
);

AOI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1309),
.A2(n_1318),
.B(n_1290),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_SL g1361 ( 
.A(n_1319),
.B(n_57),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1253),
.B(n_1260),
.Y(n_1362)
);

OAI21x1_ASAP7_75t_L g1363 ( 
.A1(n_1289),
.A2(n_129),
.B(n_127),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1297),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1319),
.B(n_1258),
.Y(n_1365)
);

BUFx10_ASAP7_75t_L g1366 ( 
.A(n_1266),
.Y(n_1366)
);

BUFx5_ASAP7_75t_L g1367 ( 
.A(n_1281),
.Y(n_1367)
);

BUFx3_ASAP7_75t_L g1368 ( 
.A(n_1270),
.Y(n_1368)
);

BUFx5_ASAP7_75t_L g1369 ( 
.A(n_1282),
.Y(n_1369)
);

AOI21xp5_ASAP7_75t_L g1370 ( 
.A1(n_1274),
.A2(n_57),
.B(n_58),
.Y(n_1370)
);

OAI21x1_ASAP7_75t_L g1371 ( 
.A1(n_1308),
.A2(n_1295),
.B(n_1254),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1285),
.B(n_58),
.Y(n_1372)
);

OAI21x1_ASAP7_75t_L g1373 ( 
.A1(n_1308),
.A2(n_131),
.B(n_130),
.Y(n_1373)
);

AOI21xp5_ASAP7_75t_L g1374 ( 
.A1(n_1258),
.A2(n_60),
.B(n_61),
.Y(n_1374)
);

AND2x4_ASAP7_75t_L g1375 ( 
.A(n_1275),
.B(n_60),
.Y(n_1375)
);

A2O1A1Ixp33_ASAP7_75t_L g1376 ( 
.A1(n_1319),
.A2(n_64),
.B(n_62),
.C(n_63),
.Y(n_1376)
);

AOI21x1_ASAP7_75t_L g1377 ( 
.A1(n_1275),
.A2(n_133),
.B(n_132),
.Y(n_1377)
);

AOI21xp5_ASAP7_75t_L g1378 ( 
.A1(n_1277),
.A2(n_62),
.B(n_63),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1285),
.B(n_64),
.Y(n_1379)
);

OAI21xp5_ASAP7_75t_L g1380 ( 
.A1(n_1299),
.A2(n_65),
.B(n_66),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1249),
.Y(n_1381)
);

INVx3_ASAP7_75t_L g1382 ( 
.A(n_1248),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1263),
.B(n_1303),
.Y(n_1383)
);

A2O1A1Ixp33_ASAP7_75t_L g1384 ( 
.A1(n_1306),
.A2(n_68),
.B(n_66),
.C(n_67),
.Y(n_1384)
);

OAI21x1_ASAP7_75t_SL g1385 ( 
.A1(n_1268),
.A2(n_67),
.B(n_68),
.Y(n_1385)
);

HB1xp67_ASAP7_75t_L g1386 ( 
.A(n_1302),
.Y(n_1386)
);

AOI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1277),
.A2(n_69),
.B(n_70),
.Y(n_1387)
);

O2A1O1Ixp33_ASAP7_75t_L g1388 ( 
.A1(n_1263),
.A2(n_71),
.B(n_69),
.C(n_70),
.Y(n_1388)
);

INVx5_ASAP7_75t_L g1389 ( 
.A(n_1264),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1294),
.B(n_71),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1294),
.B(n_72),
.Y(n_1391)
);

AND2x4_ASAP7_75t_L g1392 ( 
.A(n_1311),
.B(n_73),
.Y(n_1392)
);

OA21x2_ASAP7_75t_L g1393 ( 
.A1(n_1255),
.A2(n_73),
.B(n_74),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_1259),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1265),
.B(n_1248),
.Y(n_1395)
);

OAI22xp5_ASAP7_75t_L g1396 ( 
.A1(n_1279),
.A2(n_76),
.B1(n_74),
.B2(n_75),
.Y(n_1396)
);

CKINVDCx8_ASAP7_75t_R g1397 ( 
.A(n_1271),
.Y(n_1397)
);

OA21x2_ASAP7_75t_L g1398 ( 
.A1(n_1276),
.A2(n_77),
.B(n_78),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1302),
.Y(n_1399)
);

AOI21xp5_ASAP7_75t_L g1400 ( 
.A1(n_1269),
.A2(n_77),
.B(n_78),
.Y(n_1400)
);

OAI21x1_ASAP7_75t_L g1401 ( 
.A1(n_1302),
.A2(n_1312),
.B(n_1280),
.Y(n_1401)
);

OAI21xp5_ASAP7_75t_L g1402 ( 
.A1(n_1269),
.A2(n_79),
.B(n_80),
.Y(n_1402)
);

NOR2xp33_ASAP7_75t_L g1403 ( 
.A(n_1242),
.B(n_79),
.Y(n_1403)
);

AOI21x1_ASAP7_75t_SL g1404 ( 
.A1(n_1314),
.A2(n_80),
.B(n_81),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_L g1405 ( 
.A1(n_1291),
.A2(n_135),
.B(n_134),
.Y(n_1405)
);

OAI21x1_ASAP7_75t_L g1406 ( 
.A1(n_1291),
.A2(n_137),
.B(n_136),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1267),
.B(n_82),
.Y(n_1407)
);

BUFx2_ASAP7_75t_L g1408 ( 
.A(n_1243),
.Y(n_1408)
);

OAI21x1_ASAP7_75t_L g1409 ( 
.A1(n_1291),
.A2(n_139),
.B(n_138),
.Y(n_1409)
);

AND2x4_ASAP7_75t_L g1410 ( 
.A(n_1339),
.B(n_141),
.Y(n_1410)
);

AOI21x1_ASAP7_75t_L g1411 ( 
.A1(n_1322),
.A2(n_82),
.B(n_83),
.Y(n_1411)
);

CKINVDCx5p33_ASAP7_75t_R g1412 ( 
.A(n_1397),
.Y(n_1412)
);

BUFx2_ASAP7_75t_L g1413 ( 
.A(n_1408),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1362),
.B(n_84),
.Y(n_1414)
);

AOI21xp5_ASAP7_75t_L g1415 ( 
.A1(n_1402),
.A2(n_84),
.B(n_85),
.Y(n_1415)
);

INVx6_ASAP7_75t_L g1416 ( 
.A(n_1389),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1338),
.B(n_1342),
.Y(n_1417)
);

INVx2_ASAP7_75t_SL g1418 ( 
.A(n_1389),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1347),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1327),
.Y(n_1420)
);

AND2x4_ASAP7_75t_L g1421 ( 
.A(n_1368),
.B(n_142),
.Y(n_1421)
);

AOI21xp5_ASAP7_75t_L g1422 ( 
.A1(n_1360),
.A2(n_85),
.B(n_86),
.Y(n_1422)
);

BUFx3_ASAP7_75t_L g1423 ( 
.A(n_1341),
.Y(n_1423)
);

AOI21xp5_ASAP7_75t_L g1424 ( 
.A1(n_1325),
.A2(n_86),
.B(n_87),
.Y(n_1424)
);

AND2x2_ASAP7_75t_SL g1425 ( 
.A(n_1346),
.B(n_1403),
.Y(n_1425)
);

AOI22xp5_ASAP7_75t_L g1426 ( 
.A1(n_1332),
.A2(n_1348),
.B1(n_1340),
.B2(n_1380),
.Y(n_1426)
);

AOI21xp5_ASAP7_75t_L g1427 ( 
.A1(n_1405),
.A2(n_87),
.B(n_88),
.Y(n_1427)
);

OAI22xp5_ASAP7_75t_L g1428 ( 
.A1(n_1374),
.A2(n_88),
.B1(n_89),
.B2(n_143),
.Y(n_1428)
);

INVx3_ASAP7_75t_L g1429 ( 
.A(n_1341),
.Y(n_1429)
);

INVx3_ASAP7_75t_SL g1430 ( 
.A(n_1366),
.Y(n_1430)
);

OR2x2_ASAP7_75t_L g1431 ( 
.A(n_1335),
.B(n_144),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1407),
.B(n_147),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1321),
.B(n_148),
.Y(n_1433)
);

HB1xp67_ASAP7_75t_L g1434 ( 
.A(n_1386),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1351),
.A2(n_154),
.B1(n_152),
.B2(n_153),
.Y(n_1435)
);

NOR2xp33_ASAP7_75t_L g1436 ( 
.A(n_1375),
.B(n_156),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1364),
.Y(n_1437)
);

AO22x2_ASAP7_75t_L g1438 ( 
.A1(n_1352),
.A2(n_159),
.B1(n_157),
.B2(n_158),
.Y(n_1438)
);

AND2x4_ASAP7_75t_L g1439 ( 
.A(n_1399),
.B(n_160),
.Y(n_1439)
);

BUFx2_ASAP7_75t_L g1440 ( 
.A(n_1383),
.Y(n_1440)
);

NOR2x1_ASAP7_75t_SL g1441 ( 
.A(n_1365),
.B(n_162),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1351),
.B(n_163),
.Y(n_1442)
);

HB1xp67_ASAP7_75t_L g1443 ( 
.A(n_1371),
.Y(n_1443)
);

AOI21xp5_ASAP7_75t_L g1444 ( 
.A1(n_1406),
.A2(n_164),
.B(n_165),
.Y(n_1444)
);

AOI21xp5_ASAP7_75t_L g1445 ( 
.A1(n_1409),
.A2(n_166),
.B(n_168),
.Y(n_1445)
);

INVx3_ASAP7_75t_L g1446 ( 
.A(n_1382),
.Y(n_1446)
);

BUFx6f_ASAP7_75t_L g1447 ( 
.A(n_1401),
.Y(n_1447)
);

NOR2xp33_ASAP7_75t_L g1448 ( 
.A(n_1357),
.B(n_169),
.Y(n_1448)
);

CKINVDCx16_ASAP7_75t_R g1449 ( 
.A(n_1395),
.Y(n_1449)
);

INVx4_ASAP7_75t_L g1450 ( 
.A(n_1355),
.Y(n_1450)
);

AOI21xp5_ASAP7_75t_L g1451 ( 
.A1(n_1324),
.A2(n_170),
.B(n_171),
.Y(n_1451)
);

OAI22xp5_ASAP7_75t_SL g1452 ( 
.A1(n_1390),
.A2(n_174),
.B1(n_172),
.B2(n_173),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1381),
.Y(n_1453)
);

O2A1O1Ixp5_ASAP7_75t_SL g1454 ( 
.A1(n_1361),
.A2(n_179),
.B(n_177),
.C(n_178),
.Y(n_1454)
);

BUFx4f_ASAP7_75t_L g1455 ( 
.A(n_1356),
.Y(n_1455)
);

BUFx12f_ASAP7_75t_L g1456 ( 
.A(n_1392),
.Y(n_1456)
);

INVx1_ASAP7_75t_SL g1457 ( 
.A(n_1343),
.Y(n_1457)
);

AOI21xp5_ASAP7_75t_L g1458 ( 
.A1(n_1331),
.A2(n_180),
.B(n_182),
.Y(n_1458)
);

BUFx8_ASAP7_75t_L g1459 ( 
.A(n_1372),
.Y(n_1459)
);

CKINVDCx20_ASAP7_75t_R g1460 ( 
.A(n_1391),
.Y(n_1460)
);

AOI22xp33_ASAP7_75t_L g1461 ( 
.A1(n_1323),
.A2(n_187),
.B1(n_183),
.B2(n_186),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1328),
.B(n_190),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1394),
.Y(n_1463)
);

NAND2x1p5_ASAP7_75t_L g1464 ( 
.A(n_1326),
.B(n_191),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1337),
.B(n_192),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1379),
.B(n_193),
.Y(n_1466)
);

OR2x2_ASAP7_75t_L g1467 ( 
.A(n_1345),
.B(n_194),
.Y(n_1467)
);

BUFx3_ASAP7_75t_L g1468 ( 
.A(n_1367),
.Y(n_1468)
);

NOR2xp67_ASAP7_75t_SL g1469 ( 
.A(n_1378),
.B(n_195),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1393),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1398),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1353),
.Y(n_1472)
);

AND2x4_ASAP7_75t_L g1473 ( 
.A(n_1387),
.B(n_196),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1349),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_SL g1475 ( 
.A(n_1367),
.B(n_197),
.Y(n_1475)
);

NOR2x1_ASAP7_75t_L g1476 ( 
.A(n_1329),
.B(n_199),
.Y(n_1476)
);

AOI22xp5_ASAP7_75t_L g1477 ( 
.A1(n_1358),
.A2(n_205),
.B1(n_201),
.B2(n_202),
.Y(n_1477)
);

AND2x6_ASAP7_75t_L g1478 ( 
.A(n_1377),
.B(n_206),
.Y(n_1478)
);

AOI21xp5_ASAP7_75t_SL g1479 ( 
.A1(n_1376),
.A2(n_207),
.B(n_208),
.Y(n_1479)
);

INVx3_ASAP7_75t_L g1480 ( 
.A(n_1367),
.Y(n_1480)
);

AND2x4_ASAP7_75t_L g1481 ( 
.A(n_1400),
.B(n_209),
.Y(n_1481)
);

AOI21xp5_ASAP7_75t_L g1482 ( 
.A1(n_1344),
.A2(n_1373),
.B(n_1359),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1349),
.Y(n_1483)
);

INVx1_ASAP7_75t_SL g1484 ( 
.A(n_1367),
.Y(n_1484)
);

AOI22xp33_ASAP7_75t_L g1485 ( 
.A1(n_1334),
.A2(n_214),
.B1(n_211),
.B2(n_212),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1369),
.B(n_1384),
.Y(n_1486)
);

OR2x2_ASAP7_75t_L g1487 ( 
.A(n_1369),
.B(n_215),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1369),
.Y(n_1488)
);

BUFx2_ASAP7_75t_L g1489 ( 
.A(n_1369),
.Y(n_1489)
);

OAI21xp33_ASAP7_75t_L g1490 ( 
.A1(n_1396),
.A2(n_219),
.B(n_220),
.Y(n_1490)
);

BUFx3_ASAP7_75t_L g1491 ( 
.A(n_1385),
.Y(n_1491)
);

OR2x2_ASAP7_75t_L g1492 ( 
.A(n_1370),
.B(n_222),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1388),
.B(n_223),
.Y(n_1493)
);

INVx2_ASAP7_75t_L g1494 ( 
.A(n_1354),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1363),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_SL g1496 ( 
.A(n_1350),
.B(n_224),
.Y(n_1496)
);

NOR2xp33_ASAP7_75t_SL g1497 ( 
.A(n_1404),
.B(n_225),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1330),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1333),
.B(n_226),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1336),
.B(n_227),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1339),
.B(n_228),
.Y(n_1501)
);

AOI21xp5_ASAP7_75t_L g1502 ( 
.A1(n_1322),
.A2(n_229),
.B(n_230),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1338),
.Y(n_1503)
);

AOI21xp5_ASAP7_75t_L g1504 ( 
.A1(n_1322),
.A2(n_231),
.B(n_232),
.Y(n_1504)
);

INVx6_ASAP7_75t_L g1505 ( 
.A(n_1389),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_SL g1506 ( 
.A(n_1360),
.B(n_233),
.Y(n_1506)
);

A2O1A1Ixp33_ASAP7_75t_L g1507 ( 
.A1(n_1360),
.A2(n_236),
.B(n_234),
.C(n_235),
.Y(n_1507)
);

OAI22xp5_ASAP7_75t_L g1508 ( 
.A1(n_1403),
.A2(n_239),
.B1(n_237),
.B2(n_238),
.Y(n_1508)
);

O2A1O1Ixp5_ASAP7_75t_L g1509 ( 
.A1(n_1422),
.A2(n_248),
.B(n_240),
.C(n_241),
.Y(n_1509)
);

AOI21xp5_ASAP7_75t_SL g1510 ( 
.A1(n_1507),
.A2(n_249),
.B(n_250),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1417),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1440),
.B(n_525),
.Y(n_1512)
);

BUFx8_ASAP7_75t_L g1513 ( 
.A(n_1456),
.Y(n_1513)
);

CKINVDCx5p33_ASAP7_75t_R g1514 ( 
.A(n_1412),
.Y(n_1514)
);

O2A1O1Ixp5_ASAP7_75t_L g1515 ( 
.A1(n_1506),
.A2(n_254),
.B(n_251),
.C(n_253),
.Y(n_1515)
);

NOR2xp33_ASAP7_75t_L g1516 ( 
.A(n_1449),
.B(n_1429),
.Y(n_1516)
);

HB1xp67_ASAP7_75t_L g1517 ( 
.A(n_1434),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1413),
.B(n_524),
.Y(n_1518)
);

AOI21xp5_ASAP7_75t_L g1519 ( 
.A1(n_1502),
.A2(n_1504),
.B(n_1482),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1420),
.Y(n_1520)
);

OR2x2_ASAP7_75t_SL g1521 ( 
.A(n_1416),
.B(n_255),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1457),
.B(n_521),
.Y(n_1522)
);

OR2x6_ASAP7_75t_SL g1523 ( 
.A(n_1414),
.B(n_1442),
.Y(n_1523)
);

O2A1O1Ixp5_ASAP7_75t_L g1524 ( 
.A1(n_1415),
.A2(n_260),
.B(n_257),
.C(n_258),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1503),
.Y(n_1525)
);

CKINVDCx5p33_ASAP7_75t_R g1526 ( 
.A(n_1423),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1450),
.B(n_519),
.Y(n_1527)
);

O2A1O1Ixp5_ASAP7_75t_L g1528 ( 
.A1(n_1508),
.A2(n_264),
.B(n_262),
.C(n_263),
.Y(n_1528)
);

OR2x2_ASAP7_75t_L g1529 ( 
.A(n_1437),
.B(n_1472),
.Y(n_1529)
);

NOR2xp67_ASAP7_75t_L g1530 ( 
.A(n_1418),
.B(n_265),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1501),
.B(n_268),
.Y(n_1531)
);

A2O1A1Ixp33_ASAP7_75t_L g1532 ( 
.A1(n_1425),
.A2(n_273),
.B(n_269),
.C(n_271),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1453),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1489),
.B(n_275),
.Y(n_1534)
);

AOI21xp5_ASAP7_75t_L g1535 ( 
.A1(n_1451),
.A2(n_1486),
.B(n_1496),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1446),
.B(n_518),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1463),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1470),
.Y(n_1538)
);

HB1xp67_ASAP7_75t_L g1539 ( 
.A(n_1419),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1410),
.B(n_276),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1484),
.B(n_517),
.Y(n_1541)
);

A2O1A1Ixp33_ASAP7_75t_SL g1542 ( 
.A1(n_1469),
.A2(n_280),
.B(n_277),
.C(n_278),
.Y(n_1542)
);

AOI21xp5_ASAP7_75t_L g1543 ( 
.A1(n_1479),
.A2(n_1455),
.B(n_1490),
.Y(n_1543)
);

INVx3_ASAP7_75t_L g1544 ( 
.A(n_1416),
.Y(n_1544)
);

INVx2_ASAP7_75t_SL g1545 ( 
.A(n_1505),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1488),
.B(n_515),
.Y(n_1546)
);

OA21x2_ASAP7_75t_L g1547 ( 
.A1(n_1474),
.A2(n_281),
.B(n_284),
.Y(n_1547)
);

AND2x4_ASAP7_75t_L g1548 ( 
.A(n_1468),
.B(n_285),
.Y(n_1548)
);

CKINVDCx6p67_ASAP7_75t_R g1549 ( 
.A(n_1430),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1505),
.B(n_514),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1471),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1421),
.B(n_286),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1443),
.Y(n_1553)
);

HB1xp67_ASAP7_75t_L g1554 ( 
.A(n_1495),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1483),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1480),
.B(n_512),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1447),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1436),
.B(n_287),
.Y(n_1558)
);

OA21x2_ASAP7_75t_L g1559 ( 
.A1(n_1494),
.A2(n_288),
.B(n_291),
.Y(n_1559)
);

O2A1O1Ixp5_ASAP7_75t_L g1560 ( 
.A1(n_1428),
.A2(n_292),
.B(n_293),
.C(n_294),
.Y(n_1560)
);

INVxp67_ASAP7_75t_L g1561 ( 
.A(n_1465),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1447),
.Y(n_1562)
);

CKINVDCx16_ASAP7_75t_R g1563 ( 
.A(n_1460),
.Y(n_1563)
);

OR2x2_ASAP7_75t_L g1564 ( 
.A(n_1426),
.B(n_1431),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1411),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1498),
.Y(n_1566)
);

NOR2xp33_ASAP7_75t_SL g1567 ( 
.A(n_1448),
.B(n_295),
.Y(n_1567)
);

CKINVDCx20_ASAP7_75t_R g1568 ( 
.A(n_1459),
.Y(n_1568)
);

HB1xp67_ASAP7_75t_L g1569 ( 
.A(n_1464),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_SL g1570 ( 
.A(n_1491),
.B(n_296),
.Y(n_1570)
);

O2A1O1Ixp5_ASAP7_75t_L g1571 ( 
.A1(n_1493),
.A2(n_298),
.B(n_299),
.C(n_300),
.Y(n_1571)
);

HB1xp67_ASAP7_75t_L g1572 ( 
.A(n_1433),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1466),
.B(n_511),
.Y(n_1573)
);

INVxp67_ASAP7_75t_L g1574 ( 
.A(n_1467),
.Y(n_1574)
);

OR2x2_ASAP7_75t_L g1575 ( 
.A(n_1487),
.B(n_301),
.Y(n_1575)
);

O2A1O1Ixp33_ASAP7_75t_L g1576 ( 
.A1(n_1432),
.A2(n_302),
.B(n_305),
.C(n_308),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1438),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1438),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1441),
.B(n_309),
.Y(n_1579)
);

BUFx6f_ASAP7_75t_L g1580 ( 
.A(n_1439),
.Y(n_1580)
);

OAI22xp5_ASAP7_75t_L g1581 ( 
.A1(n_1477),
.A2(n_311),
.B1(n_312),
.B2(n_314),
.Y(n_1581)
);

O2A1O1Ixp5_ASAP7_75t_L g1582 ( 
.A1(n_1424),
.A2(n_316),
.B(n_317),
.C(n_318),
.Y(n_1582)
);

AND2x4_ASAP7_75t_SL g1583 ( 
.A(n_1481),
.B(n_319),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1462),
.B(n_320),
.Y(n_1584)
);

AOI21xp5_ASAP7_75t_L g1585 ( 
.A1(n_1475),
.A2(n_323),
.B(n_324),
.Y(n_1585)
);

AOI21xp5_ASAP7_75t_SL g1586 ( 
.A1(n_1473),
.A2(n_326),
.B(n_327),
.Y(n_1586)
);

AOI21xp5_ASAP7_75t_L g1587 ( 
.A1(n_1444),
.A2(n_1445),
.B(n_1497),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1492),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1435),
.B(n_510),
.Y(n_1589)
);

CKINVDCx5p33_ASAP7_75t_R g1590 ( 
.A(n_1452),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1476),
.B(n_328),
.Y(n_1591)
);

CKINVDCx20_ASAP7_75t_R g1592 ( 
.A(n_1499),
.Y(n_1592)
);

AOI21xp5_ASAP7_75t_L g1593 ( 
.A1(n_1458),
.A2(n_329),
.B(n_330),
.Y(n_1593)
);

A2O1A1Ixp33_ASAP7_75t_L g1594 ( 
.A1(n_1427),
.A2(n_331),
.B(n_332),
.C(n_335),
.Y(n_1594)
);

INVx1_ASAP7_75t_SL g1595 ( 
.A(n_1478),
.Y(n_1595)
);

O2A1O1Ixp5_ASAP7_75t_L g1596 ( 
.A1(n_1500),
.A2(n_336),
.B(n_337),
.C(n_338),
.Y(n_1596)
);

AOI21xp5_ASAP7_75t_L g1597 ( 
.A1(n_1485),
.A2(n_340),
.B(n_343),
.Y(n_1597)
);

AND2x6_ASAP7_75t_L g1598 ( 
.A(n_1478),
.B(n_344),
.Y(n_1598)
);

AND2x2_ASAP7_75t_SL g1599 ( 
.A(n_1461),
.B(n_345),
.Y(n_1599)
);

A2O1A1Ixp33_ASAP7_75t_SL g1600 ( 
.A1(n_1454),
.A2(n_346),
.B(n_347),
.C(n_348),
.Y(n_1600)
);

INVxp67_ASAP7_75t_L g1601 ( 
.A(n_1478),
.Y(n_1601)
);

HB1xp67_ASAP7_75t_L g1602 ( 
.A(n_1434),
.Y(n_1602)
);

AND2x4_ASAP7_75t_L g1603 ( 
.A(n_1413),
.B(n_349),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1420),
.Y(n_1604)
);

A2O1A1Ixp33_ASAP7_75t_L g1605 ( 
.A1(n_1425),
.A2(n_350),
.B(n_352),
.C(n_353),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1417),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_SL g1607 ( 
.A(n_1449),
.B(n_354),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1525),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1529),
.Y(n_1609)
);

CKINVDCx5p33_ASAP7_75t_R g1610 ( 
.A(n_1514),
.Y(n_1610)
);

HB1xp67_ASAP7_75t_L g1611 ( 
.A(n_1553),
.Y(n_1611)
);

OA21x2_ASAP7_75t_L g1612 ( 
.A1(n_1577),
.A2(n_355),
.B(n_356),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1520),
.Y(n_1613)
);

AO21x1_ASAP7_75t_SL g1614 ( 
.A1(n_1565),
.A2(n_357),
.B(n_359),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_1551),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1517),
.B(n_360),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1538),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1537),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1604),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1533),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1602),
.B(n_361),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1511),
.Y(n_1622)
);

HB1xp67_ASAP7_75t_L g1623 ( 
.A(n_1539),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1555),
.Y(n_1624)
);

OAI21xp5_ASAP7_75t_L g1625 ( 
.A1(n_1532),
.A2(n_362),
.B(n_363),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1606),
.Y(n_1626)
);

AND2x4_ASAP7_75t_L g1627 ( 
.A(n_1557),
.B(n_364),
.Y(n_1627)
);

OAI21x1_ASAP7_75t_L g1628 ( 
.A1(n_1535),
.A2(n_365),
.B(n_366),
.Y(n_1628)
);

INVxp33_ASAP7_75t_L g1629 ( 
.A(n_1516),
.Y(n_1629)
);

OR2x2_ASAP7_75t_L g1630 ( 
.A(n_1574),
.B(n_368),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1566),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1554),
.Y(n_1632)
);

AO21x2_ASAP7_75t_L g1633 ( 
.A1(n_1562),
.A2(n_369),
.B(n_370),
.Y(n_1633)
);

AO21x2_ASAP7_75t_L g1634 ( 
.A1(n_1578),
.A2(n_371),
.B(n_372),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1572),
.B(n_374),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1588),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1563),
.B(n_379),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1564),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1523),
.Y(n_1639)
);

AND2x4_ASAP7_75t_L g1640 ( 
.A(n_1601),
.B(n_380),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1592),
.Y(n_1641)
);

OA21x2_ASAP7_75t_L g1642 ( 
.A1(n_1519),
.A2(n_381),
.B(n_382),
.Y(n_1642)
);

INVx4_ASAP7_75t_L g1643 ( 
.A(n_1549),
.Y(n_1643)
);

OR2x2_ASAP7_75t_L g1644 ( 
.A(n_1561),
.B(n_384),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1547),
.Y(n_1645)
);

AO21x2_ASAP7_75t_L g1646 ( 
.A1(n_1587),
.A2(n_385),
.B(n_387),
.Y(n_1646)
);

BUFx3_ASAP7_75t_L g1647 ( 
.A(n_1513),
.Y(n_1647)
);

INVx4_ASAP7_75t_L g1648 ( 
.A(n_1544),
.Y(n_1648)
);

HB1xp67_ASAP7_75t_L g1649 ( 
.A(n_1518),
.Y(n_1649)
);

INVx3_ASAP7_75t_L g1650 ( 
.A(n_1545),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1595),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1569),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1512),
.Y(n_1653)
);

CKINVDCx20_ASAP7_75t_R g1654 ( 
.A(n_1568),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1547),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1580),
.Y(n_1656)
);

INVx3_ASAP7_75t_L g1657 ( 
.A(n_1603),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1580),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1580),
.Y(n_1659)
);

OAI21x1_ASAP7_75t_L g1660 ( 
.A1(n_1543),
.A2(n_388),
.B(n_389),
.Y(n_1660)
);

HB1xp67_ASAP7_75t_L g1661 ( 
.A(n_1534),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1546),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1559),
.Y(n_1663)
);

AOI22xp5_ASAP7_75t_SL g1664 ( 
.A1(n_1590),
.A2(n_391),
.B1(n_393),
.B2(n_394),
.Y(n_1664)
);

OAI21x1_ASAP7_75t_L g1665 ( 
.A1(n_1559),
.A2(n_395),
.B(n_396),
.Y(n_1665)
);

BUFx12f_ASAP7_75t_L g1666 ( 
.A(n_1526),
.Y(n_1666)
);

INVx3_ASAP7_75t_L g1667 ( 
.A(n_1548),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1522),
.Y(n_1668)
);

HB1xp67_ASAP7_75t_L g1669 ( 
.A(n_1541),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1575),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1521),
.Y(n_1671)
);

BUFx2_ASAP7_75t_L g1672 ( 
.A(n_1527),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1550),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1556),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1548),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_1591),
.Y(n_1676)
);

OAI21x1_ASAP7_75t_L g1677 ( 
.A1(n_1596),
.A2(n_397),
.B(n_398),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1617),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1617),
.Y(n_1679)
);

AOI22xp33_ASAP7_75t_L g1680 ( 
.A1(n_1625),
.A2(n_1599),
.B1(n_1598),
.B2(n_1581),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1661),
.B(n_1531),
.Y(n_1681)
);

HB1xp67_ASAP7_75t_L g1682 ( 
.A(n_1623),
.Y(n_1682)
);

NOR2xp67_ASAP7_75t_SL g1683 ( 
.A(n_1647),
.B(n_1586),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1611),
.Y(n_1684)
);

INVx1_ASAP7_75t_SL g1685 ( 
.A(n_1672),
.Y(n_1685)
);

INVxp67_ASAP7_75t_SL g1686 ( 
.A(n_1623),
.Y(n_1686)
);

BUFx2_ASAP7_75t_L g1687 ( 
.A(n_1661),
.Y(n_1687)
);

INVx5_ASAP7_75t_SL g1688 ( 
.A(n_1640),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1639),
.B(n_1536),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1624),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1649),
.B(n_1607),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1649),
.B(n_1552),
.Y(n_1692)
);

HB1xp67_ASAP7_75t_L g1693 ( 
.A(n_1611),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1669),
.B(n_1558),
.Y(n_1694)
);

OAI21xp5_ASAP7_75t_SL g1695 ( 
.A1(n_1625),
.A2(n_1605),
.B(n_1540),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1622),
.B(n_1579),
.Y(n_1696)
);

INVx4_ASAP7_75t_L g1697 ( 
.A(n_1647),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1624),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1669),
.B(n_1570),
.Y(n_1699)
);

AOI21xp33_ASAP7_75t_SL g1700 ( 
.A1(n_1610),
.A2(n_1584),
.B(n_1573),
.Y(n_1700)
);

AOI22xp33_ASAP7_75t_L g1701 ( 
.A1(n_1634),
.A2(n_1598),
.B1(n_1589),
.B2(n_1567),
.Y(n_1701)
);

OAI22xp33_ASAP7_75t_L g1702 ( 
.A1(n_1671),
.A2(n_1530),
.B1(n_1597),
.B2(n_1593),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1626),
.Y(n_1703)
);

INVx4_ASAP7_75t_SL g1704 ( 
.A(n_1666),
.Y(n_1704)
);

INVx2_ASAP7_75t_L g1705 ( 
.A(n_1631),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1608),
.Y(n_1706)
);

BUFx3_ASAP7_75t_L g1707 ( 
.A(n_1654),
.Y(n_1707)
);

BUFx2_ASAP7_75t_L g1708 ( 
.A(n_1648),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1613),
.Y(n_1709)
);

CKINVDCx8_ASAP7_75t_R g1710 ( 
.A(n_1610),
.Y(n_1710)
);

OR2x2_ASAP7_75t_L g1711 ( 
.A(n_1609),
.B(n_1594),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1619),
.Y(n_1712)
);

INVx4_ASAP7_75t_L g1713 ( 
.A(n_1643),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1620),
.Y(n_1714)
);

INVx4_ASAP7_75t_L g1715 ( 
.A(n_1643),
.Y(n_1715)
);

AND2x4_ASAP7_75t_L g1716 ( 
.A(n_1667),
.B(n_1598),
.Y(n_1716)
);

INVxp67_ASAP7_75t_SL g1717 ( 
.A(n_1655),
.Y(n_1717)
);

BUFx2_ASAP7_75t_L g1718 ( 
.A(n_1648),
.Y(n_1718)
);

BUFx3_ASAP7_75t_L g1719 ( 
.A(n_1654),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1652),
.B(n_1583),
.Y(n_1720)
);

BUFx2_ASAP7_75t_L g1721 ( 
.A(n_1650),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1629),
.B(n_1598),
.Y(n_1722)
);

NOR2xp33_ASAP7_75t_L g1723 ( 
.A(n_1629),
.B(n_1576),
.Y(n_1723)
);

INVx2_ASAP7_75t_SL g1724 ( 
.A(n_1650),
.Y(n_1724)
);

HB1xp67_ASAP7_75t_L g1725 ( 
.A(n_1632),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1631),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1638),
.Y(n_1727)
);

AND2x4_ASAP7_75t_L g1728 ( 
.A(n_1667),
.B(n_1585),
.Y(n_1728)
);

AND2x4_ASAP7_75t_L g1729 ( 
.A(n_1651),
.B(n_1656),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1693),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1725),
.B(n_1670),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1690),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1685),
.B(n_1641),
.Y(n_1733)
);

OR2x6_ASAP7_75t_L g1734 ( 
.A(n_1697),
.B(n_1640),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1685),
.B(n_1657),
.Y(n_1735)
);

OR2x2_ASAP7_75t_L g1736 ( 
.A(n_1687),
.B(n_1653),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1694),
.B(n_1657),
.Y(n_1737)
);

INVx4_ASAP7_75t_L g1738 ( 
.A(n_1697),
.Y(n_1738)
);

OR2x2_ASAP7_75t_L g1739 ( 
.A(n_1682),
.B(n_1662),
.Y(n_1739)
);

BUFx3_ASAP7_75t_L g1740 ( 
.A(n_1707),
.Y(n_1740)
);

NAND2x1_ASAP7_75t_L g1741 ( 
.A(n_1721),
.B(n_1675),
.Y(n_1741)
);

OAI321xp33_ASAP7_75t_L g1742 ( 
.A1(n_1680),
.A2(n_1645),
.A3(n_1635),
.B1(n_1676),
.B2(n_1663),
.C(n_1644),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1725),
.Y(n_1743)
);

HB1xp67_ASAP7_75t_L g1744 ( 
.A(n_1693),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1698),
.Y(n_1745)
);

INVx2_ASAP7_75t_L g1746 ( 
.A(n_1705),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1706),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1714),
.Y(n_1748)
);

OR2x2_ASAP7_75t_L g1749 ( 
.A(n_1727),
.B(n_1674),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1681),
.B(n_1658),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1726),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1709),
.Y(n_1752)
);

INVxp67_ASAP7_75t_SL g1753 ( 
.A(n_1723),
.Y(n_1753)
);

AND2x4_ASAP7_75t_L g1754 ( 
.A(n_1716),
.B(n_1659),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1712),
.Y(n_1755)
);

BUFx3_ASAP7_75t_L g1756 ( 
.A(n_1719),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1678),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1679),
.Y(n_1758)
);

AND2x4_ASAP7_75t_L g1759 ( 
.A(n_1716),
.B(n_1616),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1717),
.Y(n_1760)
);

INVx2_ASAP7_75t_L g1761 ( 
.A(n_1711),
.Y(n_1761)
);

AND2x4_ASAP7_75t_L g1762 ( 
.A(n_1708),
.B(n_1718),
.Y(n_1762)
);

AND2x4_ASAP7_75t_L g1763 ( 
.A(n_1729),
.B(n_1621),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1717),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1747),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1763),
.B(n_1724),
.Y(n_1766)
);

AND2x4_ASAP7_75t_L g1767 ( 
.A(n_1762),
.B(n_1692),
.Y(n_1767)
);

AND2x4_ASAP7_75t_L g1768 ( 
.A(n_1762),
.B(n_1713),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1748),
.Y(n_1769)
);

INVx1_ASAP7_75t_SL g1770 ( 
.A(n_1740),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1752),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1753),
.B(n_1684),
.Y(n_1772)
);

AND2x4_ASAP7_75t_SL g1773 ( 
.A(n_1734),
.B(n_1713),
.Y(n_1773)
);

OR2x2_ASAP7_75t_L g1774 ( 
.A(n_1731),
.B(n_1686),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1755),
.Y(n_1775)
);

OR2x2_ASAP7_75t_L g1776 ( 
.A(n_1739),
.B(n_1686),
.Y(n_1776)
);

INVxp67_ASAP7_75t_L g1777 ( 
.A(n_1733),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1763),
.B(n_1715),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1735),
.B(n_1715),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1743),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1749),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1730),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1730),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1757),
.Y(n_1784)
);

HB1xp67_ASAP7_75t_L g1785 ( 
.A(n_1744),
.Y(n_1785)
);

BUFx2_ASAP7_75t_SL g1786 ( 
.A(n_1756),
.Y(n_1786)
);

AND2x4_ASAP7_75t_L g1787 ( 
.A(n_1759),
.B(n_1704),
.Y(n_1787)
);

INVx4_ASAP7_75t_L g1788 ( 
.A(n_1738),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1737),
.B(n_1729),
.Y(n_1789)
);

INVx2_ASAP7_75t_L g1790 ( 
.A(n_1736),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1759),
.B(n_1699),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1750),
.B(n_1754),
.Y(n_1792)
);

INVx3_ASAP7_75t_L g1793 ( 
.A(n_1738),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1761),
.B(n_1703),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1757),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1754),
.B(n_1734),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1732),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1784),
.Y(n_1798)
);

AO21x2_ASAP7_75t_L g1799 ( 
.A1(n_1783),
.A2(n_1764),
.B(n_1760),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_1791),
.Y(n_1800)
);

AOI22xp5_ASAP7_75t_L g1801 ( 
.A1(n_1777),
.A2(n_1695),
.B1(n_1701),
.B2(n_1683),
.Y(n_1801)
);

AND2x2_ASAP7_75t_SL g1802 ( 
.A(n_1787),
.B(n_1722),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1765),
.Y(n_1803)
);

HB1xp67_ASAP7_75t_L g1804 ( 
.A(n_1785),
.Y(n_1804)
);

AND2x4_ASAP7_75t_L g1805 ( 
.A(n_1787),
.B(n_1704),
.Y(n_1805)
);

BUFx2_ASAP7_75t_L g1806 ( 
.A(n_1768),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1765),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1794),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1769),
.Y(n_1809)
);

OR2x2_ASAP7_75t_L g1810 ( 
.A(n_1772),
.B(n_1696),
.Y(n_1810)
);

NAND3xp33_ASAP7_75t_L g1811 ( 
.A(n_1782),
.B(n_1764),
.C(n_1760),
.Y(n_1811)
);

AO21x2_ASAP7_75t_L g1812 ( 
.A1(n_1783),
.A2(n_1700),
.B(n_1635),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1771),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1781),
.B(n_1758),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1784),
.Y(n_1815)
);

OR2x2_ASAP7_75t_L g1816 ( 
.A(n_1808),
.B(n_1804),
.Y(n_1816)
);

BUFx2_ASAP7_75t_L g1817 ( 
.A(n_1805),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1800),
.B(n_1790),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1805),
.B(n_1792),
.Y(n_1819)
);

INVx2_ASAP7_75t_L g1820 ( 
.A(n_1812),
.Y(n_1820)
);

HB1xp67_ASAP7_75t_L g1821 ( 
.A(n_1809),
.Y(n_1821)
);

NAND2x1p5_ASAP7_75t_L g1822 ( 
.A(n_1806),
.B(n_1770),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1798),
.Y(n_1823)
);

INVx2_ASAP7_75t_SL g1824 ( 
.A(n_1802),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1798),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1815),
.Y(n_1826)
);

INVx2_ASAP7_75t_SL g1827 ( 
.A(n_1814),
.Y(n_1827)
);

INVx2_ASAP7_75t_SL g1828 ( 
.A(n_1810),
.Y(n_1828)
);

NAND2x1p5_ASAP7_75t_L g1829 ( 
.A(n_1801),
.B(n_1637),
.Y(n_1829)
);

INVx2_ASAP7_75t_L g1830 ( 
.A(n_1822),
.Y(n_1830)
);

INVx2_ASAP7_75t_L g1831 ( 
.A(n_1817),
.Y(n_1831)
);

AOI211xp5_ASAP7_75t_L g1832 ( 
.A1(n_1824),
.A2(n_1811),
.B(n_1700),
.C(n_1695),
.Y(n_1832)
);

AOI22xp33_ASAP7_75t_L g1833 ( 
.A1(n_1820),
.A2(n_1799),
.B1(n_1797),
.B2(n_1646),
.Y(n_1833)
);

INVx2_ASAP7_75t_L g1834 ( 
.A(n_1819),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1828),
.B(n_1813),
.Y(n_1835)
);

OR2x2_ASAP7_75t_L g1836 ( 
.A(n_1816),
.B(n_1780),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1827),
.B(n_1786),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1821),
.B(n_1803),
.Y(n_1838)
);

AND2x2_ASAP7_75t_L g1839 ( 
.A(n_1818),
.B(n_1768),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1823),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1825),
.B(n_1807),
.Y(n_1841)
);

AND2x4_ASAP7_75t_L g1842 ( 
.A(n_1823),
.B(n_1788),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1831),
.B(n_1826),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1840),
.Y(n_1844)
);

NOR2xp33_ASAP7_75t_L g1845 ( 
.A(n_1837),
.B(n_1788),
.Y(n_1845)
);

AND2x2_ASAP7_75t_L g1846 ( 
.A(n_1830),
.B(n_1796),
.Y(n_1846)
);

HB1xp67_ASAP7_75t_L g1847 ( 
.A(n_1834),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1839),
.Y(n_1848)
);

OR2x2_ASAP7_75t_L g1849 ( 
.A(n_1835),
.B(n_1774),
.Y(n_1849)
);

HB1xp67_ASAP7_75t_L g1850 ( 
.A(n_1842),
.Y(n_1850)
);

OR2x2_ASAP7_75t_L g1851 ( 
.A(n_1836),
.B(n_1826),
.Y(n_1851)
);

OR2x2_ASAP7_75t_L g1852 ( 
.A(n_1838),
.B(n_1776),
.Y(n_1852)
);

NOR2xp33_ASAP7_75t_R g1853 ( 
.A(n_1842),
.B(n_1710),
.Y(n_1853)
);

INVxp67_ASAP7_75t_SL g1854 ( 
.A(n_1850),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1848),
.B(n_1847),
.Y(n_1855)
);

NAND2x1_ASAP7_75t_SL g1856 ( 
.A(n_1846),
.B(n_1793),
.Y(n_1856)
);

OR2x2_ASAP7_75t_L g1857 ( 
.A(n_1852),
.B(n_1841),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1853),
.B(n_1832),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1851),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1845),
.B(n_1849),
.Y(n_1860)
);

INVx2_ASAP7_75t_L g1861 ( 
.A(n_1844),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1843),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1848),
.B(n_1778),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1854),
.Y(n_1864)
);

AOI21xp5_ASAP7_75t_L g1865 ( 
.A1(n_1855),
.A2(n_1859),
.B(n_1860),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1859),
.Y(n_1866)
);

NAND3xp33_ASAP7_75t_SL g1867 ( 
.A(n_1858),
.B(n_1833),
.C(n_1829),
.Y(n_1867)
);

AOI21xp33_ASAP7_75t_L g1868 ( 
.A1(n_1857),
.A2(n_1815),
.B(n_1664),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1862),
.B(n_1775),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1861),
.Y(n_1870)
);

AOI222xp33_ASAP7_75t_L g1871 ( 
.A1(n_1863),
.A2(n_1742),
.B1(n_1795),
.B2(n_1645),
.C1(n_1702),
.C2(n_1691),
.Y(n_1871)
);

INVx1_ASAP7_75t_SL g1872 ( 
.A(n_1864),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1865),
.B(n_1856),
.Y(n_1873)
);

AOI22xp33_ASAP7_75t_L g1874 ( 
.A1(n_1867),
.A2(n_1646),
.B1(n_1612),
.B2(n_1795),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1866),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_L g1876 ( 
.A(n_1870),
.B(n_1767),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1868),
.B(n_1767),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1869),
.B(n_1779),
.Y(n_1878)
);

INVx2_ASAP7_75t_L g1879 ( 
.A(n_1871),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1865),
.B(n_1793),
.Y(n_1880)
);

OR2x2_ASAP7_75t_L g1881 ( 
.A(n_1864),
.B(n_1789),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1864),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1865),
.B(n_1773),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_SL g1884 ( 
.A(n_1873),
.B(n_1766),
.Y(n_1884)
);

NOR3xp33_ASAP7_75t_SL g1885 ( 
.A(n_1880),
.B(n_1696),
.C(n_1758),
.Y(n_1885)
);

NOR4xp25_ASAP7_75t_SL g1886 ( 
.A(n_1875),
.B(n_1688),
.C(n_1741),
.D(n_1614),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1881),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1878),
.B(n_1689),
.Y(n_1888)
);

AO22x2_ASAP7_75t_L g1889 ( 
.A1(n_1872),
.A2(n_1879),
.B1(n_1882),
.B2(n_1883),
.Y(n_1889)
);

XNOR2xp5_ASAP7_75t_L g1890 ( 
.A(n_1876),
.B(n_1877),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_SL g1891 ( 
.A(n_1874),
.B(n_1688),
.Y(n_1891)
);

BUFx2_ASAP7_75t_L g1892 ( 
.A(n_1873),
.Y(n_1892)
);

NAND4xp75_ASAP7_75t_L g1893 ( 
.A(n_1887),
.B(n_1642),
.C(n_1571),
.D(n_1524),
.Y(n_1893)
);

INVxp67_ASAP7_75t_L g1894 ( 
.A(n_1889),
.Y(n_1894)
);

INVx1_ASAP7_75t_SL g1895 ( 
.A(n_1892),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1889),
.Y(n_1896)
);

NAND4xp25_ASAP7_75t_L g1897 ( 
.A(n_1884),
.B(n_1528),
.C(n_1542),
.D(n_1560),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1888),
.B(n_1720),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1890),
.Y(n_1899)
);

AOI211xp5_ASAP7_75t_L g1900 ( 
.A1(n_1894),
.A2(n_1891),
.B(n_1885),
.C(n_1886),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1895),
.B(n_1668),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1896),
.Y(n_1902)
);

INVxp67_ASAP7_75t_L g1903 ( 
.A(n_1899),
.Y(n_1903)
);

NAND3xp33_ASAP7_75t_SL g1904 ( 
.A(n_1898),
.B(n_1630),
.C(n_1509),
.Y(n_1904)
);

NOR2xp33_ASAP7_75t_SL g1905 ( 
.A(n_1897),
.B(n_1728),
.Y(n_1905)
);

AND2x2_ASAP7_75t_L g1906 ( 
.A(n_1893),
.B(n_1728),
.Y(n_1906)
);

NOR3xp33_ASAP7_75t_L g1907 ( 
.A(n_1894),
.B(n_1582),
.C(n_1515),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_SL g1908 ( 
.A(n_1895),
.B(n_1627),
.Y(n_1908)
);

AND2x2_ASAP7_75t_L g1909 ( 
.A(n_1895),
.B(n_1745),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1896),
.Y(n_1910)
);

OAI211xp5_ASAP7_75t_SL g1911 ( 
.A1(n_1895),
.A2(n_1510),
.B(n_1600),
.C(n_1751),
.Y(n_1911)
);

XNOR2xp5_ASAP7_75t_L g1912 ( 
.A(n_1900),
.B(n_1612),
.Y(n_1912)
);

INVxp67_ASAP7_75t_L g1913 ( 
.A(n_1909),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1903),
.B(n_1642),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1901),
.Y(n_1915)
);

OAI21xp33_ASAP7_75t_L g1916 ( 
.A1(n_1905),
.A2(n_1627),
.B(n_1628),
.Y(n_1916)
);

OAI211xp5_ASAP7_75t_SL g1917 ( 
.A1(n_1902),
.A2(n_1746),
.B(n_1673),
.C(n_403),
.Y(n_1917)
);

OAI22xp5_ASAP7_75t_L g1918 ( 
.A1(n_1906),
.A2(n_1618),
.B1(n_1636),
.B2(n_1677),
.Y(n_1918)
);

OR2x2_ASAP7_75t_L g1919 ( 
.A(n_1908),
.B(n_1634),
.Y(n_1919)
);

AOI221xp5_ASAP7_75t_L g1920 ( 
.A1(n_1910),
.A2(n_1633),
.B1(n_1618),
.B2(n_1615),
.C(n_1636),
.Y(n_1920)
);

NOR2x1_ASAP7_75t_L g1921 ( 
.A(n_1904),
.B(n_1633),
.Y(n_1921)
);

AND2x2_ASAP7_75t_L g1922 ( 
.A(n_1907),
.B(n_1660),
.Y(n_1922)
);

NAND3xp33_ASAP7_75t_L g1923 ( 
.A(n_1911),
.B(n_399),
.C(n_401),
.Y(n_1923)
);

NOR3xp33_ASAP7_75t_L g1924 ( 
.A(n_1903),
.B(n_1665),
.C(n_406),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1909),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1909),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1909),
.B(n_404),
.Y(n_1927)
);

NOR2x1_ASAP7_75t_L g1928 ( 
.A(n_1915),
.B(n_408),
.Y(n_1928)
);

XOR2xp5_ASAP7_75t_SL g1929 ( 
.A(n_1921),
.B(n_409),
.Y(n_1929)
);

NOR3x1_ASAP7_75t_L g1930 ( 
.A(n_1923),
.B(n_410),
.C(n_412),
.Y(n_1930)
);

OR2x2_ASAP7_75t_L g1931 ( 
.A(n_1925),
.B(n_1615),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1926),
.Y(n_1932)
);

NAND3xp33_ASAP7_75t_SL g1933 ( 
.A(n_1927),
.B(n_413),
.C(n_415),
.Y(n_1933)
);

NOR2xp33_ASAP7_75t_L g1934 ( 
.A(n_1913),
.B(n_416),
.Y(n_1934)
);

NOR2x1_ASAP7_75t_L g1935 ( 
.A(n_1912),
.B(n_419),
.Y(n_1935)
);

NOR2xp67_ASAP7_75t_L g1936 ( 
.A(n_1914),
.B(n_420),
.Y(n_1936)
);

NOR2x1_ASAP7_75t_L g1937 ( 
.A(n_1922),
.B(n_423),
.Y(n_1937)
);

NOR2xp33_ASAP7_75t_L g1938 ( 
.A(n_1917),
.B(n_424),
.Y(n_1938)
);

NOR2xp33_ASAP7_75t_L g1939 ( 
.A(n_1919),
.B(n_426),
.Y(n_1939)
);

NOR3xp33_ASAP7_75t_L g1940 ( 
.A(n_1916),
.B(n_428),
.C(n_429),
.Y(n_1940)
);

NOR3xp33_ASAP7_75t_L g1941 ( 
.A(n_1924),
.B(n_431),
.C(n_432),
.Y(n_1941)
);

AND2x2_ASAP7_75t_SL g1942 ( 
.A(n_1920),
.B(n_433),
.Y(n_1942)
);

INVx1_ASAP7_75t_SL g1943 ( 
.A(n_1918),
.Y(n_1943)
);

NOR2x1_ASAP7_75t_L g1944 ( 
.A(n_1915),
.B(n_436),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1925),
.Y(n_1945)
);

OA21x2_ASAP7_75t_L g1946 ( 
.A1(n_1913),
.A2(n_437),
.B(n_438),
.Y(n_1946)
);

OR2x2_ASAP7_75t_L g1947 ( 
.A(n_1929),
.B(n_439),
.Y(n_1947)
);

AOI22xp5_ASAP7_75t_L g1948 ( 
.A1(n_1932),
.A2(n_440),
.B1(n_441),
.B2(n_442),
.Y(n_1948)
);

NOR2x1_ASAP7_75t_L g1949 ( 
.A(n_1945),
.B(n_445),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1928),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1944),
.Y(n_1951)
);

AOI222xp33_ASAP7_75t_L g1952 ( 
.A1(n_1936),
.A2(n_446),
.B1(n_448),
.B2(n_449),
.C1(n_451),
.C2(n_452),
.Y(n_1952)
);

OR2x2_ASAP7_75t_L g1953 ( 
.A(n_1943),
.B(n_454),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1937),
.Y(n_1954)
);

NAND2xp33_ASAP7_75t_R g1955 ( 
.A(n_1946),
.B(n_455),
.Y(n_1955)
);

INVx2_ASAP7_75t_L g1956 ( 
.A(n_1930),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1938),
.B(n_457),
.Y(n_1957)
);

XOR2x1_ASAP7_75t_L g1958 ( 
.A(n_1950),
.B(n_1946),
.Y(n_1958)
);

NAND2x1_ASAP7_75t_L g1959 ( 
.A(n_1956),
.B(n_1935),
.Y(n_1959)
);

NOR3xp33_ASAP7_75t_SL g1960 ( 
.A(n_1955),
.B(n_1939),
.C(n_1934),
.Y(n_1960)
);

AND3x4_ASAP7_75t_L g1961 ( 
.A(n_1949),
.B(n_1941),
.C(n_1940),
.Y(n_1961)
);

XOR2x2_ASAP7_75t_L g1962 ( 
.A(n_1947),
.B(n_1933),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1951),
.Y(n_1963)
);

OAI22xp5_ASAP7_75t_SL g1964 ( 
.A1(n_1954),
.A2(n_1957),
.B1(n_1953),
.B2(n_1942),
.Y(n_1964)
);

NOR2xp33_ASAP7_75t_L g1965 ( 
.A(n_1948),
.B(n_1931),
.Y(n_1965)
);

INVxp67_ASAP7_75t_L g1966 ( 
.A(n_1958),
.Y(n_1966)
);

AOI22xp5_ASAP7_75t_L g1967 ( 
.A1(n_1963),
.A2(n_1952),
.B1(n_459),
.B2(n_460),
.Y(n_1967)
);

INVx2_ASAP7_75t_L g1968 ( 
.A(n_1962),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1959),
.Y(n_1969)
);

XOR2xp5_ASAP7_75t_L g1970 ( 
.A(n_1968),
.B(n_1964),
.Y(n_1970)
);

AOI221xp5_ASAP7_75t_L g1971 ( 
.A1(n_1966),
.A2(n_1969),
.B1(n_1965),
.B2(n_1960),
.C(n_1967),
.Y(n_1971)
);

NOR2x1p5_ASAP7_75t_L g1972 ( 
.A(n_1969),
.B(n_1961),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1970),
.Y(n_1973)
);

NAND3xp33_ASAP7_75t_L g1974 ( 
.A(n_1971),
.B(n_458),
.C(n_462),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1973),
.B(n_1972),
.Y(n_1975)
);

CKINVDCx20_ASAP7_75t_R g1976 ( 
.A(n_1974),
.Y(n_1976)
);

NOR3xp33_ASAP7_75t_L g1977 ( 
.A(n_1975),
.B(n_465),
.C(n_466),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_L g1978 ( 
.A(n_1976),
.B(n_467),
.Y(n_1978)
);

HB1xp67_ASAP7_75t_L g1979 ( 
.A(n_1978),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1977),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_SL g1981 ( 
.A(n_1979),
.B(n_468),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1980),
.B(n_469),
.Y(n_1982)
);

OAI21x1_ASAP7_75t_SL g1983 ( 
.A1(n_1982),
.A2(n_470),
.B(n_473),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1981),
.Y(n_1984)
);

AOI21xp5_ASAP7_75t_L g1985 ( 
.A1(n_1981),
.A2(n_474),
.B(n_476),
.Y(n_1985)
);

OAI21xp5_ASAP7_75t_SL g1986 ( 
.A1(n_1981),
.A2(n_477),
.B(n_478),
.Y(n_1986)
);

AOI22x1_ASAP7_75t_L g1987 ( 
.A1(n_1981),
.A2(n_480),
.B1(n_481),
.B2(n_482),
.Y(n_1987)
);

INVx3_ASAP7_75t_L g1988 ( 
.A(n_1984),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1983),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1986),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1985),
.Y(n_1991)
);

OR2x6_ASAP7_75t_L g1992 ( 
.A(n_1988),
.B(n_1987),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_L g1993 ( 
.A(n_1989),
.B(n_484),
.Y(n_1993)
);

AOI221xp5_ASAP7_75t_L g1994 ( 
.A1(n_1990),
.A2(n_485),
.B1(n_486),
.B2(n_487),
.C(n_489),
.Y(n_1994)
);

AO21x2_ASAP7_75t_L g1995 ( 
.A1(n_1992),
.A2(n_1991),
.B(n_491),
.Y(n_1995)
);

AOI211xp5_ASAP7_75t_L g1996 ( 
.A1(n_1995),
.A2(n_1993),
.B(n_1994),
.C(n_493),
.Y(n_1996)
);


endmodule