module fake_jpeg_14032_n_482 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_482);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_482;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx8_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_13),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_10),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

BUFx16f_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_1),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_9),
.Y(n_52)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_9),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_7),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_11),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_17),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_57),
.B(n_65),
.Y(n_125)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_58),
.Y(n_189)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_59),
.Y(n_123)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_27),
.Y(n_60)
);

NAND2xp33_ASAP7_75t_SL g187 ( 
.A(n_60),
.B(n_95),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_61),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g140 ( 
.A(n_62),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_63),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_64),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_37),
.B(n_16),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_66),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_67),
.Y(n_181)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_68),
.Y(n_126)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_69),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_70),
.Y(n_190)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_71),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_22),
.B(n_16),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_72),
.B(n_74),
.Y(n_127)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_20),
.Y(n_73)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_73),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_22),
.B(n_16),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g133 ( 
.A(n_75),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_76),
.Y(n_191)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_28),
.Y(n_77)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_77),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_78),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_30),
.Y(n_79)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_79),
.Y(n_151)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_18),
.Y(n_80)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_80),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_42),
.Y(n_81)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_81),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_29),
.Y(n_82)
);

BUFx2_ASAP7_75t_SL g171 ( 
.A(n_82),
.Y(n_171)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_26),
.Y(n_83)
);

INVx11_ASAP7_75t_L g178 ( 
.A(n_83),
.Y(n_178)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_21),
.Y(n_84)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_84),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_50),
.B(n_15),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_85),
.B(n_96),
.Y(n_128)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_18),
.Y(n_86)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_86),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_87),
.Y(n_182)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_35),
.Y(n_88)
);

INVx3_ASAP7_75t_SL g166 ( 
.A(n_88),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

INVx8_ASAP7_75t_L g183 ( 
.A(n_89),
.Y(n_183)
);

INVx3_ASAP7_75t_SL g90 ( 
.A(n_53),
.Y(n_90)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_90),
.Y(n_138)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_21),
.Y(n_91)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_91),
.Y(n_169)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_35),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_92),
.Y(n_149)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_26),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_93),
.Y(n_164)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_18),
.Y(n_94)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_94),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_30),
.Y(n_96)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_47),
.Y(n_97)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_97),
.Y(n_153)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_30),
.Y(n_98)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_98),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_47),
.Y(n_99)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_99),
.Y(n_160)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_35),
.Y(n_100)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_100),
.Y(n_162)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_23),
.Y(n_101)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_101),
.Y(n_174)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_30),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_102),
.B(n_107),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_49),
.Y(n_103)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_103),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_19),
.B(n_15),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_104),
.B(n_111),
.Y(n_147)
);

INVx13_ASAP7_75t_L g105 ( 
.A(n_26),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_105),
.Y(n_150)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_24),
.Y(n_106)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_106),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_50),
.B(n_15),
.Y(n_107)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_24),
.Y(n_108)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_108),
.Y(n_177)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_23),
.Y(n_109)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_109),
.Y(n_176)
);

BUFx5_ASAP7_75t_L g110 ( 
.A(n_44),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_56),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_28),
.B(n_13),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_24),
.Y(n_112)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_112),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_49),
.Y(n_113)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_113),
.Y(n_179)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_24),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_114),
.B(n_116),
.Y(n_188)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_24),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_115),
.B(n_117),
.Y(n_157)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_46),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_33),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_46),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_118),
.B(n_52),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_97),
.A2(n_113),
.B1(n_103),
.B2(n_61),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_119),
.A2(n_121),
.B1(n_122),
.B2(n_144),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_63),
.A2(n_53),
.B1(n_49),
.B2(n_44),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_90),
.A2(n_38),
.B1(n_28),
.B2(n_53),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_134),
.Y(n_204)
);

OAI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_64),
.A2(n_44),
.B1(n_49),
.B2(n_38),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_137),
.A2(n_156),
.B1(n_163),
.B2(n_167),
.Y(n_218)
);

AND2x2_ASAP7_75t_SL g142 ( 
.A(n_79),
.B(n_33),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_142),
.B(n_5),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_79),
.A2(n_56),
.B1(n_33),
.B2(n_38),
.Y(n_144)
);

A2O1A1Ixp33_ASAP7_75t_L g148 ( 
.A1(n_72),
.A2(n_34),
.B(n_54),
.C(n_25),
.Y(n_148)
);

A2O1A1Ixp33_ASAP7_75t_L g253 ( 
.A1(n_148),
.A2(n_178),
.B(n_140),
.C(n_146),
.Y(n_253)
);

NOR2x1_ASAP7_75t_L g152 ( 
.A(n_60),
.B(n_34),
.Y(n_152)
);

NOR3xp33_ASAP7_75t_L g238 ( 
.A(n_152),
.B(n_171),
.C(n_131),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_96),
.A2(n_33),
.B1(n_54),
.B2(n_51),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_155),
.A2(n_159),
.B1(n_173),
.B2(n_4),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_85),
.A2(n_55),
.B1(n_19),
.B2(n_36),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_158),
.B(n_125),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_96),
.A2(n_33),
.B1(n_51),
.B2(n_48),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_67),
.A2(n_52),
.B1(n_31),
.B2(n_48),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_161),
.A2(n_192),
.B1(n_10),
.B2(n_121),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_107),
.A2(n_55),
.B1(n_41),
.B2(n_36),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_74),
.A2(n_41),
.B1(n_43),
.B2(n_40),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_88),
.B(n_43),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_168),
.B(n_175),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_102),
.A2(n_100),
.B1(n_92),
.B2(n_39),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_102),
.B(n_40),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_70),
.A2(n_39),
.B1(n_31),
.B2(n_25),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g249 ( 
.A1(n_180),
.A2(n_145),
.B1(n_181),
.B2(n_164),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_76),
.B(n_12),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_186),
.B(n_149),
.Y(n_227)
);

OAI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_78),
.A2(n_46),
.B1(n_1),
.B2(n_2),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_120),
.Y(n_193)
);

INVx5_ASAP7_75t_L g294 ( 
.A(n_193),
.Y(n_294)
);

NAND3xp33_ASAP7_75t_L g194 ( 
.A(n_147),
.B(n_12),
.C(n_2),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_194),
.B(n_205),
.Y(n_282)
);

AOI21xp33_ASAP7_75t_L g195 ( 
.A1(n_127),
.A2(n_12),
.B(n_46),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_195),
.B(n_198),
.Y(n_274)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_153),
.Y(n_196)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_196),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_148),
.B(n_0),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_197),
.B(n_200),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_132),
.B(n_81),
.C(n_99),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_199),
.B(n_219),
.C(n_217),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_127),
.B(n_2),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_169),
.B(n_4),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_201),
.B(n_206),
.Y(n_263)
);

OAI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_134),
.A2(n_87),
.B1(n_89),
.B2(n_105),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_202),
.A2(n_222),
.B1(n_231),
.B2(n_235),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_203),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_188),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_174),
.B(n_4),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_154),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_207),
.Y(n_297)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_160),
.Y(n_208)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_208),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_176),
.B(n_4),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_209),
.B(n_212),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_142),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_210),
.B(n_211),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_123),
.B(n_5),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_124),
.B(n_5),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_133),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_213),
.B(n_214),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_128),
.B(n_170),
.Y(n_214)
);

BUFx2_ASAP7_75t_L g215 ( 
.A(n_183),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_215),
.Y(n_267)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_151),
.Y(n_216)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_216),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_217),
.B(n_225),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_157),
.B(n_5),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_152),
.B(n_9),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_220),
.B(n_221),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_161),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_150),
.B(n_10),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_223),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_119),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_224),
.B(n_228),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_126),
.B(n_130),
.Y(n_225)
);

AOI21xp33_ASAP7_75t_L g226 ( 
.A1(n_187),
.A2(n_149),
.B(n_133),
.Y(n_226)
);

OR2x2_ASAP7_75t_L g303 ( 
.A(n_226),
.B(n_227),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_166),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_172),
.B(n_185),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_229),
.B(n_242),
.Y(n_298)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_138),
.Y(n_230)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_230),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_144),
.A2(n_137),
.B1(n_173),
.B2(n_155),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_179),
.Y(n_232)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_232),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_159),
.Y(n_233)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_233),
.Y(n_279)
);

AND2x4_ASAP7_75t_SL g234 ( 
.A(n_135),
.B(n_136),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_234),
.B(n_240),
.Y(n_302)
);

OAI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_192),
.A2(n_162),
.B1(n_166),
.B2(n_139),
.Y(n_235)
);

INVx5_ASAP7_75t_L g236 ( 
.A(n_151),
.Y(n_236)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_236),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_120),
.Y(n_237)
);

INVx8_ASAP7_75t_L g259 ( 
.A(n_237),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_238),
.A2(n_250),
.B(n_213),
.Y(n_264)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_165),
.Y(n_239)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_239),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_184),
.B(n_189),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_141),
.A2(n_182),
.B1(n_143),
.B2(n_191),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_241),
.A2(n_244),
.B1(n_255),
.B2(n_243),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_177),
.B(n_183),
.Y(n_242)
);

AND2x4_ASAP7_75t_L g243 ( 
.A(n_184),
.B(n_129),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_243),
.A2(n_228),
.B(n_250),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_141),
.A2(n_182),
.B1(n_143),
.B2(n_190),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_146),
.B(n_129),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_246),
.Y(n_257)
);

AO22x1_ASAP7_75t_SL g247 ( 
.A1(n_131),
.A2(n_191),
.B1(n_145),
.B2(n_190),
.Y(n_247)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_247),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_249),
.A2(n_224),
.B1(n_221),
.B2(n_204),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_140),
.B(n_178),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_140),
.Y(n_251)
);

INVx11_ASAP7_75t_L g275 ( 
.A(n_251),
.Y(n_275)
);

INVx6_ASAP7_75t_L g252 ( 
.A(n_181),
.Y(n_252)
);

INVx8_ASAP7_75t_L g299 ( 
.A(n_252),
.Y(n_299)
);

A2O1A1Ixp33_ASAP7_75t_L g276 ( 
.A1(n_253),
.A2(n_217),
.B(n_197),
.C(n_204),
.Y(n_276)
);

AO22x1_ASAP7_75t_SL g254 ( 
.A1(n_137),
.A2(n_192),
.B1(n_126),
.B2(n_130),
.Y(n_254)
);

O2A1O1Ixp33_ASAP7_75t_SL g289 ( 
.A1(n_254),
.A2(n_241),
.B(n_244),
.C(n_219),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_121),
.A2(n_119),
.B1(n_122),
.B2(n_168),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_258),
.B(n_293),
.Y(n_315)
);

BUFx5_ASAP7_75t_L g262 ( 
.A(n_193),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_264),
.A2(n_215),
.B(n_237),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_242),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_272),
.B(n_265),
.Y(n_322)
);

O2A1O1Ixp33_ASAP7_75t_L g305 ( 
.A1(n_276),
.A2(n_243),
.B(n_247),
.C(n_251),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_L g320 ( 
.A1(n_278),
.A2(n_291),
.B1(n_302),
.B2(n_280),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_218),
.A2(n_233),
.B1(n_254),
.B2(n_248),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_280),
.A2(n_283),
.B1(n_285),
.B2(n_243),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_218),
.A2(n_254),
.B1(n_255),
.B2(n_245),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_284),
.A2(n_290),
.B(n_236),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_227),
.A2(n_222),
.B1(n_231),
.B2(n_199),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_229),
.B(n_200),
.C(n_205),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_287),
.B(n_292),
.Y(n_310)
);

OA22x2_ASAP7_75t_L g337 ( 
.A1(n_289),
.A2(n_296),
.B1(n_276),
.B2(n_261),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_253),
.A2(n_219),
.B(n_201),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_234),
.B(n_230),
.C(n_206),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_234),
.B(n_212),
.C(n_209),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_271),
.A2(n_247),
.B1(n_232),
.B2(n_196),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_304),
.A2(n_329),
.B1(n_260),
.B2(n_300),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_305),
.B(n_312),
.Y(n_355)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_281),
.Y(n_306)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_306),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_307),
.A2(n_314),
.B1(n_320),
.B2(n_325),
.Y(n_353)
);

INVx13_ASAP7_75t_L g308 ( 
.A(n_275),
.Y(n_308)
);

INVx1_ASAP7_75t_SL g367 ( 
.A(n_308),
.Y(n_367)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_281),
.Y(n_309)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_309),
.Y(n_342)
);

OR2x2_ASAP7_75t_L g311 ( 
.A(n_290),
.B(n_216),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_311),
.B(n_322),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_275),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_313),
.B(n_317),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_283),
.A2(n_208),
.B1(n_239),
.B2(n_252),
.Y(n_314)
);

INVx1_ASAP7_75t_SL g316 ( 
.A(n_302),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_316),
.B(n_327),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_257),
.B(n_215),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_277),
.Y(n_318)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_318),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_319),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_286),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_321),
.B(n_324),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_257),
.B(n_301),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_323),
.B(n_326),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_256),
.B(n_274),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_285),
.A2(n_291),
.B1(n_278),
.B2(n_272),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_263),
.B(n_265),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_295),
.B(n_287),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_263),
.B(n_298),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_328),
.B(n_332),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_271),
.A2(n_296),
.B1(n_298),
.B2(n_273),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_277),
.Y(n_330)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_330),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_289),
.A2(n_279),
.B1(n_302),
.B2(n_256),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_331),
.A2(n_336),
.B1(n_282),
.B2(n_267),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_293),
.B(n_258),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_261),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_333),
.B(n_337),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_297),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_334),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_292),
.B(n_266),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_335),
.B(n_266),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_289),
.A2(n_279),
.B1(n_266),
.B2(n_284),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_260),
.Y(n_338)
);

AOI22xp33_ASAP7_75t_L g348 ( 
.A1(n_338),
.A2(n_339),
.B1(n_300),
.B2(n_268),
.Y(n_348)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_268),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_SL g373 ( 
.A(n_344),
.B(n_310),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_346),
.A2(n_350),
.B1(n_354),
.B2(n_366),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_336),
.A2(n_303),
.B(n_264),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_L g374 ( 
.A1(n_347),
.A2(n_311),
.B(n_327),
.Y(n_374)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_348),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_329),
.A2(n_303),
.B1(n_299),
.B2(n_259),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_332),
.B(n_288),
.C(n_270),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_351),
.B(n_365),
.C(n_311),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_304),
.A2(n_299),
.B1(n_259),
.B2(n_294),
.Y(n_354)
);

OA21x2_ASAP7_75t_L g358 ( 
.A1(n_307),
.A2(n_269),
.B(n_270),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_358),
.B(n_337),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_360),
.A2(n_364),
.B1(n_369),
.B2(n_305),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_325),
.A2(n_314),
.B1(n_309),
.B2(n_306),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_315),
.B(n_269),
.C(n_267),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_305),
.A2(n_262),
.B1(n_294),
.B2(n_316),
.Y(n_366)
);

MAJx2_ASAP7_75t_L g368 ( 
.A(n_315),
.B(n_310),
.C(n_335),
.Y(n_368)
);

MAJx2_ASAP7_75t_L g387 ( 
.A(n_368),
.B(n_337),
.C(n_318),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_331),
.A2(n_322),
.B1(n_312),
.B2(n_337),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_343),
.Y(n_371)
);

OAI22xp33_ASAP7_75t_SL g412 ( 
.A1(n_371),
.A2(n_367),
.B1(n_363),
.B2(n_345),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_349),
.B(n_321),
.Y(n_372)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_372),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_374),
.A2(n_355),
.B(n_341),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_349),
.B(n_328),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_375),
.B(n_376),
.C(n_380),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_368),
.B(n_326),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_361),
.B(n_352),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_377),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_378),
.A2(n_385),
.B1(n_389),
.B2(n_393),
.Y(n_399)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_379),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_344),
.B(n_359),
.C(n_365),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_381),
.B(n_384),
.C(n_386),
.Y(n_397)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_345),
.Y(n_382)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_382),
.Y(n_406)
);

CKINVDCx16_ASAP7_75t_R g383 ( 
.A(n_356),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_383),
.B(n_388),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_359),
.B(n_323),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_SL g385 ( 
.A(n_352),
.B(n_324),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_359),
.B(n_337),
.C(n_319),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_343),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_341),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_351),
.B(n_334),
.Y(n_390)
);

NAND2xp33_ASAP7_75t_R g413 ( 
.A(n_390),
.B(n_363),
.Y(n_413)
);

INVx1_ASAP7_75t_SL g391 ( 
.A(n_355),
.Y(n_391)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_391),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_340),
.B(n_339),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_378),
.A2(n_350),
.B1(n_357),
.B2(n_347),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_400),
.B(n_410),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_392),
.A2(n_353),
.B1(n_369),
.B2(n_362),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_401),
.A2(n_408),
.B1(n_386),
.B2(n_389),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_403),
.B(n_413),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_373),
.B(n_355),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_404),
.B(n_405),
.C(n_407),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_381),
.B(n_342),
.C(n_340),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_376),
.B(n_362),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_392),
.A2(n_362),
.B1(n_357),
.B2(n_358),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_384),
.B(n_342),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_409),
.B(n_380),
.C(n_374),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_379),
.A2(n_346),
.B1(n_366),
.B2(n_354),
.Y(n_410)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_412),
.Y(n_419)
);

AOI22x1_ASAP7_75t_L g436 ( 
.A1(n_414),
.A2(n_400),
.B1(n_410),
.B2(n_408),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_394),
.B(n_385),
.Y(n_415)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_415),
.Y(n_431)
);

INVx2_ASAP7_75t_SL g417 ( 
.A(n_406),
.Y(n_417)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_417),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_402),
.B(n_375),
.Y(n_418)
);

CKINVDCx16_ASAP7_75t_R g443 ( 
.A(n_418),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_395),
.B(n_388),
.Y(n_420)
);

AO221x1_ASAP7_75t_L g433 ( 
.A1(n_420),
.A2(n_382),
.B1(n_333),
.B2(n_411),
.C(n_370),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_395),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_421),
.B(n_425),
.Y(n_441)
);

CKINVDCx14_ASAP7_75t_R g424 ( 
.A(n_399),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_424),
.B(n_430),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_406),
.Y(n_425)
);

INVx1_ASAP7_75t_SL g426 ( 
.A(n_398),
.Y(n_426)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_426),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_398),
.B(n_371),
.Y(n_427)
);

HB1xp67_ASAP7_75t_L g442 ( 
.A(n_427),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_428),
.B(n_397),
.C(n_396),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_401),
.A2(n_391),
.B1(n_370),
.B2(n_387),
.Y(n_429)
);

BUFx2_ASAP7_75t_L g432 ( 
.A(n_429),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_405),
.B(n_330),
.Y(n_430)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_433),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_436),
.B(n_422),
.Y(n_446)
);

NOR2xp67_ASAP7_75t_SL g452 ( 
.A(n_438),
.B(n_423),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_423),
.B(n_397),
.C(n_396),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_439),
.B(n_438),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_421),
.B(n_409),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_SL g449 ( 
.A(n_440),
.B(n_416),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g444 ( 
.A1(n_441),
.A2(n_416),
.B(n_427),
.Y(n_444)
);

AOI21xp5_ASAP7_75t_L g454 ( 
.A1(n_444),
.A2(n_447),
.B(n_452),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_445),
.B(n_448),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_SL g460 ( 
.A1(n_446),
.A2(n_422),
.B(n_444),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_SL g447 ( 
.A1(n_439),
.A2(n_403),
.B(n_428),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_431),
.B(n_419),
.Y(n_448)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_449),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_434),
.B(n_419),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_450),
.B(n_443),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_SL g451 ( 
.A(n_432),
.B(n_404),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_451),
.B(n_429),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_451),
.B(n_414),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_455),
.B(n_457),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_456),
.B(n_461),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_446),
.B(n_432),
.C(n_436),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_460),
.B(n_441),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_453),
.B(n_442),
.Y(n_461)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_462),
.Y(n_466)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_464),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_SL g465 ( 
.A1(n_454),
.A2(n_437),
.B(n_435),
.Y(n_465)
);

AOI21xp5_ASAP7_75t_L g472 ( 
.A1(n_465),
.A2(n_467),
.B(n_457),
.Y(n_472)
);

AOI21xp33_ASAP7_75t_L g467 ( 
.A1(n_458),
.A2(n_459),
.B(n_437),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_455),
.B(n_425),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_468),
.B(n_417),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_470),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_469),
.B(n_463),
.Y(n_471)
);

INVxp33_ASAP7_75t_L g474 ( 
.A(n_471),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_472),
.B(n_466),
.C(n_464),
.Y(n_475)
);

OAI21xp5_ASAP7_75t_SL g478 ( 
.A1(n_475),
.A2(n_460),
.B(n_471),
.Y(n_478)
);

OAI21xp33_ASAP7_75t_L g477 ( 
.A1(n_474),
.A2(n_473),
.B(n_476),
.Y(n_477)
);

AOI21x1_ASAP7_75t_L g479 ( 
.A1(n_477),
.A2(n_478),
.B(n_435),
.Y(n_479)
);

AO21x1_ASAP7_75t_L g480 ( 
.A1(n_479),
.A2(n_411),
.B(n_417),
.Y(n_480)
);

AOI221xp5_ASAP7_75t_L g481 ( 
.A1(n_480),
.A2(n_313),
.B1(n_426),
.B2(n_436),
.C(n_338),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_481),
.B(n_358),
.Y(n_482)
);


endmodule