module fake_jpeg_24186_n_179 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_179);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_179;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx2_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_35),
.B(n_37),
.Y(n_64)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_39),
.Y(n_48)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_0),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_41),
.Y(n_51)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_16),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_19),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_37),
.A2(n_26),
.B1(n_32),
.B2(n_25),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_44),
.A2(n_45),
.B1(n_47),
.B2(n_50),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_35),
.A2(n_26),
.B1(n_18),
.B2(n_27),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_57),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_41),
.A2(n_25),
.B1(n_23),
.B2(n_18),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_40),
.A2(n_25),
.B1(n_23),
.B2(n_18),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_27),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_53),
.B(n_58),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_L g54 ( 
.A1(n_36),
.A2(n_18),
.B1(n_23),
.B2(n_21),
.Y(n_54)
);

OA22x2_ASAP7_75t_L g69 ( 
.A1(n_54),
.A2(n_61),
.B1(n_20),
.B2(n_16),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_55),
.B(n_62),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_40),
.A2(n_18),
.B1(n_30),
.B2(n_22),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_33),
.B(n_31),
.C(n_28),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_43),
.A2(n_31),
.B1(n_28),
.B2(n_29),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_33),
.B(n_19),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_34),
.B(n_0),
.Y(n_63)
);

A2O1A1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_63),
.A2(n_20),
.B(n_22),
.C(n_24),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_65),
.Y(n_94)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_64),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_66),
.B(n_80),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_69),
.A2(n_59),
.B1(n_56),
.B2(n_21),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_70),
.B(n_73),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_24),
.Y(n_72)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_48),
.B(n_30),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_51),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_78),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_53),
.B(n_29),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_79),
.B(n_15),
.Y(n_102)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_82),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_58),
.B(n_21),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_42),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_83),
.B(n_84),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_42),
.Y(n_84)
);

NOR3xp33_ASAP7_75t_L g86 ( 
.A(n_81),
.B(n_57),
.C(n_45),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_86),
.B(n_101),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_51),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_95),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_83),
.B(n_34),
.C(n_38),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_89),
.B(n_98),
.C(n_68),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_67),
.A2(n_56),
.B(n_46),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_90),
.A2(n_97),
.B(n_79),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_84),
.B(n_42),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_77),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_38),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_74),
.B(n_38),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_96),
.B(n_69),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_76),
.B(n_80),
.C(n_66),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_75),
.B(n_59),
.Y(n_101)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_103),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_105),
.B(n_107),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_113),
.C(n_118),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_100),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_95),
.B(n_69),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_108),
.B(n_92),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_99),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_109),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_110),
.A2(n_94),
.B1(n_91),
.B2(n_93),
.Y(n_135)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_103),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_111),
.B(n_112),
.Y(n_136)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_98),
.Y(n_112)
);

NOR4xp25_ASAP7_75t_L g114 ( 
.A(n_85),
.B(n_69),
.C(n_73),
.D(n_70),
.Y(n_114)
);

A2O1A1O1Ixp25_ASAP7_75t_L g134 ( 
.A1(n_114),
.A2(n_117),
.B(n_102),
.C(n_60),
.D(n_49),
.Y(n_134)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_88),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_116),
.B(n_120),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_96),
.A2(n_34),
.B(n_77),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_65),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_119),
.B(n_94),
.Y(n_131)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_121),
.A2(n_134),
.B(n_135),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_116),
.B(n_85),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_125),
.B(n_129),
.Y(n_148)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_104),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_126),
.B(n_133),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_118),
.B(n_89),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_127),
.B(n_128),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_104),
.B(n_90),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_112),
.B(n_87),
.Y(n_129)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_131),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_87),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_1),
.Y(n_145)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_109),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_108),
.B(n_93),
.Y(n_137)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_137),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_137),
.A2(n_113),
.B1(n_120),
.B2(n_108),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_138),
.A2(n_78),
.B1(n_71),
.B2(n_4),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_135),
.A2(n_110),
.B1(n_115),
.B2(n_107),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_139),
.A2(n_136),
.B1(n_130),
.B2(n_121),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_123),
.A2(n_133),
.B(n_126),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_141),
.A2(n_124),
.B(n_129),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_145),
.B(n_128),
.Y(n_150)
);

BUFx2_ASAP7_75t_L g146 ( 
.A(n_122),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g151 ( 
.A(n_146),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_149),
.A2(n_155),
.B(n_156),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_150),
.B(n_153),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_152),
.A2(n_138),
.B1(n_148),
.B2(n_139),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_143),
.B(n_127),
.C(n_130),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_143),
.B(n_132),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_154),
.B(n_157),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_142),
.B(n_121),
.C(n_91),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_144),
.B(n_65),
.C(n_78),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_156),
.A2(n_147),
.B(n_144),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_158),
.A2(n_155),
.B(n_140),
.Y(n_166)
);

MAJx2_ASAP7_75t_L g160 ( 
.A(n_154),
.B(n_145),
.C(n_148),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_160),
.B(n_162),
.C(n_150),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_149),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_163),
.B(n_159),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_165),
.B(n_168),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_166),
.B(n_167),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_164),
.B(n_153),
.C(n_152),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_161),
.B(n_146),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_169),
.B(n_170),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_161),
.B(n_151),
.C(n_3),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_165),
.A2(n_2),
.B1(n_3),
.B2(n_6),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_172),
.B(n_174),
.C(n_171),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_175),
.B(n_176),
.C(n_173),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_171),
.B(n_7),
.C(n_8),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_177),
.A2(n_9),
.B(n_10),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_178),
.B(n_10),
.Y(n_179)
);


endmodule