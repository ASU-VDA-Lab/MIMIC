module real_aes_807_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_547;
wire n_454;
wire n_122;
wire n_443;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_527;
wire n_502;
wire n_434;
wire n_505;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_87;
wire n_171;
wire n_531;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_501;
wire n_488;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_536;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_456;
wire n_359;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
NAND2xp5_ASAP7_75t_SL g294 ( .A(n_0), .B(n_221), .Y(n_294) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_1), .A2(n_229), .B(n_234), .Y(n_228) );
AOI22xp33_ASAP7_75t_SL g124 ( .A1(n_2), .A2(n_4), .B1(n_125), .B2(n_130), .Y(n_124) );
AO22x2_ASAP7_75t_L g96 ( .A1(n_3), .A2(n_55), .B1(n_93), .B2(n_97), .Y(n_96) );
NAND2xp5_ASAP7_75t_SL g275 ( .A(n_5), .B(n_236), .Y(n_275) );
INVx1_ASAP7_75t_L g202 ( .A(n_6), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_7), .B(n_236), .Y(n_326) );
AO22x2_ASAP7_75t_L g92 ( .A1(n_8), .A2(n_25), .B1(n_93), .B2(n_94), .Y(n_92) );
AOI22xp33_ASAP7_75t_L g135 ( .A1(n_9), .A2(n_40), .B1(n_136), .B2(n_140), .Y(n_135) );
NAND2xp33_ASAP7_75t_L g318 ( .A(n_10), .B(n_238), .Y(n_318) );
INVx2_ASAP7_75t_L g218 ( .A(n_11), .Y(n_218) );
AOI221x1_ASAP7_75t_L g260 ( .A1(n_12), .A2(n_20), .B1(n_221), .B2(n_229), .C(n_261), .Y(n_260) );
INVx1_ASAP7_75t_L g549 ( .A(n_12), .Y(n_549) );
NAND2xp5_ASAP7_75t_SL g314 ( .A(n_13), .B(n_221), .Y(n_314) );
AO21x2_ASAP7_75t_L g311 ( .A1(n_14), .A2(n_312), .B(n_313), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_15), .B(n_240), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_16), .B(n_236), .Y(n_249) );
AO21x1_ASAP7_75t_L g270 ( .A1(n_17), .A2(n_221), .B(n_271), .Y(n_270) );
INVx1_ASAP7_75t_L g180 ( .A(n_18), .Y(n_180) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_19), .Y(n_122) );
OAI22xp5_ASAP7_75t_SL g183 ( .A1(n_21), .A2(n_184), .B1(n_187), .B2(n_188), .Y(n_183) );
INVx1_ASAP7_75t_L g188 ( .A(n_21), .Y(n_188) );
NAND2x1_ASAP7_75t_L g292 ( .A(n_22), .B(n_236), .Y(n_292) );
NAND2x1_ASAP7_75t_L g325 ( .A(n_23), .B(n_238), .Y(n_325) );
AOI22xp33_ASAP7_75t_L g153 ( .A1(n_24), .A2(n_74), .B1(n_154), .B2(n_158), .Y(n_153) );
OAI221xp5_ASAP7_75t_L g194 ( .A1(n_25), .A2(n_55), .B1(n_62), .B2(n_195), .C(n_197), .Y(n_194) );
OA21x2_ASAP7_75t_L g217 ( .A1(n_26), .A2(n_68), .B(n_218), .Y(n_217) );
OR2x2_ASAP7_75t_L g242 ( .A(n_26), .B(n_68), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_27), .B(n_238), .Y(n_237) );
INVx3_ASAP7_75t_L g93 ( .A(n_28), .Y(n_93) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_29), .B(n_236), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_30), .B(n_238), .Y(n_274) );
AOI22xp33_ASAP7_75t_L g146 ( .A1(n_31), .A2(n_57), .B1(n_147), .B2(n_149), .Y(n_146) );
AOI21xp5_ASAP7_75t_L g280 ( .A1(n_32), .A2(n_229), .B(n_281), .Y(n_280) );
INVx1_ASAP7_75t_SL g101 ( .A(n_33), .Y(n_101) );
INVx1_ASAP7_75t_L g204 ( .A(n_34), .Y(n_204) );
AND2x2_ASAP7_75t_L g227 ( .A(n_34), .B(n_202), .Y(n_227) );
AND2x2_ASAP7_75t_L g230 ( .A(n_34), .B(n_231), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g284 ( .A(n_35), .B(n_221), .Y(n_284) );
CKINVDCx20_ASAP7_75t_R g253 ( .A(n_36), .Y(n_253) );
OAI22xp5_ASAP7_75t_L g184 ( .A1(n_37), .A2(n_69), .B1(n_185), .B2(n_186), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_37), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_37), .B(n_238), .Y(n_282) );
AOI22xp5_ASAP7_75t_L g80 ( .A1(n_38), .A2(n_81), .B1(n_82), .B2(n_174), .Y(n_80) );
CKINVDCx16_ASAP7_75t_R g174 ( .A(n_38), .Y(n_174) );
AOI22xp33_ASAP7_75t_L g169 ( .A1(n_39), .A2(n_47), .B1(n_170), .B2(n_173), .Y(n_169) );
AOI21xp5_ASAP7_75t_L g323 ( .A1(n_41), .A2(n_229), .B(n_324), .Y(n_323) );
AO22x2_ASAP7_75t_L g104 ( .A1(n_42), .A2(n_62), .B1(n_93), .B2(n_105), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_43), .B(n_238), .Y(n_293) );
INVx1_ASAP7_75t_L g224 ( .A(n_44), .Y(n_224) );
INVx1_ASAP7_75t_L g233 ( .A(n_44), .Y(n_233) );
INVx1_ASAP7_75t_L g102 ( .A(n_45), .Y(n_102) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_46), .B(n_236), .Y(n_263) );
AOI22xp5_ASAP7_75t_L g176 ( .A1(n_48), .A2(n_177), .B1(n_178), .B2(n_182), .Y(n_176) );
INVx1_ASAP7_75t_L g182 ( .A(n_48), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g290 ( .A1(n_49), .A2(n_229), .B(n_291), .Y(n_290) );
OAI22xp5_ASAP7_75t_SL g178 ( .A1(n_50), .A2(n_179), .B1(n_180), .B2(n_181), .Y(n_178) );
INVx1_ASAP7_75t_L g181 ( .A(n_50), .Y(n_181) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_51), .Y(n_115) );
AO21x1_ASAP7_75t_L g272 ( .A1(n_52), .A2(n_229), .B(n_273), .Y(n_272) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_53), .B(n_221), .Y(n_220) );
NAND2xp5_ASAP7_75t_SL g327 ( .A(n_54), .B(n_221), .Y(n_327) );
INVxp33_ASAP7_75t_L g199 ( .A(n_55), .Y(n_199) );
AOI22xp33_ASAP7_75t_L g162 ( .A1(n_56), .A2(n_63), .B1(n_163), .B2(n_166), .Y(n_162) );
AND2x2_ASAP7_75t_L g286 ( .A(n_58), .B(n_241), .Y(n_286) );
AOI22xp5_ASAP7_75t_L g536 ( .A1(n_59), .A2(n_81), .B1(n_82), .B2(n_537), .Y(n_536) );
CKINVDCx20_ASAP7_75t_R g537 ( .A(n_59), .Y(n_537) );
INVx1_ASAP7_75t_L g226 ( .A(n_60), .Y(n_226) );
INVx1_ASAP7_75t_L g231 ( .A(n_60), .Y(n_231) );
AND2x2_ASAP7_75t_L g329 ( .A(n_61), .B(n_215), .Y(n_329) );
INVxp67_ASAP7_75t_L g198 ( .A(n_62), .Y(n_198) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_64), .Y(n_106) );
AND2x2_ASAP7_75t_L g214 ( .A(n_65), .B(n_215), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g251 ( .A(n_66), .B(n_221), .Y(n_251) );
AND2x2_ASAP7_75t_L g271 ( .A(n_67), .B(n_245), .Y(n_271) );
INVx1_ASAP7_75t_L g186 ( .A(n_69), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_69), .B(n_238), .Y(n_250) );
AND2x2_ASAP7_75t_L g295 ( .A(n_70), .B(n_215), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_71), .B(n_236), .Y(n_283) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_72), .A2(n_229), .B(n_248), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_73), .B(n_238), .Y(n_262) );
AOI22xp5_ASAP7_75t_L g528 ( .A1(n_73), .A2(n_81), .B1(n_82), .B2(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_73), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_75), .B(n_236), .Y(n_235) );
BUFx2_ASAP7_75t_SL g196 ( .A(n_76), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g315 ( .A1(n_77), .A2(n_229), .B(n_316), .Y(n_315) );
AOI221xp5_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_191), .B1(n_205), .B2(n_525), .C(n_527), .Y(n_78) );
XNOR2xp5_ASAP7_75t_L g79 ( .A(n_80), .B(n_175), .Y(n_79) );
CKINVDCx16_ASAP7_75t_R g81 ( .A(n_82), .Y(n_81) );
HB1xp67_ASAP7_75t_L g82 ( .A(n_83), .Y(n_82) );
NAND2xp5_ASAP7_75t_SL g83 ( .A(n_84), .B(n_144), .Y(n_83) );
NOR2x1_ASAP7_75t_L g84 ( .A(n_85), .B(n_123), .Y(n_84) );
OAI222xp33_ASAP7_75t_L g85 ( .A1(n_86), .A2(n_106), .B1(n_107), .B2(n_115), .C1(n_116), .C2(n_122), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
HB1xp67_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
INVx2_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
INVx2_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
AND2x2_ASAP7_75t_L g90 ( .A(n_91), .B(n_98), .Y(n_90) );
AND2x4_ASAP7_75t_L g137 ( .A(n_91), .B(n_138), .Y(n_137) );
AND2x4_ASAP7_75t_L g168 ( .A(n_91), .B(n_152), .Y(n_168) );
AND2x4_ASAP7_75t_L g91 ( .A(n_92), .B(n_95), .Y(n_91) );
INVx1_ASAP7_75t_L g114 ( .A(n_92), .Y(n_114) );
AND2x2_ASAP7_75t_L g120 ( .A(n_92), .B(n_96), .Y(n_120) );
INVx1_ASAP7_75t_L g129 ( .A(n_92), .Y(n_129) );
INVx2_ASAP7_75t_L g94 ( .A(n_93), .Y(n_94) );
INVx1_ASAP7_75t_L g97 ( .A(n_93), .Y(n_97) );
OAI22x1_ASAP7_75t_L g99 ( .A1(n_93), .A2(n_100), .B1(n_101), .B2(n_102), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_93), .Y(n_100) );
INVx1_ASAP7_75t_L g105 ( .A(n_93), .Y(n_105) );
AND2x4_ASAP7_75t_L g113 ( .A(n_95), .B(n_114), .Y(n_113) );
INVxp67_ASAP7_75t_L g143 ( .A(n_95), .Y(n_143) );
INVx2_ASAP7_75t_L g95 ( .A(n_96), .Y(n_95) );
AND2x2_ASAP7_75t_L g128 ( .A(n_96), .B(n_129), .Y(n_128) );
AND2x2_ASAP7_75t_L g127 ( .A(n_98), .B(n_128), .Y(n_127) );
AND2x4_ASAP7_75t_L g172 ( .A(n_98), .B(n_113), .Y(n_172) );
AND2x2_ASAP7_75t_L g98 ( .A(n_99), .B(n_103), .Y(n_98) );
AND2x2_ASAP7_75t_L g112 ( .A(n_99), .B(n_104), .Y(n_112) );
HB1xp67_ASAP7_75t_L g121 ( .A(n_99), .Y(n_121) );
INVx2_ASAP7_75t_L g139 ( .A(n_99), .Y(n_139) );
AND2x4_ASAP7_75t_L g152 ( .A(n_103), .B(n_139), .Y(n_152) );
INVx2_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
AND2x2_ASAP7_75t_L g138 ( .A(n_104), .B(n_139), .Y(n_138) );
BUFx2_ASAP7_75t_L g160 ( .A(n_104), .Y(n_160) );
INVx3_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
BUFx6f_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx3_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
INVx6_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
AND2x2_ASAP7_75t_L g111 ( .A(n_112), .B(n_113), .Y(n_111) );
AND2x4_ASAP7_75t_L g132 ( .A(n_112), .B(n_133), .Y(n_132) );
AND2x4_ASAP7_75t_L g142 ( .A(n_112), .B(n_143), .Y(n_142) );
AND2x2_ASAP7_75t_L g148 ( .A(n_113), .B(n_138), .Y(n_148) );
AND2x4_ASAP7_75t_L g165 ( .A(n_113), .B(n_152), .Y(n_165) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
BUFx3_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
BUFx12f_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
AND2x2_ASAP7_75t_L g119 ( .A(n_120), .B(n_121), .Y(n_119) );
AND2x4_ASAP7_75t_L g159 ( .A(n_120), .B(n_160), .Y(n_159) );
AND2x4_ASAP7_75t_L g173 ( .A(n_120), .B(n_152), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_124), .B(n_135), .Y(n_123) );
BUFx6f_ASAP7_75t_SL g125 ( .A(n_126), .Y(n_125) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
AND2x4_ASAP7_75t_L g151 ( .A(n_128), .B(n_152), .Y(n_151) );
AND2x2_ASAP7_75t_L g157 ( .A(n_128), .B(n_138), .Y(n_157) );
HB1xp67_ASAP7_75t_L g134 ( .A(n_129), .Y(n_134) );
INVx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx2_ASAP7_75t_SL g140 ( .A(n_141), .Y(n_140) );
INVx6_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
NOR2xp33_ASAP7_75t_L g144 ( .A(n_145), .B(n_161), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_146), .B(n_153), .Y(n_145) );
BUFx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx8_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
BUFx3_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_162), .B(n_169), .Y(n_161) );
INVx3_ASAP7_75t_SL g163 ( .A(n_164), .Y(n_163) );
INVx8_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
HB1xp67_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx3_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx6_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
OAI22xp5_ASAP7_75t_SL g175 ( .A1(n_176), .A2(n_183), .B1(n_189), .B2(n_190), .Y(n_175) );
CKINVDCx20_ASAP7_75t_R g189 ( .A(n_176), .Y(n_189) );
CKINVDCx16_ASAP7_75t_R g177 ( .A(n_178), .Y(n_177) );
INVx1_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
CKINVDCx20_ASAP7_75t_R g190 ( .A(n_183), .Y(n_190) );
CKINVDCx16_ASAP7_75t_R g187 ( .A(n_184), .Y(n_187) );
CKINVDCx20_ASAP7_75t_R g191 ( .A(n_192), .Y(n_191) );
CKINVDCx20_ASAP7_75t_R g192 ( .A(n_193), .Y(n_192) );
AND3x1_ASAP7_75t_SL g193 ( .A(n_194), .B(n_200), .C(n_203), .Y(n_193) );
INVxp67_ASAP7_75t_L g535 ( .A(n_194), .Y(n_535) );
CKINVDCx8_ASAP7_75t_R g195 ( .A(n_196), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_198), .B(n_199), .Y(n_197) );
CKINVDCx16_ASAP7_75t_R g533 ( .A(n_200), .Y(n_533) );
OAI21xp5_ASAP7_75t_L g542 ( .A1(n_200), .A2(n_543), .B(n_546), .Y(n_542) );
INVx1_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
OR2x2_ASAP7_75t_SL g540 ( .A(n_201), .B(n_203), .Y(n_540) );
AND2x2_ASAP7_75t_L g547 ( .A(n_201), .B(n_548), .Y(n_547) );
HB1xp67_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
AND2x2_ASAP7_75t_L g232 ( .A(n_202), .B(n_233), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_203), .B(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
HB1xp67_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
INVx3_ASAP7_75t_SL g206 ( .A(n_207), .Y(n_206) );
NOR2x2_ASAP7_75t_L g207 ( .A(n_208), .B(n_412), .Y(n_207) );
AO211x2_ASAP7_75t_L g208 ( .A1(n_209), .A2(n_254), .B(n_305), .C(n_380), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
INVxp67_ASAP7_75t_SL g210 ( .A(n_211), .Y(n_210) );
AND3x2_ASAP7_75t_L g461 ( .A(n_211), .B(n_342), .C(n_358), .Y(n_461) );
AND2x4_ASAP7_75t_L g464 ( .A(n_211), .B(n_465), .Y(n_464) );
AND2x2_ASAP7_75t_L g211 ( .A(n_212), .B(n_243), .Y(n_211) );
NAND2x1p5_ASAP7_75t_L g319 ( .A(n_212), .B(n_320), .Y(n_319) );
INVx4_ASAP7_75t_L g373 ( .A(n_212), .Y(n_373) );
AND2x2_ASAP7_75t_SL g458 ( .A(n_212), .B(n_367), .Y(n_458) );
AND2x2_ASAP7_75t_L g501 ( .A(n_212), .B(n_321), .Y(n_501) );
INVx5_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
BUFx2_ASAP7_75t_L g350 ( .A(n_213), .Y(n_350) );
AND2x2_ASAP7_75t_L g369 ( .A(n_213), .B(n_311), .Y(n_369) );
AND2x2_ASAP7_75t_L g387 ( .A(n_213), .B(n_321), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_213), .B(n_320), .Y(n_447) );
NOR2x1_ASAP7_75t_SL g474 ( .A(n_213), .B(n_243), .Y(n_474) );
OR2x6_ASAP7_75t_L g213 ( .A(n_214), .B(n_219), .Y(n_213) );
INVx3_ASAP7_75t_L g285 ( .A(n_215), .Y(n_285) );
INVx4_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
INVx3_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
BUFx4f_ASAP7_75t_L g312 ( .A(n_217), .Y(n_312) );
AND2x2_ASAP7_75t_SL g241 ( .A(n_218), .B(n_242), .Y(n_241) );
AND2x4_ASAP7_75t_L g245 ( .A(n_218), .B(n_242), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_228), .B(n_240), .Y(n_219) );
AND2x4_ASAP7_75t_L g221 ( .A(n_222), .B(n_227), .Y(n_221) );
AND2x4_ASAP7_75t_L g222 ( .A(n_223), .B(n_225), .Y(n_222) );
AND2x6_ASAP7_75t_L g238 ( .A(n_223), .B(n_231), .Y(n_238) );
INVx2_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
AND2x4_ASAP7_75t_L g236 ( .A(n_225), .B(n_233), .Y(n_236) );
INVx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
INVx5_ASAP7_75t_L g239 ( .A(n_227), .Y(n_239) );
HB1xp67_ASAP7_75t_L g526 ( .A(n_229), .Y(n_526) );
AND2x6_ASAP7_75t_L g229 ( .A(n_230), .B(n_232), .Y(n_229) );
BUFx3_ASAP7_75t_L g545 ( .A(n_230), .Y(n_545) );
INVx2_ASAP7_75t_L g548 ( .A(n_233), .Y(n_548) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_237), .B(n_239), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_239), .A2(n_249), .B(n_250), .Y(n_248) );
AOI21xp5_ASAP7_75t_L g261 ( .A1(n_239), .A2(n_262), .B(n_263), .Y(n_261) );
AOI21xp5_ASAP7_75t_L g273 ( .A1(n_239), .A2(n_274), .B(n_275), .Y(n_273) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_239), .A2(n_282), .B(n_283), .Y(n_281) );
AOI21xp5_ASAP7_75t_L g291 ( .A1(n_239), .A2(n_292), .B(n_293), .Y(n_291) );
AOI21xp5_ASAP7_75t_L g316 ( .A1(n_239), .A2(n_317), .B(n_318), .Y(n_316) );
AOI21xp5_ASAP7_75t_L g324 ( .A1(n_239), .A2(n_325), .B(n_326), .Y(n_324) );
OA21x2_ASAP7_75t_L g259 ( .A1(n_240), .A2(n_260), .B(n_264), .Y(n_259) );
CKINVDCx5p33_ASAP7_75t_R g328 ( .A(n_240), .Y(n_328) );
OA21x2_ASAP7_75t_L g333 ( .A1(n_240), .A2(n_260), .B(n_264), .Y(n_333) );
BUFx6f_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_243), .B(n_311), .Y(n_310) );
AO21x2_ASAP7_75t_L g243 ( .A1(n_244), .A2(n_246), .B(n_252), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g252 ( .A(n_244), .B(n_253), .Y(n_252) );
AO21x2_ASAP7_75t_L g346 ( .A1(n_244), .A2(n_246), .B(n_252), .Y(n_346) );
INVx1_ASAP7_75t_SL g244 ( .A(n_245), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_245), .B(n_277), .Y(n_276) );
AOI21xp5_ASAP7_75t_L g313 ( .A1(n_245), .A2(n_314), .B(n_315), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_247), .B(n_251), .Y(n_246) );
AO21x1_ASAP7_75t_L g254 ( .A1(n_255), .A2(n_287), .B(n_296), .Y(n_254) );
INVx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
OAI22xp33_ASAP7_75t_L g355 ( .A1(n_256), .A2(n_356), .B1(n_360), .B2(n_361), .Y(n_355) );
OR2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_265), .Y(n_256) );
AND2x2_ASAP7_75t_L g416 ( .A(n_257), .B(n_302), .Y(n_416) );
BUFx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
AND2x4_ASAP7_75t_L g349 ( .A(n_258), .B(n_332), .Y(n_349) );
AND2x2_ASAP7_75t_L g421 ( .A(n_258), .B(n_304), .Y(n_421) );
AND2x2_ASAP7_75t_L g440 ( .A(n_258), .B(n_406), .Y(n_440) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
INVx2_ASAP7_75t_L g297 ( .A(n_259), .Y(n_297) );
HB1xp67_ASAP7_75t_L g427 ( .A(n_259), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_265), .B(n_410), .Y(n_409) );
INVx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g400 ( .A(n_266), .B(n_299), .Y(n_400) );
AND2x4_ASAP7_75t_L g266 ( .A(n_267), .B(n_278), .Y(n_266) );
AND2x2_ASAP7_75t_L g302 ( .A(n_267), .B(n_303), .Y(n_302) );
OR2x2_ASAP7_75t_L g337 ( .A(n_267), .B(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_SL g397 ( .A(n_267), .B(n_333), .Y(n_397) );
INVx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
BUFx2_ASAP7_75t_L g490 ( .A(n_268), .Y(n_490) );
INVx2_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
INVx2_ASAP7_75t_L g332 ( .A(n_269), .Y(n_332) );
OAI21x1_ASAP7_75t_SL g269 ( .A1(n_270), .A2(n_272), .B(n_276), .Y(n_269) );
INVx1_ASAP7_75t_L g277 ( .A(n_271), .Y(n_277) );
INVx2_ASAP7_75t_L g338 ( .A(n_278), .Y(n_338) );
HB1xp67_ASAP7_75t_L g438 ( .A(n_278), .Y(n_438) );
AO21x2_ASAP7_75t_L g278 ( .A1(n_279), .A2(n_285), .B(n_286), .Y(n_278) );
AO21x2_ASAP7_75t_L g304 ( .A1(n_279), .A2(n_285), .B(n_286), .Y(n_304) );
NAND2xp5_ASAP7_75t_SL g279 ( .A(n_280), .B(n_284), .Y(n_279) );
AO21x2_ASAP7_75t_L g288 ( .A1(n_285), .A2(n_289), .B(n_295), .Y(n_288) );
AO21x2_ASAP7_75t_L g301 ( .A1(n_285), .A2(n_289), .B(n_295), .Y(n_301) );
INVx2_ASAP7_75t_L g334 ( .A(n_287), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_287), .B(n_466), .Y(n_492) );
AND2x2_ASAP7_75t_L g511 ( .A(n_287), .B(n_501), .Y(n_511) );
BUFx2_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x4_ASAP7_75t_SL g379 ( .A(n_288), .B(n_338), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_290), .B(n_294), .Y(n_289) );
AND2x2_ASAP7_75t_SL g296 ( .A(n_297), .B(n_298), .Y(n_296) );
AND2x2_ASAP7_75t_L g378 ( .A(n_297), .B(n_379), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_297), .B(n_348), .Y(n_383) );
INVx1_ASAP7_75t_SL g510 ( .A(n_297), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_298), .B(n_461), .Y(n_460) );
AND2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_302), .Y(n_298) );
INVx1_ASAP7_75t_L g336 ( .A(n_299), .Y(n_336) );
AND2x2_ASAP7_75t_L g522 ( .A(n_299), .B(n_523), .Y(n_522) );
BUFx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g398 ( .A(n_300), .B(n_303), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_300), .B(n_411), .Y(n_410) );
AND2x2_ASAP7_75t_L g452 ( .A(n_300), .B(n_304), .Y(n_452) );
AND2x2_ASAP7_75t_L g483 ( .A(n_300), .B(n_484), .Y(n_483) );
INVx2_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g348 ( .A(n_301), .B(n_304), .Y(n_348) );
INVxp67_ASAP7_75t_L g365 ( .A(n_301), .Y(n_365) );
BUFx3_ASAP7_75t_L g406 ( .A(n_301), .Y(n_406) );
AND2x2_ASAP7_75t_L g426 ( .A(n_302), .B(n_427), .Y(n_426) );
NAND2xp33_ASAP7_75t_L g439 ( .A(n_302), .B(n_440), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_303), .B(n_332), .Y(n_395) );
AND2x2_ASAP7_75t_L g484 ( .A(n_303), .B(n_333), .Y(n_484) );
INVx2_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g411 ( .A(n_304), .B(n_333), .Y(n_411) );
OR3x1_ASAP7_75t_L g305 ( .A(n_306), .B(n_355), .C(n_370), .Y(n_305) );
OAI321xp33_ASAP7_75t_L g306 ( .A1(n_307), .A2(n_319), .A3(n_330), .B1(n_335), .B2(n_339), .C(n_347), .Y(n_306) );
INVx1_ASAP7_75t_SL g307 ( .A(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVxp67_ASAP7_75t_SL g386 ( .A(n_310), .Y(n_386) );
INVxp67_ASAP7_75t_SL g404 ( .A(n_310), .Y(n_404) );
OR2x2_ASAP7_75t_L g408 ( .A(n_310), .B(n_319), .Y(n_408) );
BUFx3_ASAP7_75t_L g342 ( .A(n_311), .Y(n_342) );
AND2x2_ASAP7_75t_L g359 ( .A(n_311), .B(n_345), .Y(n_359) );
INVx1_ASAP7_75t_L g376 ( .A(n_311), .Y(n_376) );
INVx2_ASAP7_75t_L g392 ( .A(n_311), .Y(n_392) );
OR2x2_ASAP7_75t_L g431 ( .A(n_311), .B(n_320), .Y(n_431) );
INVx2_ASAP7_75t_L g419 ( .A(n_319), .Y(n_419) );
AND2x2_ASAP7_75t_L g343 ( .A(n_320), .B(n_344), .Y(n_343) );
INVx2_ASAP7_75t_L g358 ( .A(n_320), .Y(n_358) );
AND2x4_ASAP7_75t_L g367 ( .A(n_320), .B(n_368), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_320), .B(n_344), .Y(n_390) );
AND2x2_ASAP7_75t_L g497 ( .A(n_320), .B(n_392), .Y(n_497) );
INVx4_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
HB1xp67_ASAP7_75t_L g456 ( .A(n_321), .Y(n_456) );
AO21x2_ASAP7_75t_L g321 ( .A1(n_322), .A2(n_328), .B(n_329), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_323), .B(n_327), .Y(n_322) );
INVx1_ASAP7_75t_L g384 ( .A(n_330), .Y(n_384) );
NAND2xp5_ASAP7_75t_SL g330 ( .A(n_331), .B(n_334), .Y(n_330) );
AND2x2_ASAP7_75t_L g471 ( .A(n_331), .B(n_398), .Y(n_471) );
INVx1_ASAP7_75t_SL g488 ( .A(n_331), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_331), .B(n_464), .Y(n_517) );
AND2x4_ASAP7_75t_L g331 ( .A(n_332), .B(n_333), .Y(n_331) );
OR2x2_ASAP7_75t_L g360 ( .A(n_332), .B(n_333), .Y(n_360) );
AND2x2_ASAP7_75t_L g453 ( .A(n_334), .B(n_349), .Y(n_453) );
OR2x2_ASAP7_75t_L g335 ( .A(n_336), .B(n_337), .Y(n_335) );
NAND2xp5_ASAP7_75t_SL g476 ( .A(n_338), .B(n_349), .Y(n_476) );
INVx2_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_340), .A2(n_489), .B1(n_494), .B2(n_496), .Y(n_493) );
AND2x4_ASAP7_75t_L g340 ( .A(n_341), .B(n_343), .Y(n_340) );
AND2x2_ASAP7_75t_L g418 ( .A(n_341), .B(n_419), .Y(n_418) );
OR2x2_ASAP7_75t_L g513 ( .A(n_341), .B(n_514), .Y(n_513) );
INVx2_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g469 ( .A(n_342), .B(n_387), .Y(n_469) );
AND2x4_ASAP7_75t_L g423 ( .A(n_343), .B(n_369), .Y(n_423) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
HB1xp67_ASAP7_75t_L g521 ( .A(n_345), .Y(n_521) );
INVx2_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g354 ( .A(n_346), .Y(n_354) );
INVx1_ASAP7_75t_L g368 ( .A(n_346), .Y(n_368) );
NAND4xp25_ASAP7_75t_L g347 ( .A(n_348), .B(n_349), .C(n_350), .D(n_351), .Y(n_347) );
AND2x2_ASAP7_75t_L g505 ( .A(n_348), .B(n_490), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_348), .B(n_516), .Y(n_515) );
NOR2xp33_ASAP7_75t_L g424 ( .A(n_349), .B(n_425), .Y(n_424) );
OAI322xp33_ASAP7_75t_L g432 ( .A1(n_349), .A2(n_433), .A3(n_437), .B1(n_439), .B2(n_441), .C1(n_443), .C2(n_448), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_349), .B(n_398), .Y(n_448) );
INVx1_ASAP7_75t_L g516 ( .A(n_349), .Y(n_516) );
INVx2_ASAP7_75t_L g362 ( .A(n_350), .Y(n_362) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_353), .B(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_354), .B(n_373), .Y(n_430) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_357), .B(n_400), .Y(n_399) );
AND2x2_ASAP7_75t_L g357 ( .A(n_358), .B(n_359), .Y(n_357) );
INVx1_ASAP7_75t_L g403 ( .A(n_358), .Y(n_403) );
AND2x2_ASAP7_75t_L g475 ( .A(n_358), .B(n_386), .Y(n_475) );
AOI31xp33_ASAP7_75t_L g361 ( .A1(n_359), .A2(n_362), .A3(n_363), .B(n_366), .Y(n_361) );
AND2x2_ASAP7_75t_L g372 ( .A(n_359), .B(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g500 ( .A(n_359), .B(n_501), .Y(n_500) );
AND2x2_ASAP7_75t_SL g507 ( .A(n_359), .B(n_387), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_359), .Y(n_508) );
INVx1_ASAP7_75t_SL g466 ( .A(n_360), .Y(n_466) );
NAND3xp33_ASAP7_75t_SL g494 ( .A(n_360), .B(n_488), .C(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
OR2x2_ASAP7_75t_L g394 ( .A(n_365), .B(n_395), .Y(n_394) );
AND2x2_ASAP7_75t_L g366 ( .A(n_367), .B(n_369), .Y(n_366) );
AND2x2_ASAP7_75t_L g375 ( .A(n_367), .B(n_376), .Y(n_375) );
INVx2_ASAP7_75t_L g436 ( .A(n_367), .Y(n_436) );
AOI322xp5_ASAP7_75t_L g518 ( .A1(n_367), .A2(n_397), .A3(n_400), .B1(n_519), .B2(n_520), .C1(n_522), .C2(n_524), .Y(n_518) );
AND2x2_ASAP7_75t_L g524 ( .A(n_367), .B(n_373), .Y(n_524) );
AOI21xp5_ASAP7_75t_L g370 ( .A1(n_371), .A2(n_374), .B(n_377), .Y(n_370) );
INVx1_ASAP7_75t_SL g371 ( .A(n_372), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_373), .B(n_392), .Y(n_391) );
AND2x4_ASAP7_75t_L g519 ( .A(n_373), .B(n_406), .Y(n_519) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g445 ( .A(n_376), .Y(n_445) );
AND2x2_ASAP7_75t_L g473 ( .A(n_376), .B(n_474), .Y(n_473) );
AND2x2_ASAP7_75t_L g520 ( .A(n_376), .B(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g425 ( .A(n_379), .Y(n_425) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
O2A1O1Ixp5_ASAP7_75t_L g381 ( .A1(n_382), .A2(n_384), .B(n_385), .C(n_388), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
AND2x2_ASAP7_75t_L g385 ( .A(n_386), .B(n_387), .Y(n_385) );
AND2x2_ASAP7_75t_L g442 ( .A(n_387), .B(n_392), .Y(n_442) );
OAI211xp5_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_393), .B(n_399), .C(n_401), .Y(n_388) );
OAI221xp5_ASAP7_75t_L g414 ( .A1(n_389), .A2(n_415), .B1(n_417), .B2(n_420), .C(n_422), .Y(n_414) );
OR2x2_ASAP7_75t_L g389 ( .A(n_390), .B(n_391), .Y(n_389) );
INVx1_ASAP7_75t_L g434 ( .A(n_391), .Y(n_434) );
OR2x2_ASAP7_75t_L g454 ( .A(n_391), .B(n_455), .Y(n_454) );
AND2x2_ASAP7_75t_L g393 ( .A(n_394), .B(n_396), .Y(n_393) );
INVx1_ASAP7_75t_L g499 ( .A(n_394), .Y(n_499) );
INVx1_ASAP7_75t_L g523 ( .A(n_395), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g396 ( .A(n_397), .B(n_398), .Y(n_396) );
AND2x2_ASAP7_75t_L g405 ( .A(n_397), .B(n_406), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_397), .B(n_467), .Y(n_479) );
INVx1_ASAP7_75t_L g459 ( .A(n_398), .Y(n_459) );
AOI22xp5_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_405), .B1(n_407), .B2(n_409), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_403), .B(n_404), .Y(n_402) );
INVx1_ASAP7_75t_SL g467 ( .A(n_406), .Y(n_467) );
INVx2_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
NAND4xp75_ASAP7_75t_L g412 ( .A(n_413), .B(n_449), .C(n_477), .D(n_502), .Y(n_412) );
NOR2xp67_ASAP7_75t_L g413 ( .A(n_414), .B(n_432), .Y(n_413) );
INVx1_ASAP7_75t_SL g415 ( .A(n_416), .Y(n_415) );
INVx2_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
AND2x2_ASAP7_75t_SL g489 ( .A(n_421), .B(n_490), .Y(n_489) );
AOI22xp5_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_424), .B1(n_426), .B2(n_428), .Y(n_422) );
NOR2xp33_ASAP7_75t_L g487 ( .A(n_425), .B(n_488), .Y(n_487) );
INVx2_ASAP7_75t_SL g428 ( .A(n_429), .Y(n_428) );
OR2x2_ASAP7_75t_L g429 ( .A(n_430), .B(n_431), .Y(n_429) );
INVx2_ASAP7_75t_L g465 ( .A(n_431), .Y(n_465) );
OR2x2_ASAP7_75t_L g480 ( .A(n_431), .B(n_481), .Y(n_480) );
NAND2xp5_ASAP7_75t_SL g433 ( .A(n_434), .B(n_435), .Y(n_433) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g495 ( .A(n_440), .Y(n_495) );
INVx1_ASAP7_75t_SL g441 ( .A(n_442), .Y(n_441) );
OAI21xp5_ASAP7_75t_SL g486 ( .A1(n_442), .A2(n_487), .B(n_489), .Y(n_486) );
INVxp67_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_445), .B(n_446), .Y(n_444) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
NOR2x1_ASAP7_75t_L g449 ( .A(n_450), .B(n_462), .Y(n_449) );
OAI221xp5_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_454), .B1(n_457), .B2(n_459), .C(n_460), .Y(n_450) );
NOR2xp33_ASAP7_75t_L g451 ( .A(n_452), .B(n_453), .Y(n_451) );
OAI21xp33_ASAP7_75t_L g498 ( .A1(n_452), .A2(n_499), .B(n_500), .Y(n_498) );
INVx3_ASAP7_75t_SL g457 ( .A(n_458), .Y(n_457) );
OAI322xp33_ASAP7_75t_L g462 ( .A1(n_463), .A2(n_466), .A3(n_467), .B1(n_468), .B2(n_470), .C1(n_472), .C2(n_476), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_SL g470 ( .A(n_471), .Y(n_470) );
NOR2x1_ASAP7_75t_L g472 ( .A(n_473), .B(n_475), .Y(n_472) );
INVx1_ASAP7_75t_L g485 ( .A(n_473), .Y(n_485) );
INVx1_ASAP7_75t_L g481 ( .A(n_474), .Y(n_481) );
AND2x2_ASAP7_75t_L g496 ( .A(n_474), .B(n_497), .Y(n_496) );
NOR2x1_ASAP7_75t_L g477 ( .A(n_478), .B(n_491), .Y(n_477) );
OAI221xp5_ASAP7_75t_L g478 ( .A1(n_479), .A2(n_480), .B1(n_482), .B2(n_485), .C(n_486), .Y(n_478) );
INVx1_ASAP7_75t_SL g482 ( .A(n_483), .Y(n_482) );
OAI211xp5_ASAP7_75t_SL g491 ( .A1(n_485), .A2(n_492), .B(n_493), .C(n_498), .Y(n_491) );
INVx2_ASAP7_75t_SL g514 ( .A(n_501), .Y(n_514) );
NOR2x1_ASAP7_75t_L g502 ( .A(n_503), .B(n_512), .Y(n_502) );
OAI22xp33_ASAP7_75t_L g503 ( .A1(n_504), .A2(n_506), .B1(n_508), .B2(n_509), .Y(n_503) );
INVx1_ASAP7_75t_SL g504 ( .A(n_505), .Y(n_504) );
INVx2_ASAP7_75t_SL g506 ( .A(n_507), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_510), .B(n_511), .Y(n_509) );
OAI211xp5_ASAP7_75t_SL g512 ( .A1(n_513), .A2(n_515), .B(n_517), .C(n_518), .Y(n_512) );
HB1xp67_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
OAI222xp33_ASAP7_75t_L g527 ( .A1(n_528), .A2(n_530), .B1(n_536), .B2(n_538), .C1(n_541), .C2(n_549), .Y(n_527) );
CKINVDCx20_ASAP7_75t_R g530 ( .A(n_531), .Y(n_530) );
CKINVDCx20_ASAP7_75t_R g531 ( .A(n_532), .Y(n_531) );
OR2x2_ASAP7_75t_L g532 ( .A(n_533), .B(n_534), .Y(n_532) );
CKINVDCx20_ASAP7_75t_R g538 ( .A(n_539), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
CKINVDCx16_ASAP7_75t_R g541 ( .A(n_542), .Y(n_541) );
INVxp67_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
endmodule