module real_jpeg_8767_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_247;
wire n_146;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_131;
wire n_47;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_255;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_195;
wire n_61;
wire n_110;
wire n_258;
wire n_205;
wire n_117;
wire n_193;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_150;
wire n_32;
wire n_20;
wire n_74;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_52;
wire n_58;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_128;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_0),
.A2(n_38),
.B1(n_39),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_0),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_0),
.A2(n_27),
.B1(n_30),
.B2(n_49),
.Y(n_95)
);

BUFx24_ASAP7_75t_L g61 ( 
.A(n_1),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_2),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_2),
.A2(n_29),
.B1(n_59),
.B2(n_60),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_2),
.A2(n_29),
.B1(n_38),
.B2(n_39),
.Y(n_90)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_4),
.A2(n_54),
.B1(n_63),
.B2(n_64),
.Y(n_62)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_4),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_4),
.A2(n_59),
.B1(n_60),
.B2(n_64),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_4),
.A2(n_27),
.B1(n_30),
.B2(n_64),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_4),
.A2(n_38),
.B1(n_39),
.B2(n_64),
.Y(n_224)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

BUFx6f_ASAP7_75t_SL g72 ( 
.A(n_8),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_10),
.A2(n_54),
.B1(n_63),
.B2(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_10),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_10),
.A2(n_59),
.B1(n_60),
.B2(n_104),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_10),
.A2(n_27),
.B1(n_30),
.B2(n_104),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_10),
.A2(n_38),
.B1(n_39),
.B2(n_104),
.Y(n_216)
);

OAI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_11),
.A2(n_27),
.B1(n_30),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_11),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_11),
.A2(n_35),
.B1(n_54),
.B2(n_63),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_11),
.A2(n_35),
.B1(n_59),
.B2(n_60),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_11),
.A2(n_35),
.B1(n_38),
.B2(n_39),
.Y(n_153)
);

BUFx10_ASAP7_75t_L g54 ( 
.A(n_12),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_13),
.A2(n_54),
.B1(n_63),
.B2(n_123),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_13),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_13),
.A2(n_59),
.B1(n_60),
.B2(n_123),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_13),
.A2(n_38),
.B1(n_39),
.B2(n_123),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_13),
.A2(n_27),
.B1(n_30),
.B2(n_123),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_14),
.A2(n_38),
.B1(n_39),
.B2(n_42),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_14),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_14),
.A2(n_42),
.B1(n_59),
.B2(n_60),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_14),
.A2(n_27),
.B1(n_30),
.B2(n_42),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_15),
.Y(n_127)
);

AOI21xp33_ASAP7_75t_L g128 ( 
.A1(n_15),
.A2(n_56),
.B(n_60),
.Y(n_128)
);

OAI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_15),
.A2(n_54),
.B1(n_63),
.B2(n_127),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_15),
.B(n_67),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_15),
.A2(n_38),
.B(n_192),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_15),
.B(n_38),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_15),
.A2(n_84),
.B1(n_85),
.B2(n_203),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_133),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_131),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_108),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_19),
.B(n_108),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_92),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_80),
.B2(n_81),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_50),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_36),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_24),
.B(n_36),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_33),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_25),
.A2(n_85),
.B(n_130),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_31),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_26),
.B(n_32),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_27),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_27),
.A2(n_30),
.B1(n_44),
.B2(n_47),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_27),
.A2(n_195),
.B1(n_196),
.B2(n_197),
.Y(n_194)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_30),
.B(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_30),
.B(n_47),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_30),
.B(n_207),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_31),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_31),
.A2(n_32),
.B1(n_184),
.B2(n_186),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_32),
.B(n_34),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_32),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_33),
.A2(n_84),
.B(n_187),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_34),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_43),
.B1(n_46),
.B2(n_48),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_37),
.A2(n_46),
.B(n_98),
.Y(n_97)
);

A2O1A1Ixp33_ASAP7_75t_SL g43 ( 
.A1(n_38),
.A2(n_44),
.B(n_45),
.C(n_46),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_44),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_38),
.A2(n_39),
.B1(n_71),
.B2(n_72),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_38),
.B(n_71),
.Y(n_231)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_39),
.A2(n_76),
.B1(n_226),
.B2(n_231),
.Y(n_230)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_43),
.A2(n_48),
.B(n_88),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_43),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_43),
.A2(n_46),
.B1(n_191),
.B2(n_193),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_43),
.A2(n_46),
.B1(n_193),
.B2(n_216),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_43),
.A2(n_46),
.B1(n_216),
.B2(n_224),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_43),
.A2(n_224),
.B(n_247),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_44),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_45),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_46),
.B(n_90),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_46),
.B(n_127),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_46),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_52),
.B1(n_68),
.B2(n_79),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_53),
.A2(n_62),
.B(n_65),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_53),
.A2(n_58),
.B1(n_62),
.B2(n_103),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_53),
.A2(n_58),
.B1(n_103),
.B2(n_122),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_53),
.Y(n_149)
);

A2O1A1Ixp33_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_55),
.B(n_57),
.C(n_58),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_54),
.B(n_55),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_54),
.Y(n_63)
);

A2O1A1Ixp33_ASAP7_75t_L g126 ( 
.A1(n_54),
.A2(n_55),
.B(n_127),
.C(n_128),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_55),
.A2(n_56),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

O2A1O1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_60),
.A2(n_70),
.B(n_71),
.C(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_60),
.B(n_71),
.Y(n_76)
);

HAxp5_ASAP7_75t_SL g226 ( 
.A(n_60),
.B(n_127),
.CON(n_226),
.SN(n_226)
);

BUFx10_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_66),
.B(n_67),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_67),
.A2(n_149),
.B1(n_150),
.B2(n_151),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_68),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_73),
.B(n_74),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_69),
.B(n_78),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_69),
.A2(n_117),
.B1(n_118),
.B2(n_147),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_69),
.A2(n_117),
.B1(n_147),
.B2(n_170),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_69),
.B(n_127),
.Y(n_214)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_70),
.B(n_106),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_70),
.A2(n_75),
.B1(n_171),
.B2(n_226),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_77),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_75),
.A2(n_106),
.B(n_107),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_75),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_83),
.B1(n_87),
.B2(n_91),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_85),
.B(n_86),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_84),
.A2(n_95),
.B(n_96),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_84),
.A2(n_85),
.B1(n_95),
.B2(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_84),
.A2(n_85),
.B1(n_185),
.B2(n_203),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_84),
.A2(n_86),
.B(n_96),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_85),
.B(n_127),
.Y(n_207)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_87),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_89),
.A2(n_100),
.B(n_153),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_90),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_101),
.C(n_105),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_97),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_94),
.B(n_97),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_100),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_101),
.A2(n_102),
.B1(n_105),
.B2(n_111),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_105),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_112),
.C(n_113),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_109),
.B(n_112),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_113),
.A2(n_114),
.B1(n_155),
.B2(n_156),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_120),
.C(n_124),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_115),
.A2(n_116),
.B1(n_120),
.B2(n_121),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_117),
.A2(n_118),
.B(n_119),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_122),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_124),
.B(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_129),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_125),
.A2(n_126),
.B1(n_129),
.B2(n_165),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_129),
.Y(n_165)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_176),
.Y(n_133)
);

INVxp33_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_157),
.B(n_175),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

NOR3xp33_ASAP7_75t_L g176 ( 
.A(n_137),
.B(n_177),
.C(n_258),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_154),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_138),
.B(n_154),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_141),
.C(n_143),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_139),
.B(n_159),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_141),
.A2(n_142),
.B1(n_143),
.B2(n_144),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_148),
.C(n_152),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_145),
.A2(n_146),
.B1(n_152),
.B2(n_163),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_148),
.B(n_162),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_152),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_153),
.B(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_155),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_160),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_158),
.B(n_160),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_164),
.C(n_166),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_161),
.B(n_255),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_164),
.A2(n_166),
.B1(n_167),
.B2(n_256),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_164),
.Y(n_256)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_172),
.C(n_173),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_168),
.A2(n_169),
.B1(n_240),
.B2(n_241),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_172),
.A2(n_173),
.B1(n_174),
.B2(n_242),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_172),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_252),
.B(n_257),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_179),
.A2(n_235),
.B(n_251),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_219),
.B(n_234),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_181),
.A2(n_210),
.B(n_218),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_199),
.B(n_209),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_188),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_183),
.B(n_188),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_189),
.A2(n_190),
.B1(n_194),
.B2(n_198),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_189),
.B(n_198),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_192),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_194),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_204),
.B(n_208),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_201),
.B(n_202),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_211),
.B(n_212),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_213),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_213),
.B(n_220),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_213),
.B(n_220),
.Y(n_234)
);

FAx1_ASAP7_75t_SL g213 ( 
.A(n_214),
.B(n_215),
.CI(n_217),
.CON(n_213),
.SN(n_213)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_222),
.B1(n_229),
.B2(n_233),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_225),
.B1(n_227),
.B2(n_228),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_223),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_225),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_225),
.B(n_228),
.C(n_233),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_229),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_232),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_230),
.B(n_232),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_236),
.B(n_237),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_238),
.A2(n_239),
.B1(n_243),
.B2(n_244),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_238),
.B(n_246),
.C(n_249),
.Y(n_253)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_245),
.A2(n_246),
.B1(n_249),
.B2(n_250),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_245),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_246),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_253),
.B(n_254),
.Y(n_257)
);


endmodule