module real_jpeg_4540_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_202;
wire n_128;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx8_ASAP7_75t_L g74 ( 
.A(n_0),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_1),
.A2(n_81),
.B1(n_83),
.B2(n_84),
.Y(n_80)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_1),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_1),
.A2(n_83),
.B1(n_156),
.B2(n_158),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_1),
.A2(n_83),
.B1(n_184),
.B2(n_186),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_1),
.A2(n_23),
.B1(n_83),
.B2(n_194),
.Y(n_193)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_2),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_2),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_2),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_3),
.A2(n_139),
.B1(n_140),
.B2(n_143),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_3),
.Y(n_139)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_4),
.Y(n_59)
);

INVx8_ASAP7_75t_L g148 ( 
.A(n_5),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_5),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_5),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_5),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_5),
.Y(n_280)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_7),
.A2(n_22),
.B1(n_117),
.B2(n_120),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_7),
.B(n_39),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_7),
.A2(n_22),
.B1(n_169),
.B2(n_170),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_7),
.A2(n_22),
.B1(n_45),
.B2(n_202),
.Y(n_201)
);

O2A1O1Ixp33_ASAP7_75t_L g215 ( 
.A1(n_7),
.A2(n_216),
.B(n_219),
.C(n_223),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_7),
.B(n_102),
.C(n_144),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_7),
.B(n_91),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_7),
.B(n_280),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_7),
.B(n_107),
.Y(n_284)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_9),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g195 ( 
.A(n_9),
.Y(n_195)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_10),
.Y(n_101)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_10),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_10),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_11),
.A2(n_49),
.B1(n_50),
.B2(n_51),
.Y(n_48)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_11),
.A2(n_50),
.B1(n_87),
.B2(n_90),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_11),
.A2(n_50),
.B1(n_233),
.B2(n_236),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_L g254 ( 
.A1(n_11),
.A2(n_50),
.B1(n_111),
.B2(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);

OAI22xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_205),
.B1(n_308),
.B2(n_309),
.Y(n_13)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_14),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_204),
.Y(n_14)
);

INVxp67_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_174),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_17),
.B(n_174),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_123),
.C(n_159),
.Y(n_17)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_18),
.B(n_208),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_52),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_19),
.B(n_53),
.C(n_93),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_47),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_30),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B(n_26),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_22),
.B(n_27),
.Y(n_26)
);

OAI21xp33_ASAP7_75t_L g219 ( 
.A1(n_22),
.A2(n_220),
.B(n_221),
.Y(n_219)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVxp33_ASAP7_75t_L g132 ( 
.A(n_26),
.Y(n_132)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_30),
.B(n_48),
.Y(n_196)
);

NOR2x1_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_39),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_34),
.B1(n_35),
.B2(n_38),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp33_ASAP7_75t_SL g133 ( 
.A(n_35),
.B(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

AO22x2_ASAP7_75t_L g39 ( 
.A1(n_36),
.A2(n_40),
.B1(n_41),
.B2(n_45),
.Y(n_39)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_39),
.B(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_40),
.Y(n_129)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_43),
.Y(n_203)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_44),
.Y(n_128)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_45),
.Y(n_223)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_46),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_92),
.B1(n_93),
.B2(n_122),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_53),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_54),
.B(n_85),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_56),
.B(n_79),
.Y(n_55)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_56),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_69),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_60),
.B1(n_62),
.B2(n_66),
.Y(n_57)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_59),
.Y(n_218)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_69),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_69),
.B(n_200),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_71),
.B1(n_75),
.B2(n_78),
.Y(n_69)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_74),
.Y(n_77)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_74),
.Y(n_99)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_74),
.Y(n_121)
);

BUFx5_ASAP7_75t_L g236 ( 
.A(n_74),
.Y(n_236)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_76),
.Y(n_106)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_77),
.Y(n_119)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_77),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_77),
.Y(n_235)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_80),
.B(n_91),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_81),
.Y(n_90)
);

INVx6_ASAP7_75t_SL g81 ( 
.A(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_85),
.B(n_296),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_91),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_86),
.B(n_163),
.Y(n_162)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_114),
.B(n_115),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_95),
.B(n_116),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_95),
.B(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_95),
.B(n_183),
.Y(n_294)
);

NOR2x1_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_107),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_100),
.B1(n_102),
.B2(n_105),
.Y(n_96)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_98),
.Y(n_222)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_99),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_107),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_107),
.B(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_107),
.B(n_232),
.Y(n_247)
);

AO22x1_ASAP7_75t_SL g107 ( 
.A1(n_108),
.A2(n_109),
.B1(n_111),
.B2(n_113),
.Y(n_107)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_108),
.Y(n_113)
);

INVx8_ASAP7_75t_L g142 ( 
.A(n_109),
.Y(n_142)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_109),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx3_ASAP7_75t_SL g169 ( 
.A(n_111),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx5_ASAP7_75t_L g144 ( 
.A(n_112),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_114),
.B(n_115),
.Y(n_230)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_123),
.A2(n_124),
.B1(n_159),
.B2(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_137),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_125),
.B(n_137),
.Y(n_189)
);

AOI32xp33_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_129),
.A3(n_130),
.B1(n_132),
.B2(n_133),
.Y(n_125)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_145),
.B(n_149),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_138),
.A2(n_171),
.B(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_145),
.B(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_148),
.Y(n_173)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_149),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_155),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_150),
.B(n_168),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_150),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_150),
.A2(n_168),
.B(n_225),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_150),
.B(n_254),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_153),
.Y(n_150)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_151),
.Y(n_278)
);

BUFx5_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_152),
.Y(n_157)
);

BUFx8_ASAP7_75t_L g170 ( 
.A(n_152),
.Y(n_170)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_152),
.Y(n_258)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_155),
.B(n_172),
.Y(n_171)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_159),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_164),
.C(n_166),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_160),
.B(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_162),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_162),
.B(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_163),
.B(n_201),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_164),
.A2(n_165),
.B1(n_166),
.B2(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_166),
.Y(n_213)
);

OR2x2_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_171),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_167),
.B(n_270),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_168),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_171),
.B(n_253),
.Y(n_283)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_188),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_180),
.Y(n_177)
);

AND2x2_ASAP7_75t_SL g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_181),
.B(n_247),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_182),
.B(n_231),
.Y(n_260)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx5_ASAP7_75t_L g244 ( 
.A(n_185),
.Y(n_244)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g188 ( 
.A(n_189),
.B(n_190),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_197),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_196),
.Y(n_191)
);

INVx8_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVxp67_ASAP7_75t_SL g200 ( 
.A(n_201),
.Y(n_200)
);

INVx6_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_205),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_237),
.B(n_307),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_210),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_207),
.B(n_210),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_214),
.C(n_227),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_211),
.B(n_303),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_214),
.A2(n_227),
.B1(n_228),
.B2(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_214),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_224),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_215),
.A2(n_224),
.B1(n_298),
.B2(n_299),
.Y(n_297)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_215),
.Y(n_299)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_216),
.Y(n_220)
);

INVx8_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_224),
.Y(n_298)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_231),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx11_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_301),
.B(n_306),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_239),
.A2(n_288),
.B(n_300),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_264),
.B(n_287),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_248),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_241),
.B(n_248),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_246),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_242),
.A2(n_243),
.B1(n_246),
.B2(n_267),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_243),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_246),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_247),
.B(n_294),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_259),
.Y(n_248)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_249),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_252),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_254),
.B(n_271),
.Y(n_270)
);

BUFx2_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_260),
.A2(n_261),
.B1(n_262),
.B2(n_263),
.Y(n_259)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_260),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_261),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_261),
.B(n_262),
.C(n_290),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_265),
.A2(n_274),
.B(n_286),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_266),
.B(n_268),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_266),
.B(n_268),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_273),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_282),
.B(n_285),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_281),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_279),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_278),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_283),
.B(n_284),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_291),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_289),
.B(n_291),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_297),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_295),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_293),
.B(n_295),
.C(n_297),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_302),
.B(n_305),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_302),
.B(n_305),
.Y(n_306)
);


endmodule