module fake_jpeg_4325_n_216 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_216);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_216;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx3_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_13),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_7),
.B(n_1),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_31),
.B(n_44),
.Y(n_59)
);

INVx6_ASAP7_75t_SL g32 ( 
.A(n_29),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_33),
.A2(n_28),
.B1(n_30),
.B2(n_26),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_24),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_34),
.B(n_12),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_18),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_35),
.A2(n_39),
.B(n_42),
.Y(n_52)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_20),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_37),
.A2(n_17),
.B1(n_22),
.B2(n_27),
.Y(n_57)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_24),
.B(n_2),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_16),
.B(n_3),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_16),
.B(n_3),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_45),
.A2(n_8),
.B(n_9),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

CKINVDCx12_ASAP7_75t_R g47 ( 
.A(n_28),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_14),
.Y(n_69)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_48),
.B(n_49),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_17),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_50),
.B(n_54),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_35),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_51),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g53 ( 
.A1(n_39),
.A2(n_15),
.B(n_18),
.Y(n_53)
);

AO21x1_ASAP7_75t_L g95 ( 
.A1(n_53),
.A2(n_69),
.B(n_85),
.Y(n_95)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_55),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_57),
.A2(n_66),
.B1(n_79),
.B2(n_80),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_31),
.A2(n_15),
.B1(n_27),
.B2(n_19),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_60),
.A2(n_11),
.B1(n_76),
.B2(n_64),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_34),
.B(n_45),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_61),
.B(n_63),
.Y(n_109)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_22),
.Y(n_63)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_65),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_19),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_82),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_32),
.Y(n_70)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_33),
.B(n_28),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_71),
.Y(n_97)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_73),
.Y(n_102)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_74),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_46),
.B(n_6),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_75),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_77),
.Y(n_108)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_33),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_42),
.B(n_6),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_36),
.A2(n_25),
.B1(n_26),
.B2(n_30),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_83),
.A2(n_10),
.B1(n_11),
.B2(n_66),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_34),
.B(n_28),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_8),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_64),
.A2(n_30),
.B1(n_25),
.B2(n_14),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_88),
.A2(n_110),
.B1(n_104),
.B2(n_90),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_52),
.B(n_59),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_94),
.B(n_96),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_72),
.B(n_25),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_55),
.A2(n_25),
.B1(n_9),
.B2(n_10),
.Y(n_98)
);

OAI22x1_ASAP7_75t_L g124 ( 
.A1(n_98),
.A2(n_105),
.B1(n_49),
.B2(n_77),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_100),
.B(n_58),
.Y(n_114)
);

OAI32xp33_ASAP7_75t_L g104 ( 
.A1(n_78),
.A2(n_8),
.A3(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_111),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_72),
.B(n_78),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_106),
.B(n_65),
.Y(n_113)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_113),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_114),
.B(n_115),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_91),
.B(n_83),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_101),
.B(n_80),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_116),
.B(n_117),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_101),
.B(n_109),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_91),
.B(n_67),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_119),
.B(n_121),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_95),
.A2(n_67),
.B1(n_81),
.B2(n_70),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_120),
.Y(n_150)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_86),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_94),
.B(n_70),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_122),
.B(n_126),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_89),
.A2(n_56),
.B(n_81),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_123),
.A2(n_124),
.B(n_115),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_87),
.B(n_58),
.Y(n_125)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_125),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_111),
.B(n_77),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_96),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_127),
.B(n_128),
.Y(n_147)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_110),
.Y(n_128)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_129),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_87),
.B(n_107),
.Y(n_130)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_130),
.Y(n_155)
);

BUFx8_ASAP7_75t_L g131 ( 
.A(n_108),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_99),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_132),
.B(n_134),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_97),
.B(n_95),
.Y(n_133)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_133),
.Y(n_156)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_99),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_100),
.B(n_93),
.Y(n_135)
);

NAND2xp33_ASAP7_75t_SL g154 ( 
.A(n_135),
.B(n_124),
.Y(n_154)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_102),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_136),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_112),
.A2(n_90),
.B1(n_92),
.B2(n_103),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_137),
.A2(n_140),
.B1(n_129),
.B2(n_135),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_112),
.A2(n_92),
.B1(n_103),
.B2(n_108),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_118),
.B(n_122),
.C(n_126),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_146),
.B(n_148),
.C(n_151),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_118),
.B(n_102),
.C(n_127),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_149),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_119),
.B(n_120),
.C(n_133),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_154),
.B(n_136),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_123),
.B(n_117),
.C(n_128),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_157),
.B(n_132),
.C(n_134),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_138),
.A2(n_116),
.B(n_114),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_158),
.A2(n_167),
.B(n_169),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_147),
.B(n_135),
.Y(n_159)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_159),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_149),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_162),
.B(n_165),
.Y(n_178)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_163),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_147),
.B(n_121),
.Y(n_164)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_164),
.Y(n_181)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_153),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_166),
.B(n_168),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_146),
.B(n_131),
.C(n_148),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_156),
.A2(n_131),
.B(n_157),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_153),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_170),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_152),
.A2(n_131),
.B1(n_137),
.B2(n_140),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_171),
.A2(n_156),
.B1(n_152),
.B2(n_142),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_142),
.Y(n_172)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_172),
.Y(n_182)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_175),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_172),
.B(n_151),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_176),
.B(n_184),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_164),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_180),
.B(n_185),
.Y(n_186)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_171),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_159),
.B(n_139),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_183),
.A2(n_167),
.B(n_161),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_188),
.A2(n_189),
.B(n_176),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_183),
.A2(n_169),
.B(n_166),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_181),
.B(n_155),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_190),
.B(n_181),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_174),
.B(n_168),
.C(n_160),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_191),
.B(n_192),
.C(n_193),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_174),
.B(n_160),
.C(n_145),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_173),
.B(n_145),
.C(n_163),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_186),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_195),
.B(n_199),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_193),
.B(n_194),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_197),
.B(n_175),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_198),
.B(n_179),
.Y(n_205)
);

NOR3xp33_ASAP7_75t_SL g199 ( 
.A(n_187),
.B(n_154),
.C(n_158),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_200),
.B(n_201),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_186),
.B(n_143),
.Y(n_201)
);

AOI322xp5_ASAP7_75t_L g208 ( 
.A1(n_202),
.A2(n_205),
.A3(n_177),
.B1(n_197),
.B2(n_173),
.C1(n_170),
.C2(n_182),
.Y(n_208)
);

AO22x1_ASAP7_75t_L g206 ( 
.A1(n_199),
.A2(n_178),
.B1(n_184),
.B2(n_179),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_206),
.A2(n_143),
.B1(n_155),
.B2(n_144),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_204),
.B(n_165),
.Y(n_207)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_207),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_208),
.B(n_209),
.Y(n_213)
);

AOI322xp5_ASAP7_75t_L g209 ( 
.A1(n_203),
.A2(n_177),
.A3(n_196),
.B1(n_141),
.B2(n_182),
.C1(n_150),
.C2(n_139),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_210),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_211),
.B(n_196),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_214),
.A2(n_215),
.B(n_213),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_212),
.A2(n_207),
.B1(n_204),
.B2(n_144),
.Y(n_215)
);


endmodule