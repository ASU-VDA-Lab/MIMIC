module real_aes_2884_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_769;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_617;
wire n_552;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_728;
wire n_598;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_753;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g229 ( .A(n_0), .B(n_144), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_1), .B(n_740), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_2), .B(n_128), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_3), .B(n_146), .Y(n_451) );
INVx1_ASAP7_75t_L g135 ( .A(n_4), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_5), .B(n_128), .Y(n_127) );
NAND2xp33_ASAP7_75t_SL g214 ( .A(n_6), .B(n_134), .Y(n_214) );
INVx1_ASAP7_75t_L g205 ( .A(n_7), .Y(n_205) );
CKINVDCx16_ASAP7_75t_R g740 ( .A(n_8), .Y(n_740) );
AND2x2_ASAP7_75t_L g122 ( .A(n_9), .B(n_123), .Y(n_122) );
AOI221xp5_ASAP7_75t_L g103 ( .A1(n_10), .A2(n_104), .B1(n_733), .B2(n_744), .C(n_753), .Y(n_103) );
AND2x2_ASAP7_75t_L g453 ( .A(n_10), .B(n_175), .Y(n_453) );
OAI22xp5_ASAP7_75t_SL g759 ( .A1(n_10), .A2(n_69), .B1(n_760), .B2(n_761), .Y(n_759) );
CKINVDCx20_ASAP7_75t_R g760 ( .A(n_10), .Y(n_760) );
AND2x2_ASAP7_75t_L g461 ( .A(n_11), .B(n_211), .Y(n_461) );
INVx2_ASAP7_75t_L g124 ( .A(n_12), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_13), .B(n_146), .Y(n_469) );
CKINVDCx16_ASAP7_75t_R g108 ( .A(n_14), .Y(n_108) );
AOI221x1_ASAP7_75t_L g208 ( .A1(n_15), .A2(n_137), .B1(n_209), .B2(n_211), .C(n_213), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_16), .B(n_128), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g493 ( .A(n_17), .B(n_128), .Y(n_493) );
INVx1_ASAP7_75t_L g111 ( .A(n_18), .Y(n_111) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_19), .A2(n_92), .B1(n_128), .B2(n_179), .Y(n_522) );
AOI22xp5_ASAP7_75t_L g756 ( .A1(n_20), .A2(n_73), .B1(n_757), .B2(n_758), .Y(n_756) );
CKINVDCx20_ASAP7_75t_R g758 ( .A(n_20), .Y(n_758) );
AOI21xp5_ASAP7_75t_L g136 ( .A1(n_21), .A2(n_137), .B(n_142), .Y(n_136) );
AOI221xp5_ASAP7_75t_SL g219 ( .A1(n_22), .A2(n_36), .B1(n_128), .B2(n_137), .C(n_220), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_23), .B(n_144), .Y(n_143) );
OR2x2_ASAP7_75t_L g125 ( .A(n_24), .B(n_91), .Y(n_125) );
OA21x2_ASAP7_75t_L g176 ( .A1(n_24), .A2(n_91), .B(n_124), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_25), .B(n_146), .Y(n_199) );
INVxp67_ASAP7_75t_L g207 ( .A(n_26), .Y(n_207) );
AND2x2_ASAP7_75t_L g168 ( .A(n_27), .B(n_158), .Y(n_168) );
AOI22xp5_ASAP7_75t_SL g721 ( .A1(n_28), .A2(n_722), .B1(n_723), .B2(n_724), .Y(n_721) );
CKINVDCx20_ASAP7_75t_R g722 ( .A(n_28), .Y(n_722) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_29), .A2(n_137), .B(n_228), .Y(n_227) );
AO21x2_ASAP7_75t_L g464 ( .A1(n_30), .A2(n_211), .B(n_465), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_31), .B(n_146), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g448 ( .A1(n_32), .A2(n_137), .B(n_449), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_33), .B(n_146), .Y(n_477) );
AND2x2_ASAP7_75t_L g134 ( .A(n_34), .B(n_135), .Y(n_134) );
AND2x2_ASAP7_75t_L g138 ( .A(n_34), .B(n_139), .Y(n_138) );
INVx1_ASAP7_75t_L g187 ( .A(n_34), .Y(n_187) );
OR2x6_ASAP7_75t_L g109 ( .A(n_35), .B(n_110), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_37), .B(n_128), .Y(n_452) );
AOI22xp5_ASAP7_75t_L g184 ( .A1(n_38), .A2(n_84), .B1(n_137), .B2(n_185), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_39), .B(n_146), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_40), .B(n_128), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_41), .B(n_144), .Y(n_166) );
AOI21xp5_ASAP7_75t_L g456 ( .A1(n_42), .A2(n_137), .B(n_457), .Y(n_456) );
AND2x2_ASAP7_75t_L g232 ( .A(n_43), .B(n_158), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_44), .B(n_144), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_45), .B(n_158), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g466 ( .A(n_46), .B(n_128), .Y(n_466) );
AOI22xp33_ASAP7_75t_L g727 ( .A1(n_47), .A2(n_720), .B1(n_728), .B2(n_731), .Y(n_727) );
INVx1_ASAP7_75t_L g131 ( .A(n_48), .Y(n_131) );
INVx1_ASAP7_75t_L g141 ( .A(n_48), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_49), .B(n_146), .Y(n_459) );
AND2x2_ASAP7_75t_L g484 ( .A(n_50), .B(n_158), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_51), .B(n_769), .Y(n_768) );
NAND2xp5_ASAP7_75t_SL g167 ( .A(n_52), .B(n_128), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_53), .B(n_144), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_54), .B(n_144), .Y(n_476) );
AND2x2_ASAP7_75t_L g159 ( .A(n_55), .B(n_158), .Y(n_159) );
NAND2xp5_ASAP7_75t_SL g460 ( .A(n_56), .B(n_128), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_57), .B(n_146), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g486 ( .A(n_58), .B(n_128), .Y(n_486) );
AOI21xp5_ASAP7_75t_L g474 ( .A1(n_59), .A2(n_137), .B(n_475), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_60), .B(n_144), .Y(n_155) );
AND2x2_ASAP7_75t_SL g200 ( .A(n_61), .B(n_123), .Y(n_200) );
AND2x2_ASAP7_75t_L g499 ( .A(n_62), .B(n_123), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g163 ( .A1(n_63), .A2(n_137), .B(n_164), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_64), .B(n_146), .Y(n_145) );
AND2x2_ASAP7_75t_SL g190 ( .A(n_65), .B(n_175), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_66), .B(n_144), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_67), .B(n_144), .Y(n_470) );
AOI22xp5_ASAP7_75t_L g523 ( .A1(n_68), .A2(n_95), .B1(n_137), .B2(n_185), .Y(n_523) );
INVx1_ASAP7_75t_L g761 ( .A(n_69), .Y(n_761) );
OAI22xp5_ASAP7_75t_SL g724 ( .A1(n_70), .A2(n_80), .B1(n_725), .B2(n_726), .Y(n_724) );
CKINVDCx14_ASAP7_75t_R g726 ( .A(n_70), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_71), .B(n_146), .Y(n_496) );
INVx1_ASAP7_75t_L g133 ( .A(n_72), .Y(n_133) );
INVx1_ASAP7_75t_L g139 ( .A(n_72), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g757 ( .A(n_73), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_74), .B(n_144), .Y(n_450) );
XNOR2xp5_ASAP7_75t_L g720 ( .A(n_75), .B(n_721), .Y(n_720) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_76), .A2(n_137), .B(n_488), .Y(n_487) );
AOI21xp5_ASAP7_75t_L g439 ( .A1(n_77), .A2(n_137), .B(n_440), .Y(n_439) );
AOI21xp5_ASAP7_75t_L g467 ( .A1(n_78), .A2(n_137), .B(n_468), .Y(n_467) );
AND2x2_ASAP7_75t_L g479 ( .A(n_79), .B(n_123), .Y(n_479) );
CKINVDCx20_ASAP7_75t_R g725 ( .A(n_80), .Y(n_725) );
NAND2xp5_ASAP7_75t_SL g520 ( .A(n_81), .B(n_158), .Y(n_520) );
NAND2xp5_ASAP7_75t_SL g156 ( .A(n_82), .B(n_128), .Y(n_156) );
AOI22xp5_ASAP7_75t_L g178 ( .A1(n_83), .A2(n_86), .B1(n_128), .B2(n_179), .Y(n_178) );
INVx1_ASAP7_75t_L g112 ( .A(n_85), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_87), .B(n_144), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_88), .B(n_144), .Y(n_222) );
AND2x2_ASAP7_75t_L g443 ( .A(n_89), .B(n_175), .Y(n_443) );
AOI21xp5_ASAP7_75t_L g152 ( .A1(n_90), .A2(n_137), .B(n_153), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_93), .B(n_146), .Y(n_154) );
AOI21xp5_ASAP7_75t_L g494 ( .A1(n_94), .A2(n_137), .B(n_495), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_96), .B(n_146), .Y(n_441) );
INVxp67_ASAP7_75t_L g210 ( .A(n_97), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_98), .B(n_128), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_99), .B(n_146), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g196 ( .A1(n_100), .A2(n_137), .B(n_197), .Y(n_196) );
BUFx2_ASAP7_75t_L g498 ( .A(n_101), .Y(n_498) );
BUFx2_ASAP7_75t_L g741 ( .A(n_102), .Y(n_741) );
BUFx2_ASAP7_75t_SL g750 ( .A(n_102), .Y(n_750) );
OAI21xp5_ASAP7_75t_SL g104 ( .A1(n_105), .A2(n_720), .B(n_727), .Y(n_104) );
INVxp67_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
AO22x2_ASAP7_75t_L g106 ( .A1(n_107), .A2(n_113), .B1(n_426), .B2(n_429), .Y(n_106) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_107), .B(n_114), .Y(n_730) );
AND2x6_ASAP7_75t_SL g107 ( .A(n_108), .B(n_109), .Y(n_107) );
OR2x6_ASAP7_75t_SL g427 ( .A(n_108), .B(n_428), .Y(n_427) );
OR2x2_ASAP7_75t_L g732 ( .A(n_108), .B(n_109), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_108), .B(n_428), .Y(n_743) );
CKINVDCx5p33_ASAP7_75t_R g428 ( .A(n_109), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_111), .B(n_112), .Y(n_110) );
INVx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
XNOR2xp5_ASAP7_75t_L g755 ( .A(n_114), .B(n_756), .Y(n_755) );
AND2x2_ASAP7_75t_L g114 ( .A(n_115), .B(n_348), .Y(n_114) );
NOR3xp33_ASAP7_75t_SL g115 ( .A(n_116), .B(n_272), .C(n_322), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_117), .B(n_252), .Y(n_116) );
AOI21xp5_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_191), .B(n_233), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
NOR2xp33_ASAP7_75t_L g119 ( .A(n_120), .B(n_169), .Y(n_119) );
INVx1_ASAP7_75t_SL g358 ( .A(n_120), .Y(n_358) );
AOI32xp33_ASAP7_75t_L g389 ( .A1(n_120), .A2(n_371), .A3(n_390), .B1(n_391), .B2(n_392), .Y(n_389) );
AND2x2_ASAP7_75t_L g391 ( .A(n_120), .B(n_248), .Y(n_391) );
AND2x4_ASAP7_75t_SL g120 ( .A(n_121), .B(n_149), .Y(n_120) );
HB1xp67_ASAP7_75t_L g170 ( .A(n_121), .Y(n_170) );
INVx5_ASAP7_75t_L g251 ( .A(n_121), .Y(n_251) );
OR2x2_ASAP7_75t_L g258 ( .A(n_121), .B(n_250), .Y(n_258) );
INVx2_ASAP7_75t_L g263 ( .A(n_121), .Y(n_263) );
AND2x2_ASAP7_75t_L g275 ( .A(n_121), .B(n_150), .Y(n_275) );
AND2x2_ASAP7_75t_L g280 ( .A(n_121), .B(n_160), .Y(n_280) );
OR2x2_ASAP7_75t_L g287 ( .A(n_121), .B(n_172), .Y(n_287) );
AND2x4_ASAP7_75t_L g296 ( .A(n_121), .B(n_161), .Y(n_296) );
O2A1O1Ixp33_ASAP7_75t_SL g338 ( .A1(n_121), .A2(n_254), .B(n_289), .C(n_327), .Y(n_338) );
OR2x6_ASAP7_75t_L g121 ( .A(n_122), .B(n_126), .Y(n_121) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_123), .Y(n_158) );
AND2x2_ASAP7_75t_SL g123 ( .A(n_124), .B(n_125), .Y(n_123) );
AND2x4_ASAP7_75t_L g148 ( .A(n_124), .B(n_125), .Y(n_148) );
AOI21xp5_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_136), .B(n_148), .Y(n_126) );
AND2x4_ASAP7_75t_L g128 ( .A(n_129), .B(n_134), .Y(n_128) );
INVx1_ASAP7_75t_L g215 ( .A(n_129), .Y(n_215) );
AND2x4_ASAP7_75t_L g129 ( .A(n_130), .B(n_132), .Y(n_129) );
AND2x6_ASAP7_75t_L g144 ( .A(n_130), .B(n_139), .Y(n_144) );
INVx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
AND2x4_ASAP7_75t_L g146 ( .A(n_132), .B(n_141), .Y(n_146) );
INVx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx5_ASAP7_75t_L g147 ( .A(n_134), .Y(n_147) );
AND2x2_ASAP7_75t_L g140 ( .A(n_135), .B(n_141), .Y(n_140) );
HB1xp67_ASAP7_75t_L g182 ( .A(n_135), .Y(n_182) );
AND2x6_ASAP7_75t_L g137 ( .A(n_138), .B(n_140), .Y(n_137) );
BUFx3_ASAP7_75t_L g183 ( .A(n_138), .Y(n_183) );
INVx2_ASAP7_75t_L g189 ( .A(n_139), .Y(n_189) );
AND2x4_ASAP7_75t_L g185 ( .A(n_140), .B(n_186), .Y(n_185) );
INVx2_ASAP7_75t_L g181 ( .A(n_141), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_145), .B(n_147), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_144), .B(n_498), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g153 ( .A1(n_147), .A2(n_154), .B(n_155), .Y(n_153) );
AOI21xp5_ASAP7_75t_L g164 ( .A1(n_147), .A2(n_165), .B(n_166), .Y(n_164) );
AOI21xp5_ASAP7_75t_L g197 ( .A1(n_147), .A2(n_198), .B(n_199), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_147), .A2(n_221), .B(n_222), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_147), .A2(n_229), .B(n_230), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g440 ( .A1(n_147), .A2(n_441), .B(n_442), .Y(n_440) );
AOI21xp5_ASAP7_75t_L g449 ( .A1(n_147), .A2(n_450), .B(n_451), .Y(n_449) );
AOI21xp5_ASAP7_75t_L g457 ( .A1(n_147), .A2(n_458), .B(n_459), .Y(n_457) );
AOI21xp5_ASAP7_75t_L g468 ( .A1(n_147), .A2(n_469), .B(n_470), .Y(n_468) );
AOI21xp5_ASAP7_75t_L g475 ( .A1(n_147), .A2(n_476), .B(n_477), .Y(n_475) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_147), .A2(n_489), .B(n_490), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_147), .A2(n_496), .B(n_497), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g204 ( .A(n_148), .B(n_205), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g206 ( .A(n_148), .B(n_207), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_148), .B(n_210), .Y(n_209) );
NOR3xp33_ASAP7_75t_L g213 ( .A(n_148), .B(n_214), .C(n_215), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g465 ( .A1(n_148), .A2(n_466), .B(n_467), .Y(n_465) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_148), .A2(n_486), .B(n_487), .Y(n_485) );
INVx3_ASAP7_75t_SL g288 ( .A(n_149), .Y(n_288) );
AND2x2_ASAP7_75t_L g334 ( .A(n_149), .B(n_251), .Y(n_334) );
AND2x4_ASAP7_75t_L g149 ( .A(n_150), .B(n_160), .Y(n_149) );
AND2x2_ASAP7_75t_L g171 ( .A(n_150), .B(n_172), .Y(n_171) );
OR2x2_ASAP7_75t_L g265 ( .A(n_150), .B(n_161), .Y(n_265) );
AND2x2_ASAP7_75t_L g269 ( .A(n_150), .B(n_248), .Y(n_269) );
INVx1_ASAP7_75t_L g295 ( .A(n_150), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_150), .B(n_161), .Y(n_317) );
INVx2_ASAP7_75t_L g321 ( .A(n_150), .Y(n_321) );
HB1xp67_ASAP7_75t_L g331 ( .A(n_150), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_150), .B(n_251), .Y(n_398) );
AO21x2_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_157), .B(n_159), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_152), .B(n_156), .Y(n_151) );
AO21x2_ASAP7_75t_L g161 ( .A1(n_157), .A2(n_162), .B(n_168), .Y(n_161) );
AO21x2_ASAP7_75t_L g250 ( .A1(n_157), .A2(n_162), .B(n_168), .Y(n_250) );
AOI21x1_ASAP7_75t_L g446 ( .A1(n_157), .A2(n_447), .B(n_453), .Y(n_446) );
CKINVDCx5p33_ASAP7_75t_R g157 ( .A(n_158), .Y(n_157) );
OA21x2_ASAP7_75t_L g218 ( .A1(n_158), .A2(n_219), .B(n_223), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g437 ( .A1(n_158), .A2(n_438), .B(n_439), .Y(n_437) );
AO21x2_ASAP7_75t_L g521 ( .A1(n_158), .A2(n_522), .B(n_523), .Y(n_521) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
AND2x2_ASAP7_75t_L g332 ( .A(n_161), .B(n_172), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_163), .B(n_167), .Y(n_162) );
AND2x2_ASAP7_75t_L g169 ( .A(n_170), .B(n_171), .Y(n_169) );
INVx1_ASAP7_75t_L g342 ( .A(n_170), .Y(n_342) );
NAND2xp33_ASAP7_75t_SL g367 ( .A(n_170), .B(n_259), .Y(n_367) );
AND2x2_ASAP7_75t_L g409 ( .A(n_171), .B(n_251), .Y(n_409) );
AND2x2_ASAP7_75t_L g320 ( .A(n_172), .B(n_321), .Y(n_320) );
BUFx2_ASAP7_75t_L g383 ( .A(n_172), .Y(n_383) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
BUFx6f_ASAP7_75t_L g248 ( .A(n_173), .Y(n_248) );
AOI21x1_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_177), .B(n_190), .Y(n_173) );
INVx2_ASAP7_75t_SL g174 ( .A(n_175), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_175), .A2(n_195), .B(n_196), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_175), .A2(n_493), .B(n_494), .Y(n_492) );
BUFx4f_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx3_ASAP7_75t_L g212 ( .A(n_176), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_178), .B(n_184), .Y(n_177) );
AOI22xp5_ASAP7_75t_L g203 ( .A1(n_179), .A2(n_185), .B1(n_204), .B2(n_206), .Y(n_203) );
AND2x4_ASAP7_75t_L g179 ( .A(n_180), .B(n_183), .Y(n_179) );
AND2x2_ASAP7_75t_L g180 ( .A(n_181), .B(n_182), .Y(n_180) );
NOR2x1p5_ASAP7_75t_L g186 ( .A(n_187), .B(n_188), .Y(n_186) );
INVx3_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
AOI22xp5_ASAP7_75t_L g413 ( .A1(n_191), .A2(n_274), .B1(n_376), .B2(n_414), .Y(n_413) );
AND2x2_ASAP7_75t_L g191 ( .A(n_192), .B(n_216), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_192), .B(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_192), .B(n_299), .Y(n_298) );
AND2x4_ASAP7_75t_L g192 ( .A(n_193), .B(n_201), .Y(n_192) );
INVx2_ASAP7_75t_L g239 ( .A(n_193), .Y(n_239) );
OR2x2_ASAP7_75t_L g243 ( .A(n_193), .B(n_244), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_193), .B(n_256), .Y(n_261) );
AND2x4_ASAP7_75t_SL g271 ( .A(n_193), .B(n_202), .Y(n_271) );
OR2x2_ASAP7_75t_L g278 ( .A(n_193), .B(n_218), .Y(n_278) );
OR2x2_ASAP7_75t_L g290 ( .A(n_193), .B(n_202), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_193), .B(n_218), .Y(n_304) );
INVx1_ASAP7_75t_L g309 ( .A(n_193), .Y(n_309) );
HB1xp67_ASAP7_75t_L g327 ( .A(n_193), .Y(n_327) );
AND2x2_ASAP7_75t_L g390 ( .A(n_193), .B(n_310), .Y(n_390) );
INVx2_ASAP7_75t_L g394 ( .A(n_193), .Y(n_394) );
OR2x2_ASAP7_75t_L g401 ( .A(n_193), .B(n_291), .Y(n_401) );
OR2x2_ASAP7_75t_L g423 ( .A(n_193), .B(n_424), .Y(n_423) );
OR2x6_ASAP7_75t_L g193 ( .A(n_194), .B(n_200), .Y(n_193) );
AND2x2_ASAP7_75t_L g240 ( .A(n_201), .B(n_241), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_201), .B(n_224), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_201), .B(n_300), .Y(n_362) );
INVx3_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx1_ASAP7_75t_L g259 ( .A(n_202), .Y(n_259) );
AND2x4_ASAP7_75t_L g310 ( .A(n_202), .B(n_311), .Y(n_310) );
NOR2xp33_ASAP7_75t_L g324 ( .A(n_202), .B(n_255), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_202), .B(n_356), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_202), .B(n_244), .Y(n_403) );
AND2x4_ASAP7_75t_L g202 ( .A(n_203), .B(n_208), .Y(n_202) );
INVx3_ASAP7_75t_L g472 ( .A(n_211), .Y(n_472) );
INVx4_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
AOI21x1_ASAP7_75t_L g225 ( .A1(n_212), .A2(n_226), .B(n_232), .Y(n_225) );
AO21x2_ASAP7_75t_L g454 ( .A1(n_212), .A2(n_455), .B(n_461), .Y(n_454) );
AND2x2_ASAP7_75t_L g270 ( .A(n_216), .B(n_271), .Y(n_270) );
AO221x1_ASAP7_75t_L g344 ( .A1(n_216), .A2(n_259), .B1(n_290), .B2(n_345), .C(n_346), .Y(n_344) );
OAI322xp33_ASAP7_75t_L g396 ( .A1(n_216), .A2(n_316), .A3(n_397), .B1(n_399), .B2(n_400), .C1(n_401), .C2(n_402), .Y(n_396) );
AND2x2_ASAP7_75t_L g216 ( .A(n_217), .B(n_224), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
BUFx3_ASAP7_75t_L g238 ( .A(n_218), .Y(n_238) );
INVx2_ASAP7_75t_L g244 ( .A(n_218), .Y(n_244) );
AND2x2_ASAP7_75t_L g256 ( .A(n_218), .B(n_224), .Y(n_256) );
INVx1_ASAP7_75t_L g301 ( .A(n_218), .Y(n_301) );
HB1xp67_ASAP7_75t_L g357 ( .A(n_218), .Y(n_357) );
INVx1_ASAP7_75t_L g241 ( .A(n_224), .Y(n_241) );
OR2x2_ASAP7_75t_L g291 ( .A(n_224), .B(n_244), .Y(n_291) );
INVx2_ASAP7_75t_L g311 ( .A(n_224), .Y(n_311) );
INVx1_ASAP7_75t_L g364 ( .A(n_224), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_224), .B(n_394), .Y(n_393) );
INVx3_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_227), .B(n_231), .Y(n_226) );
INVx1_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
OAI21xp33_ASAP7_75t_SL g234 ( .A1(n_235), .A2(n_242), .B(n_245), .Y(n_234) );
AOI221xp5_ASAP7_75t_L g273 ( .A1(n_235), .A2(n_274), .B1(n_276), .B2(n_280), .C(n_281), .Y(n_273) );
INVx1_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_237), .B(n_240), .Y(n_236) );
NOR2x1p5_ASAP7_75t_L g237 ( .A(n_238), .B(n_239), .Y(n_237) );
INVx1_ASAP7_75t_L g360 ( .A(n_239), .Y(n_360) );
INVx1_ASAP7_75t_SL g279 ( .A(n_240), .Y(n_279) );
OAI21xp5_ASAP7_75t_L g384 ( .A1(n_240), .A2(n_385), .B(n_387), .Y(n_384) );
HB1xp67_ASAP7_75t_L g284 ( .A(n_241), .Y(n_284) );
INVx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
HB1xp67_ASAP7_75t_L g347 ( .A(n_244), .Y(n_347) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_247), .B(n_249), .Y(n_246) );
OAI211xp5_ASAP7_75t_L g322 ( .A1(n_247), .A2(n_323), .B(n_328), .C(n_339), .Y(n_322) );
OR2x2_ASAP7_75t_L g412 ( .A(n_247), .B(n_317), .Y(n_412) );
AND2x2_ASAP7_75t_L g414 ( .A(n_247), .B(n_280), .Y(n_414) );
INVx2_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
OR2x2_ASAP7_75t_L g254 ( .A(n_248), .B(n_255), .Y(n_254) );
OR2x2_ASAP7_75t_L g316 ( .A(n_248), .B(n_317), .Y(n_316) );
AND2x4_ASAP7_75t_L g354 ( .A(n_248), .B(n_321), .Y(n_354) );
OA33x2_ASAP7_75t_L g361 ( .A1(n_248), .A2(n_278), .A3(n_362), .B1(n_363), .B2(n_365), .B3(n_367), .Y(n_361) );
OR2x2_ASAP7_75t_L g372 ( .A(n_248), .B(n_357), .Y(n_372) );
NAND2xp5_ASAP7_75t_SL g386 ( .A(n_248), .B(n_296), .Y(n_386) );
AND2x4_ASAP7_75t_L g249 ( .A(n_250), .B(n_251), .Y(n_249) );
AND2x2_ASAP7_75t_L g274 ( .A(n_250), .B(n_275), .Y(n_274) );
AOI22xp33_ASAP7_75t_SL g323 ( .A1(n_250), .A2(n_280), .B1(n_324), .B2(n_325), .Y(n_323) );
NAND3xp33_ASAP7_75t_L g363 ( .A(n_251), .B(n_331), .C(n_364), .Y(n_363) );
AOI322xp5_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_257), .A3(n_259), .B1(n_260), .B2(n_262), .C1(n_266), .C2(n_270), .Y(n_252) );
INVx3_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
OR2x2_ASAP7_75t_L g359 ( .A(n_255), .B(n_360), .Y(n_359) );
INVx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
A2O1A1Ixp33_ASAP7_75t_L g314 ( .A1(n_256), .A2(n_271), .B(n_315), .C(n_318), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_257), .B(n_320), .Y(n_319) );
INVx1_ASAP7_75t_SL g257 ( .A(n_258), .Y(n_257) );
NAND4xp25_ASAP7_75t_SL g378 ( .A(n_258), .B(n_287), .C(n_379), .D(n_381), .Y(n_378) );
INVx1_ASAP7_75t_SL g260 ( .A(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
INVx2_ASAP7_75t_L g268 ( .A(n_263), .Y(n_268) );
OR2x2_ASAP7_75t_L g313 ( .A(n_263), .B(n_265), .Y(n_313) );
AND2x2_ASAP7_75t_L g382 ( .A(n_264), .B(n_383), .Y(n_382) );
INVx2_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_268), .B(n_269), .Y(n_267) );
AND2x2_ASAP7_75t_L g387 ( .A(n_268), .B(n_382), .Y(n_387) );
BUFx2_ASAP7_75t_L g380 ( .A(n_269), .Y(n_380) );
INVx1_ASAP7_75t_SL g410 ( .A(n_270), .Y(n_410) );
AND2x4_ASAP7_75t_L g346 ( .A(n_271), .B(n_347), .Y(n_346) );
INVx1_ASAP7_75t_SL g399 ( .A(n_271), .Y(n_399) );
NAND3xp33_ASAP7_75t_L g272 ( .A(n_273), .B(n_292), .C(n_314), .Y(n_272) );
INVx1_ASAP7_75t_SL g276 ( .A(n_277), .Y(n_276) );
OR2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
INVx1_ASAP7_75t_SL g336 ( .A(n_278), .Y(n_336) );
OAI211xp5_ASAP7_75t_L g404 ( .A1(n_278), .A2(n_405), .B(n_406), .C(n_415), .Y(n_404) );
OR2x2_ASAP7_75t_L g326 ( .A(n_279), .B(n_327), .Y(n_326) );
OAI22xp33_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_285), .B1(n_288), .B2(n_289), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_283), .B(n_366), .Y(n_365) );
INVxp67_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_286), .B(n_288), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_286), .B(n_343), .Y(n_425) );
INVx1_ASAP7_75t_SL g286 ( .A(n_287), .Y(n_286) );
OR2x2_ASAP7_75t_L g400 ( .A(n_287), .B(n_288), .Y(n_400) );
OR2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
INVx1_ASAP7_75t_L g345 ( .A(n_291), .Y(n_345) );
AOI222xp33_ASAP7_75t_L g292 ( .A1(n_293), .A2(n_297), .B1(n_302), .B2(n_306), .C1(n_307), .C2(n_312), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
HB1xp67_ASAP7_75t_L g306 ( .A(n_295), .Y(n_306) );
AND2x2_ASAP7_75t_L g353 ( .A(n_296), .B(n_354), .Y(n_353) );
AOI22xp5_ASAP7_75t_L g368 ( .A1(n_296), .A2(n_369), .B1(n_374), .B2(n_378), .Y(n_368) );
INVx2_ASAP7_75t_SL g421 ( .A(n_296), .Y(n_421) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVxp67_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
HB1xp67_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g377 ( .A(n_301), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_301), .B(n_364), .Y(n_424) );
INVx2_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
OR2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_305), .Y(n_303) );
INVx1_ASAP7_75t_L g337 ( .A(n_305), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_307), .B(n_371), .Y(n_370) );
INVx1_ASAP7_75t_SL g307 ( .A(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
INVx1_ASAP7_75t_L g375 ( .A(n_309), .Y(n_375) );
AND2x2_ASAP7_75t_SL g376 ( .A(n_310), .B(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_L g418 ( .A(n_310), .B(n_347), .Y(n_418) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx1_ASAP7_75t_SL g315 ( .A(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g343 ( .A(n_317), .Y(n_343) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g422 ( .A(n_320), .Y(n_422) );
HB1xp67_ASAP7_75t_L g366 ( .A(n_321), .Y(n_366) );
INVx1_ASAP7_75t_SL g325 ( .A(n_326), .Y(n_325) );
O2A1O1Ixp33_ASAP7_75t_L g328 ( .A1(n_329), .A2(n_333), .B(n_335), .C(n_338), .Y(n_328) );
AND2x2_ASAP7_75t_SL g329 ( .A(n_330), .B(n_332), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
HB1xp67_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g373 ( .A(n_335), .Y(n_373) );
AND2x2_ASAP7_75t_L g335 ( .A(n_336), .B(n_337), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_340), .B(n_344), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
NAND2xp5_ASAP7_75t_SL g341 ( .A(n_342), .B(n_343), .Y(n_341) );
NOR3xp33_ASAP7_75t_L g348 ( .A(n_349), .B(n_388), .C(n_404), .Y(n_348) );
NAND3xp33_ASAP7_75t_L g349 ( .A(n_350), .B(n_368), .C(n_384), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
OAI221xp5_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_355), .B1(n_358), .B2(n_359), .C(n_361), .Y(n_351) );
INVx1_ASAP7_75t_SL g352 ( .A(n_353), .Y(n_352) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
NAND2xp5_ASAP7_75t_SL g369 ( .A(n_370), .B(n_373), .Y(n_369) );
INVx1_ASAP7_75t_SL g371 ( .A(n_372), .Y(n_371) );
AND2x2_ASAP7_75t_L g374 ( .A(n_375), .B(n_376), .Y(n_374) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx2_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
OR2x2_ASAP7_75t_L g397 ( .A(n_383), .B(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g405 ( .A(n_387), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_389), .B(n_395), .Y(n_388) );
INVx2_ASAP7_75t_L g411 ( .A(n_390), .Y(n_411) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
OR2x2_ASAP7_75t_L g402 ( .A(n_393), .B(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
OAI221xp5_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_410), .B1(n_411), .B2(n_412), .C(n_413), .Y(n_407) );
INVxp67_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
OAI22xp5_ASAP7_75t_L g416 ( .A1(n_417), .A2(n_419), .B1(n_423), .B2(n_425), .Y(n_416) );
INVx1_ASAP7_75t_SL g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
NOR2xp33_ASAP7_75t_L g420 ( .A(n_421), .B(n_422), .Y(n_420) );
INVx1_ASAP7_75t_SL g729 ( .A(n_426), .Y(n_729) );
CKINVDCx11_ASAP7_75t_R g426 ( .A(n_427), .Y(n_426) );
OAI21x1_ASAP7_75t_SL g728 ( .A1(n_429), .A2(n_729), .B(n_730), .Y(n_728) );
INVx4_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
AND2x4_ASAP7_75t_L g430 ( .A(n_431), .B(n_628), .Y(n_430) );
NOR3xp33_ASAP7_75t_SL g431 ( .A(n_432), .B(n_551), .C(n_586), .Y(n_431) );
OAI211xp5_ASAP7_75t_L g432 ( .A1(n_433), .A2(n_462), .B(n_513), .C(n_541), .Y(n_432) );
INVx1_ASAP7_75t_SL g433 ( .A(n_434), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_435), .B(n_444), .Y(n_434) );
AND2x2_ASAP7_75t_L g534 ( .A(n_435), .B(n_535), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_435), .B(n_540), .Y(n_574) );
AND2x2_ASAP7_75t_L g599 ( .A(n_435), .B(n_554), .Y(n_599) );
INVx4_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
BUFx2_ASAP7_75t_L g516 ( .A(n_436), .Y(n_516) );
OR2x2_ASAP7_75t_L g537 ( .A(n_436), .B(n_538), .Y(n_537) );
AND2x2_ASAP7_75t_L g545 ( .A(n_436), .B(n_454), .Y(n_545) );
AND2x2_ASAP7_75t_L g553 ( .A(n_436), .B(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g580 ( .A(n_436), .B(n_581), .Y(n_580) );
NOR2x1_ASAP7_75t_L g591 ( .A(n_436), .B(n_583), .Y(n_591) );
AND2x4_ASAP7_75t_L g608 ( .A(n_436), .B(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g646 ( .A(n_436), .Y(n_646) );
AND2x4_ASAP7_75t_SL g651 ( .A(n_436), .B(n_445), .Y(n_651) );
OR2x6_ASAP7_75t_L g436 ( .A(n_437), .B(n_443), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_444), .B(n_534), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_444), .B(n_685), .Y(n_684) );
AND2x2_ASAP7_75t_L g444 ( .A(n_445), .B(n_454), .Y(n_444) );
HB1xp67_ASAP7_75t_L g546 ( .A(n_445), .Y(n_546) );
INVx2_ASAP7_75t_L g582 ( .A(n_445), .Y(n_582) );
INVx1_ASAP7_75t_L g609 ( .A(n_445), .Y(n_609) );
AND2x2_ASAP7_75t_L g708 ( .A(n_445), .B(n_618), .Y(n_708) );
INVx3_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
HB1xp67_ASAP7_75t_L g540 ( .A(n_446), .Y(n_540) );
AND2x2_ASAP7_75t_L g554 ( .A(n_446), .B(n_454), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_448), .B(n_452), .Y(n_447) );
INVx2_ASAP7_75t_L g583 ( .A(n_454), .Y(n_583) );
INVx2_ASAP7_75t_L g618 ( .A(n_454), .Y(n_618) );
OR2x2_ASAP7_75t_L g703 ( .A(n_454), .B(n_535), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_456), .B(n_460), .Y(n_455) );
AOI211xp5_ASAP7_75t_L g462 ( .A1(n_463), .A2(n_480), .B(n_500), .C(n_507), .Y(n_462) );
INVx2_ASAP7_75t_SL g592 ( .A(n_463), .Y(n_592) );
AND2x2_ASAP7_75t_L g598 ( .A(n_463), .B(n_481), .Y(n_598) );
AND2x2_ASAP7_75t_L g463 ( .A(n_464), .B(n_471), .Y(n_463) );
INVx1_ASAP7_75t_L g504 ( .A(n_464), .Y(n_504) );
INVx1_ASAP7_75t_L g510 ( .A(n_464), .Y(n_510) );
INVx2_ASAP7_75t_L g525 ( .A(n_464), .Y(n_525) );
AND2x2_ASAP7_75t_L g549 ( .A(n_464), .B(n_483), .Y(n_549) );
HB1xp67_ASAP7_75t_L g578 ( .A(n_464), .Y(n_578) );
OR2x2_ASAP7_75t_L g658 ( .A(n_464), .B(n_491), .Y(n_658) );
AND2x2_ASAP7_75t_L g524 ( .A(n_471), .B(n_525), .Y(n_524) );
NOR2x1_ASAP7_75t_SL g556 ( .A(n_471), .B(n_491), .Y(n_556) );
AO21x1_ASAP7_75t_SL g471 ( .A1(n_472), .A2(n_473), .B(n_479), .Y(n_471) );
AO21x2_ASAP7_75t_L g506 ( .A1(n_472), .A2(n_473), .B(n_479), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_474), .B(n_478), .Y(n_473) );
INVxp67_ASAP7_75t_SL g480 ( .A(n_481), .Y(n_480) );
AND2x2_ASAP7_75t_L g570 ( .A(n_481), .B(n_503), .Y(n_570) );
AND2x2_ASAP7_75t_L g481 ( .A(n_482), .B(n_491), .Y(n_481) );
OR2x2_ASAP7_75t_L g512 ( .A(n_482), .B(n_491), .Y(n_512) );
BUFx2_ASAP7_75t_L g526 ( .A(n_482), .Y(n_526) );
NOR2xp67_ASAP7_75t_L g577 ( .A(n_482), .B(n_578), .Y(n_577) );
INVx4_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
HB1xp67_ASAP7_75t_L g529 ( .A(n_483), .Y(n_529) );
AND2x2_ASAP7_75t_L g555 ( .A(n_483), .B(n_556), .Y(n_555) );
INVx2_ASAP7_75t_L g565 ( .A(n_483), .Y(n_565) );
NAND2x1_ASAP7_75t_L g603 ( .A(n_483), .B(n_491), .Y(n_603) );
OR2x2_ASAP7_75t_L g678 ( .A(n_483), .B(n_505), .Y(n_678) );
OR2x6_ASAP7_75t_L g483 ( .A(n_484), .B(n_485), .Y(n_483) );
INVx2_ASAP7_75t_SL g501 ( .A(n_491), .Y(n_501) );
AND2x2_ASAP7_75t_L g550 ( .A(n_491), .B(n_505), .Y(n_550) );
AND2x2_ASAP7_75t_L g621 ( .A(n_491), .B(n_622), .Y(n_621) );
BUFx2_ASAP7_75t_L g642 ( .A(n_491), .Y(n_642) );
OR2x6_ASAP7_75t_L g491 ( .A(n_492), .B(n_499), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g500 ( .A(n_501), .B(n_502), .Y(n_500) );
INVx1_ASAP7_75t_SL g502 ( .A(n_503), .Y(n_502) );
AND2x2_ASAP7_75t_L g564 ( .A(n_503), .B(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g503 ( .A(n_504), .B(n_505), .Y(n_503) );
BUFx2_ASAP7_75t_L g559 ( .A(n_504), .Y(n_559) );
AND2x2_ASAP7_75t_L g531 ( .A(n_505), .B(n_532), .Y(n_531) );
INVx2_ASAP7_75t_L g622 ( .A(n_505), .Y(n_622) );
INVx3_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_509), .B(n_511), .Y(n_508) );
OR2x2_ASAP7_75t_L g568 ( .A(n_509), .B(n_569), .Y(n_568) );
AND2x4_ASAP7_75t_SL g610 ( .A(n_509), .B(n_611), .Y(n_610) );
AOI322xp5_ASAP7_75t_L g647 ( .A1(n_509), .A2(n_526), .A3(n_648), .B1(n_650), .B2(n_653), .C1(n_655), .C2(n_657), .Y(n_647) );
AND2x2_ASAP7_75t_L g712 ( .A(n_509), .B(n_713), .Y(n_712) );
INVx3_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_510), .B(n_526), .Y(n_536) );
AOI322xp5_ASAP7_75t_L g587 ( .A1(n_511), .A2(n_588), .A3(n_592), .B1(n_593), .B2(n_596), .C1(n_598), .C2(n_599), .Y(n_587) );
INVx2_ASAP7_75t_SL g511 ( .A(n_512), .Y(n_511) );
OR2x2_ASAP7_75t_L g639 ( .A(n_512), .B(n_592), .Y(n_639) );
OAI22xp5_ASAP7_75t_L g698 ( .A1(n_512), .A2(n_699), .B1(n_701), .B2(n_704), .Y(n_698) );
OR2x2_ASAP7_75t_L g716 ( .A(n_512), .B(n_665), .Y(n_716) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_514), .A2(n_526), .B(n_527), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_515), .B(n_517), .Y(n_514) );
AOI221xp5_ASAP7_75t_SL g566 ( .A1(n_515), .A2(n_542), .B1(n_567), .B2(n_570), .C(n_571), .Y(n_566) );
AND2x2_ASAP7_75t_L g593 ( .A(n_515), .B(n_594), .Y(n_593) );
INVx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_516), .B(n_633), .Y(n_632) );
OR2x2_ASAP7_75t_L g635 ( .A(n_516), .B(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g664 ( .A(n_517), .Y(n_664) );
AND2x2_ASAP7_75t_L g517 ( .A(n_518), .B(n_524), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_518), .B(n_539), .Y(n_538) );
INVx2_ASAP7_75t_L g606 ( .A(n_518), .Y(n_606) );
OR2x2_ASAP7_75t_L g613 ( .A(n_518), .B(n_614), .Y(n_613) );
INVx3_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
AND2x2_ASAP7_75t_L g656 ( .A(n_519), .B(n_618), .Y(n_656) );
AND2x4_ASAP7_75t_L g519 ( .A(n_520), .B(n_521), .Y(n_519) );
AND2x4_ASAP7_75t_L g535 ( .A(n_520), .B(n_521), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_524), .B(n_585), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_524), .B(n_565), .Y(n_661) );
INVx1_ASAP7_75t_L g665 ( .A(n_524), .Y(n_665) );
INVx1_ASAP7_75t_L g532 ( .A(n_525), .Y(n_532) );
OAI22xp5_ASAP7_75t_L g527 ( .A1(n_528), .A2(n_533), .B1(n_536), .B2(n_537), .Y(n_527) );
OR2x2_ASAP7_75t_L g528 ( .A(n_529), .B(n_530), .Y(n_528) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
BUFx2_ASAP7_75t_SL g643 ( .A(n_531), .Y(n_643) );
AND2x2_ASAP7_75t_L g700 ( .A(n_532), .B(n_556), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_534), .B(n_563), .Y(n_562) );
NOR2xp33_ASAP7_75t_SL g572 ( .A(n_534), .B(n_573), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_534), .B(n_693), .Y(n_692) );
BUFx3_ASAP7_75t_L g560 ( .A(n_535), .Y(n_560) );
INVx2_ASAP7_75t_L g590 ( .A(n_535), .Y(n_590) );
AND2x2_ASAP7_75t_L g633 ( .A(n_535), .B(n_617), .Y(n_633) );
INVx1_ASAP7_75t_L g547 ( .A(n_537), .Y(n_547) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
OAI21xp5_ASAP7_75t_SL g541 ( .A1(n_542), .A2(n_547), .B(n_548), .Y(n_541) );
INVx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_545), .B(n_546), .Y(n_544) );
INVx1_ASAP7_75t_L g626 ( .A(n_545), .Y(n_626) );
INVx2_ASAP7_75t_L g614 ( .A(n_546), .Y(n_614) );
AND2x2_ASAP7_75t_L g548 ( .A(n_549), .B(n_550), .Y(n_548) );
AND2x2_ASAP7_75t_L g611 ( .A(n_550), .B(n_565), .Y(n_611) );
OAI21xp5_ASAP7_75t_L g671 ( .A1(n_550), .A2(n_648), .B(n_672), .Y(n_671) );
NAND2xp5_ASAP7_75t_SL g551 ( .A(n_552), .B(n_566), .Y(n_551) );
AOI32xp33_ASAP7_75t_L g552 ( .A1(n_553), .A2(n_555), .A3(n_557), .B1(n_561), .B2(n_564), .Y(n_552) );
HB1xp67_ASAP7_75t_L g627 ( .A(n_553), .Y(n_627) );
AOI221xp5_ASAP7_75t_L g659 ( .A1(n_553), .A2(n_642), .B1(n_660), .B2(n_662), .C(n_668), .Y(n_659) );
AND2x2_ASAP7_75t_L g679 ( .A(n_553), .B(n_560), .Y(n_679) );
BUFx2_ASAP7_75t_L g563 ( .A(n_554), .Y(n_563) );
INVx1_ASAP7_75t_L g688 ( .A(n_554), .Y(n_688) );
INVx1_ASAP7_75t_L g693 ( .A(n_554), .Y(n_693) );
INVx1_ASAP7_75t_SL g686 ( .A(n_555), .Y(n_686) );
INVx2_ASAP7_75t_L g569 ( .A(n_556), .Y(n_569) );
AND2x2_ASAP7_75t_L g681 ( .A(n_557), .B(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
OR2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_560), .Y(n_558) );
AND2x2_ASAP7_75t_L g653 ( .A(n_559), .B(n_654), .Y(n_653) );
OR2x2_ASAP7_75t_L g625 ( .A(n_560), .B(n_626), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_560), .B(n_651), .Y(n_673) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx2_ASAP7_75t_L g585 ( .A(n_565), .Y(n_585) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
OR2x2_ASAP7_75t_L g575 ( .A(n_569), .B(n_576), .Y(n_575) );
OR2x2_ASAP7_75t_L g584 ( .A(n_569), .B(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g689 ( .A(n_570), .Y(n_689) );
OAI22xp5_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_575), .B1(n_579), .B2(n_584), .Y(n_571) );
INVx2_ASAP7_75t_SL g663 ( .A(n_573), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_573), .B(n_702), .Y(n_704) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
AOI21xp5_ASAP7_75t_L g668 ( .A1(n_575), .A2(n_669), .B(n_670), .Y(n_668) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g620 ( .A(n_577), .B(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g648 ( .A(n_580), .B(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g595 ( .A(n_581), .Y(n_595) );
AND2x2_ASAP7_75t_L g581 ( .A(n_582), .B(n_583), .Y(n_581) );
INVx1_ASAP7_75t_L g637 ( .A(n_583), .Y(n_637) );
INVx1_ASAP7_75t_L g682 ( .A(n_584), .Y(n_682) );
NAND3xp33_ASAP7_75t_L g586 ( .A(n_587), .B(n_600), .C(n_623), .Y(n_586) );
AND2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_591), .Y(n_588) );
INVx2_ASAP7_75t_L g649 ( .A(n_589), .Y(n_649) );
AND2x2_ASAP7_75t_L g667 ( .A(n_589), .B(n_608), .Y(n_667) );
OR2x2_ASAP7_75t_L g706 ( .A(n_589), .B(n_707), .Y(n_706) );
INVx2_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_590), .B(n_637), .Y(n_636) );
OR2x2_ASAP7_75t_L g602 ( .A(n_592), .B(n_603), .Y(n_602) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
OR2x2_ASAP7_75t_L g669 ( .A(n_595), .B(n_606), .Y(n_669) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_598), .B(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g710 ( .A(n_598), .Y(n_710) );
AOI221xp5_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_604), .B1(n_608), .B2(n_610), .C(n_612), .Y(n_600) );
OAI21xp5_ASAP7_75t_L g623 ( .A1(n_601), .A2(n_624), .B(n_627), .Y(n_623) );
INVx2_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx3_ASAP7_75t_L g654 ( .A(n_603), .Y(n_654) );
NOR2xp33_ASAP7_75t_L g696 ( .A(n_603), .B(n_697), .Y(n_696) );
INVxp33_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
OR2x2_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .Y(n_605) );
INVx2_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g615 ( .A(n_611), .Y(n_615) );
OAI22xp33_ASAP7_75t_L g612 ( .A1(n_613), .A2(n_615), .B1(n_616), .B2(n_619), .Y(n_612) );
INVx2_ASAP7_75t_L g718 ( .A(n_614), .Y(n_718) );
BUFx2_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVxp67_ASAP7_75t_L g697 ( .A(n_622), .Y(n_697) );
INVx1_ASAP7_75t_SL g624 ( .A(n_625), .Y(n_624) );
NOR2x1_ASAP7_75t_L g628 ( .A(n_629), .B(n_674), .Y(n_628) );
NAND4xp25_ASAP7_75t_L g629 ( .A(n_630), .B(n_647), .C(n_659), .D(n_671), .Y(n_629) );
O2A1O1Ixp33_ASAP7_75t_L g630 ( .A1(n_631), .A2(n_634), .B(n_638), .C(n_640), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g670 ( .A(n_633), .Y(n_670) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
OAI21xp5_ASAP7_75t_L g640 ( .A1(n_635), .A2(n_641), .B(n_644), .Y(n_640) );
INVx2_ASAP7_75t_L g719 ( .A(n_636), .Y(n_719) );
NOR2xp33_ASAP7_75t_L g645 ( .A(n_637), .B(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g652 ( .A(n_637), .Y(n_652) );
INVx2_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_642), .B(n_643), .Y(n_641) );
OR2x2_ASAP7_75t_L g714 ( .A(n_642), .B(n_678), .Y(n_714) );
INVxp67_ASAP7_75t_SL g685 ( .A(n_649), .Y(n_685) );
AND2x2_ASAP7_75t_SL g650 ( .A(n_651), .B(n_652), .Y(n_650) );
AND2x2_ASAP7_75t_L g655 ( .A(n_651), .B(n_656), .Y(n_655) );
AOI21xp5_ASAP7_75t_L g680 ( .A1(n_651), .A2(n_681), .B(n_683), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_651), .B(n_702), .Y(n_701) );
INVx2_ASAP7_75t_SL g709 ( .A(n_651), .Y(n_709) );
INVxp67_ASAP7_75t_SL g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
OAI22xp33_ASAP7_75t_SL g662 ( .A1(n_663), .A2(n_664), .B1(n_665), .B2(n_666), .Y(n_662) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
NAND4xp25_ASAP7_75t_L g674 ( .A(n_675), .B(n_680), .C(n_690), .D(n_711), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_676), .B(n_679), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
HB1xp67_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
OAI22xp5_ASAP7_75t_L g683 ( .A1(n_684), .A2(n_686), .B1(n_687), .B2(n_689), .Y(n_683) );
HB1xp67_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
AOI211xp5_ASAP7_75t_SL g690 ( .A1(n_691), .A2(n_694), .B(n_698), .C(n_705), .Y(n_690) );
INVxp67_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx2_ASAP7_75t_SL g702 ( .A(n_703), .Y(n_702) );
AOI21xp33_ASAP7_75t_L g705 ( .A1(n_706), .A2(n_709), .B(n_710), .Y(n_705) );
INVx1_ASAP7_75t_SL g707 ( .A(n_708), .Y(n_707) );
OAI21xp5_ASAP7_75t_SL g711 ( .A1(n_712), .A2(n_715), .B(n_717), .Y(n_711) );
INVx1_ASAP7_75t_SL g713 ( .A(n_714), .Y(n_713) );
INVx2_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
AND2x2_ASAP7_75t_L g717 ( .A(n_718), .B(n_719), .Y(n_717) );
INVxp67_ASAP7_75t_SL g723 ( .A(n_724), .Y(n_723) );
INVx2_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
CKINVDCx20_ASAP7_75t_R g733 ( .A(n_734), .Y(n_733) );
INVx2_ASAP7_75t_SL g734 ( .A(n_735), .Y(n_734) );
AND2x2_ASAP7_75t_L g735 ( .A(n_736), .B(n_742), .Y(n_735) );
INVxp67_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
NAND2xp5_ASAP7_75t_SL g737 ( .A(n_738), .B(n_741), .Y(n_737) );
INVx2_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
AOI21xp5_ASAP7_75t_L g747 ( .A1(n_739), .A2(n_748), .B(n_751), .Y(n_747) );
OR2x2_ASAP7_75t_SL g770 ( .A(n_739), .B(n_741), .Y(n_770) );
INVx1_ASAP7_75t_L g769 ( .A(n_742), .Y(n_769) );
BUFx2_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
BUFx2_ASAP7_75t_L g752 ( .A(n_743), .Y(n_752) );
BUFx3_ASAP7_75t_L g767 ( .A(n_743), .Y(n_767) );
INVx1_ASAP7_75t_SL g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_SL g746 ( .A(n_747), .Y(n_746) );
CKINVDCx11_ASAP7_75t_R g748 ( .A(n_749), .Y(n_748) );
CKINVDCx8_ASAP7_75t_R g749 ( .A(n_750), .Y(n_749) );
INVx2_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
O2A1O1Ixp33_ASAP7_75t_R g753 ( .A1(n_754), .A2(n_764), .B(n_768), .C(n_770), .Y(n_753) );
AOI22xp5_ASAP7_75t_L g754 ( .A1(n_755), .A2(n_759), .B1(n_762), .B2(n_763), .Y(n_754) );
INVx2_ASAP7_75t_L g762 ( .A(n_755), .Y(n_762) );
INVx1_ASAP7_75t_L g763 ( .A(n_759), .Y(n_763) );
CKINVDCx20_ASAP7_75t_R g764 ( .A(n_765), .Y(n_764) );
CKINVDCx11_ASAP7_75t_R g765 ( .A(n_766), .Y(n_765) );
CKINVDCx20_ASAP7_75t_R g766 ( .A(n_767), .Y(n_766) );
endmodule