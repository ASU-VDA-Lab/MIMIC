module fake_netlist_1_4934_n_586 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_586);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_586;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_461;
wire n_305;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_540;
wire n_563;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_554;
wire n_447;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_420;
wire n_446;
wire n_423;
wire n_342;
wire n_165;
wire n_370;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_357;
wire n_90;
wire n_245;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g82 ( .A(n_21), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_51), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_36), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_10), .Y(n_85) );
BUFx6f_ASAP7_75t_L g86 ( .A(n_16), .Y(n_86) );
INVxp67_ASAP7_75t_L g87 ( .A(n_11), .Y(n_87) );
BUFx3_ASAP7_75t_L g88 ( .A(n_76), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_47), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_41), .Y(n_90) );
INVx2_ASAP7_75t_L g91 ( .A(n_33), .Y(n_91) );
INVxp33_ASAP7_75t_L g92 ( .A(n_64), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_57), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_34), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_44), .Y(n_95) );
INVxp33_ASAP7_75t_SL g96 ( .A(n_24), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_1), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_59), .Y(n_98) );
INVx2_ASAP7_75t_L g99 ( .A(n_67), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_66), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_16), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_2), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_29), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_70), .Y(n_104) );
BUFx2_ASAP7_75t_SL g105 ( .A(n_81), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_55), .Y(n_106) );
INVx2_ASAP7_75t_L g107 ( .A(n_43), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_53), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_12), .Y(n_109) );
XOR2xp5_ASAP7_75t_L g110 ( .A(n_11), .B(n_45), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_35), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_30), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_46), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_17), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_12), .Y(n_115) );
INVxp67_ASAP7_75t_SL g116 ( .A(n_62), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_4), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_1), .Y(n_118) );
CKINVDCx16_ASAP7_75t_R g119 ( .A(n_63), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_13), .Y(n_120) );
INVxp67_ASAP7_75t_L g121 ( .A(n_54), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_39), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_27), .Y(n_123) );
AND2x4_ASAP7_75t_L g124 ( .A(n_117), .B(n_85), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_85), .B(n_0), .Y(n_125) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_88), .Y(n_126) );
HB1xp67_ASAP7_75t_L g127 ( .A(n_97), .Y(n_127) );
AND2x2_ASAP7_75t_L g128 ( .A(n_92), .B(n_0), .Y(n_128) );
HB1xp67_ASAP7_75t_L g129 ( .A(n_97), .Y(n_129) );
AND2x4_ASAP7_75t_L g130 ( .A(n_117), .B(n_2), .Y(n_130) );
AND2x4_ASAP7_75t_L g131 ( .A(n_101), .B(n_3), .Y(n_131) );
AND2x4_ASAP7_75t_L g132 ( .A(n_101), .B(n_3), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_119), .Y(n_133) );
HB1xp67_ASAP7_75t_L g134 ( .A(n_109), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_109), .B(n_4), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_114), .B(n_5), .Y(n_136) );
BUFx2_ASAP7_75t_L g137 ( .A(n_87), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_96), .Y(n_138) );
OAI22xp5_ASAP7_75t_L g139 ( .A1(n_110), .A2(n_5), .B1(n_6), .B2(n_7), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_114), .B(n_6), .Y(n_140) );
AND2x2_ASAP7_75t_L g141 ( .A(n_115), .B(n_7), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_82), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_93), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_82), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_91), .Y(n_145) );
CKINVDCx20_ASAP7_75t_R g146 ( .A(n_110), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_84), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_126), .Y(n_148) );
BUFx2_ASAP7_75t_L g149 ( .A(n_143), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_126), .Y(n_150) );
AND2x2_ASAP7_75t_L g151 ( .A(n_127), .B(n_115), .Y(n_151) );
AO22x2_ASAP7_75t_L g152 ( .A1(n_139), .A2(n_108), .B1(n_84), .B2(n_89), .Y(n_152) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_126), .Y(n_153) );
INVx4_ASAP7_75t_SL g154 ( .A(n_131), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_126), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_145), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_145), .Y(n_157) );
NAND2xp5_ASAP7_75t_SL g158 ( .A(n_142), .B(n_121), .Y(n_158) );
NOR2xp33_ASAP7_75t_L g159 ( .A(n_138), .B(n_83), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_142), .B(n_91), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_145), .Y(n_161) );
BUFx3_ASAP7_75t_L g162 ( .A(n_126), .Y(n_162) );
NOR2xp33_ASAP7_75t_L g163 ( .A(n_137), .B(n_104), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_137), .B(n_106), .Y(n_164) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_126), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_126), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_131), .Y(n_167) );
INVx2_ASAP7_75t_SL g168 ( .A(n_144), .Y(n_168) );
AND2x2_ASAP7_75t_L g169 ( .A(n_127), .B(n_120), .Y(n_169) );
AOI22xp33_ASAP7_75t_L g170 ( .A1(n_131), .A2(n_120), .B1(n_118), .B2(n_102), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_131), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_144), .B(n_99), .Y(n_172) );
BUFx3_ASAP7_75t_L g173 ( .A(n_124), .Y(n_173) );
INVx4_ASAP7_75t_SL g174 ( .A(n_132), .Y(n_174) );
BUFx3_ASAP7_75t_L g175 ( .A(n_124), .Y(n_175) );
INVx1_ASAP7_75t_SL g176 ( .A(n_154), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_168), .B(n_128), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_156), .Y(n_178) );
INVx2_ASAP7_75t_SL g179 ( .A(n_154), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_168), .B(n_128), .Y(n_180) );
AOI22xp33_ASAP7_75t_L g181 ( .A1(n_173), .A2(n_132), .B1(n_130), .B2(n_141), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_168), .B(n_129), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_173), .B(n_129), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_156), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_162), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_151), .B(n_134), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_162), .Y(n_187) );
INVx2_ASAP7_75t_SL g188 ( .A(n_154), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_157), .Y(n_189) );
OAI22xp33_ASAP7_75t_L g190 ( .A1(n_149), .A2(n_139), .B1(n_133), .B2(n_134), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_162), .Y(n_191) );
AOI22xp33_ASAP7_75t_L g192 ( .A1(n_173), .A2(n_132), .B1(n_130), .B2(n_141), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_153), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_154), .B(n_132), .Y(n_194) );
AOI22xp33_ASAP7_75t_L g195 ( .A1(n_175), .A2(n_130), .B1(n_141), .B2(n_147), .Y(n_195) );
O2A1O1Ixp33_ASAP7_75t_L g196 ( .A1(n_151), .A2(n_135), .B(n_125), .C(n_140), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_154), .B(n_174), .Y(n_197) );
AOI22xp5_ASAP7_75t_L g198 ( .A1(n_152), .A2(n_130), .B1(n_147), .B2(n_124), .Y(n_198) );
AND2x2_ASAP7_75t_L g199 ( .A(n_169), .B(n_124), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_157), .Y(n_200) );
AOI22xp33_ASAP7_75t_L g201 ( .A1(n_175), .A2(n_140), .B1(n_136), .B2(n_135), .Y(n_201) );
NAND2x1_ASAP7_75t_L g202 ( .A(n_167), .B(n_99), .Y(n_202) );
INVx3_ASAP7_75t_L g203 ( .A(n_175), .Y(n_203) );
AND2x2_ASAP7_75t_L g204 ( .A(n_169), .B(n_125), .Y(n_204) );
A2O1A1Ixp33_ASAP7_75t_L g205 ( .A1(n_167), .A2(n_136), .B(n_112), .C(n_111), .Y(n_205) );
BUFx2_ASAP7_75t_L g206 ( .A(n_149), .Y(n_206) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_174), .B(n_123), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_163), .B(n_103), .Y(n_208) );
BUFx4f_ASAP7_75t_L g209 ( .A(n_171), .Y(n_209) );
AND2x4_ASAP7_75t_L g210 ( .A(n_174), .B(n_118), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_171), .B(n_116), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_161), .Y(n_212) );
HB1xp67_ASAP7_75t_L g213 ( .A(n_206), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_204), .B(n_170), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_178), .Y(n_215) );
O2A1O1Ixp33_ASAP7_75t_L g216 ( .A1(n_196), .A2(n_164), .B(n_172), .C(n_160), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g217 ( .A(n_186), .B(n_159), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_178), .Y(n_218) );
BUFx12f_ASAP7_75t_L g219 ( .A(n_206), .Y(n_219) );
INVx3_ASAP7_75t_L g220 ( .A(n_203), .Y(n_220) );
AND2x2_ASAP7_75t_L g221 ( .A(n_204), .B(n_152), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_182), .B(n_174), .Y(n_222) );
INVxp67_ASAP7_75t_L g223 ( .A(n_186), .Y(n_223) );
AND2x4_ASAP7_75t_L g224 ( .A(n_198), .B(n_174), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_182), .B(n_160), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_209), .B(n_94), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_201), .B(n_172), .Y(n_227) );
INVxp67_ASAP7_75t_L g228 ( .A(n_199), .Y(n_228) );
HB1xp67_ASAP7_75t_L g229 ( .A(n_210), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g230 ( .A(n_199), .B(n_158), .Y(n_230) );
OAI22xp5_ASAP7_75t_L g231 ( .A1(n_198), .A2(n_152), .B1(n_146), .B2(n_161), .Y(n_231) );
BUFx12f_ASAP7_75t_L g232 ( .A(n_210), .Y(n_232) );
OAI22x1_ASAP7_75t_L g233 ( .A1(n_210), .A2(n_152), .B1(n_89), .B2(n_112), .Y(n_233) );
INVx4_ASAP7_75t_L g234 ( .A(n_179), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_194), .A2(n_166), .B(n_155), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_184), .Y(n_236) );
OAI22x1_ASAP7_75t_L g237 ( .A1(n_210), .A2(n_152), .B1(n_90), .B2(n_122), .Y(n_237) );
BUFx2_ASAP7_75t_L g238 ( .A(n_209), .Y(n_238) );
AOI22xp5_ASAP7_75t_L g239 ( .A1(n_177), .A2(n_108), .B1(n_90), .B2(n_98), .Y(n_239) );
XNOR2xp5_ASAP7_75t_SL g240 ( .A(n_181), .B(n_8), .Y(n_240) );
AND2x2_ASAP7_75t_L g241 ( .A(n_177), .B(n_122), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_184), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_189), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_189), .Y(n_244) );
INVx3_ASAP7_75t_L g245 ( .A(n_203), .Y(n_245) );
AND2x4_ASAP7_75t_L g246 ( .A(n_203), .B(n_98), .Y(n_246) );
INVx1_ASAP7_75t_SL g247 ( .A(n_176), .Y(n_247) );
AND2x2_ASAP7_75t_L g248 ( .A(n_180), .B(n_100), .Y(n_248) );
INVx2_ASAP7_75t_SL g249 ( .A(n_232), .Y(n_249) );
AO21x2_ASAP7_75t_L g250 ( .A1(n_227), .A2(n_205), .B(n_166), .Y(n_250) );
OAI21x1_ASAP7_75t_L g251 ( .A1(n_235), .A2(n_202), .B(n_193), .Y(n_251) );
OAI21x1_ASAP7_75t_L g252 ( .A1(n_218), .A2(n_202), .B(n_193), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_218), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_218), .Y(n_254) );
INVx1_ASAP7_75t_SL g255 ( .A(n_219), .Y(n_255) );
OAI21xp5_ASAP7_75t_L g256 ( .A1(n_215), .A2(n_209), .B(n_180), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_244), .Y(n_257) );
OAI22xp5_ASAP7_75t_L g258 ( .A1(n_225), .A2(n_192), .B1(n_195), .B2(n_212), .Y(n_258) );
BUFx4f_ASAP7_75t_L g259 ( .A(n_232), .Y(n_259) );
OAI21xp5_ASAP7_75t_L g260 ( .A1(n_215), .A2(n_209), .B(n_200), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_244), .Y(n_261) );
OAI21x1_ASAP7_75t_L g262 ( .A1(n_244), .A2(n_193), .B(n_166), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_236), .Y(n_263) );
INVx2_ASAP7_75t_L g264 ( .A(n_236), .Y(n_264) );
OAI22xp5_ASAP7_75t_L g265 ( .A1(n_224), .A2(n_200), .B1(n_212), .B2(n_211), .Y(n_265) );
CKINVDCx16_ASAP7_75t_R g266 ( .A(n_219), .Y(n_266) );
INVxp67_ASAP7_75t_L g267 ( .A(n_213), .Y(n_267) );
OAI21xp5_ASAP7_75t_L g268 ( .A1(n_242), .A2(n_211), .B(n_187), .Y(n_268) );
BUFx2_ASAP7_75t_L g269 ( .A(n_232), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_242), .Y(n_270) );
OAI21xp5_ASAP7_75t_L g271 ( .A1(n_243), .A2(n_191), .B(n_185), .Y(n_271) );
A2O1A1Ixp33_ASAP7_75t_L g272 ( .A1(n_216), .A2(n_203), .B(n_183), .C(n_208), .Y(n_272) );
AND2x4_ASAP7_75t_L g273 ( .A(n_224), .B(n_179), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g274 ( .A(n_223), .B(n_190), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_243), .Y(n_275) );
HB1xp67_ASAP7_75t_L g276 ( .A(n_219), .Y(n_276) );
OAI21x1_ASAP7_75t_SL g277 ( .A1(n_234), .A2(n_188), .B(n_100), .Y(n_277) );
AND2x4_ASAP7_75t_L g278 ( .A(n_224), .B(n_188), .Y(n_278) );
A2O1A1Ixp33_ASAP7_75t_SL g279 ( .A1(n_274), .A2(n_217), .B(n_230), .C(n_228), .Y(n_279) );
OA21x2_ASAP7_75t_L g280 ( .A1(n_262), .A2(n_150), .B(n_155), .Y(n_280) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_272), .A2(n_222), .B(n_224), .Y(n_281) );
INVx3_ASAP7_75t_L g282 ( .A(n_253), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_261), .Y(n_283) );
AND2x2_ASAP7_75t_L g284 ( .A(n_253), .B(n_221), .Y(n_284) );
INVx3_ASAP7_75t_L g285 ( .A(n_253), .Y(n_285) );
AOI21xp5_ASAP7_75t_L g286 ( .A1(n_254), .A2(n_248), .B(n_241), .Y(n_286) );
INVx8_ASAP7_75t_L g287 ( .A(n_273), .Y(n_287) );
CKINVDCx5p33_ASAP7_75t_R g288 ( .A(n_266), .Y(n_288) );
AOI21xp5_ASAP7_75t_L g289 ( .A1(n_254), .A2(n_248), .B(n_241), .Y(n_289) );
CKINVDCx11_ASAP7_75t_R g290 ( .A(n_266), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_254), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_257), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_257), .Y(n_293) );
OAI221xp5_ASAP7_75t_L g294 ( .A1(n_267), .A2(n_231), .B1(n_214), .B2(n_239), .C(n_221), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_263), .B(n_239), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_261), .Y(n_296) );
OR2x2_ASAP7_75t_L g297 ( .A(n_257), .B(n_246), .Y(n_297) );
AOI22xp5_ASAP7_75t_L g298 ( .A1(n_265), .A2(n_237), .B1(n_233), .B2(n_240), .Y(n_298) );
AOI22xp33_ASAP7_75t_SL g299 ( .A1(n_265), .A2(n_240), .B1(n_238), .B2(n_246), .Y(n_299) );
OAI222xp33_ASAP7_75t_L g300 ( .A1(n_255), .A2(n_111), .B1(n_238), .B2(n_247), .C1(n_246), .C2(n_237), .Y(n_300) );
OR2x2_ASAP7_75t_L g301 ( .A(n_264), .B(n_246), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_263), .B(n_233), .Y(n_302) );
OR2x2_ASAP7_75t_L g303 ( .A(n_264), .B(n_247), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_264), .Y(n_304) );
AND2x2_ASAP7_75t_L g305 ( .A(n_304), .B(n_275), .Y(n_305) );
BUFx2_ASAP7_75t_L g306 ( .A(n_282), .Y(n_306) );
OR2x2_ASAP7_75t_L g307 ( .A(n_304), .B(n_275), .Y(n_307) );
INVx5_ASAP7_75t_L g308 ( .A(n_282), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_283), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_279), .B(n_267), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_299), .B(n_255), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_284), .B(n_275), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_283), .Y(n_313) );
BUFx2_ASAP7_75t_L g314 ( .A(n_282), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_296), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_296), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_291), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_284), .B(n_295), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_291), .Y(n_319) );
AND2x2_ASAP7_75t_L g320 ( .A(n_292), .B(n_270), .Y(n_320) );
AOI21xp5_ASAP7_75t_L g321 ( .A1(n_286), .A2(n_260), .B(n_277), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_292), .B(n_270), .Y(n_322) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_297), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_293), .Y(n_324) );
AO31x2_ASAP7_75t_L g325 ( .A1(n_281), .A2(n_258), .A3(n_155), .B(n_148), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_293), .Y(n_326) );
INVx4_ASAP7_75t_SL g327 ( .A(n_298), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_285), .Y(n_328) );
OR2x2_ASAP7_75t_L g329 ( .A(n_303), .B(n_276), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_309), .B(n_302), .Y(n_330) );
AOI22xp33_ASAP7_75t_L g331 ( .A1(n_327), .A2(n_298), .B1(n_294), .B2(n_287), .Y(n_331) );
OAI22xp33_ASAP7_75t_L g332 ( .A1(n_311), .A2(n_259), .B1(n_287), .B2(n_288), .Y(n_332) );
AND2x4_ASAP7_75t_SL g333 ( .A(n_305), .B(n_285), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_327), .B(n_285), .Y(n_334) );
AOI221xp5_ASAP7_75t_L g335 ( .A1(n_318), .A2(n_258), .B1(n_289), .B2(n_86), .C(n_300), .Y(n_335) );
INVxp67_ASAP7_75t_SL g336 ( .A(n_307), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_317), .Y(n_337) );
OR2x2_ASAP7_75t_L g338 ( .A(n_307), .B(n_303), .Y(n_338) );
AND2x2_ASAP7_75t_L g339 ( .A(n_327), .B(n_297), .Y(n_339) );
INVx2_ASAP7_75t_SL g340 ( .A(n_308), .Y(n_340) );
BUFx2_ASAP7_75t_L g341 ( .A(n_306), .Y(n_341) );
OR2x2_ASAP7_75t_L g342 ( .A(n_329), .B(n_301), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_317), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_327), .B(n_301), .Y(n_344) );
NAND2xp5_ASAP7_75t_SL g345 ( .A(n_308), .B(n_288), .Y(n_345) );
AOI31xp33_ASAP7_75t_L g346 ( .A1(n_323), .A2(n_276), .A3(n_249), .B(n_290), .Y(n_346) );
OR2x2_ASAP7_75t_L g347 ( .A(n_329), .B(n_287), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_305), .B(n_250), .Y(n_348) );
OR2x2_ASAP7_75t_L g349 ( .A(n_309), .B(n_287), .Y(n_349) );
INVx1_ASAP7_75t_SL g350 ( .A(n_306), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_313), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_312), .B(n_250), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_312), .B(n_250), .Y(n_353) );
INVx4_ASAP7_75t_L g354 ( .A(n_308), .Y(n_354) );
OR2x2_ASAP7_75t_L g355 ( .A(n_313), .B(n_250), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_324), .B(n_280), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_315), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_315), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_319), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_324), .B(n_280), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_352), .B(n_325), .Y(n_361) );
OR2x2_ASAP7_75t_L g362 ( .A(n_336), .B(n_326), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_337), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_352), .B(n_325), .Y(n_364) );
INVx6_ASAP7_75t_L g365 ( .A(n_354), .Y(n_365) );
INVx4_ASAP7_75t_L g366 ( .A(n_354), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_351), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_351), .Y(n_368) );
OAI33xp33_ASAP7_75t_L g369 ( .A1(n_357), .A2(n_310), .A3(n_316), .B1(n_107), .B2(n_326), .B3(n_14), .Y(n_369) );
OR2x6_ASAP7_75t_L g370 ( .A(n_354), .B(n_314), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_353), .B(n_325), .Y(n_371) );
NOR3xp33_ASAP7_75t_SL g372 ( .A(n_332), .B(n_113), .C(n_95), .Y(n_372) );
AOI21xp5_ASAP7_75t_L g373 ( .A1(n_335), .A2(n_321), .B(n_314), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_353), .B(n_325), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_357), .Y(n_375) );
OR2x2_ASAP7_75t_L g376 ( .A(n_336), .B(n_325), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_348), .B(n_316), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_338), .B(n_320), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_338), .B(n_320), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_348), .B(n_319), .Y(n_380) );
OR2x2_ASAP7_75t_L g381 ( .A(n_355), .B(n_322), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_358), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_358), .Y(n_383) );
AND2x4_ASAP7_75t_L g384 ( .A(n_334), .B(n_308), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_356), .B(n_328), .Y(n_385) );
INVx1_ASAP7_75t_SL g386 ( .A(n_333), .Y(n_386) );
OAI211xp5_ASAP7_75t_SL g387 ( .A1(n_331), .A2(n_107), .B(n_249), .C(n_226), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_342), .B(n_322), .Y(n_388) );
HB1xp67_ASAP7_75t_L g389 ( .A(n_341), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_356), .B(n_328), .Y(n_390) );
OR2x2_ASAP7_75t_L g391 ( .A(n_355), .B(n_86), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_342), .B(n_308), .Y(n_392) );
OR2x2_ASAP7_75t_L g393 ( .A(n_341), .B(n_86), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_360), .B(n_308), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_360), .B(n_337), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_337), .B(n_280), .Y(n_396) );
BUFx2_ASAP7_75t_L g397 ( .A(n_354), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_330), .B(n_86), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_343), .Y(n_399) );
OR2x2_ASAP7_75t_L g400 ( .A(n_350), .B(n_86), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_343), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_343), .B(n_280), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_359), .B(n_105), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_359), .B(n_105), .Y(n_404) );
NAND2xp5_ASAP7_75t_SL g405 ( .A(n_346), .B(n_259), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_368), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_368), .Y(n_407) );
OR2x2_ASAP7_75t_L g408 ( .A(n_391), .B(n_350), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_377), .B(n_330), .Y(n_409) );
NAND2x1_ASAP7_75t_L g410 ( .A(n_366), .B(n_346), .Y(n_410) );
INVx1_ASAP7_75t_SL g411 ( .A(n_365), .Y(n_411) );
AOI21xp5_ASAP7_75t_L g412 ( .A1(n_373), .A2(n_335), .B(n_340), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_361), .B(n_359), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_361), .B(n_334), .Y(n_414) );
INVxp33_ASAP7_75t_L g415 ( .A(n_397), .Y(n_415) );
OR2x2_ASAP7_75t_L g416 ( .A(n_391), .B(n_347), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_377), .B(n_333), .Y(n_417) );
OR2x2_ASAP7_75t_L g418 ( .A(n_381), .B(n_347), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_378), .B(n_333), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_364), .B(n_344), .Y(n_420) );
NAND2x1_ASAP7_75t_SL g421 ( .A(n_366), .B(n_344), .Y(n_421) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_400), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_375), .Y(n_423) );
NAND3xp33_ASAP7_75t_SL g424 ( .A(n_405), .B(n_345), .C(n_269), .Y(n_424) );
NAND2x1p5_ASAP7_75t_SL g425 ( .A(n_394), .B(n_340), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_379), .B(n_339), .Y(n_426) );
OR2x2_ASAP7_75t_L g427 ( .A(n_381), .B(n_349), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_375), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_382), .Y(n_429) );
OR2x2_ASAP7_75t_L g430 ( .A(n_362), .B(n_349), .Y(n_430) );
NOR2xp33_ASAP7_75t_L g431 ( .A(n_369), .B(n_339), .Y(n_431) );
OR2x2_ASAP7_75t_L g432 ( .A(n_362), .B(n_340), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_364), .B(n_88), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_382), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_388), .B(n_8), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_371), .B(n_153), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_367), .B(n_9), .Y(n_437) );
NOR3xp33_ASAP7_75t_SL g438 ( .A(n_387), .B(n_256), .C(n_260), .Y(n_438) );
INVx1_ASAP7_75t_SL g439 ( .A(n_365), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_371), .B(n_153), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_383), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_380), .B(n_9), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_383), .B(n_10), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_380), .B(n_13), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_393), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_393), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_398), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_363), .Y(n_448) );
XNOR2xp5_ASAP7_75t_L g449 ( .A(n_392), .B(n_269), .Y(n_449) );
INVx1_ASAP7_75t_SL g450 ( .A(n_365), .Y(n_450) );
NOR2xp33_ASAP7_75t_L g451 ( .A(n_389), .B(n_14), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_395), .B(n_15), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_374), .B(n_153), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_374), .B(n_153), .Y(n_454) );
OR2x2_ASAP7_75t_L g455 ( .A(n_395), .B(n_15), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_385), .B(n_153), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_403), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_385), .B(n_17), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_390), .B(n_18), .Y(n_459) );
OAI22xp33_ASAP7_75t_L g460 ( .A1(n_410), .A2(n_366), .B1(n_397), .B2(n_370), .Y(n_460) );
OAI21xp5_ASAP7_75t_L g461 ( .A1(n_424), .A2(n_372), .B(n_400), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_406), .Y(n_462) );
NAND3xp33_ASAP7_75t_L g463 ( .A(n_431), .B(n_404), .C(n_403), .Y(n_463) );
NAND3xp33_ASAP7_75t_SL g464 ( .A(n_412), .B(n_386), .C(n_404), .Y(n_464) );
AOI22xp5_ASAP7_75t_L g465 ( .A1(n_431), .A2(n_365), .B1(n_394), .B2(n_390), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_433), .B(n_376), .Y(n_466) );
OR2x2_ASAP7_75t_L g467 ( .A(n_427), .B(n_376), .Y(n_467) );
NAND2xp33_ASAP7_75t_L g468 ( .A(n_415), .B(n_384), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_433), .B(n_401), .Y(n_469) );
NAND3xp33_ASAP7_75t_L g470 ( .A(n_451), .B(n_370), .C(n_401), .Y(n_470) );
INVx1_ASAP7_75t_SL g471 ( .A(n_421), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_409), .B(n_363), .Y(n_472) );
OAI21xp33_ASAP7_75t_L g473 ( .A1(n_415), .A2(n_370), .B(n_399), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_407), .Y(n_474) );
NAND2x1_ASAP7_75t_L g475 ( .A(n_425), .B(n_370), .Y(n_475) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_435), .B(n_384), .Y(n_476) );
NAND2xp5_ASAP7_75t_SL g477 ( .A(n_411), .B(n_384), .Y(n_477) );
OAI221xp5_ASAP7_75t_L g478 ( .A1(n_451), .A2(n_249), .B1(n_399), .B2(n_259), .C(n_256), .Y(n_478) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_455), .B(n_18), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_423), .Y(n_480) );
NAND2xp5_ASAP7_75t_SL g481 ( .A(n_439), .B(n_402), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_428), .Y(n_482) );
HB1xp67_ASAP7_75t_L g483 ( .A(n_422), .Y(n_483) );
OAI22xp5_ASAP7_75t_L g484 ( .A1(n_449), .A2(n_402), .B1(n_396), .B2(n_259), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_422), .B(n_396), .Y(n_485) );
AOI22xp5_ASAP7_75t_L g486 ( .A1(n_445), .A2(n_278), .B1(n_273), .B2(n_268), .Y(n_486) );
OAI21xp33_ASAP7_75t_L g487 ( .A1(n_420), .A2(n_414), .B(n_413), .Y(n_487) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_450), .A2(n_277), .B(n_271), .Y(n_488) );
AOI22xp5_ASAP7_75t_L g489 ( .A1(n_446), .A2(n_278), .B1(n_273), .B2(n_268), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_429), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_413), .B(n_19), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_434), .B(n_19), .Y(n_492) );
OAI311xp33_ASAP7_75t_L g493 ( .A1(n_452), .A2(n_271), .A3(n_245), .B1(n_220), .C1(n_25), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_458), .B(n_278), .Y(n_494) );
OR2x2_ASAP7_75t_L g495 ( .A(n_430), .B(n_148), .Y(n_495) );
AND2x4_ASAP7_75t_L g496 ( .A(n_436), .B(n_278), .Y(n_496) );
AND2x4_ASAP7_75t_L g497 ( .A(n_436), .B(n_273), .Y(n_497) );
AOI22xp5_ASAP7_75t_L g498 ( .A1(n_442), .A2(n_252), .B1(n_251), .B2(n_165), .Y(n_498) );
AOI21xp33_ASAP7_75t_SL g499 ( .A1(n_425), .A2(n_20), .B(n_22), .Y(n_499) );
INVx1_ASAP7_75t_SL g500 ( .A(n_432), .Y(n_500) );
OAI22xp5_ASAP7_75t_L g501 ( .A1(n_418), .A2(n_229), .B1(n_220), .B2(n_245), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_441), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_448), .Y(n_503) );
OAI22xp33_ASAP7_75t_L g504 ( .A1(n_416), .A2(n_234), .B1(n_220), .B2(n_245), .Y(n_504) );
OAI221xp5_ASAP7_75t_L g505 ( .A1(n_459), .A2(n_148), .B1(n_150), .B2(n_165), .C(n_245), .Y(n_505) );
OAI32xp33_ASAP7_75t_L g506 ( .A1(n_417), .A2(n_176), .A3(n_150), .B1(n_234), .B2(n_197), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_426), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_483), .Y(n_508) );
OAI221xp5_ASAP7_75t_L g509 ( .A1(n_465), .A2(n_437), .B1(n_443), .B2(n_419), .C(n_447), .Y(n_509) );
INVx1_ASAP7_75t_SL g510 ( .A(n_500), .Y(n_510) );
NAND3xp33_ASAP7_75t_L g511 ( .A(n_463), .B(n_454), .C(n_453), .Y(n_511) );
XNOR2x1_ASAP7_75t_L g512 ( .A(n_484), .B(n_444), .Y(n_512) );
AOI211xp5_ASAP7_75t_L g513 ( .A1(n_460), .A2(n_420), .B(n_414), .C(n_408), .Y(n_513) );
INVxp67_ASAP7_75t_L g514 ( .A(n_464), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_503), .Y(n_515) );
INVx1_ASAP7_75t_SL g516 ( .A(n_471), .Y(n_516) );
AOI21xp33_ASAP7_75t_L g517 ( .A1(n_470), .A2(n_454), .B(n_453), .Y(n_517) );
OAI21xp5_ASAP7_75t_L g518 ( .A1(n_470), .A2(n_438), .B(n_440), .Y(n_518) );
AOI22xp5_ASAP7_75t_L g519 ( .A1(n_476), .A2(n_440), .B1(n_457), .B2(n_456), .Y(n_519) );
INVxp67_ASAP7_75t_L g520 ( .A(n_491), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_462), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_507), .B(n_456), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_474), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_473), .B(n_448), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_487), .B(n_438), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_480), .Y(n_526) );
NOR3x1_ASAP7_75t_L g527 ( .A(n_475), .B(n_251), .C(n_252), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_481), .Y(n_528) );
AOI22xp5_ASAP7_75t_L g529 ( .A1(n_479), .A2(n_251), .B1(n_252), .B2(n_165), .Y(n_529) );
XNOR2xp5_ASAP7_75t_L g530 ( .A(n_467), .B(n_23), .Y(n_530) );
OAI21xp5_ASAP7_75t_SL g531 ( .A1(n_461), .A2(n_165), .B(n_207), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_482), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_490), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_485), .B(n_165), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_478), .B(n_26), .Y(n_535) );
O2A1O1Ixp33_ASAP7_75t_L g536 ( .A1(n_493), .A2(n_220), .B(n_31), .C(n_32), .Y(n_536) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_499), .B(n_165), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_472), .B(n_262), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_502), .Y(n_539) );
OAI22xp5_ASAP7_75t_L g540 ( .A1(n_513), .A2(n_477), .B1(n_466), .B2(n_469), .Y(n_540) );
INVx2_ASAP7_75t_SL g541 ( .A(n_510), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_508), .Y(n_542) );
AOI322xp5_ASAP7_75t_L g543 ( .A1(n_514), .A2(n_468), .A3(n_492), .B1(n_494), .B2(n_497), .C1(n_496), .C2(n_486), .Y(n_543) );
OAI22xp5_ASAP7_75t_L g544 ( .A1(n_514), .A2(n_498), .B1(n_496), .B2(n_497), .Y(n_544) );
NOR2xp33_ASAP7_75t_L g545 ( .A(n_516), .B(n_495), .Y(n_545) );
INVx1_ASAP7_75t_SL g546 ( .A(n_530), .Y(n_546) );
OAI21xp5_ASAP7_75t_L g547 ( .A1(n_536), .A2(n_488), .B(n_505), .Y(n_547) );
AOI21xp5_ASAP7_75t_L g548 ( .A1(n_537), .A2(n_506), .B(n_504), .Y(n_548) );
OAI21xp33_ASAP7_75t_L g549 ( .A1(n_525), .A2(n_489), .B(n_501), .Y(n_549) );
AOI21xp33_ASAP7_75t_SL g550 ( .A1(n_512), .A2(n_28), .B(n_37), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_522), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_528), .B(n_38), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_521), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_523), .Y(n_554) );
NAND3xp33_ASAP7_75t_L g555 ( .A(n_531), .B(n_234), .C(n_191), .Y(n_555) );
NOR3x1_ASAP7_75t_L g556 ( .A(n_518), .B(n_262), .C(n_42), .Y(n_556) );
AOI21xp5_ASAP7_75t_L g557 ( .A1(n_536), .A2(n_191), .B(n_187), .Y(n_557) );
OAI21xp33_ASAP7_75t_SL g558 ( .A1(n_517), .A2(n_40), .B(n_48), .Y(n_558) );
OAI211xp5_ASAP7_75t_L g559 ( .A1(n_558), .A2(n_520), .B(n_511), .C(n_509), .Y(n_559) );
OAI21xp5_ASAP7_75t_L g560 ( .A1(n_543), .A2(n_520), .B(n_535), .Y(n_560) );
OAI211xp5_ASAP7_75t_SL g561 ( .A1(n_549), .A2(n_529), .B(n_519), .C(n_535), .Y(n_561) );
NOR3xp33_ASAP7_75t_L g562 ( .A(n_547), .B(n_534), .C(n_524), .Y(n_562) );
INVxp67_ASAP7_75t_L g563 ( .A(n_541), .Y(n_563) );
A2O1A1Ixp33_ASAP7_75t_L g564 ( .A1(n_550), .A2(n_539), .B(n_533), .C(n_532), .Y(n_564) );
AOI21xp5_ASAP7_75t_L g565 ( .A1(n_540), .A2(n_557), .B(n_548), .Y(n_565) );
NOR3xp33_ASAP7_75t_L g566 ( .A(n_544), .B(n_526), .C(n_538), .Y(n_566) );
OAI211xp5_ASAP7_75t_SL g567 ( .A1(n_546), .A2(n_515), .B(n_527), .C(n_52), .Y(n_567) );
OA211x2_ASAP7_75t_L g568 ( .A1(n_545), .A2(n_49), .B(n_50), .C(n_56), .Y(n_568) );
NOR3xp33_ASAP7_75t_L g569 ( .A(n_557), .B(n_185), .C(n_187), .Y(n_569) );
NOR2x1_ASAP7_75t_L g570 ( .A(n_565), .B(n_555), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_563), .B(n_551), .Y(n_571) );
NOR2xp67_ASAP7_75t_L g572 ( .A(n_559), .B(n_542), .Y(n_572) );
NOR4xp75_ASAP7_75t_SL g573 ( .A(n_560), .B(n_556), .C(n_548), .D(n_553), .Y(n_573) );
NOR3xp33_ASAP7_75t_L g574 ( .A(n_567), .B(n_552), .C(n_554), .Y(n_574) );
AOI211xp5_ASAP7_75t_L g575 ( .A1(n_561), .A2(n_58), .B(n_60), .C(n_61), .Y(n_575) );
AND3x4_ASAP7_75t_L g576 ( .A(n_570), .B(n_566), .C(n_562), .Y(n_576) );
AND2x2_ASAP7_75t_SL g577 ( .A(n_574), .B(n_569), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_572), .A2(n_568), .B1(n_564), .B2(n_185), .Y(n_578) );
INVx2_ASAP7_75t_L g579 ( .A(n_576), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_577), .B(n_571), .Y(n_580) );
AOI22x1_ASAP7_75t_L g581 ( .A1(n_579), .A2(n_573), .B1(n_578), .B2(n_575), .Y(n_581) );
NOR3xp33_ASAP7_75t_L g582 ( .A(n_580), .B(n_65), .C(n_68), .Y(n_582) );
AOI22xp5_ASAP7_75t_L g583 ( .A1(n_582), .A2(n_69), .B1(n_71), .B2(n_72), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_583), .A2(n_581), .B1(n_74), .B2(n_75), .Y(n_584) );
AOI22x1_ASAP7_75t_L g585 ( .A1(n_584), .A2(n_73), .B1(n_77), .B2(n_78), .Y(n_585) );
AOI21xp5_ASAP7_75t_L g586 ( .A1(n_585), .A2(n_79), .B(n_80), .Y(n_586) );
endmodule