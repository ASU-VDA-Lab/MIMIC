module fake_netlist_6_4274_n_2408 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_235, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_223, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_226, n_228, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_227, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_233, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_234, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_236, n_38, n_110, n_151, n_61, n_112, n_172, n_237, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_231, n_65, n_230, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_229, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_232, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_2408);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_235;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_223;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_226;
input n_228;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_227;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_233;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_234;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_236;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_237;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_231;
input n_65;
input n_230;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_229;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_232;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_2408;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_2332;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_1854;
wire n_2324;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_2405;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_2179;
wire n_2386;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_2382;
wire n_2291;
wire n_415;
wire n_830;
wire n_2299;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_1590;
wire n_1532;
wire n_2313;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_2365;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_522;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2094;
wire n_2018;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_2212;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_2256;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_405;
wire n_538;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_2394;
wire n_2108;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_381;
wire n_2378;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_2155;
wire n_1445;
wire n_2364;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_2370;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_2214;
wire n_913;
wire n_407;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_2300;
wire n_564;
wire n_2397;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_577;
wire n_1843;
wire n_619;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_2093;
wire n_483;
wire n_2207;
wire n_1970;
wire n_608;
wire n_261;
wire n_2101;
wire n_630;
wire n_2059;
wire n_2198;
wire n_541;
wire n_512;
wire n_2073;
wire n_2273;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_2355;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2245;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_2192;
wire n_2254;
wire n_2345;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2350;
wire n_286;
wire n_254;
wire n_2193;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_850;
wire n_690;
wire n_1886;
wire n_1801;
wire n_2092;
wire n_2347;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2206;
wire n_604;
wire n_2319;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_2377;
wire n_701;
wire n_295;
wire n_2178;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_1825;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_2194;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_2279;
wire n_1052;
wire n_462;
wire n_1033;
wire n_1296;
wire n_1990;
wire n_2391;
wire n_304;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_595;
wire n_627;
wire n_297;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2349;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_2230;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_963;
wire n_320;
wire n_639;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_851;
wire n_682;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_2316;
wire n_631;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_2407;
wire n_1277;
wire n_797;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_2307;
wire n_2362;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_2231;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_2251;
wire n_1384;
wire n_2238;
wire n_293;
wire n_2368;
wire n_1070;
wire n_458;
wire n_2403;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_2338;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_2354;
wire n_1395;
wire n_2199;
wire n_2110;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_1021;
wire n_931;
wire n_527;
wire n_474;
wire n_811;
wire n_683;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_2294;
wire n_1363;
wire n_1334;
wire n_1966;
wire n_1942;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_399;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1736;
wire n_1564;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2330;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_1141;
wire n_562;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_556;
wire n_2209;
wire n_2301;
wire n_2387;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_2357;
wire n_1125;
wire n_970;
wire n_2224;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_441;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_2115;
wire n_1053;
wire n_2374;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_2384;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_2204;
wire n_1520;
wire n_496;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2289;
wire n_1077;
wire n_1733;
wire n_2315;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_2276;
wire n_663;
wire n_856;
wire n_2100;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_2379;
wire n_435;
wire n_1905;
wire n_2016;
wire n_2343;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_2219;
wire n_1203;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_952;
wire n_725;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_732;
wire n_974;
wire n_2240;
wire n_392;
wire n_2278;
wire n_724;
wire n_2375;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2381;
wire n_1847;
wire n_2052;
wire n_248;
wire n_2302;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_2177;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_2337;
wire n_2401;
wire n_1356;
wire n_1589;
wire n_2309;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_2264;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_2220;
wire n_1262;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_239;
wire n_2037;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_2169;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_2244;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2200;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_2376;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_2346;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_1524;
wire n_543;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_2406;
wire n_533;
wire n_2390;
wire n_806;
wire n_879;
wire n_959;
wire n_2310;
wire n_584;
wire n_2141;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_2383;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2196;
wire n_273;
wire n_1633;
wire n_2195;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_550;
wire n_2322;
wire n_275;
wire n_652;
wire n_2154;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_2283;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_2361;
wire n_306;
wire n_1292;
wire n_1373;
wire n_2266;
wire n_346;
wire n_1029;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_2189;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2348;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_2366;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_2400;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_1074;
wire n_698;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_246;
wire n_1338;
wire n_1097;
wire n_2395;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_2380;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_2295;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_2020;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_2048;
wire n_300;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_2175;
wire n_601;
wire n_2182;
wire n_338;
wire n_1283;
wire n_2385;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1848;
wire n_763;
wire n_1147;
wire n_1785;
wire n_360;
wire n_1754;
wire n_2149;
wire n_2396;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2284;
wire n_387;
wire n_2287;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2081;
wire n_2168;
wire n_2022;
wire n_2203;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_472;
wire n_270;
wire n_2265;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_2267;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_854;
wire n_1058;
wire n_2312;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_390;
wire n_1148;
wire n_2188;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_2318;
wire n_1149;
wire n_265;
wire n_1184;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_859;
wire n_570;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_985;
wire n_2233;
wire n_481;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2360;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_436;
wire n_2334;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_2303;
wire n_1619;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_2367;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_973;
wire n_359;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2217;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_2215;
wire n_404;
wire n_271;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_588;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2223;
wire n_2091;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_2116;
wire n_336;
wire n_2320;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_53),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_160),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_35),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_207),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_20),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_20),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_15),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_152),
.Y(n_245)
);

INVx2_ASAP7_75t_SL g246 ( 
.A(n_201),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_216),
.Y(n_247)
);

BUFx5_ASAP7_75t_L g248 ( 
.A(n_74),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_204),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_107),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_89),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_199),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_42),
.Y(n_253)
);

INVx2_ASAP7_75t_SL g254 ( 
.A(n_145),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_33),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_5),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_86),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_69),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_136),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_158),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_105),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_54),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_237),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_156),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_134),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_223),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_162),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_13),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_132),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_92),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_49),
.Y(n_271)
);

BUFx3_ASAP7_75t_L g272 ( 
.A(n_141),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_53),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_173),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_55),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_22),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_159),
.Y(n_277)
);

BUFx2_ASAP7_75t_L g278 ( 
.A(n_46),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_78),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_22),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_52),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_17),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_83),
.Y(n_283)
);

INVx2_ASAP7_75t_SL g284 ( 
.A(n_234),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_210),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_17),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_174),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_24),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_38),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_79),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_4),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_56),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_144),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_90),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_33),
.Y(n_295)
);

CKINVDCx14_ASAP7_75t_R g296 ( 
.A(n_124),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_198),
.Y(n_297)
);

BUFx5_ASAP7_75t_L g298 ( 
.A(n_4),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_61),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_24),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_93),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_167),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_236),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_25),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_35),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_78),
.Y(n_306)
);

BUFx3_ASAP7_75t_L g307 ( 
.A(n_73),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_83),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_79),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_157),
.Y(n_310)
);

BUFx10_ASAP7_75t_L g311 ( 
.A(n_56),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_50),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_125),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_222),
.Y(n_314)
);

BUFx10_ASAP7_75t_L g315 ( 
.A(n_138),
.Y(n_315)
);

BUFx10_ASAP7_75t_L g316 ( 
.A(n_225),
.Y(n_316)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_85),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_166),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_58),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_30),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_171),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_193),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_101),
.Y(n_323)
);

BUFx2_ASAP7_75t_L g324 ( 
.A(n_179),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_70),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_154),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_96),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_66),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_123),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_137),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_172),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_98),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_71),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_175),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_34),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_72),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_191),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_14),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_215),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_19),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_235),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_110),
.Y(n_342)
);

INVx1_ASAP7_75t_SL g343 ( 
.A(n_0),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_133),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_211),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_30),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_66),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_185),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_6),
.Y(n_349)
);

INVx1_ASAP7_75t_SL g350 ( 
.A(n_214),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_41),
.Y(n_351)
);

BUFx2_ASAP7_75t_L g352 ( 
.A(n_106),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_95),
.Y(n_353)
);

BUFx3_ASAP7_75t_L g354 ( 
.A(n_109),
.Y(n_354)
);

INVx2_ASAP7_75t_SL g355 ( 
.A(n_40),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_97),
.Y(n_356)
);

BUFx10_ASAP7_75t_L g357 ( 
.A(n_87),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_59),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_92),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_227),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_41),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_25),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_102),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_205),
.Y(n_364)
);

BUFx2_ASAP7_75t_L g365 ( 
.A(n_170),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_44),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_183),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_5),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_232),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_189),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_190),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_65),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_163),
.Y(n_373)
);

CKINVDCx14_ASAP7_75t_R g374 ( 
.A(n_203),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_202),
.Y(n_375)
);

INVx1_ASAP7_75t_SL g376 ( 
.A(n_31),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_87),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_187),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_9),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_27),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_72),
.Y(n_381)
);

BUFx3_ASAP7_75t_L g382 ( 
.A(n_32),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_64),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_139),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_47),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_176),
.Y(n_386)
);

INVx1_ASAP7_75t_SL g387 ( 
.A(n_192),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_12),
.Y(n_388)
);

CKINVDCx16_ASAP7_75t_R g389 ( 
.A(n_181),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_67),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_45),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_90),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_231),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_217),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_117),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_149),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_142),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_93),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_81),
.Y(n_399)
);

INVx1_ASAP7_75t_SL g400 ( 
.A(n_70),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_102),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_2),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_208),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_37),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_130),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_91),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_42),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_31),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_28),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_120),
.Y(n_410)
);

INVx1_ASAP7_75t_SL g411 ( 
.A(n_151),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_165),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_122),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_10),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_177),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_127),
.Y(n_416)
);

INVx2_ASAP7_75t_SL g417 ( 
.A(n_48),
.Y(n_417)
);

CKINVDCx16_ASAP7_75t_R g418 ( 
.A(n_80),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_61),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_63),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_91),
.Y(n_421)
);

BUFx10_ASAP7_75t_L g422 ( 
.A(n_221),
.Y(n_422)
);

CKINVDCx16_ASAP7_75t_R g423 ( 
.A(n_180),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_150),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_114),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_64),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_1),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_219),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_135),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_28),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_101),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_43),
.Y(n_432)
);

INVx1_ASAP7_75t_SL g433 ( 
.A(n_197),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_196),
.Y(n_434)
);

CKINVDCx14_ASAP7_75t_R g435 ( 
.A(n_51),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_81),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_129),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_100),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_86),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_213),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_103),
.Y(n_441)
);

INVx1_ASAP7_75t_SL g442 ( 
.A(n_98),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_40),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_108),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_34),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_12),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_113),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_54),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_186),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_2),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_8),
.Y(n_451)
);

BUFx10_ASAP7_75t_L g452 ( 
.A(n_218),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_96),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_209),
.Y(n_454)
);

BUFx3_ASAP7_75t_L g455 ( 
.A(n_228),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_131),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_229),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_46),
.Y(n_458)
);

INVxp67_ASAP7_75t_L g459 ( 
.A(n_111),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_164),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_188),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_0),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_32),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_65),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_39),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_248),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_239),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_248),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_248),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_247),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_248),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_249),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_250),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_248),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_248),
.Y(n_475)
);

INVxp33_ASAP7_75t_SL g476 ( 
.A(n_278),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_261),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_248),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_248),
.Y(n_479)
);

INVxp67_ASAP7_75t_L g480 ( 
.A(n_278),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_264),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_324),
.B(n_1),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_248),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_298),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_252),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_259),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_260),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_263),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_265),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_318),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_267),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_269),
.Y(n_492)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_338),
.Y(n_493)
);

INVxp67_ASAP7_75t_SL g494 ( 
.A(n_324),
.Y(n_494)
);

INVxp67_ASAP7_75t_SL g495 ( 
.A(n_352),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_298),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_298),
.Y(n_497)
);

HB1xp67_ASAP7_75t_L g498 ( 
.A(n_255),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_274),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_344),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_285),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_287),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_410),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_298),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_352),
.B(n_3),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_298),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_298),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_425),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_298),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_298),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_444),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_298),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_338),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_454),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_338),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_389),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_338),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_338),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_338),
.Y(n_519)
);

INVxp67_ASAP7_75t_SL g520 ( 
.A(n_365),
.Y(n_520)
);

BUFx6f_ASAP7_75t_SL g521 ( 
.A(n_315),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_349),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_349),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_293),
.Y(n_524)
);

CKINVDCx16_ASAP7_75t_R g525 ( 
.A(n_435),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_349),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_349),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_303),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_349),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_325),
.Y(n_530)
);

CKINVDCx16_ASAP7_75t_R g531 ( 
.A(n_255),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_310),
.Y(n_532)
);

INVxp33_ASAP7_75t_SL g533 ( 
.A(n_238),
.Y(n_533)
);

HB1xp67_ASAP7_75t_L g534 ( 
.A(n_312),
.Y(n_534)
);

CKINVDCx20_ASAP7_75t_R g535 ( 
.A(n_389),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_325),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_423),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g538 ( 
.A(n_423),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_296),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g540 ( 
.A(n_374),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_313),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_365),
.B(n_3),
.Y(n_542)
);

INVxp67_ASAP7_75t_L g543 ( 
.A(n_251),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_321),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_322),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_329),
.Y(n_546)
);

BUFx2_ASAP7_75t_SL g547 ( 
.A(n_246),
.Y(n_547)
);

CKINVDCx20_ASAP7_75t_R g548 ( 
.A(n_331),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_334),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_380),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_380),
.Y(n_551)
);

INVxp67_ASAP7_75t_SL g552 ( 
.A(n_272),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g553 ( 
.A(n_337),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_246),
.B(n_6),
.Y(n_554)
);

CKINVDCx20_ASAP7_75t_R g555 ( 
.A(n_339),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_341),
.Y(n_556)
);

CKINVDCx20_ASAP7_75t_R g557 ( 
.A(n_342),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_383),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_383),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_345),
.Y(n_560)
);

CKINVDCx20_ASAP7_75t_R g561 ( 
.A(n_348),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_398),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_398),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_427),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_254),
.B(n_7),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_427),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_360),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_443),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_443),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_462),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_254),
.B(n_7),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_462),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_364),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_367),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g575 ( 
.A(n_369),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_251),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_253),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_371),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_375),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_378),
.Y(n_580)
);

INVxp33_ASAP7_75t_SL g581 ( 
.A(n_240),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_384),
.Y(n_582)
);

CKINVDCx20_ASAP7_75t_R g583 ( 
.A(n_386),
.Y(n_583)
);

INVxp67_ASAP7_75t_L g584 ( 
.A(n_253),
.Y(n_584)
);

INVxp67_ASAP7_75t_L g585 ( 
.A(n_257),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_257),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_258),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_258),
.Y(n_588)
);

CKINVDCx20_ASAP7_75t_R g589 ( 
.A(n_393),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_395),
.Y(n_590)
);

AND2x2_ASAP7_75t_L g591 ( 
.A(n_307),
.B(n_8),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_266),
.Y(n_592)
);

NOR2xp67_ASAP7_75t_L g593 ( 
.A(n_414),
.B(n_9),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_515),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_466),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_515),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_591),
.B(n_552),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_466),
.Y(n_598)
);

NAND2xp33_ASAP7_75t_SL g599 ( 
.A(n_542),
.B(n_355),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_468),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_565),
.B(n_284),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_571),
.B(n_284),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_517),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_517),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_547),
.B(n_312),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_518),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_518),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_493),
.Y(n_608)
);

INVxp67_ASAP7_75t_L g609 ( 
.A(n_498),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_522),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_468),
.Y(n_611)
);

OAI21x1_ASAP7_75t_L g612 ( 
.A1(n_469),
.A2(n_456),
.B(n_245),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_469),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_522),
.Y(n_614)
);

BUFx2_ASAP7_75t_L g615 ( 
.A(n_516),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_523),
.Y(n_616)
);

OAI22xp5_ASAP7_75t_SL g617 ( 
.A1(n_476),
.A2(n_275),
.B1(n_340),
.B2(n_262),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_523),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_526),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_526),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_591),
.B(n_272),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_527),
.B(n_397),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_471),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_471),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_474),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_527),
.B(n_403),
.Y(n_626)
);

AND2x4_ASAP7_75t_L g627 ( 
.A(n_493),
.B(n_354),
.Y(n_627)
);

BUFx3_ASAP7_75t_L g628 ( 
.A(n_493),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_513),
.Y(n_629)
);

OAI22xp5_ASAP7_75t_L g630 ( 
.A1(n_480),
.A2(n_418),
.B1(n_421),
.B2(n_358),
.Y(n_630)
);

INVxp67_ASAP7_75t_L g631 ( 
.A(n_534),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_547),
.B(n_418),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_592),
.B(n_354),
.Y(n_633)
);

BUFx6f_ASAP7_75t_L g634 ( 
.A(n_474),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_554),
.B(n_459),
.Y(n_635)
);

BUFx6f_ASAP7_75t_L g636 ( 
.A(n_475),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_475),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_513),
.Y(n_638)
);

INVx3_ASAP7_75t_L g639 ( 
.A(n_519),
.Y(n_639)
);

HB1xp67_ASAP7_75t_L g640 ( 
.A(n_593),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_519),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_478),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_478),
.Y(n_643)
);

AOI22xp5_ASAP7_75t_L g644 ( 
.A1(n_482),
.A2(n_432),
.B1(n_450),
.B2(n_431),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_529),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_529),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_592),
.B(n_455),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_530),
.B(n_455),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_479),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_525),
.B(n_315),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_479),
.Y(n_651)
);

BUFx6f_ASAP7_75t_L g652 ( 
.A(n_483),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_483),
.Y(n_653)
);

HB1xp67_ASAP7_75t_L g654 ( 
.A(n_543),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_484),
.Y(n_655)
);

INVx3_ASAP7_75t_L g656 ( 
.A(n_484),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_530),
.Y(n_657)
);

INVx4_ASAP7_75t_L g658 ( 
.A(n_568),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_496),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_568),
.Y(n_660)
);

BUFx8_ASAP7_75t_L g661 ( 
.A(n_521),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_496),
.Y(n_662)
);

HB1xp67_ASAP7_75t_L g663 ( 
.A(n_584),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_576),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_497),
.Y(n_665)
);

BUFx6f_ASAP7_75t_L g666 ( 
.A(n_497),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_576),
.Y(n_667)
);

BUFx6f_ASAP7_75t_L g668 ( 
.A(n_504),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_504),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_506),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_506),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_507),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_507),
.Y(n_673)
);

BUFx2_ASAP7_75t_L g674 ( 
.A(n_535),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_548),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_509),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_509),
.Y(n_677)
);

OA22x2_ASAP7_75t_SL g678 ( 
.A1(n_494),
.A2(n_270),
.B1(n_271),
.B2(n_268),
.Y(n_678)
);

INVx3_ASAP7_75t_L g679 ( 
.A(n_510),
.Y(n_679)
);

AND2x4_ASAP7_75t_L g680 ( 
.A(n_510),
.B(n_245),
.Y(n_680)
);

BUFx12f_ASAP7_75t_L g681 ( 
.A(n_467),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_512),
.Y(n_682)
);

BUFx6f_ASAP7_75t_L g683 ( 
.A(n_512),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_536),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_536),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_550),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_550),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_551),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_495),
.B(n_307),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_551),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_558),
.Y(n_691)
);

AOI22xp5_ASAP7_75t_L g692 ( 
.A1(n_635),
.A2(n_505),
.B1(n_520),
.B2(n_317),
.Y(n_692)
);

NAND2xp33_ASAP7_75t_L g693 ( 
.A(n_601),
.B(n_602),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_597),
.B(n_470),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_595),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_595),
.Y(n_696)
);

INVx2_ASAP7_75t_SL g697 ( 
.A(n_597),
.Y(n_697)
);

BUFx10_ASAP7_75t_L g698 ( 
.A(n_605),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_670),
.Y(n_699)
);

INVx3_ASAP7_75t_L g700 ( 
.A(n_600),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_601),
.B(n_533),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_605),
.B(n_525),
.Y(n_702)
);

INVx2_ASAP7_75t_SL g703 ( 
.A(n_597),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_595),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_602),
.B(n_581),
.Y(n_705)
);

OR2x2_ASAP7_75t_L g706 ( 
.A(n_609),
.B(n_531),
.Y(n_706)
);

INVx4_ASAP7_75t_SL g707 ( 
.A(n_600),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_670),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_595),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_635),
.B(n_622),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_632),
.B(n_472),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_670),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_632),
.B(n_473),
.Y(n_713)
);

BUFx4f_ASAP7_75t_L g714 ( 
.A(n_600),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_673),
.Y(n_715)
);

BUFx2_ASAP7_75t_L g716 ( 
.A(n_609),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_621),
.B(n_558),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_650),
.B(n_485),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_673),
.Y(n_719)
);

BUFx6f_ASAP7_75t_L g720 ( 
.A(n_628),
.Y(n_720)
);

INVx3_ASAP7_75t_L g721 ( 
.A(n_600),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_598),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_673),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_598),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_598),
.Y(n_725)
);

INVx3_ASAP7_75t_L g726 ( 
.A(n_600),
.Y(n_726)
);

BUFx3_ASAP7_75t_L g727 ( 
.A(n_628),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_676),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_661),
.B(n_486),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_621),
.B(n_559),
.Y(n_730)
);

OR2x2_ASAP7_75t_L g731 ( 
.A(n_631),
.B(n_487),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_598),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_622),
.B(n_488),
.Y(n_733)
);

INVx2_ASAP7_75t_SL g734 ( 
.A(n_621),
.Y(n_734)
);

AOI21x1_ASAP7_75t_L g735 ( 
.A1(n_680),
.A2(n_277),
.B(n_266),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_676),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_611),
.Y(n_737)
);

INVx2_ASAP7_75t_SL g738 ( 
.A(n_689),
.Y(n_738)
);

AO22x2_ASAP7_75t_L g739 ( 
.A1(n_630),
.A2(n_417),
.B1(n_355),
.B2(n_270),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_611),
.Y(n_740)
);

CKINVDCx20_ASAP7_75t_R g741 ( 
.A(n_675),
.Y(n_741)
);

OR2x6_ASAP7_75t_L g742 ( 
.A(n_681),
.B(n_277),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_611),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_676),
.Y(n_744)
);

AOI22xp33_ASAP7_75t_L g745 ( 
.A1(n_599),
.A2(n_417),
.B1(n_382),
.B2(n_268),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_656),
.Y(n_746)
);

INVx4_ASAP7_75t_L g747 ( 
.A(n_600),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_611),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_613),
.Y(n_749)
);

AOI22xp33_ASAP7_75t_L g750 ( 
.A1(n_599),
.A2(n_382),
.B1(n_271),
.B2(n_288),
.Y(n_750)
);

NAND3xp33_ASAP7_75t_L g751 ( 
.A(n_680),
.B(n_585),
.C(n_302),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_661),
.B(n_489),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_661),
.B(n_491),
.Y(n_753)
);

BUFx3_ASAP7_75t_L g754 ( 
.A(n_628),
.Y(n_754)
);

INVx2_ASAP7_75t_SL g755 ( 
.A(n_689),
.Y(n_755)
);

INVx1_ASAP7_75t_SL g756 ( 
.A(n_675),
.Y(n_756)
);

INVx3_ASAP7_75t_L g757 ( 
.A(n_600),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_656),
.Y(n_758)
);

AND2x6_ASAP7_75t_L g759 ( 
.A(n_680),
.B(n_396),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_613),
.Y(n_760)
);

INVx4_ASAP7_75t_L g761 ( 
.A(n_600),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_661),
.B(n_492),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_681),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_613),
.Y(n_764)
);

XNOR2xp5_ASAP7_75t_L g765 ( 
.A(n_617),
.B(n_477),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_661),
.B(n_499),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_613),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_623),
.Y(n_768)
);

CKINVDCx20_ASAP7_75t_R g769 ( 
.A(n_681),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_661),
.B(n_501),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_656),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_623),
.Y(n_772)
);

OAI22xp33_ASAP7_75t_L g773 ( 
.A1(n_650),
.A2(n_343),
.B1(n_376),
.B2(n_281),
.Y(n_773)
);

INVx3_ASAP7_75t_L g774 ( 
.A(n_634),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_656),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_631),
.B(n_502),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_626),
.B(n_524),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_626),
.B(n_528),
.Y(n_778)
);

AOI22xp33_ASAP7_75t_L g779 ( 
.A1(n_689),
.A2(n_280),
.B1(n_300),
.B2(n_288),
.Y(n_779)
);

INVx3_ASAP7_75t_L g780 ( 
.A(n_634),
.Y(n_780)
);

INVx3_ASAP7_75t_L g781 ( 
.A(n_634),
.Y(n_781)
);

INVx3_ASAP7_75t_L g782 ( 
.A(n_634),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_640),
.B(n_532),
.Y(n_783)
);

BUFx6f_ASAP7_75t_L g784 ( 
.A(n_628),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_627),
.B(n_541),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_623),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_656),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_679),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_640),
.B(n_544),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_623),
.Y(n_790)
);

BUFx4f_ASAP7_75t_L g791 ( 
.A(n_634),
.Y(n_791)
);

BUFx6f_ASAP7_75t_L g792 ( 
.A(n_634),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_679),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_679),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_654),
.B(n_545),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_SL g796 ( 
.A(n_681),
.B(n_537),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_627),
.B(n_679),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_679),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_627),
.B(n_546),
.Y(n_799)
);

AOI22xp33_ASAP7_75t_L g800 ( 
.A1(n_680),
.A2(n_280),
.B1(n_323),
.B2(n_300),
.Y(n_800)
);

INVx3_ASAP7_75t_L g801 ( 
.A(n_634),
.Y(n_801)
);

INVx4_ASAP7_75t_L g802 ( 
.A(n_634),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_624),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_627),
.B(n_556),
.Y(n_804)
);

CKINVDCx16_ASAP7_75t_R g805 ( 
.A(n_615),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_L g806 ( 
.A(n_654),
.B(n_560),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_615),
.Y(n_807)
);

OR2x6_ASAP7_75t_L g808 ( 
.A(n_627),
.B(n_297),
.Y(n_808)
);

OR2x6_ASAP7_75t_L g809 ( 
.A(n_627),
.B(n_297),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_633),
.B(n_567),
.Y(n_810)
);

AND2x2_ASAP7_75t_L g811 ( 
.A(n_648),
.B(n_559),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_663),
.B(n_573),
.Y(n_812)
);

BUFx3_ASAP7_75t_L g813 ( 
.A(n_648),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_624),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_624),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_624),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_625),
.Y(n_817)
);

OR2x2_ASAP7_75t_L g818 ( 
.A(n_663),
.B(n_574),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_625),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_625),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_625),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_637),
.Y(n_822)
);

NAND3xp33_ASAP7_75t_L g823 ( 
.A(n_680),
.B(n_314),
.C(n_302),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_633),
.B(n_578),
.Y(n_824)
);

INVx4_ASAP7_75t_L g825 ( 
.A(n_636),
.Y(n_825)
);

NAND2xp33_ASAP7_75t_L g826 ( 
.A(n_633),
.B(n_579),
.Y(n_826)
);

AOI22xp33_ASAP7_75t_L g827 ( 
.A1(n_680),
.A2(n_647),
.B1(n_648),
.B2(n_658),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_664),
.B(n_580),
.Y(n_828)
);

OR2x2_ASAP7_75t_L g829 ( 
.A(n_630),
.B(n_582),
.Y(n_829)
);

OR2x2_ASAP7_75t_L g830 ( 
.A(n_644),
.B(n_590),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_637),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_637),
.Y(n_832)
);

AOI22xp33_ASAP7_75t_L g833 ( 
.A1(n_647),
.A2(n_327),
.B1(n_328),
.B2(n_323),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_637),
.Y(n_834)
);

AND2x4_ASAP7_75t_L g835 ( 
.A(n_647),
.B(n_314),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_644),
.B(n_539),
.Y(n_836)
);

INVx4_ASAP7_75t_L g837 ( 
.A(n_636),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_643),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_643),
.Y(n_839)
);

INVx3_ASAP7_75t_L g840 ( 
.A(n_636),
.Y(n_840)
);

OAI22xp33_ASAP7_75t_L g841 ( 
.A1(n_664),
.A2(n_442),
.B1(n_400),
.B2(n_242),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_643),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_643),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_649),
.Y(n_844)
);

CKINVDCx12_ASAP7_75t_R g845 ( 
.A(n_617),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_649),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_649),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_649),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_651),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_651),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_658),
.B(n_350),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_651),
.Y(n_852)
);

AND3x2_ASAP7_75t_L g853 ( 
.A(n_615),
.B(n_456),
.C(n_330),
.Y(n_853)
);

INVx2_ASAP7_75t_SL g854 ( 
.A(n_813),
.Y(n_854)
);

AOI22xp5_ASAP7_75t_L g855 ( 
.A1(n_701),
.A2(n_549),
.B1(n_555),
.B2(n_553),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_710),
.B(n_636),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_813),
.B(n_636),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_813),
.B(n_636),
.Y(n_858)
);

INVx2_ASAP7_75t_SL g859 ( 
.A(n_717),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_705),
.B(n_557),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_711),
.B(n_561),
.Y(n_861)
);

HB1xp67_ASAP7_75t_L g862 ( 
.A(n_738),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_693),
.B(n_636),
.Y(n_863)
);

AOI22x1_ASAP7_75t_SL g864 ( 
.A1(n_769),
.A2(n_538),
.B1(n_490),
.B2(n_500),
.Y(n_864)
);

OAI221xp5_ASAP7_75t_L g865 ( 
.A1(n_779),
.A2(n_678),
.B1(n_697),
.B2(n_703),
.C(n_800),
.Y(n_865)
);

INVx1_ASAP7_75t_SL g866 ( 
.A(n_716),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_827),
.B(n_636),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_734),
.B(n_642),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_L g869 ( 
.A(n_713),
.B(n_575),
.Y(n_869)
);

INVxp67_ASAP7_75t_SL g870 ( 
.A(n_792),
.Y(n_870)
);

A2O1A1Ixp33_ASAP7_75t_L g871 ( 
.A1(n_697),
.A2(n_612),
.B(n_327),
.C(n_333),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_699),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_703),
.B(n_642),
.Y(n_873)
);

BUFx6f_ASAP7_75t_L g874 ( 
.A(n_720),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_734),
.B(n_642),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_733),
.B(n_642),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_738),
.B(n_642),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_783),
.B(n_806),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_699),
.Y(n_879)
);

INVx8_ASAP7_75t_L g880 ( 
.A(n_808),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_777),
.B(n_583),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_811),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_708),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_708),
.Y(n_884)
);

AOI22xp5_ASAP7_75t_L g885 ( 
.A1(n_755),
.A2(n_589),
.B1(n_503),
.B2(n_508),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_L g886 ( 
.A(n_778),
.B(n_540),
.Y(n_886)
);

NAND2xp33_ASAP7_75t_L g887 ( 
.A(n_797),
.B(n_396),
.Y(n_887)
);

AOI22xp33_ASAP7_75t_L g888 ( 
.A1(n_755),
.A2(n_653),
.B1(n_655),
.B2(n_651),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_712),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_694),
.B(n_828),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_712),
.B(n_642),
.Y(n_891)
);

INVx8_ASAP7_75t_L g892 ( 
.A(n_808),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_SL g893 ( 
.A(n_718),
.B(n_642),
.Y(n_893)
);

INVxp67_ASAP7_75t_L g894 ( 
.A(n_716),
.Y(n_894)
);

AOI22xp5_ASAP7_75t_L g895 ( 
.A1(n_826),
.A2(n_511),
.B1(n_514),
.B2(n_481),
.Y(n_895)
);

INVx2_ASAP7_75t_SL g896 ( 
.A(n_811),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_776),
.B(n_674),
.Y(n_897)
);

BUFx6f_ASAP7_75t_L g898 ( 
.A(n_720),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_717),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_810),
.B(n_674),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_730),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_715),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_730),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_715),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_773),
.B(n_642),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_719),
.Y(n_906)
);

O2A1O1Ixp5_ASAP7_75t_L g907 ( 
.A1(n_719),
.A2(n_655),
.B(n_659),
.C(n_653),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_723),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_L g909 ( 
.A(n_824),
.B(n_674),
.Y(n_909)
);

INVx3_ASAP7_75t_L g910 ( 
.A(n_727),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_818),
.B(n_667),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_698),
.B(n_652),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_723),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_728),
.B(n_652),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_SL g915 ( 
.A(n_698),
.B(n_652),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_728),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_736),
.B(n_652),
.Y(n_917)
);

AOI22xp5_ASAP7_75t_L g918 ( 
.A1(n_702),
.A2(n_799),
.B1(n_804),
.B2(n_785),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_736),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_744),
.B(n_652),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_744),
.Y(n_921)
);

BUFx6f_ASAP7_75t_L g922 ( 
.A(n_720),
.Y(n_922)
);

AND2x4_ASAP7_75t_SL g923 ( 
.A(n_742),
.B(n_315),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_SL g924 ( 
.A(n_698),
.B(n_720),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_746),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_818),
.B(n_521),
.Y(n_926)
);

INVx2_ASAP7_75t_SL g927 ( 
.A(n_853),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_763),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_SL g929 ( 
.A(n_698),
.B(n_652),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_741),
.Y(n_930)
);

NAND2xp33_ASAP7_75t_L g931 ( 
.A(n_759),
.B(n_396),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_SL g932 ( 
.A(n_720),
.B(n_652),
.Y(n_932)
);

OAI22xp5_ASAP7_75t_L g933 ( 
.A1(n_692),
.A2(n_326),
.B1(n_370),
.B2(n_330),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_731),
.B(n_521),
.Y(n_934)
);

BUFx6f_ASAP7_75t_SL g935 ( 
.A(n_742),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_746),
.Y(n_936)
);

OR2x2_ASAP7_75t_L g937 ( 
.A(n_706),
.B(n_667),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_722),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_722),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_851),
.B(n_652),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_758),
.B(n_662),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_758),
.Y(n_942)
);

BUFx3_ASAP7_75t_L g943 ( 
.A(n_727),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_771),
.B(n_662),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_771),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_775),
.B(n_662),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_SL g947 ( 
.A(n_720),
.B(n_662),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_722),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_775),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_787),
.B(n_662),
.Y(n_950)
);

OR2x2_ASAP7_75t_L g951 ( 
.A(n_706),
.B(n_577),
.Y(n_951)
);

INVx1_ASAP7_75t_SL g952 ( 
.A(n_756),
.Y(n_952)
);

BUFx6f_ASAP7_75t_L g953 ( 
.A(n_784),
.Y(n_953)
);

AOI22xp33_ASAP7_75t_L g954 ( 
.A1(n_835),
.A2(n_655),
.B1(n_659),
.B2(n_653),
.Y(n_954)
);

INVx8_ASAP7_75t_L g955 ( 
.A(n_808),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_784),
.B(n_787),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_740),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_740),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_788),
.B(n_662),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_784),
.B(n_662),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_788),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_740),
.Y(n_962)
);

AND2x2_ASAP7_75t_L g963 ( 
.A(n_731),
.B(n_311),
.Y(n_963)
);

AOI22xp5_ASAP7_75t_L g964 ( 
.A1(n_835),
.A2(n_411),
.B1(n_433),
.B2(n_387),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_793),
.B(n_662),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_743),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_793),
.Y(n_967)
);

NAND2xp33_ASAP7_75t_L g968 ( 
.A(n_759),
.B(n_396),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_L g969 ( 
.A(n_795),
.B(n_243),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_743),
.Y(n_970)
);

AOI22xp33_ASAP7_75t_L g971 ( 
.A1(n_835),
.A2(n_655),
.B1(n_659),
.B2(n_653),
.Y(n_971)
);

OAI22xp5_ASAP7_75t_L g972 ( 
.A1(n_692),
.A2(n_326),
.B1(n_373),
.B2(n_370),
.Y(n_972)
);

BUFx3_ASAP7_75t_L g973 ( 
.A(n_727),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_794),
.B(n_798),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_SL g975 ( 
.A(n_784),
.B(n_666),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_743),
.Y(n_976)
);

INVxp67_ASAP7_75t_L g977 ( 
.A(n_812),
.Y(n_977)
);

AOI22xp5_ASAP7_75t_L g978 ( 
.A1(n_835),
.A2(n_809),
.B1(n_808),
.B2(n_752),
.Y(n_978)
);

AOI22xp5_ASAP7_75t_L g979 ( 
.A1(n_808),
.A2(n_412),
.B1(n_413),
.B2(n_405),
.Y(n_979)
);

NOR3xp33_ASAP7_75t_L g980 ( 
.A(n_836),
.B(n_256),
.C(n_244),
.Y(n_980)
);

NAND2xp33_ASAP7_75t_L g981 ( 
.A(n_759),
.B(n_396),
.Y(n_981)
);

NOR3xp33_ASAP7_75t_L g982 ( 
.A(n_805),
.B(n_276),
.C(n_273),
.Y(n_982)
);

BUFx3_ASAP7_75t_L g983 ( 
.A(n_754),
.Y(n_983)
);

INVx2_ASAP7_75t_SL g984 ( 
.A(n_789),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_SL g985 ( 
.A(n_784),
.B(n_666),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_794),
.B(n_666),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_798),
.B(n_754),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_754),
.Y(n_988)
);

NAND2xp33_ASAP7_75t_L g989 ( 
.A(n_759),
.B(n_396),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_700),
.B(n_666),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_SL g991 ( 
.A(n_784),
.B(n_666),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_700),
.B(n_666),
.Y(n_992)
);

INVxp67_ASAP7_75t_L g993 ( 
.A(n_829),
.Y(n_993)
);

NOR2xp67_ASAP7_75t_L g994 ( 
.A(n_729),
.B(n_658),
.Y(n_994)
);

AOI22xp5_ASAP7_75t_L g995 ( 
.A1(n_809),
.A2(n_428),
.B1(n_429),
.B2(n_416),
.Y(n_995)
);

NOR2xp33_ASAP7_75t_L g996 ( 
.A(n_829),
.B(n_279),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_748),
.Y(n_997)
);

INVxp67_ASAP7_75t_L g998 ( 
.A(n_830),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_814),
.Y(n_999)
);

AOI22xp5_ASAP7_75t_L g1000 ( 
.A1(n_809),
.A2(n_437),
.B1(n_461),
.B2(n_434),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_L g1001 ( 
.A(n_830),
.B(n_282),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_792),
.B(n_666),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_700),
.B(n_721),
.Y(n_1003)
);

BUFx8_ASAP7_75t_L g1004 ( 
.A(n_805),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_814),
.Y(n_1005)
);

INVx2_ASAP7_75t_SL g1006 ( 
.A(n_809),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_SL g1007 ( 
.A(n_792),
.B(n_666),
.Y(n_1007)
);

AOI22xp33_ASAP7_75t_SL g1008 ( 
.A1(n_796),
.A2(n_316),
.B1(n_422),
.B2(n_315),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_748),
.Y(n_1009)
);

BUFx6f_ASAP7_75t_L g1010 ( 
.A(n_792),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_748),
.Y(n_1011)
);

NOR2xp33_ASAP7_75t_L g1012 ( 
.A(n_753),
.B(n_283),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_700),
.B(n_721),
.Y(n_1013)
);

AOI22xp5_ASAP7_75t_L g1014 ( 
.A1(n_809),
.A2(n_394),
.B1(n_415),
.B2(n_373),
.Y(n_1014)
);

BUFx3_ASAP7_75t_L g1015 ( 
.A(n_742),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_721),
.B(n_668),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_721),
.B(n_668),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_749),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_749),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_726),
.B(n_668),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_749),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_726),
.B(n_668),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_760),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_820),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_760),
.Y(n_1025)
);

NAND3xp33_ASAP7_75t_L g1026 ( 
.A(n_745),
.B(n_289),
.C(n_286),
.Y(n_1026)
);

A2O1A1Ixp33_ASAP7_75t_L g1027 ( 
.A1(n_751),
.A2(n_612),
.B(n_333),
.C(n_336),
.Y(n_1027)
);

OAI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_867),
.A2(n_791),
.B(n_714),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_890),
.B(n_726),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_SL g1030 ( 
.A(n_928),
.B(n_807),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_878),
.B(n_726),
.Y(n_1031)
);

AND2x2_ASAP7_75t_L g1032 ( 
.A(n_911),
.B(n_739),
.Y(n_1032)
);

INVx3_ASAP7_75t_L g1033 ( 
.A(n_943),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_893),
.A2(n_791),
.B(n_714),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_854),
.B(n_757),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_893),
.A2(n_791),
.B(n_714),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_854),
.B(n_757),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_876),
.A2(n_761),
.B(n_747),
.Y(n_1038)
);

OAI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_856),
.A2(n_822),
.B(n_820),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_SL g1040 ( 
.A(n_918),
.B(n_757),
.Y(n_1040)
);

NOR2xp67_ASAP7_75t_L g1041 ( 
.A(n_885),
.B(n_762),
.Y(n_1041)
);

AND2x2_ASAP7_75t_L g1042 ( 
.A(n_866),
.B(n_739),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_940),
.A2(n_761),
.B(n_747),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_872),
.Y(n_1044)
);

A2O1A1Ixp33_ASAP7_75t_L g1045 ( 
.A1(n_996),
.A2(n_751),
.B(n_770),
.C(n_766),
.Y(n_1045)
);

O2A1O1Ixp33_ASAP7_75t_L g1046 ( 
.A1(n_933),
.A2(n_841),
.B(n_823),
.C(n_831),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_896),
.B(n_757),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_879),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_857),
.A2(n_761),
.B(n_747),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_SL g1050 ( 
.A(n_928),
.B(n_742),
.Y(n_1050)
);

NOR2x1p5_ASAP7_75t_SL g1051 ( 
.A(n_938),
.B(n_939),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_879),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_963),
.B(n_739),
.Y(n_1053)
);

OAI22xp5_ASAP7_75t_L g1054 ( 
.A1(n_978),
.A2(n_742),
.B1(n_833),
.B2(n_823),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_858),
.A2(n_761),
.B(n_747),
.Y(n_1055)
);

BUFx6f_ASAP7_75t_L g1056 ( 
.A(n_1010),
.Y(n_1056)
);

AND2x4_ASAP7_75t_L g1057 ( 
.A(n_859),
.B(n_750),
.Y(n_1057)
);

O2A1O1Ixp33_ASAP7_75t_SL g1058 ( 
.A1(n_871),
.A2(n_1027),
.B(n_905),
.C(n_972),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_896),
.B(n_774),
.Y(n_1059)
);

OR2x2_ASAP7_75t_L g1060 ( 
.A(n_952),
.B(n_765),
.Y(n_1060)
);

OAI21xp33_ASAP7_75t_L g1061 ( 
.A1(n_1001),
.A2(n_739),
.B(n_291),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_862),
.B(n_774),
.Y(n_1062)
);

AND2x2_ASAP7_75t_L g1063 ( 
.A(n_897),
.B(n_765),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_904),
.B(n_774),
.Y(n_1064)
);

AOI21x1_ASAP7_75t_L g1065 ( 
.A1(n_912),
.A2(n_831),
.B(n_822),
.Y(n_1065)
);

AND2x2_ASAP7_75t_SL g1066 ( 
.A(n_923),
.B(n_394),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_870),
.A2(n_825),
.B(n_802),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_863),
.A2(n_825),
.B(n_802),
.Y(n_1068)
);

AOI22xp33_ASAP7_75t_L g1069 ( 
.A1(n_899),
.A2(n_328),
.B1(n_346),
.B2(n_336),
.Y(n_1069)
);

BUFx6f_ASAP7_75t_L g1070 ( 
.A(n_1010),
.Y(n_1070)
);

AOI22xp5_ASAP7_75t_L g1071 ( 
.A1(n_881),
.A2(n_759),
.B1(n_780),
.B2(n_774),
.Y(n_1071)
);

NOR2xp33_ASAP7_75t_SL g1072 ( 
.A(n_860),
.B(n_316),
.Y(n_1072)
);

AND2x2_ASAP7_75t_L g1073 ( 
.A(n_900),
.B(n_311),
.Y(n_1073)
);

O2A1O1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_865),
.A2(n_834),
.B(n_838),
.C(n_832),
.Y(n_1074)
);

A2O1A1Ixp33_ASAP7_75t_L g1075 ( 
.A1(n_1012),
.A2(n_424),
.B(n_440),
.C(n_415),
.Y(n_1075)
);

NOR3xp33_ASAP7_75t_L g1076 ( 
.A(n_861),
.B(n_440),
.C(n_424),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_SL g1077 ( 
.A(n_883),
.B(n_780),
.Y(n_1077)
);

INVx2_ASAP7_75t_SL g1078 ( 
.A(n_937),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_L g1079 ( 
.A(n_993),
.B(n_845),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_916),
.B(n_919),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_868),
.A2(n_825),
.B(n_802),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_921),
.B(n_780),
.Y(n_1082)
);

BUFx6f_ASAP7_75t_L g1083 ( 
.A(n_1010),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_882),
.B(n_901),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_875),
.A2(n_825),
.B(n_802),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_910),
.A2(n_837),
.B(n_792),
.Y(n_1086)
);

OR2x6_ASAP7_75t_L g1087 ( 
.A(n_880),
.B(n_441),
.Y(n_1087)
);

O2A1O1Ixp33_ASAP7_75t_L g1088 ( 
.A1(n_905),
.A2(n_834),
.B(n_838),
.C(n_832),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_910),
.A2(n_837),
.B(n_792),
.Y(n_1089)
);

NOR2xp33_ASAP7_75t_SL g1090 ( 
.A(n_869),
.B(n_316),
.Y(n_1090)
);

A2O1A1Ixp33_ASAP7_75t_L g1091 ( 
.A1(n_903),
.A2(n_612),
.B(n_353),
.C(n_362),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_883),
.B(n_780),
.Y(n_1092)
);

O2A1O1Ixp33_ASAP7_75t_L g1093 ( 
.A1(n_1027),
.A2(n_843),
.B(n_847),
.C(n_839),
.Y(n_1093)
);

INVx4_ASAP7_75t_L g1094 ( 
.A(n_943),
.Y(n_1094)
);

OAI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_1006),
.A2(n_441),
.B1(n_449),
.B2(n_447),
.Y(n_1095)
);

AND2x2_ASAP7_75t_L g1096 ( 
.A(n_909),
.B(n_311),
.Y(n_1096)
);

OAI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_907),
.A2(n_843),
.B(n_839),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_884),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_910),
.A2(n_837),
.B(n_782),
.Y(n_1099)
);

OAI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_873),
.A2(n_848),
.B(n_847),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_884),
.B(n_781),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_889),
.B(n_781),
.Y(n_1102)
);

NOR2xp67_ASAP7_75t_L g1103 ( 
.A(n_977),
.B(n_735),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_SL g1104 ( 
.A(n_930),
.B(n_316),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_930),
.Y(n_1105)
);

OR2x2_ASAP7_75t_L g1106 ( 
.A(n_951),
.B(n_577),
.Y(n_1106)
);

OAI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_873),
.A2(n_849),
.B(n_848),
.Y(n_1107)
);

BUFx6f_ASAP7_75t_L g1108 ( 
.A(n_1010),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_987),
.A2(n_837),
.B(n_782),
.Y(n_1109)
);

AND2x4_ASAP7_75t_L g1110 ( 
.A(n_973),
.B(n_586),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_1003),
.A2(n_782),
.B(n_781),
.Y(n_1111)
);

OAI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_974),
.A2(n_849),
.B(n_852),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_889),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_1013),
.A2(n_782),
.B(n_781),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_877),
.A2(n_840),
.B(n_801),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_902),
.Y(n_1116)
);

OAI22x1_ASAP7_75t_L g1117 ( 
.A1(n_855),
.A2(n_845),
.B1(n_678),
.B2(n_292),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_SL g1118 ( 
.A(n_902),
.B(n_801),
.Y(n_1118)
);

A2O1A1Ixp33_ASAP7_75t_L g1119 ( 
.A1(n_969),
.A2(n_353),
.B(n_362),
.C(n_346),
.Y(n_1119)
);

A2O1A1Ixp33_ASAP7_75t_L g1120 ( 
.A1(n_886),
.A2(n_449),
.B(n_457),
.C(n_447),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_877),
.A2(n_840),
.B(n_801),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_SL g1122 ( 
.A(n_906),
.B(n_801),
.Y(n_1122)
);

NOR2xp33_ASAP7_75t_L g1123 ( 
.A(n_998),
.B(n_840),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_906),
.B(n_840),
.Y(n_1124)
);

CKINVDCx8_ASAP7_75t_R g1125 ( 
.A(n_880),
.Y(n_1125)
);

OAI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_891),
.A2(n_696),
.B(n_695),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_912),
.A2(n_696),
.B(n_695),
.Y(n_1127)
);

AND2x4_ASAP7_75t_L g1128 ( 
.A(n_973),
.B(n_586),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_915),
.A2(n_709),
.B(n_704),
.Y(n_1129)
);

BUFx2_ASAP7_75t_SL g1130 ( 
.A(n_935),
.Y(n_1130)
);

INVx3_ASAP7_75t_L g1131 ( 
.A(n_983),
.Y(n_1131)
);

OAI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_914),
.A2(n_852),
.B(n_709),
.Y(n_1132)
);

BUFx4f_ASAP7_75t_L g1133 ( 
.A(n_984),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_915),
.A2(n_724),
.B(n_704),
.Y(n_1134)
);

INVx5_ASAP7_75t_L g1135 ( 
.A(n_874),
.Y(n_1135)
);

A2O1A1Ixp33_ASAP7_75t_L g1136 ( 
.A1(n_964),
.A2(n_460),
.B(n_457),
.C(n_724),
.Y(n_1136)
);

INVx3_ASAP7_75t_L g1137 ( 
.A(n_983),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_908),
.Y(n_1138)
);

NOR2xp33_ASAP7_75t_R g1139 ( 
.A(n_1004),
.B(n_735),
.Y(n_1139)
);

NOR2x1p5_ASAP7_75t_SL g1140 ( 
.A(n_938),
.B(n_760),
.Y(n_1140)
);

NOR2xp33_ASAP7_75t_L g1141 ( 
.A(n_894),
.B(n_725),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_908),
.B(n_725),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_929),
.A2(n_737),
.B(n_732),
.Y(n_1143)
);

OAI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_917),
.A2(n_850),
.B(n_737),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_913),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_913),
.B(n_732),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_929),
.A2(n_768),
.B(n_767),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_925),
.B(n_850),
.Y(n_1148)
);

BUFx8_ASAP7_75t_L g1149 ( 
.A(n_935),
.Y(n_1149)
);

OAI22xp5_ASAP7_75t_L g1150 ( 
.A1(n_1006),
.A2(n_460),
.B1(n_768),
.B2(n_767),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_956),
.A2(n_786),
.B(n_772),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_SL g1152 ( 
.A(n_994),
.B(n_707),
.Y(n_1152)
);

AOI21xp33_ASAP7_75t_L g1153 ( 
.A1(n_934),
.A2(n_294),
.B(n_290),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_SL g1154 ( 
.A(n_954),
.B(n_707),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_956),
.A2(n_786),
.B(n_772),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_936),
.Y(n_1156)
);

OAI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_920),
.A2(n_846),
.B(n_815),
.Y(n_1157)
);

OAI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_871),
.A2(n_846),
.B(n_815),
.Y(n_1158)
);

OAI21x1_ASAP7_75t_L g1159 ( 
.A1(n_990),
.A2(n_1016),
.B(n_992),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_1017),
.A2(n_816),
.B(n_803),
.Y(n_1160)
);

BUFx4f_ASAP7_75t_L g1161 ( 
.A(n_927),
.Y(n_1161)
);

INVx3_ASAP7_75t_L g1162 ( 
.A(n_874),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1020),
.A2(n_816),
.B(n_803),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_942),
.B(n_844),
.Y(n_1164)
);

INVx3_ASAP7_75t_L g1165 ( 
.A(n_874),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1022),
.A2(n_819),
.B(n_817),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_932),
.A2(n_819),
.B(n_817),
.Y(n_1167)
);

NOR2xp33_ASAP7_75t_L g1168 ( 
.A(n_895),
.B(n_842),
.Y(n_1168)
);

OAI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_945),
.A2(n_844),
.B(n_842),
.Y(n_1169)
);

AOI21x1_ASAP7_75t_L g1170 ( 
.A1(n_932),
.A2(n_790),
.B(n_764),
.Y(n_1170)
);

OAI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_949),
.A2(n_790),
.B(n_764),
.Y(n_1171)
);

INVx3_ASAP7_75t_L g1172 ( 
.A(n_874),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_961),
.B(n_764),
.Y(n_1173)
);

O2A1O1Ixp33_ASAP7_75t_L g1174 ( 
.A1(n_967),
.A2(n_1005),
.B(n_1024),
.C(n_999),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_939),
.Y(n_1175)
);

O2A1O1Ixp33_ASAP7_75t_L g1176 ( 
.A1(n_924),
.A2(n_821),
.B(n_790),
.C(n_665),
.Y(n_1176)
);

NOR2xp33_ASAP7_75t_L g1177 ( 
.A(n_926),
.B(n_821),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_948),
.Y(n_1178)
);

AND2x2_ASAP7_75t_L g1179 ( 
.A(n_980),
.B(n_311),
.Y(n_1179)
);

O2A1O1Ixp5_ASAP7_75t_L g1180 ( 
.A1(n_924),
.A2(n_821),
.B(n_646),
.C(n_645),
.Y(n_1180)
);

AOI21xp33_ASAP7_75t_L g1181 ( 
.A1(n_1008),
.A2(n_299),
.B(n_295),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_988),
.B(n_659),
.Y(n_1182)
);

NOR2xp67_ASAP7_75t_L g1183 ( 
.A(n_1026),
.B(n_587),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_888),
.B(n_665),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_948),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_947),
.A2(n_669),
.B(n_665),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_SL g1187 ( 
.A(n_971),
.B(n_707),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_957),
.B(n_665),
.Y(n_1188)
);

INVxp67_ASAP7_75t_SL g1189 ( 
.A(n_898),
.Y(n_1189)
);

NAND2xp33_ASAP7_75t_SL g1190 ( 
.A(n_935),
.B(n_377),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_SL g1191 ( 
.A(n_898),
.B(n_707),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_SL g1192 ( 
.A(n_898),
.B(n_707),
.Y(n_1192)
);

INVx2_ASAP7_75t_L g1193 ( 
.A(n_958),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_947),
.A2(n_975),
.B(n_960),
.Y(n_1194)
);

OAI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_941),
.A2(n_671),
.B(n_669),
.Y(n_1195)
);

AOI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_880),
.A2(n_759),
.B1(n_669),
.B2(n_671),
.Y(n_1196)
);

INVx1_ASAP7_75t_SL g1197 ( 
.A(n_864),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_958),
.B(n_669),
.Y(n_1198)
);

AO21x1_ASAP7_75t_L g1199 ( 
.A1(n_887),
.A2(n_379),
.B(n_377),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_960),
.A2(n_672),
.B(n_671),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_SL g1201 ( 
.A(n_922),
.B(n_668),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_962),
.B(n_671),
.Y(n_1202)
);

INVxp67_ASAP7_75t_SL g1203 ( 
.A(n_922),
.Y(n_1203)
);

NAND3xp33_ASAP7_75t_L g1204 ( 
.A(n_982),
.B(n_304),
.C(n_301),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_966),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_975),
.A2(n_677),
.B(n_672),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_966),
.B(n_672),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_985),
.A2(n_677),
.B(n_672),
.Y(n_1208)
);

AOI21x1_ASAP7_75t_L g1209 ( 
.A1(n_985),
.A2(n_682),
.B(n_677),
.Y(n_1209)
);

OAI22xp5_ASAP7_75t_L g1210 ( 
.A1(n_1015),
.A2(n_241),
.B1(n_610),
.B2(n_614),
.Y(n_1210)
);

INVx1_ASAP7_75t_SL g1211 ( 
.A(n_923),
.Y(n_1211)
);

A2O1A1Ixp33_ASAP7_75t_L g1212 ( 
.A1(n_1014),
.A2(n_448),
.B(n_391),
.C(n_399),
.Y(n_1212)
);

NAND2xp33_ASAP7_75t_L g1213 ( 
.A(n_880),
.B(n_241),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_970),
.B(n_677),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_970),
.B(n_682),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_976),
.Y(n_1216)
);

AOI22xp5_ASAP7_75t_L g1217 ( 
.A1(n_892),
.A2(n_682),
.B1(n_658),
.B2(n_608),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_991),
.A2(n_682),
.B(n_668),
.Y(n_1218)
);

BUFx6f_ASAP7_75t_L g1219 ( 
.A(n_1056),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_1185),
.Y(n_1220)
);

A2O1A1Ixp33_ASAP7_75t_L g1221 ( 
.A1(n_1045),
.A2(n_1168),
.B(n_1076),
.C(n_1061),
.Y(n_1221)
);

O2A1O1Ixp33_ASAP7_75t_L g1222 ( 
.A1(n_1076),
.A2(n_887),
.B(n_1015),
.C(n_379),
.Y(n_1222)
);

OAI22xp5_ASAP7_75t_L g1223 ( 
.A1(n_1069),
.A2(n_955),
.B1(n_892),
.B2(n_979),
.Y(n_1223)
);

O2A1O1Ixp33_ASAP7_75t_L g1224 ( 
.A1(n_1120),
.A2(n_391),
.B(n_407),
.C(n_399),
.Y(n_1224)
);

OAI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1074),
.A2(n_946),
.B(n_944),
.Y(n_1225)
);

INVxp67_ASAP7_75t_L g1226 ( 
.A(n_1078),
.Y(n_1226)
);

BUFx8_ASAP7_75t_L g1227 ( 
.A(n_1042),
.Y(n_1227)
);

AO22x1_ASAP7_75t_L g1228 ( 
.A1(n_1063),
.A2(n_1004),
.B1(n_305),
.B2(n_308),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1135),
.A2(n_953),
.B(n_922),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1141),
.B(n_892),
.Y(n_1230)
);

AND2x2_ASAP7_75t_L g1231 ( 
.A(n_1073),
.B(n_1096),
.Y(n_1231)
);

OAI22xp5_ASAP7_75t_L g1232 ( 
.A1(n_1069),
.A2(n_955),
.B1(n_892),
.B2(n_995),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1135),
.A2(n_953),
.B(n_991),
.Y(n_1233)
);

A2O1A1Ixp33_ASAP7_75t_L g1234 ( 
.A1(n_1168),
.A2(n_1000),
.B(n_955),
.C(n_959),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1141),
.B(n_955),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1031),
.B(n_976),
.Y(n_1236)
);

O2A1O1Ixp33_ASAP7_75t_L g1237 ( 
.A1(n_1119),
.A2(n_407),
.B(n_426),
.C(n_430),
.Y(n_1237)
);

O2A1O1Ixp33_ASAP7_75t_L g1238 ( 
.A1(n_1119),
.A2(n_438),
.B(n_464),
.C(n_453),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1213),
.A2(n_1007),
.B(n_1002),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1044),
.Y(n_1240)
);

NAND2xp33_ASAP7_75t_SL g1241 ( 
.A(n_1053),
.B(n_1004),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1057),
.B(n_997),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_1105),
.Y(n_1243)
);

OAI22xp5_ASAP7_75t_SL g1244 ( 
.A1(n_1060),
.A2(n_351),
.B1(n_306),
.B2(n_309),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1067),
.A2(n_1007),
.B(n_968),
.Y(n_1245)
);

NOR3xp33_ASAP7_75t_SL g1246 ( 
.A(n_1079),
.B(n_320),
.C(n_319),
.Y(n_1246)
);

OAI22x1_ASAP7_75t_L g1247 ( 
.A1(n_1079),
.A2(n_332),
.B1(n_335),
.B2(n_347),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1052),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_SL g1249 ( 
.A(n_1041),
.B(n_997),
.Y(n_1249)
);

A2O1A1Ixp33_ASAP7_75t_L g1250 ( 
.A1(n_1046),
.A2(n_965),
.B(n_986),
.C(n_950),
.Y(n_1250)
);

A2O1A1Ixp33_ASAP7_75t_L g1251 ( 
.A1(n_1090),
.A2(n_1025),
.B(n_1023),
.C(n_1021),
.Y(n_1251)
);

A2O1A1Ixp33_ASAP7_75t_L g1252 ( 
.A1(n_1054),
.A2(n_1025),
.B(n_1023),
.C(n_1021),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_SL g1253 ( 
.A(n_1066),
.B(n_1009),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_1193),
.Y(n_1254)
);

INVx1_ASAP7_75t_SL g1255 ( 
.A(n_1030),
.Y(n_1255)
);

NOR2xp33_ASAP7_75t_L g1256 ( 
.A(n_1072),
.B(n_1009),
.Y(n_1256)
);

INVx3_ASAP7_75t_L g1257 ( 
.A(n_1056),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1098),
.Y(n_1258)
);

INVx3_ASAP7_75t_SL g1259 ( 
.A(n_1197),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1116),
.Y(n_1260)
);

OAI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1028),
.A2(n_1018),
.B(n_1011),
.Y(n_1261)
);

BUFx6f_ASAP7_75t_L g1262 ( 
.A(n_1056),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1145),
.Y(n_1263)
);

OAI21xp33_ASAP7_75t_SL g1264 ( 
.A1(n_1154),
.A2(n_1018),
.B(n_1011),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1038),
.A2(n_968),
.B(n_931),
.Y(n_1265)
);

HB1xp67_ASAP7_75t_L g1266 ( 
.A(n_1110),
.Y(n_1266)
);

OR2x2_ASAP7_75t_L g1267 ( 
.A(n_1106),
.B(n_1019),
.Y(n_1267)
);

A2O1A1Ixp33_ASAP7_75t_L g1268 ( 
.A1(n_1080),
.A2(n_1019),
.B(n_989),
.C(n_981),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1034),
.A2(n_981),
.B(n_931),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1057),
.B(n_658),
.Y(n_1270)
);

BUFx2_ASAP7_75t_L g1271 ( 
.A(n_1110),
.Y(n_1271)
);

A2O1A1Ixp33_ASAP7_75t_L g1272 ( 
.A1(n_1123),
.A2(n_989),
.B(n_451),
.C(n_448),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_1048),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1113),
.Y(n_1274)
);

A2O1A1Ixp33_ASAP7_75t_L g1275 ( 
.A1(n_1123),
.A2(n_1177),
.B(n_1174),
.C(n_1075),
.Y(n_1275)
);

A2O1A1Ixp33_ASAP7_75t_SL g1276 ( 
.A1(n_1177),
.A2(n_610),
.B(n_619),
.C(n_618),
.Y(n_1276)
);

OAI22xp5_ASAP7_75t_L g1277 ( 
.A1(n_1066),
.A2(n_464),
.B1(n_453),
.B2(n_451),
.Y(n_1277)
);

AOI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1036),
.A2(n_683),
.B(n_668),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1138),
.Y(n_1279)
);

BUFx6f_ASAP7_75t_L g1280 ( 
.A(n_1056),
.Y(n_1280)
);

BUFx6f_ASAP7_75t_L g1281 ( 
.A(n_1070),
.Y(n_1281)
);

NOR2xp33_ASAP7_75t_L g1282 ( 
.A(n_1153),
.B(n_356),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_SL g1283 ( 
.A(n_1050),
.B(n_422),
.Y(n_1283)
);

INVx4_ASAP7_75t_L g1284 ( 
.A(n_1070),
.Y(n_1284)
);

OAI22xp5_ASAP7_75t_L g1285 ( 
.A1(n_1084),
.A2(n_446),
.B1(n_439),
.B2(n_438),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1032),
.B(n_685),
.Y(n_1286)
);

INVx4_ASAP7_75t_L g1287 ( 
.A(n_1070),
.Y(n_1287)
);

AOI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1029),
.A2(n_683),
.B(n_668),
.Y(n_1288)
);

INVxp67_ASAP7_75t_L g1289 ( 
.A(n_1104),
.Y(n_1289)
);

AOI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1068),
.A2(n_683),
.B(n_241),
.Y(n_1290)
);

NOR2xp33_ASAP7_75t_L g1291 ( 
.A(n_1211),
.B(n_359),
.Y(n_1291)
);

NOR2xp33_ASAP7_75t_L g1292 ( 
.A(n_1179),
.B(n_361),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_SL g1293 ( 
.A(n_1133),
.B(n_1094),
.Y(n_1293)
);

AOI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1086),
.A2(n_683),
.B(n_241),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_1175),
.Y(n_1295)
);

NAND3xp33_ASAP7_75t_SL g1296 ( 
.A(n_1204),
.B(n_366),
.C(n_363),
.Y(n_1296)
);

AOI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1089),
.A2(n_683),
.B(n_241),
.Y(n_1297)
);

AOI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1043),
.A2(n_683),
.B(n_608),
.Y(n_1298)
);

NOR2xp33_ASAP7_75t_L g1299 ( 
.A(n_1181),
.B(n_368),
.Y(n_1299)
);

OAI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1040),
.A2(n_596),
.B(n_594),
.Y(n_1300)
);

O2A1O1Ixp33_ASAP7_75t_L g1301 ( 
.A1(n_1136),
.A2(n_446),
.B(n_439),
.C(n_436),
.Y(n_1301)
);

INVxp67_ASAP7_75t_SL g1302 ( 
.A(n_1070),
.Y(n_1302)
);

INVx1_ASAP7_75t_SL g1303 ( 
.A(n_1128),
.Y(n_1303)
);

O2A1O1Ixp5_ASAP7_75t_L g1304 ( 
.A1(n_1040),
.A2(n_691),
.B(n_690),
.C(n_688),
.Y(n_1304)
);

O2A1O1Ixp5_ASAP7_75t_L g1305 ( 
.A1(n_1152),
.A2(n_691),
.B(n_690),
.C(n_688),
.Y(n_1305)
);

NOR2xp67_ASAP7_75t_L g1306 ( 
.A(n_1117),
.B(n_104),
.Y(n_1306)
);

NOR2xp33_ASAP7_75t_L g1307 ( 
.A(n_1133),
.B(n_372),
.Y(n_1307)
);

BUFx8_ASAP7_75t_L g1308 ( 
.A(n_1128),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_SL g1309 ( 
.A(n_1094),
.B(n_422),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_SL g1310 ( 
.A(n_1033),
.B(n_422),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1156),
.Y(n_1311)
);

AOI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1039),
.A2(n_683),
.B(n_608),
.Y(n_1312)
);

INVx2_ASAP7_75t_SL g1313 ( 
.A(n_1161),
.Y(n_1313)
);

AOI221xp5_ASAP7_75t_L g1314 ( 
.A1(n_1095),
.A2(n_408),
.B1(n_381),
.B2(n_385),
.C(n_388),
.Y(n_1314)
);

AOI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1049),
.A2(n_1055),
.B(n_1081),
.Y(n_1315)
);

BUFx6f_ASAP7_75t_L g1316 ( 
.A(n_1083),
.Y(n_1316)
);

AND2x4_ASAP7_75t_L g1317 ( 
.A(n_1033),
.B(n_587),
.Y(n_1317)
);

OAI22xp5_ASAP7_75t_L g1318 ( 
.A1(n_1125),
.A2(n_426),
.B1(n_430),
.B2(n_436),
.Y(n_1318)
);

BUFx2_ASAP7_75t_L g1319 ( 
.A(n_1087),
.Y(n_1319)
);

NOR2xp33_ASAP7_75t_L g1320 ( 
.A(n_1062),
.B(n_1131),
.Y(n_1320)
);

AOI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1085),
.A2(n_683),
.B(n_596),
.Y(n_1321)
);

AOI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1152),
.A2(n_596),
.B(n_594),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1178),
.Y(n_1323)
);

O2A1O1Ixp33_ASAP7_75t_L g1324 ( 
.A1(n_1058),
.A2(n_588),
.B(n_620),
.C(n_616),
.Y(n_1324)
);

O2A1O1Ixp33_ASAP7_75t_L g1325 ( 
.A1(n_1058),
.A2(n_588),
.B(n_620),
.C(n_616),
.Y(n_1325)
);

AOI21x1_ASAP7_75t_L g1326 ( 
.A1(n_1065),
.A2(n_603),
.B(n_594),
.Y(n_1326)
);

OAI22xp5_ASAP7_75t_L g1327 ( 
.A1(n_1184),
.A2(n_409),
.B1(n_465),
.B2(n_463),
.Y(n_1327)
);

OAI22xp5_ASAP7_75t_L g1328 ( 
.A1(n_1189),
.A2(n_406),
.B1(n_458),
.B2(n_445),
.Y(n_1328)
);

AOI22x1_ASAP7_75t_L g1329 ( 
.A1(n_1194),
.A2(n_646),
.B1(n_645),
.B2(n_614),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1131),
.B(n_685),
.Y(n_1330)
);

HB1xp67_ASAP7_75t_L g1331 ( 
.A(n_1183),
.Y(n_1331)
);

AOI22xp5_ASAP7_75t_L g1332 ( 
.A1(n_1190),
.A2(n_452),
.B1(n_619),
.B2(n_618),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1137),
.B(n_1189),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1161),
.B(n_357),
.Y(n_1334)
);

NOR2xp33_ASAP7_75t_L g1335 ( 
.A(n_1137),
.B(n_390),
.Y(n_1335)
);

NAND3xp33_ASAP7_75t_SL g1336 ( 
.A(n_1139),
.B(n_402),
.C(n_420),
.Y(n_1336)
);

AOI21x1_ASAP7_75t_L g1337 ( 
.A1(n_1170),
.A2(n_607),
.B(n_603),
.Y(n_1337)
);

O2A1O1Ixp33_ASAP7_75t_SL g1338 ( 
.A1(n_1091),
.A2(n_607),
.B(n_603),
.C(n_604),
.Y(n_1338)
);

AOI21xp33_ASAP7_75t_L g1339 ( 
.A1(n_1093),
.A2(n_691),
.B(n_690),
.Y(n_1339)
);

INVx8_ASAP7_75t_L g1340 ( 
.A(n_1083),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1203),
.B(n_685),
.Y(n_1341)
);

NOR3xp33_ASAP7_75t_L g1342 ( 
.A(n_1212),
.B(n_401),
.C(n_419),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1203),
.B(n_686),
.Y(n_1343)
);

NOR2xp33_ASAP7_75t_L g1344 ( 
.A(n_1047),
.B(n_392),
.Y(n_1344)
);

NOR2xp33_ASAP7_75t_L g1345 ( 
.A(n_1059),
.B(n_404),
.Y(n_1345)
);

AOI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1154),
.A2(n_607),
.B(n_606),
.Y(n_1346)
);

OAI22xp5_ASAP7_75t_L g1347 ( 
.A1(n_1187),
.A2(n_688),
.B1(n_686),
.B2(n_562),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1205),
.B(n_686),
.Y(n_1348)
);

O2A1O1Ixp33_ASAP7_75t_L g1349 ( 
.A1(n_1212),
.A2(n_1150),
.B(n_1091),
.C(n_1082),
.Y(n_1349)
);

BUFx6f_ASAP7_75t_L g1350 ( 
.A(n_1083),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1216),
.B(n_657),
.Y(n_1351)
);

CKINVDCx5p33_ASAP7_75t_R g1352 ( 
.A(n_1149),
.Y(n_1352)
);

CKINVDCx20_ASAP7_75t_R g1353 ( 
.A(n_1149),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1148),
.Y(n_1354)
);

O2A1O1Ixp33_ASAP7_75t_L g1355 ( 
.A1(n_1064),
.A2(n_646),
.B(n_645),
.C(n_606),
.Y(n_1355)
);

AND2x2_ASAP7_75t_SL g1356 ( 
.A(n_1083),
.B(n_562),
.Y(n_1356)
);

HB1xp67_ASAP7_75t_L g1357 ( 
.A(n_1087),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_SL g1358 ( 
.A(n_1108),
.B(n_1139),
.Y(n_1358)
);

BUFx4f_ASAP7_75t_L g1359 ( 
.A(n_1087),
.Y(n_1359)
);

BUFx6f_ASAP7_75t_L g1360 ( 
.A(n_1108),
.Y(n_1360)
);

AOI22xp5_ASAP7_75t_L g1361 ( 
.A1(n_1071),
.A2(n_452),
.B1(n_660),
.B2(n_657),
.Y(n_1361)
);

OAI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1158),
.A2(n_604),
.B(n_606),
.Y(n_1362)
);

INVxp67_ASAP7_75t_SL g1363 ( 
.A(n_1108),
.Y(n_1363)
);

AND2x4_ASAP7_75t_L g1364 ( 
.A(n_1162),
.B(n_563),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1164),
.Y(n_1365)
);

AOI21xp5_ASAP7_75t_L g1366 ( 
.A1(n_1187),
.A2(n_604),
.B(n_639),
.Y(n_1366)
);

NOR2x1_ASAP7_75t_L g1367 ( 
.A(n_1130),
.B(n_660),
.Y(n_1367)
);

O2A1O1Ixp33_ASAP7_75t_L g1368 ( 
.A1(n_1077),
.A2(n_570),
.B(n_563),
.C(n_564),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_SL g1369 ( 
.A(n_1108),
.B(n_452),
.Y(n_1369)
);

OAI22xp5_ASAP7_75t_L g1370 ( 
.A1(n_1196),
.A2(n_572),
.B1(n_564),
.B2(n_566),
.Y(n_1370)
);

AOI21xp5_ASAP7_75t_L g1371 ( 
.A1(n_1099),
.A2(n_639),
.B(n_641),
.Y(n_1371)
);

O2A1O1Ixp33_ASAP7_75t_L g1372 ( 
.A1(n_1077),
.A2(n_566),
.B(n_569),
.C(n_570),
.Y(n_1372)
);

INVx4_ASAP7_75t_L g1373 ( 
.A(n_1162),
.Y(n_1373)
);

INVx3_ASAP7_75t_L g1374 ( 
.A(n_1165),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1142),
.B(n_1146),
.Y(n_1375)
);

OAI22x1_ASAP7_75t_L g1376 ( 
.A1(n_1191),
.A2(n_569),
.B1(n_357),
.B2(n_13),
.Y(n_1376)
);

AOI21xp5_ASAP7_75t_L g1377 ( 
.A1(n_1035),
.A2(n_639),
.B(n_641),
.Y(n_1377)
);

AOI21xp5_ASAP7_75t_L g1378 ( 
.A1(n_1037),
.A2(n_639),
.B(n_641),
.Y(n_1378)
);

A2O1A1Ixp33_ASAP7_75t_SL g1379 ( 
.A1(n_1165),
.A2(n_687),
.B(n_684),
.C(n_638),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1173),
.Y(n_1380)
);

AOI21xp5_ASAP7_75t_L g1381 ( 
.A1(n_1109),
.A2(n_639),
.B(n_638),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1231),
.B(n_357),
.Y(n_1382)
);

AND2x4_ASAP7_75t_L g1383 ( 
.A(n_1271),
.B(n_1172),
.Y(n_1383)
);

NAND3xp33_ASAP7_75t_SL g1384 ( 
.A(n_1282),
.B(n_1199),
.C(n_1217),
.Y(n_1384)
);

AO31x2_ASAP7_75t_L g1385 ( 
.A1(n_1221),
.A2(n_1210),
.A3(n_1127),
.B(n_1134),
.Y(n_1385)
);

AO22x2_ASAP7_75t_L g1386 ( 
.A1(n_1277),
.A2(n_1191),
.B1(n_1192),
.B2(n_1118),
.Y(n_1386)
);

AOI21xp5_ASAP7_75t_SL g1387 ( 
.A1(n_1234),
.A2(n_1112),
.B(n_1088),
.Y(n_1387)
);

NOR2xp33_ASAP7_75t_L g1388 ( 
.A(n_1292),
.B(n_1118),
.Y(n_1388)
);

OAI21x1_ASAP7_75t_L g1389 ( 
.A1(n_1337),
.A2(n_1159),
.B(n_1209),
.Y(n_1389)
);

AOI21xp5_ASAP7_75t_L g1390 ( 
.A1(n_1315),
.A2(n_1195),
.B(n_1171),
.Y(n_1390)
);

AO31x2_ASAP7_75t_L g1391 ( 
.A1(n_1275),
.A2(n_1147),
.A3(n_1129),
.B(n_1143),
.Y(n_1391)
);

AOI21xp5_ASAP7_75t_L g1392 ( 
.A1(n_1265),
.A2(n_1101),
.B(n_1092),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1354),
.B(n_1172),
.Y(n_1393)
);

A2O1A1Ixp33_ASAP7_75t_L g1394 ( 
.A1(n_1299),
.A2(n_1103),
.B(n_1180),
.C(n_1051),
.Y(n_1394)
);

BUFx6f_ASAP7_75t_L g1395 ( 
.A(n_1219),
.Y(n_1395)
);

OAI21x1_ASAP7_75t_L g1396 ( 
.A1(n_1278),
.A2(n_1097),
.B(n_1111),
.Y(n_1396)
);

INVx1_ASAP7_75t_SL g1397 ( 
.A(n_1303),
.Y(n_1397)
);

NOR2x1_ASAP7_75t_SL g1398 ( 
.A(n_1230),
.B(n_1235),
.Y(n_1398)
);

AO31x2_ASAP7_75t_L g1399 ( 
.A1(n_1251),
.A2(n_1114),
.A3(n_1160),
.B(n_1163),
.Y(n_1399)
);

A2O1A1Ixp33_ASAP7_75t_L g1400 ( 
.A1(n_1222),
.A2(n_1140),
.B(n_1176),
.C(n_1121),
.Y(n_1400)
);

AO31x2_ASAP7_75t_L g1401 ( 
.A1(n_1252),
.A2(n_1166),
.A3(n_1151),
.B(n_1155),
.Y(n_1401)
);

AOI21xp5_ASAP7_75t_L g1402 ( 
.A1(n_1375),
.A2(n_1102),
.B(n_1124),
.Y(n_1402)
);

AO31x2_ASAP7_75t_L g1403 ( 
.A1(n_1250),
.A2(n_1218),
.A3(n_1167),
.B(n_1115),
.Y(n_1403)
);

OAI21x1_ASAP7_75t_L g1404 ( 
.A1(n_1326),
.A2(n_1132),
.B(n_1144),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_L g1405 ( 
.A1(n_1298),
.A2(n_1157),
.B(n_1126),
.Y(n_1405)
);

OAI21x1_ASAP7_75t_L g1406 ( 
.A1(n_1321),
.A2(n_1186),
.B(n_1200),
.Y(n_1406)
);

BUFx12f_ASAP7_75t_L g1407 ( 
.A(n_1352),
.Y(n_1407)
);

O2A1O1Ixp33_ASAP7_75t_L g1408 ( 
.A1(n_1277),
.A2(n_1122),
.B(n_1182),
.C(n_1201),
.Y(n_1408)
);

AOI21xp5_ASAP7_75t_L g1409 ( 
.A1(n_1375),
.A2(n_1169),
.B(n_1214),
.Y(n_1409)
);

O2A1O1Ixp33_ASAP7_75t_L g1410 ( 
.A1(n_1289),
.A2(n_1122),
.B(n_1201),
.C(n_1100),
.Y(n_1410)
);

OAI21xp5_ASAP7_75t_L g1411 ( 
.A1(n_1269),
.A2(n_1208),
.B(n_1206),
.Y(n_1411)
);

OR2x2_ASAP7_75t_L g1412 ( 
.A(n_1267),
.B(n_1188),
.Y(n_1412)
);

AOI22xp5_ASAP7_75t_SL g1413 ( 
.A1(n_1247),
.A2(n_357),
.B1(n_1107),
.B2(n_452),
.Y(n_1413)
);

BUFx2_ASAP7_75t_L g1414 ( 
.A(n_1227),
.Y(n_1414)
);

OAI21x1_ASAP7_75t_L g1415 ( 
.A1(n_1261),
.A2(n_1215),
.B(n_1207),
.Y(n_1415)
);

INVx2_ASAP7_75t_SL g1416 ( 
.A(n_1313),
.Y(n_1416)
);

AOI21x1_ASAP7_75t_L g1417 ( 
.A1(n_1312),
.A2(n_1202),
.B(n_1198),
.Y(n_1417)
);

NOR2xp33_ASAP7_75t_L g1418 ( 
.A(n_1255),
.B(n_10),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1365),
.B(n_684),
.Y(n_1419)
);

O2A1O1Ixp33_ASAP7_75t_SL g1420 ( 
.A1(n_1253),
.A2(n_638),
.B(n_629),
.C(n_687),
.Y(n_1420)
);

AO31x2_ASAP7_75t_L g1421 ( 
.A1(n_1290),
.A2(n_687),
.A3(n_684),
.B(n_629),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1311),
.Y(n_1422)
);

AO31x2_ASAP7_75t_L g1423 ( 
.A1(n_1268),
.A2(n_629),
.A3(n_14),
.B(n_15),
.Y(n_1423)
);

A2O1A1Ixp33_ASAP7_75t_L g1424 ( 
.A1(n_1306),
.A2(n_11),
.B(n_16),
.C(n_18),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1323),
.Y(n_1425)
);

AOI21x1_ASAP7_75t_L g1426 ( 
.A1(n_1249),
.A2(n_233),
.B(n_230),
.Y(n_1426)
);

AO32x2_ASAP7_75t_L g1427 ( 
.A1(n_1285),
.A2(n_11),
.A3(n_16),
.B1(n_18),
.B2(n_19),
.Y(n_1427)
);

AOI21xp5_ASAP7_75t_L g1428 ( 
.A1(n_1245),
.A2(n_226),
.B(n_224),
.Y(n_1428)
);

AOI21xp5_ASAP7_75t_L g1429 ( 
.A1(n_1239),
.A2(n_220),
.B(n_212),
.Y(n_1429)
);

OAI21x1_ASAP7_75t_L g1430 ( 
.A1(n_1329),
.A2(n_206),
.B(n_200),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1266),
.B(n_21),
.Y(n_1431)
);

NAND2x1p5_ASAP7_75t_L g1432 ( 
.A(n_1284),
.B(n_112),
.Y(n_1432)
);

OAI21x1_ASAP7_75t_L g1433 ( 
.A1(n_1288),
.A2(n_195),
.B(n_194),
.Y(n_1433)
);

NOR2x2_ASAP7_75t_L g1434 ( 
.A(n_1273),
.B(n_21),
.Y(n_1434)
);

AO21x2_ASAP7_75t_L g1435 ( 
.A1(n_1362),
.A2(n_184),
.B(n_182),
.Y(n_1435)
);

AO21x1_ASAP7_75t_L g1436 ( 
.A1(n_1324),
.A2(n_1325),
.B(n_1349),
.Y(n_1436)
);

BUFx6f_ASAP7_75t_L g1437 ( 
.A(n_1219),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1380),
.B(n_1286),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1344),
.B(n_23),
.Y(n_1439)
);

BUFx2_ASAP7_75t_L g1440 ( 
.A(n_1227),
.Y(n_1440)
);

O2A1O1Ixp33_ASAP7_75t_SL g1441 ( 
.A1(n_1272),
.A2(n_178),
.B(n_169),
.C(n_168),
.Y(n_1441)
);

AO32x2_ASAP7_75t_L g1442 ( 
.A1(n_1285),
.A2(n_23),
.A3(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_1442)
);

INVx2_ASAP7_75t_SL g1443 ( 
.A(n_1308),
.Y(n_1443)
);

AOI21xp5_ASAP7_75t_L g1444 ( 
.A1(n_1236),
.A2(n_161),
.B(n_155),
.Y(n_1444)
);

AO21x2_ASAP7_75t_L g1445 ( 
.A1(n_1362),
.A2(n_153),
.B(n_148),
.Y(n_1445)
);

OAI22xp5_ASAP7_75t_L g1446 ( 
.A1(n_1356),
.A2(n_26),
.B1(n_29),
.B2(n_36),
.Y(n_1446)
);

BUFx2_ASAP7_75t_L g1447 ( 
.A(n_1226),
.Y(n_1447)
);

AOI21xp5_ASAP7_75t_L g1448 ( 
.A1(n_1223),
.A2(n_147),
.B(n_146),
.Y(n_1448)
);

A2O1A1Ixp33_ASAP7_75t_L g1449 ( 
.A1(n_1256),
.A2(n_36),
.B(n_37),
.C(n_38),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1345),
.B(n_39),
.Y(n_1450)
);

NOR2xp67_ASAP7_75t_SL g1451 ( 
.A(n_1243),
.B(n_43),
.Y(n_1451)
);

HB1xp67_ASAP7_75t_L g1452 ( 
.A(n_1317),
.Y(n_1452)
);

INVx2_ASAP7_75t_SL g1453 ( 
.A(n_1308),
.Y(n_1453)
);

O2A1O1Ixp33_ASAP7_75t_L g1454 ( 
.A1(n_1283),
.A2(n_44),
.B(n_45),
.C(n_47),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1240),
.Y(n_1455)
);

NOR2xp33_ASAP7_75t_SL g1456 ( 
.A(n_1223),
.B(n_48),
.Y(n_1456)
);

NOR2xp33_ASAP7_75t_L g1457 ( 
.A(n_1307),
.B(n_1291),
.Y(n_1457)
);

AOI21x1_ASAP7_75t_L g1458 ( 
.A1(n_1300),
.A2(n_1381),
.B(n_1346),
.Y(n_1458)
);

AO31x2_ASAP7_75t_L g1459 ( 
.A1(n_1347),
.A2(n_49),
.A3(n_50),
.B(n_51),
.Y(n_1459)
);

AO32x2_ASAP7_75t_L g1460 ( 
.A1(n_1347),
.A2(n_52),
.A3(n_55),
.B1(n_57),
.B2(n_58),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_SL g1461 ( 
.A(n_1359),
.B(n_57),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1248),
.Y(n_1462)
);

BUFx2_ASAP7_75t_L g1463 ( 
.A(n_1357),
.Y(n_1463)
);

OAI22x1_ASAP7_75t_L g1464 ( 
.A1(n_1319),
.A2(n_59),
.B1(n_60),
.B2(n_62),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1295),
.Y(n_1465)
);

INVx5_ASAP7_75t_L g1466 ( 
.A(n_1340),
.Y(n_1466)
);

NOR2xp33_ASAP7_75t_L g1467 ( 
.A(n_1335),
.B(n_60),
.Y(n_1467)
);

AO31x2_ASAP7_75t_L g1468 ( 
.A1(n_1294),
.A2(n_1297),
.A3(n_1376),
.B(n_1320),
.Y(n_1468)
);

OAI21x1_ASAP7_75t_L g1469 ( 
.A1(n_1371),
.A2(n_143),
.B(n_140),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1317),
.B(n_62),
.Y(n_1470)
);

AOI21xp5_ASAP7_75t_L g1471 ( 
.A1(n_1232),
.A2(n_128),
.B(n_126),
.Y(n_1471)
);

O2A1O1Ixp33_ASAP7_75t_SL g1472 ( 
.A1(n_1358),
.A2(n_121),
.B(n_119),
.C(n_118),
.Y(n_1472)
);

NOR2xp33_ASAP7_75t_SL g1473 ( 
.A(n_1232),
.B(n_63),
.Y(n_1473)
);

CKINVDCx5p33_ASAP7_75t_R g1474 ( 
.A(n_1353),
.Y(n_1474)
);

OAI21x1_ASAP7_75t_L g1475 ( 
.A1(n_1300),
.A2(n_116),
.B(n_115),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_SL g1476 ( 
.A(n_1359),
.B(n_67),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1334),
.B(n_1364),
.Y(n_1477)
);

OAI21x1_ASAP7_75t_L g1478 ( 
.A1(n_1304),
.A2(n_68),
.B(n_69),
.Y(n_1478)
);

AOI21xp5_ASAP7_75t_L g1479 ( 
.A1(n_1225),
.A2(n_68),
.B(n_71),
.Y(n_1479)
);

INVxp67_ASAP7_75t_SL g1480 ( 
.A(n_1333),
.Y(n_1480)
);

AO31x2_ASAP7_75t_L g1481 ( 
.A1(n_1322),
.A2(n_73),
.A3(n_74),
.B(n_75),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_L g1482 ( 
.A1(n_1342),
.A2(n_75),
.B1(n_76),
.B2(n_77),
.Y(n_1482)
);

O2A1O1Ixp33_ASAP7_75t_L g1483 ( 
.A1(n_1318),
.A2(n_76),
.B(n_77),
.C(n_80),
.Y(n_1483)
);

AO31x2_ASAP7_75t_L g1484 ( 
.A1(n_1366),
.A2(n_1370),
.A3(n_1378),
.B(n_1377),
.Y(n_1484)
);

AOI221x1_ASAP7_75t_L g1485 ( 
.A1(n_1241),
.A2(n_82),
.B1(n_84),
.B2(n_85),
.C(n_88),
.Y(n_1485)
);

O2A1O1Ixp33_ASAP7_75t_L g1486 ( 
.A1(n_1318),
.A2(n_82),
.B(n_84),
.C(n_88),
.Y(n_1486)
);

AOI21xp5_ASAP7_75t_L g1487 ( 
.A1(n_1225),
.A2(n_89),
.B(n_94),
.Y(n_1487)
);

AOI21xp5_ASAP7_75t_L g1488 ( 
.A1(n_1229),
.A2(n_94),
.B(n_95),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_SL g1489 ( 
.A(n_1331),
.B(n_1246),
.Y(n_1489)
);

INVxp67_ASAP7_75t_L g1490 ( 
.A(n_1244),
.Y(n_1490)
);

OAI21x1_ASAP7_75t_L g1491 ( 
.A1(n_1233),
.A2(n_97),
.B(n_99),
.Y(n_1491)
);

OAI21xp5_ASAP7_75t_L g1492 ( 
.A1(n_1264),
.A2(n_99),
.B(n_100),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1242),
.B(n_1270),
.Y(n_1493)
);

OAI21x1_ASAP7_75t_L g1494 ( 
.A1(n_1305),
.A2(n_1348),
.B(n_1355),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1258),
.Y(n_1495)
);

OR2x2_ASAP7_75t_L g1496 ( 
.A(n_1327),
.B(n_1328),
.Y(n_1496)
);

AND2x4_ASAP7_75t_L g1497 ( 
.A(n_1293),
.B(n_1367),
.Y(n_1497)
);

AOI22xp5_ASAP7_75t_L g1498 ( 
.A1(n_1336),
.A2(n_1327),
.B1(n_1296),
.B2(n_1364),
.Y(n_1498)
);

OAI21x1_ASAP7_75t_L g1499 ( 
.A1(n_1341),
.A2(n_1343),
.B(n_1351),
.Y(n_1499)
);

OR2x2_ASAP7_75t_L g1500 ( 
.A(n_1328),
.B(n_1279),
.Y(n_1500)
);

BUFx6f_ASAP7_75t_L g1501 ( 
.A(n_1219),
.Y(n_1501)
);

A2O1A1Ixp33_ASAP7_75t_L g1502 ( 
.A1(n_1224),
.A2(n_1237),
.B(n_1238),
.C(n_1301),
.Y(n_1502)
);

OA21x2_ASAP7_75t_L g1503 ( 
.A1(n_1339),
.A2(n_1361),
.B(n_1330),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1260),
.B(n_1263),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1274),
.B(n_1220),
.Y(n_1505)
);

O2A1O1Ixp5_ASAP7_75t_L g1506 ( 
.A1(n_1309),
.A2(n_1369),
.B(n_1310),
.C(n_1276),
.Y(n_1506)
);

INVx2_ASAP7_75t_SL g1507 ( 
.A(n_1259),
.Y(n_1507)
);

AO32x2_ASAP7_75t_L g1508 ( 
.A1(n_1370),
.A2(n_1373),
.A3(n_1287),
.B1(n_1284),
.B2(n_1338),
.Y(n_1508)
);

BUFx6f_ASAP7_75t_L g1509 ( 
.A(n_1262),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1254),
.Y(n_1510)
);

INVx5_ASAP7_75t_L g1511 ( 
.A(n_1340),
.Y(n_1511)
);

NAND3xp33_ASAP7_75t_L g1512 ( 
.A(n_1314),
.B(n_1332),
.C(n_1228),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1374),
.B(n_1257),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1374),
.B(n_1257),
.Y(n_1514)
);

OR2x6_ASAP7_75t_L g1515 ( 
.A(n_1340),
.B(n_1262),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1373),
.Y(n_1516)
);

AO21x2_ASAP7_75t_L g1517 ( 
.A1(n_1339),
.A2(n_1379),
.B(n_1302),
.Y(n_1517)
);

NOR2xp33_ASAP7_75t_L g1518 ( 
.A(n_1363),
.B(n_1287),
.Y(n_1518)
);

OR2x6_ASAP7_75t_L g1519 ( 
.A(n_1262),
.B(n_1280),
.Y(n_1519)
);

OAI21xp5_ASAP7_75t_L g1520 ( 
.A1(n_1368),
.A2(n_1372),
.B(n_1281),
.Y(n_1520)
);

OAI21x1_ASAP7_75t_L g1521 ( 
.A1(n_1280),
.A2(n_1281),
.B(n_1316),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1360),
.B(n_1316),
.Y(n_1522)
);

INVx3_ASAP7_75t_L g1523 ( 
.A(n_1350),
.Y(n_1523)
);

OAI21xp5_ASAP7_75t_L g1524 ( 
.A1(n_1350),
.A2(n_1221),
.B(n_1250),
.Y(n_1524)
);

OAI21x1_ASAP7_75t_L g1525 ( 
.A1(n_1350),
.A2(n_1337),
.B(n_1278),
.Y(n_1525)
);

AND2x4_ASAP7_75t_L g1526 ( 
.A(n_1360),
.B(n_1271),
.Y(n_1526)
);

BUFx4f_ASAP7_75t_SL g1527 ( 
.A(n_1360),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1231),
.B(n_911),
.Y(n_1528)
);

CKINVDCx11_ASAP7_75t_R g1529 ( 
.A(n_1353),
.Y(n_1529)
);

AOI21xp5_ASAP7_75t_L g1530 ( 
.A1(n_1315),
.A2(n_1213),
.B(n_1135),
.Y(n_1530)
);

AOI21xp5_ASAP7_75t_L g1531 ( 
.A1(n_1315),
.A2(n_1213),
.B(n_1135),
.Y(n_1531)
);

AOI21xp5_ASAP7_75t_L g1532 ( 
.A1(n_1315),
.A2(n_1213),
.B(n_1135),
.Y(n_1532)
);

CKINVDCx5p33_ASAP7_75t_R g1533 ( 
.A(n_1243),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1354),
.B(n_1365),
.Y(n_1534)
);

INVx6_ASAP7_75t_L g1535 ( 
.A(n_1308),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1354),
.B(n_1365),
.Y(n_1536)
);

AND2x4_ASAP7_75t_L g1537 ( 
.A(n_1271),
.B(n_1293),
.Y(n_1537)
);

A2O1A1Ixp33_ASAP7_75t_L g1538 ( 
.A1(n_1221),
.A2(n_878),
.B(n_1282),
.C(n_1299),
.Y(n_1538)
);

A2O1A1Ixp33_ASAP7_75t_L g1539 ( 
.A1(n_1221),
.A2(n_878),
.B(n_1282),
.C(n_1299),
.Y(n_1539)
);

AOI21xp5_ASAP7_75t_L g1540 ( 
.A1(n_1315),
.A2(n_1213),
.B(n_1135),
.Y(n_1540)
);

INVx3_ASAP7_75t_L g1541 ( 
.A(n_1373),
.Y(n_1541)
);

AOI21xp5_ASAP7_75t_L g1542 ( 
.A1(n_1315),
.A2(n_1213),
.B(n_1135),
.Y(n_1542)
);

AO31x2_ASAP7_75t_L g1543 ( 
.A1(n_1221),
.A2(n_1275),
.A3(n_1315),
.B(n_1251),
.Y(n_1543)
);

AO21x1_ASAP7_75t_L g1544 ( 
.A1(n_1282),
.A2(n_878),
.B(n_1076),
.Y(n_1544)
);

NOR2xp33_ASAP7_75t_L g1545 ( 
.A(n_1231),
.B(n_878),
.Y(n_1545)
);

INVx1_ASAP7_75t_SL g1546 ( 
.A(n_1303),
.Y(n_1546)
);

O2A1O1Ixp33_ASAP7_75t_L g1547 ( 
.A1(n_1221),
.A2(n_878),
.B(n_860),
.C(n_1076),
.Y(n_1547)
);

O2A1O1Ixp33_ASAP7_75t_L g1548 ( 
.A1(n_1221),
.A2(n_878),
.B(n_860),
.C(n_1076),
.Y(n_1548)
);

AOI22xp5_ASAP7_75t_L g1549 ( 
.A1(n_1282),
.A2(n_878),
.B1(n_1063),
.B2(n_1076),
.Y(n_1549)
);

AO31x2_ASAP7_75t_L g1550 ( 
.A1(n_1221),
.A2(n_1275),
.A3(n_1315),
.B(n_1251),
.Y(n_1550)
);

AOI21xp5_ASAP7_75t_L g1551 ( 
.A1(n_1315),
.A2(n_1213),
.B(n_1135),
.Y(n_1551)
);

AOI21xp5_ASAP7_75t_L g1552 ( 
.A1(n_1315),
.A2(n_1213),
.B(n_1135),
.Y(n_1552)
);

O2A1O1Ixp33_ASAP7_75t_SL g1553 ( 
.A1(n_1221),
.A2(n_1045),
.B(n_1075),
.C(n_1275),
.Y(n_1553)
);

AOI21xp5_ASAP7_75t_L g1554 ( 
.A1(n_1315),
.A2(n_1213),
.B(n_1135),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1545),
.B(n_1457),
.Y(n_1555)
);

AOI22x1_ASAP7_75t_SL g1556 ( 
.A1(n_1474),
.A2(n_1533),
.B1(n_1397),
.B2(n_1546),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1528),
.B(n_1534),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1477),
.B(n_1382),
.Y(n_1558)
);

CKINVDCx20_ASAP7_75t_R g1559 ( 
.A(n_1529),
.Y(n_1559)
);

CKINVDCx5p33_ASAP7_75t_R g1560 ( 
.A(n_1407),
.Y(n_1560)
);

BUFx8_ASAP7_75t_L g1561 ( 
.A(n_1414),
.Y(n_1561)
);

INVx4_ASAP7_75t_L g1562 ( 
.A(n_1466),
.Y(n_1562)
);

INVx3_ASAP7_75t_L g1563 ( 
.A(n_1466),
.Y(n_1563)
);

BUFx10_ASAP7_75t_L g1564 ( 
.A(n_1535),
.Y(n_1564)
);

AOI22xp33_ASAP7_75t_L g1565 ( 
.A1(n_1549),
.A2(n_1473),
.B1(n_1456),
.B2(n_1467),
.Y(n_1565)
);

AOI22xp33_ASAP7_75t_SL g1566 ( 
.A1(n_1456),
.A2(n_1473),
.B1(n_1446),
.B2(n_1413),
.Y(n_1566)
);

AOI22xp33_ASAP7_75t_SL g1567 ( 
.A1(n_1446),
.A2(n_1413),
.B1(n_1496),
.B2(n_1439),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1452),
.B(n_1431),
.Y(n_1568)
);

OAI21xp33_ASAP7_75t_L g1569 ( 
.A1(n_1549),
.A2(n_1539),
.B(n_1538),
.Y(n_1569)
);

AOI22xp33_ASAP7_75t_L g1570 ( 
.A1(n_1544),
.A2(n_1450),
.B1(n_1512),
.B2(n_1487),
.Y(n_1570)
);

INVx1_ASAP7_75t_SL g1571 ( 
.A(n_1447),
.Y(n_1571)
);

BUFx3_ASAP7_75t_L g1572 ( 
.A(n_1527),
.Y(n_1572)
);

OAI22xp5_ASAP7_75t_L g1573 ( 
.A1(n_1547),
.A2(n_1548),
.B1(n_1536),
.B2(n_1534),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1490),
.B(n_1397),
.Y(n_1574)
);

AOI22xp33_ASAP7_75t_SL g1575 ( 
.A1(n_1512),
.A2(n_1479),
.B1(n_1388),
.B2(n_1524),
.Y(n_1575)
);

AOI22xp5_ASAP7_75t_L g1576 ( 
.A1(n_1489),
.A2(n_1498),
.B1(n_1537),
.B2(n_1476),
.Y(n_1576)
);

INVx6_ASAP7_75t_L g1577 ( 
.A(n_1466),
.Y(n_1577)
);

AOI22xp33_ASAP7_75t_L g1578 ( 
.A1(n_1482),
.A2(n_1464),
.B1(n_1461),
.B2(n_1384),
.Y(n_1578)
);

AOI22xp33_ASAP7_75t_L g1579 ( 
.A1(n_1492),
.A2(n_1436),
.B1(n_1524),
.B2(n_1438),
.Y(n_1579)
);

INVx4_ASAP7_75t_L g1580 ( 
.A(n_1511),
.Y(n_1580)
);

BUFx2_ASAP7_75t_L g1581 ( 
.A(n_1526),
.Y(n_1581)
);

CKINVDCx5p33_ASAP7_75t_R g1582 ( 
.A(n_1507),
.Y(n_1582)
);

INVx1_ASAP7_75t_SL g1583 ( 
.A(n_1546),
.Y(n_1583)
);

BUFx2_ASAP7_75t_L g1584 ( 
.A(n_1526),
.Y(n_1584)
);

BUFx2_ASAP7_75t_L g1585 ( 
.A(n_1463),
.Y(n_1585)
);

BUFx2_ASAP7_75t_L g1586 ( 
.A(n_1537),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1504),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1504),
.Y(n_1588)
);

AOI22xp33_ASAP7_75t_L g1589 ( 
.A1(n_1492),
.A2(n_1438),
.B1(n_1536),
.B2(n_1448),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1480),
.B(n_1412),
.Y(n_1590)
);

AOI22xp5_ASAP7_75t_L g1591 ( 
.A1(n_1498),
.A2(n_1497),
.B1(n_1418),
.B2(n_1451),
.Y(n_1591)
);

BUFx10_ASAP7_75t_L g1592 ( 
.A(n_1535),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1425),
.Y(n_1593)
);

BUFx6f_ASAP7_75t_L g1594 ( 
.A(n_1515),
.Y(n_1594)
);

AOI22xp33_ASAP7_75t_SL g1595 ( 
.A1(n_1485),
.A2(n_1445),
.B1(n_1435),
.B2(n_1440),
.Y(n_1595)
);

AOI22xp5_ASAP7_75t_SL g1596 ( 
.A1(n_1497),
.A2(n_1470),
.B1(n_1443),
.B2(n_1453),
.Y(n_1596)
);

BUFx12f_ASAP7_75t_L g1597 ( 
.A(n_1416),
.Y(n_1597)
);

INVx1_ASAP7_75t_SL g1598 ( 
.A(n_1434),
.Y(n_1598)
);

CKINVDCx11_ASAP7_75t_R g1599 ( 
.A(n_1395),
.Y(n_1599)
);

INVx3_ASAP7_75t_L g1600 ( 
.A(n_1511),
.Y(n_1600)
);

AOI22xp33_ASAP7_75t_L g1601 ( 
.A1(n_1471),
.A2(n_1435),
.B1(n_1445),
.B2(n_1500),
.Y(n_1601)
);

INVx6_ASAP7_75t_L g1602 ( 
.A(n_1511),
.Y(n_1602)
);

AOI22xp5_ASAP7_75t_L g1603 ( 
.A1(n_1383),
.A2(n_1553),
.B1(n_1424),
.B2(n_1493),
.Y(n_1603)
);

CKINVDCx6p67_ASAP7_75t_R g1604 ( 
.A(n_1515),
.Y(n_1604)
);

INVx1_ASAP7_75t_SL g1605 ( 
.A(n_1383),
.Y(n_1605)
);

BUFx3_ASAP7_75t_L g1606 ( 
.A(n_1515),
.Y(n_1606)
);

CKINVDCx11_ASAP7_75t_R g1607 ( 
.A(n_1395),
.Y(n_1607)
);

BUFx3_ASAP7_75t_L g1608 ( 
.A(n_1395),
.Y(n_1608)
);

AOI22xp33_ASAP7_75t_L g1609 ( 
.A1(n_1488),
.A2(n_1462),
.B1(n_1495),
.B2(n_1455),
.Y(n_1609)
);

INVx6_ASAP7_75t_L g1610 ( 
.A(n_1437),
.Y(n_1610)
);

BUFx10_ASAP7_75t_L g1611 ( 
.A(n_1437),
.Y(n_1611)
);

AOI22xp33_ASAP7_75t_SL g1612 ( 
.A1(n_1427),
.A2(n_1442),
.B1(n_1460),
.B2(n_1386),
.Y(n_1612)
);

OAI21xp5_ASAP7_75t_SL g1613 ( 
.A1(n_1483),
.A2(n_1486),
.B(n_1449),
.Y(n_1613)
);

INVx1_ASAP7_75t_SL g1614 ( 
.A(n_1522),
.Y(n_1614)
);

CKINVDCx11_ASAP7_75t_R g1615 ( 
.A(n_1437),
.Y(n_1615)
);

NAND2x1p5_ASAP7_75t_L g1616 ( 
.A(n_1541),
.B(n_1521),
.Y(n_1616)
);

INVx1_ASAP7_75t_SL g1617 ( 
.A(n_1513),
.Y(n_1617)
);

INVx2_ASAP7_75t_SL g1618 ( 
.A(n_1501),
.Y(n_1618)
);

INVx6_ASAP7_75t_L g1619 ( 
.A(n_1501),
.Y(n_1619)
);

OAI22xp5_ASAP7_75t_L g1620 ( 
.A1(n_1393),
.A2(n_1387),
.B1(n_1394),
.B2(n_1505),
.Y(n_1620)
);

NAND2x1p5_ASAP7_75t_L g1621 ( 
.A(n_1541),
.B(n_1516),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1505),
.Y(n_1622)
);

CKINVDCx11_ASAP7_75t_R g1623 ( 
.A(n_1501),
.Y(n_1623)
);

BUFx3_ASAP7_75t_L g1624 ( 
.A(n_1509),
.Y(n_1624)
);

AOI22xp33_ASAP7_75t_SL g1625 ( 
.A1(n_1427),
.A2(n_1442),
.B1(n_1460),
.B2(n_1386),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1510),
.Y(n_1626)
);

AOI22xp33_ASAP7_75t_SL g1627 ( 
.A1(n_1427),
.A2(n_1442),
.B1(n_1460),
.B2(n_1432),
.Y(n_1627)
);

CKINVDCx20_ASAP7_75t_R g1628 ( 
.A(n_1509),
.Y(n_1628)
);

AOI22xp33_ASAP7_75t_L g1629 ( 
.A1(n_1503),
.A2(n_1444),
.B1(n_1419),
.B2(n_1393),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1514),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1514),
.Y(n_1631)
);

AOI22xp33_ASAP7_75t_SL g1632 ( 
.A1(n_1503),
.A2(n_1398),
.B1(n_1491),
.B2(n_1390),
.Y(n_1632)
);

AOI22xp33_ASAP7_75t_L g1633 ( 
.A1(n_1429),
.A2(n_1428),
.B1(n_1402),
.B2(n_1499),
.Y(n_1633)
);

INVx5_ASAP7_75t_L g1634 ( 
.A(n_1519),
.Y(n_1634)
);

CKINVDCx11_ASAP7_75t_R g1635 ( 
.A(n_1509),
.Y(n_1635)
);

CKINVDCx11_ASAP7_75t_R g1636 ( 
.A(n_1519),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1518),
.B(n_1454),
.Y(n_1637)
);

HB1xp67_ASAP7_75t_L g1638 ( 
.A(n_1543),
.Y(n_1638)
);

BUFx2_ASAP7_75t_L g1639 ( 
.A(n_1523),
.Y(n_1639)
);

INVx6_ASAP7_75t_L g1640 ( 
.A(n_1519),
.Y(n_1640)
);

BUFx5_ASAP7_75t_L g1641 ( 
.A(n_1391),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1481),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1481),
.Y(n_1643)
);

OAI22xp5_ASAP7_75t_L g1644 ( 
.A1(n_1502),
.A2(n_1400),
.B1(n_1410),
.B2(n_1520),
.Y(n_1644)
);

OAI21xp5_ASAP7_75t_L g1645 ( 
.A1(n_1506),
.A2(n_1409),
.B(n_1408),
.Y(n_1645)
);

BUFx6f_ASAP7_75t_L g1646 ( 
.A(n_1426),
.Y(n_1646)
);

BUFx2_ASAP7_75t_SL g1647 ( 
.A(n_1530),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1481),
.Y(n_1648)
);

CKINVDCx11_ASAP7_75t_R g1649 ( 
.A(n_1472),
.Y(n_1649)
);

AOI22xp33_ASAP7_75t_L g1650 ( 
.A1(n_1478),
.A2(n_1475),
.B1(n_1517),
.B2(n_1520),
.Y(n_1650)
);

AOI22xp33_ASAP7_75t_L g1651 ( 
.A1(n_1517),
.A2(n_1411),
.B1(n_1433),
.B2(n_1405),
.Y(n_1651)
);

OAI22xp5_ASAP7_75t_L g1652 ( 
.A1(n_1531),
.A2(n_1554),
.B1(n_1552),
.B2(n_1551),
.Y(n_1652)
);

CKINVDCx20_ASAP7_75t_R g1653 ( 
.A(n_1411),
.Y(n_1653)
);

OAI22xp5_ASAP7_75t_L g1654 ( 
.A1(n_1532),
.A2(n_1542),
.B1(n_1540),
.B2(n_1458),
.Y(n_1654)
);

BUFx2_ASAP7_75t_SL g1655 ( 
.A(n_1392),
.Y(n_1655)
);

BUFx6f_ASAP7_75t_L g1656 ( 
.A(n_1508),
.Y(n_1656)
);

OAI22xp5_ASAP7_75t_L g1657 ( 
.A1(n_1417),
.A2(n_1550),
.B1(n_1543),
.B2(n_1468),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1543),
.B(n_1550),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1459),
.B(n_1423),
.Y(n_1659)
);

AOI22xp33_ASAP7_75t_SL g1660 ( 
.A1(n_1430),
.A2(n_1459),
.B1(n_1469),
.B2(n_1550),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1459),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1420),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1468),
.B(n_1385),
.Y(n_1663)
);

OAI22xp33_ASAP7_75t_L g1664 ( 
.A1(n_1441),
.A2(n_1508),
.B1(n_1468),
.B2(n_1385),
.Y(n_1664)
);

BUFx12f_ASAP7_75t_L g1665 ( 
.A(n_1403),
.Y(n_1665)
);

INVx1_ASAP7_75t_SL g1666 ( 
.A(n_1525),
.Y(n_1666)
);

AOI22xp5_ASAP7_75t_L g1667 ( 
.A1(n_1494),
.A2(n_1396),
.B1(n_1415),
.B2(n_1404),
.Y(n_1667)
);

INVx6_ASAP7_75t_L g1668 ( 
.A(n_1508),
.Y(n_1668)
);

OAI22xp5_ASAP7_75t_L g1669 ( 
.A1(n_1385),
.A2(n_1484),
.B1(n_1391),
.B2(n_1403),
.Y(n_1669)
);

INVx11_ASAP7_75t_L g1670 ( 
.A(n_1403),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1391),
.B(n_1421),
.Y(n_1671)
);

INVx4_ASAP7_75t_L g1672 ( 
.A(n_1421),
.Y(n_1672)
);

BUFx3_ASAP7_75t_L g1673 ( 
.A(n_1484),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1401),
.Y(n_1674)
);

AOI22xp33_ASAP7_75t_SL g1675 ( 
.A1(n_1406),
.A2(n_1389),
.B1(n_1401),
.B2(n_1399),
.Y(n_1675)
);

BUFx10_ASAP7_75t_L g1676 ( 
.A(n_1399),
.Y(n_1676)
);

AOI22xp33_ASAP7_75t_L g1677 ( 
.A1(n_1401),
.A2(n_1549),
.B1(n_1456),
.B2(n_1473),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1399),
.Y(n_1678)
);

BUFx3_ASAP7_75t_L g1679 ( 
.A(n_1447),
.Y(n_1679)
);

AOI22xp33_ASAP7_75t_L g1680 ( 
.A1(n_1549),
.A2(n_1456),
.B1(n_1473),
.B2(n_1467),
.Y(n_1680)
);

AOI22xp33_ASAP7_75t_L g1681 ( 
.A1(n_1549),
.A2(n_1456),
.B1(n_1473),
.B2(n_1467),
.Y(n_1681)
);

AOI22xp33_ASAP7_75t_L g1682 ( 
.A1(n_1549),
.A2(n_1456),
.B1(n_1473),
.B2(n_1467),
.Y(n_1682)
);

BUFx12f_ASAP7_75t_L g1683 ( 
.A(n_1529),
.Y(n_1683)
);

CKINVDCx11_ASAP7_75t_R g1684 ( 
.A(n_1529),
.Y(n_1684)
);

INVx5_ASAP7_75t_L g1685 ( 
.A(n_1515),
.Y(n_1685)
);

AOI22xp33_ASAP7_75t_L g1686 ( 
.A1(n_1549),
.A2(n_1456),
.B1(n_1473),
.B2(n_1467),
.Y(n_1686)
);

AOI22xp33_ASAP7_75t_SL g1687 ( 
.A1(n_1456),
.A2(n_1473),
.B1(n_1090),
.B2(n_1072),
.Y(n_1687)
);

BUFx12f_ASAP7_75t_L g1688 ( 
.A(n_1529),
.Y(n_1688)
);

OAI22xp33_ASAP7_75t_L g1689 ( 
.A1(n_1456),
.A2(n_1473),
.B1(n_1549),
.B2(n_1090),
.Y(n_1689)
);

INVx1_ASAP7_75t_SL g1690 ( 
.A(n_1447),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1528),
.B(n_1545),
.Y(n_1691)
);

INVx6_ASAP7_75t_L g1692 ( 
.A(n_1466),
.Y(n_1692)
);

BUFx12f_ASAP7_75t_L g1693 ( 
.A(n_1529),
.Y(n_1693)
);

INVx6_ASAP7_75t_L g1694 ( 
.A(n_1466),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1545),
.B(n_878),
.Y(n_1695)
);

BUFx10_ASAP7_75t_L g1696 ( 
.A(n_1533),
.Y(n_1696)
);

AOI22xp33_ASAP7_75t_L g1697 ( 
.A1(n_1549),
.A2(n_1456),
.B1(n_1473),
.B2(n_1467),
.Y(n_1697)
);

AOI22xp33_ASAP7_75t_SL g1698 ( 
.A1(n_1456),
.A2(n_1473),
.B1(n_1090),
.B2(n_1072),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1465),
.Y(n_1699)
);

CKINVDCx5p33_ASAP7_75t_R g1700 ( 
.A(n_1533),
.Y(n_1700)
);

CKINVDCx6p67_ASAP7_75t_R g1701 ( 
.A(n_1529),
.Y(n_1701)
);

AOI22xp33_ASAP7_75t_L g1702 ( 
.A1(n_1549),
.A2(n_1456),
.B1(n_1473),
.B2(n_1467),
.Y(n_1702)
);

CKINVDCx20_ASAP7_75t_R g1703 ( 
.A(n_1529),
.Y(n_1703)
);

OAI22xp5_ASAP7_75t_L g1704 ( 
.A1(n_1549),
.A2(n_878),
.B1(n_860),
.B2(n_869),
.Y(n_1704)
);

HB1xp67_ASAP7_75t_L g1705 ( 
.A(n_1524),
.Y(n_1705)
);

INVx4_ASAP7_75t_L g1706 ( 
.A(n_1466),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1545),
.B(n_878),
.Y(n_1707)
);

AOI22xp33_ASAP7_75t_L g1708 ( 
.A1(n_1549),
.A2(n_1456),
.B1(n_1473),
.B2(n_1467),
.Y(n_1708)
);

INVx1_ASAP7_75t_SL g1709 ( 
.A(n_1447),
.Y(n_1709)
);

CKINVDCx6p67_ASAP7_75t_R g1710 ( 
.A(n_1529),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1465),
.Y(n_1711)
);

AOI22xp5_ASAP7_75t_L g1712 ( 
.A1(n_1457),
.A2(n_860),
.B1(n_869),
.B2(n_861),
.Y(n_1712)
);

AOI22xp33_ASAP7_75t_SL g1713 ( 
.A1(n_1456),
.A2(n_1473),
.B1(n_1090),
.B2(n_1072),
.Y(n_1713)
);

AOI22xp5_ASAP7_75t_L g1714 ( 
.A1(n_1457),
.A2(n_860),
.B1(n_869),
.B2(n_861),
.Y(n_1714)
);

AOI22xp33_ASAP7_75t_SL g1715 ( 
.A1(n_1456),
.A2(n_1473),
.B1(n_1090),
.B2(n_1072),
.Y(n_1715)
);

AOI22xp33_ASAP7_75t_L g1716 ( 
.A1(n_1549),
.A2(n_1456),
.B1(n_1473),
.B2(n_1467),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1545),
.B(n_878),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1528),
.B(n_1545),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1545),
.B(n_878),
.Y(n_1719)
);

INVx2_ASAP7_75t_L g1720 ( 
.A(n_1465),
.Y(n_1720)
);

OAI21xp5_ASAP7_75t_SL g1721 ( 
.A1(n_1549),
.A2(n_860),
.B(n_1457),
.Y(n_1721)
);

BUFx4f_ASAP7_75t_L g1722 ( 
.A(n_1535),
.Y(n_1722)
);

OAI21xp33_ASAP7_75t_L g1723 ( 
.A1(n_1549),
.A2(n_878),
.B(n_860),
.Y(n_1723)
);

INVx5_ASAP7_75t_L g1724 ( 
.A(n_1515),
.Y(n_1724)
);

AOI22x1_ASAP7_75t_SL g1725 ( 
.A1(n_1474),
.A2(n_769),
.B1(n_1352),
.B2(n_1353),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1422),
.Y(n_1726)
);

OAI22xp5_ASAP7_75t_L g1727 ( 
.A1(n_1549),
.A2(n_878),
.B1(n_860),
.B2(n_869),
.Y(n_1727)
);

AOI22xp33_ASAP7_75t_L g1728 ( 
.A1(n_1549),
.A2(n_1456),
.B1(n_1473),
.B2(n_1467),
.Y(n_1728)
);

BUFx2_ASAP7_75t_L g1729 ( 
.A(n_1447),
.Y(n_1729)
);

INVx6_ASAP7_75t_L g1730 ( 
.A(n_1466),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1465),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1422),
.Y(n_1732)
);

BUFx6f_ASAP7_75t_L g1733 ( 
.A(n_1515),
.Y(n_1733)
);

OR2x2_ASAP7_75t_L g1734 ( 
.A(n_1534),
.B(n_1536),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1422),
.Y(n_1735)
);

INVx3_ASAP7_75t_L g1736 ( 
.A(n_1466),
.Y(n_1736)
);

INVx6_ASAP7_75t_L g1737 ( 
.A(n_1466),
.Y(n_1737)
);

OAI22xp33_ASAP7_75t_L g1738 ( 
.A1(n_1456),
.A2(n_1473),
.B1(n_1549),
.B2(n_1090),
.Y(n_1738)
);

BUFx2_ASAP7_75t_L g1739 ( 
.A(n_1447),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1528),
.B(n_1545),
.Y(n_1740)
);

INVx4_ASAP7_75t_L g1741 ( 
.A(n_1466),
.Y(n_1741)
);

BUFx4f_ASAP7_75t_SL g1742 ( 
.A(n_1407),
.Y(n_1742)
);

BUFx2_ASAP7_75t_L g1743 ( 
.A(n_1665),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1642),
.Y(n_1744)
);

OR2x2_ASAP7_75t_L g1745 ( 
.A(n_1658),
.B(n_1663),
.Y(n_1745)
);

INVx2_ASAP7_75t_L g1746 ( 
.A(n_1674),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_1678),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1643),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1648),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1641),
.Y(n_1750)
);

NOR2xp33_ASAP7_75t_L g1751 ( 
.A(n_1712),
.B(n_1714),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1661),
.Y(n_1752)
);

AO21x2_ASAP7_75t_L g1753 ( 
.A1(n_1645),
.A2(n_1654),
.B(n_1652),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_1641),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1734),
.B(n_1590),
.Y(n_1755)
);

INVx2_ASAP7_75t_L g1756 ( 
.A(n_1630),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1659),
.B(n_1705),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1638),
.Y(n_1758)
);

BUFx3_ASAP7_75t_L g1759 ( 
.A(n_1640),
.Y(n_1759)
);

OA21x2_ASAP7_75t_L g1760 ( 
.A1(n_1650),
.A2(n_1651),
.B(n_1601),
.Y(n_1760)
);

BUFx2_ASAP7_75t_L g1761 ( 
.A(n_1653),
.Y(n_1761)
);

BUFx6f_ASAP7_75t_L g1762 ( 
.A(n_1673),
.Y(n_1762)
);

OAI21x1_ASAP7_75t_L g1763 ( 
.A1(n_1633),
.A2(n_1667),
.B(n_1669),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1705),
.B(n_1638),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_1631),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1677),
.B(n_1575),
.Y(n_1766)
);

HB1xp67_ASAP7_75t_L g1767 ( 
.A(n_1583),
.Y(n_1767)
);

BUFx3_ASAP7_75t_L g1768 ( 
.A(n_1640),
.Y(n_1768)
);

HB1xp67_ASAP7_75t_L g1769 ( 
.A(n_1617),
.Y(n_1769)
);

INVx3_ASAP7_75t_L g1770 ( 
.A(n_1670),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1671),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1656),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1656),
.Y(n_1773)
);

INVxp67_ASAP7_75t_SL g1774 ( 
.A(n_1587),
.Y(n_1774)
);

HB1xp67_ASAP7_75t_L g1775 ( 
.A(n_1585),
.Y(n_1775)
);

OAI22xp5_ASAP7_75t_L g1776 ( 
.A1(n_1687),
.A2(n_1715),
.B1(n_1698),
.B2(n_1713),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1656),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1656),
.Y(n_1778)
);

OR2x2_ASAP7_75t_L g1779 ( 
.A(n_1673),
.B(n_1657),
.Y(n_1779)
);

OA21x2_ASAP7_75t_L g1780 ( 
.A1(n_1601),
.A2(n_1629),
.B(n_1569),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1668),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1557),
.B(n_1695),
.Y(n_1782)
);

OA21x2_ASAP7_75t_L g1783 ( 
.A1(n_1629),
.A2(n_1579),
.B(n_1570),
.Y(n_1783)
);

BUFx3_ASAP7_75t_L g1784 ( 
.A(n_1640),
.Y(n_1784)
);

OAI21x1_ASAP7_75t_L g1785 ( 
.A1(n_1644),
.A2(n_1620),
.B(n_1616),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1676),
.Y(n_1786)
);

OR2x6_ASAP7_75t_L g1787 ( 
.A(n_1655),
.B(n_1647),
.Y(n_1787)
);

BUFx3_ASAP7_75t_L g1788 ( 
.A(n_1634),
.Y(n_1788)
);

AO21x2_ASAP7_75t_L g1789 ( 
.A1(n_1664),
.A2(n_1738),
.B(n_1689),
.Y(n_1789)
);

INVx2_ASAP7_75t_SL g1790 ( 
.A(n_1634),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1672),
.Y(n_1791)
);

AND2x4_ASAP7_75t_L g1792 ( 
.A(n_1685),
.B(n_1724),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_1666),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_1593),
.Y(n_1794)
);

HB1xp67_ASAP7_75t_L g1795 ( 
.A(n_1586),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1726),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1732),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1735),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1612),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1677),
.B(n_1575),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1612),
.B(n_1625),
.Y(n_1801)
);

INVxp67_ASAP7_75t_L g1802 ( 
.A(n_1729),
.Y(n_1802)
);

INVx2_ASAP7_75t_L g1803 ( 
.A(n_1626),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1625),
.B(n_1579),
.Y(n_1804)
);

AND2x4_ASAP7_75t_L g1805 ( 
.A(n_1685),
.B(n_1724),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1573),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1627),
.B(n_1588),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1664),
.Y(n_1808)
);

INVxp33_ASAP7_75t_L g1809 ( 
.A(n_1691),
.Y(n_1809)
);

AND2x4_ASAP7_75t_L g1810 ( 
.A(n_1685),
.B(n_1724),
.Y(n_1810)
);

INVx2_ASAP7_75t_L g1811 ( 
.A(n_1622),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1675),
.Y(n_1812)
);

AO21x1_ASAP7_75t_SL g1813 ( 
.A1(n_1565),
.A2(n_1716),
.B(n_1708),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1675),
.Y(n_1814)
);

HB1xp67_ASAP7_75t_SL g1815 ( 
.A(n_1561),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1627),
.B(n_1570),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1632),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1632),
.Y(n_1818)
);

INVx4_ASAP7_75t_SL g1819 ( 
.A(n_1577),
.Y(n_1819)
);

INVx2_ASAP7_75t_SL g1820 ( 
.A(n_1634),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1699),
.Y(n_1821)
);

OAI211xp5_ASAP7_75t_SL g1822 ( 
.A1(n_1721),
.A2(n_1723),
.B(n_1704),
.C(n_1727),
.Y(n_1822)
);

INVxp67_ASAP7_75t_SL g1823 ( 
.A(n_1621),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1711),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1720),
.Y(n_1825)
);

CKINVDCx5p33_ASAP7_75t_R g1826 ( 
.A(n_1684),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1731),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1660),
.Y(n_1828)
);

AND2x4_ASAP7_75t_L g1829 ( 
.A(n_1724),
.B(n_1634),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1660),
.Y(n_1830)
);

AO21x2_ASAP7_75t_L g1831 ( 
.A1(n_1689),
.A2(n_1738),
.B(n_1662),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1609),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1609),
.Y(n_1833)
);

INVx3_ASAP7_75t_L g1834 ( 
.A(n_1646),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1589),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1589),
.Y(n_1836)
);

INVx2_ASAP7_75t_L g1837 ( 
.A(n_1639),
.Y(n_1837)
);

INVx2_ASAP7_75t_L g1838 ( 
.A(n_1614),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1603),
.Y(n_1839)
);

INVx2_ASAP7_75t_L g1840 ( 
.A(n_1594),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1595),
.Y(n_1841)
);

AO21x2_ASAP7_75t_L g1842 ( 
.A1(n_1613),
.A2(n_1637),
.B(n_1576),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1595),
.Y(n_1843)
);

AND2x4_ASAP7_75t_L g1844 ( 
.A(n_1606),
.B(n_1594),
.Y(n_1844)
);

INVx3_ASAP7_75t_L g1845 ( 
.A(n_1562),
.Y(n_1845)
);

NOR2xp33_ASAP7_75t_L g1846 ( 
.A(n_1555),
.B(n_1707),
.Y(n_1846)
);

INVx2_ASAP7_75t_L g1847 ( 
.A(n_1733),
.Y(n_1847)
);

OAI21xp5_ASAP7_75t_L g1848 ( 
.A1(n_1687),
.A2(n_1698),
.B(n_1713),
.Y(n_1848)
);

HB1xp67_ASAP7_75t_L g1849 ( 
.A(n_1739),
.Y(n_1849)
);

AOI21x1_ASAP7_75t_L g1850 ( 
.A1(n_1581),
.A2(n_1584),
.B(n_1717),
.Y(n_1850)
);

OAI22xp5_ASAP7_75t_SL g1851 ( 
.A1(n_1715),
.A2(n_1566),
.B1(n_1680),
.B2(n_1697),
.Y(n_1851)
);

OAI21x1_ASAP7_75t_L g1852 ( 
.A1(n_1563),
.A2(n_1600),
.B(n_1736),
.Y(n_1852)
);

HB1xp67_ASAP7_75t_L g1853 ( 
.A(n_1679),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1567),
.Y(n_1854)
);

O2A1O1Ixp5_ASAP7_75t_L g1855 ( 
.A1(n_1719),
.A2(n_1580),
.B(n_1741),
.C(n_1706),
.Y(n_1855)
);

INVx2_ASAP7_75t_L g1856 ( 
.A(n_1733),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1567),
.Y(n_1857)
);

INVx3_ASAP7_75t_L g1858 ( 
.A(n_1562),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1566),
.Y(n_1859)
);

INVx3_ASAP7_75t_L g1860 ( 
.A(n_1580),
.Y(n_1860)
);

OAI21x1_ASAP7_75t_L g1861 ( 
.A1(n_1563),
.A2(n_1600),
.B(n_1736),
.Y(n_1861)
);

AND2x2_ASAP7_75t_L g1862 ( 
.A(n_1718),
.B(n_1740),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1606),
.Y(n_1863)
);

INVx4_ASAP7_75t_SL g1864 ( 
.A(n_1577),
.Y(n_1864)
);

AOI22xp33_ASAP7_75t_L g1865 ( 
.A1(n_1565),
.A2(n_1708),
.B1(n_1702),
.B2(n_1728),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1577),
.Y(n_1866)
);

OR2x2_ASAP7_75t_L g1867 ( 
.A(n_1680),
.B(n_1702),
.Y(n_1867)
);

BUFx12f_ASAP7_75t_L g1868 ( 
.A(n_1683),
.Y(n_1868)
);

INVx2_ASAP7_75t_L g1869 ( 
.A(n_1602),
.Y(n_1869)
);

BUFx6f_ASAP7_75t_L g1870 ( 
.A(n_1649),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1602),
.Y(n_1871)
);

BUFx2_ASAP7_75t_SL g1872 ( 
.A(n_1628),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1602),
.Y(n_1873)
);

OAI21x1_ASAP7_75t_L g1874 ( 
.A1(n_1681),
.A2(n_1686),
.B(n_1697),
.Y(n_1874)
);

AND2x4_ASAP7_75t_L g1875 ( 
.A(n_1706),
.B(n_1741),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1692),
.Y(n_1876)
);

INVx3_ASAP7_75t_L g1877 ( 
.A(n_1692),
.Y(n_1877)
);

INVx2_ASAP7_75t_L g1878 ( 
.A(n_1692),
.Y(n_1878)
);

INVx2_ASAP7_75t_L g1879 ( 
.A(n_1694),
.Y(n_1879)
);

HB1xp67_ASAP7_75t_L g1880 ( 
.A(n_1679),
.Y(n_1880)
);

NOR2xp33_ASAP7_75t_L g1881 ( 
.A(n_1571),
.B(n_1709),
.Y(n_1881)
);

AOI22xp33_ASAP7_75t_L g1882 ( 
.A1(n_1681),
.A2(n_1728),
.B1(n_1682),
.B2(n_1686),
.Y(n_1882)
);

AND2x2_ASAP7_75t_L g1883 ( 
.A(n_1682),
.B(n_1716),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1694),
.Y(n_1884)
);

INVx2_ASAP7_75t_L g1885 ( 
.A(n_1730),
.Y(n_1885)
);

OAI21x1_ASAP7_75t_L g1886 ( 
.A1(n_1578),
.A2(n_1591),
.B(n_1568),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1730),
.Y(n_1887)
);

OR2x2_ASAP7_75t_L g1888 ( 
.A(n_1690),
.B(n_1558),
.Y(n_1888)
);

INVx2_ASAP7_75t_L g1889 ( 
.A(n_1730),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1737),
.Y(n_1890)
);

NOR4xp25_ASAP7_75t_SL g1891 ( 
.A(n_1582),
.B(n_1700),
.C(n_1560),
.D(n_1596),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1737),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1737),
.Y(n_1893)
);

AO32x1_ASAP7_75t_L g1894 ( 
.A1(n_1776),
.A2(n_1574),
.A3(n_1618),
.B1(n_1578),
.B2(n_1556),
.Y(n_1894)
);

AOI22xp33_ASAP7_75t_L g1895 ( 
.A1(n_1751),
.A2(n_1598),
.B1(n_1710),
.B2(n_1701),
.Y(n_1895)
);

O2A1O1Ixp33_ASAP7_75t_SL g1896 ( 
.A1(n_1848),
.A2(n_1605),
.B(n_1703),
.C(n_1559),
.Y(n_1896)
);

O2A1O1Ixp33_ASAP7_75t_SL g1897 ( 
.A1(n_1822),
.A2(n_1867),
.B(n_1857),
.C(n_1854),
.Y(n_1897)
);

AND2x2_ASAP7_75t_L g1898 ( 
.A(n_1862),
.B(n_1608),
.Y(n_1898)
);

NOR2x1p5_ASAP7_75t_L g1899 ( 
.A(n_1868),
.B(n_1688),
.Y(n_1899)
);

A2O1A1Ixp33_ASAP7_75t_L g1900 ( 
.A1(n_1874),
.A2(n_1722),
.B(n_1572),
.C(n_1624),
.Y(n_1900)
);

HB1xp67_ASAP7_75t_L g1901 ( 
.A(n_1758),
.Y(n_1901)
);

AND2x4_ASAP7_75t_L g1902 ( 
.A(n_1770),
.B(n_1624),
.Y(n_1902)
);

OR2x2_ASAP7_75t_L g1903 ( 
.A(n_1757),
.B(n_1604),
.Y(n_1903)
);

OR2x2_ASAP7_75t_L g1904 ( 
.A(n_1757),
.B(n_1608),
.Y(n_1904)
);

OR2x2_ASAP7_75t_L g1905 ( 
.A(n_1755),
.B(n_1572),
.Y(n_1905)
);

AND2x4_ASAP7_75t_L g1906 ( 
.A(n_1770),
.B(n_1636),
.Y(n_1906)
);

AND2x2_ASAP7_75t_L g1907 ( 
.A(n_1862),
.B(n_1615),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1806),
.B(n_1619),
.Y(n_1908)
);

NOR2xp33_ASAP7_75t_L g1909 ( 
.A(n_1842),
.B(n_1619),
.Y(n_1909)
);

NOR2x1_ASAP7_75t_SL g1910 ( 
.A(n_1787),
.B(n_1693),
.Y(n_1910)
);

AND2x4_ASAP7_75t_L g1911 ( 
.A(n_1770),
.B(n_1599),
.Y(n_1911)
);

OR2x2_ASAP7_75t_L g1912 ( 
.A(n_1745),
.B(n_1696),
.Y(n_1912)
);

OR2x2_ASAP7_75t_L g1913 ( 
.A(n_1745),
.B(n_1771),
.Y(n_1913)
);

AND2x2_ASAP7_75t_L g1914 ( 
.A(n_1761),
.B(n_1837),
.Y(n_1914)
);

AO32x1_ASAP7_75t_L g1915 ( 
.A1(n_1816),
.A2(n_1883),
.A3(n_1800),
.B1(n_1766),
.B2(n_1804),
.Y(n_1915)
);

AND2x2_ASAP7_75t_L g1916 ( 
.A(n_1761),
.B(n_1635),
.Y(n_1916)
);

NOR2xp33_ASAP7_75t_L g1917 ( 
.A(n_1842),
.B(n_1610),
.Y(n_1917)
);

A2O1A1Ixp33_ASAP7_75t_L g1918 ( 
.A1(n_1874),
.A2(n_1722),
.B(n_1725),
.C(n_1623),
.Y(n_1918)
);

AOI221xp5_ASAP7_75t_L g1919 ( 
.A1(n_1851),
.A2(n_1564),
.B1(n_1592),
.B2(n_1561),
.C(n_1597),
.Y(n_1919)
);

AND2x2_ASAP7_75t_L g1920 ( 
.A(n_1837),
.B(n_1607),
.Y(n_1920)
);

AND2x2_ASAP7_75t_L g1921 ( 
.A(n_1809),
.B(n_1696),
.Y(n_1921)
);

AND2x2_ASAP7_75t_L g1922 ( 
.A(n_1853),
.B(n_1610),
.Y(n_1922)
);

CKINVDCx16_ASAP7_75t_R g1923 ( 
.A(n_1815),
.Y(n_1923)
);

AND2x4_ASAP7_75t_L g1924 ( 
.A(n_1770),
.B(n_1564),
.Y(n_1924)
);

NOR2x1_ASAP7_75t_SL g1925 ( 
.A(n_1787),
.B(n_1742),
.Y(n_1925)
);

A2O1A1Ixp33_ASAP7_75t_L g1926 ( 
.A1(n_1865),
.A2(n_1592),
.B(n_1611),
.C(n_1742),
.Y(n_1926)
);

AND2x2_ASAP7_75t_L g1927 ( 
.A(n_1880),
.B(n_1619),
.Y(n_1927)
);

AND2x2_ASAP7_75t_L g1928 ( 
.A(n_1766),
.B(n_1800),
.Y(n_1928)
);

AOI21xp5_ASAP7_75t_L g1929 ( 
.A1(n_1753),
.A2(n_1787),
.B(n_1780),
.Y(n_1929)
);

OAI21xp5_ASAP7_75t_L g1930 ( 
.A1(n_1882),
.A2(n_1806),
.B(n_1835),
.Y(n_1930)
);

A2O1A1Ixp33_ASAP7_75t_L g1931 ( 
.A1(n_1867),
.A2(n_1883),
.B(n_1886),
.C(n_1854),
.Y(n_1931)
);

AND2x2_ASAP7_75t_L g1932 ( 
.A(n_1807),
.B(n_1838),
.Y(n_1932)
);

AOI22xp5_ASAP7_75t_L g1933 ( 
.A1(n_1842),
.A2(n_1857),
.B1(n_1789),
.B2(n_1859),
.Y(n_1933)
);

INVx4_ASAP7_75t_L g1934 ( 
.A(n_1877),
.Y(n_1934)
);

INVx2_ASAP7_75t_SL g1935 ( 
.A(n_1767),
.Y(n_1935)
);

OA21x2_ASAP7_75t_L g1936 ( 
.A1(n_1763),
.A2(n_1785),
.B(n_1817),
.Y(n_1936)
);

AO32x2_ASAP7_75t_L g1937 ( 
.A1(n_1790),
.A2(n_1820),
.A3(n_1801),
.B1(n_1799),
.B2(n_1816),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1774),
.B(n_1799),
.Y(n_1938)
);

NAND2xp33_ASAP7_75t_L g1939 ( 
.A(n_1870),
.B(n_1826),
.Y(n_1939)
);

OR2x6_ASAP7_75t_L g1940 ( 
.A(n_1787),
.B(n_1743),
.Y(n_1940)
);

AND2x2_ASAP7_75t_L g1941 ( 
.A(n_1847),
.B(n_1856),
.Y(n_1941)
);

AND2x2_ASAP7_75t_L g1942 ( 
.A(n_1769),
.B(n_1859),
.Y(n_1942)
);

INVx3_ASAP7_75t_L g1943 ( 
.A(n_1844),
.Y(n_1943)
);

OAI22xp5_ASAP7_75t_L g1944 ( 
.A1(n_1870),
.A2(n_1804),
.B1(n_1782),
.B2(n_1846),
.Y(n_1944)
);

BUFx4f_ASAP7_75t_L g1945 ( 
.A(n_1868),
.Y(n_1945)
);

AND2x2_ASAP7_75t_L g1946 ( 
.A(n_1743),
.B(n_1795),
.Y(n_1946)
);

OA21x2_ASAP7_75t_L g1947 ( 
.A1(n_1817),
.A2(n_1818),
.B(n_1808),
.Y(n_1947)
);

OR2x6_ASAP7_75t_L g1948 ( 
.A(n_1787),
.B(n_1792),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1863),
.B(n_1886),
.Y(n_1949)
);

O2A1O1Ixp33_ASAP7_75t_L g1950 ( 
.A1(n_1839),
.A2(n_1836),
.B(n_1835),
.C(n_1789),
.Y(n_1950)
);

O2A1O1Ixp33_ASAP7_75t_SL g1951 ( 
.A1(n_1839),
.A2(n_1841),
.B(n_1843),
.C(n_1836),
.Y(n_1951)
);

AOI22xp5_ASAP7_75t_L g1952 ( 
.A1(n_1789),
.A2(n_1831),
.B1(n_1881),
.B2(n_1833),
.Y(n_1952)
);

AOI22xp5_ASAP7_75t_L g1953 ( 
.A1(n_1831),
.A2(n_1833),
.B1(n_1832),
.B2(n_1870),
.Y(n_1953)
);

AOI22xp5_ASAP7_75t_L g1954 ( 
.A1(n_1831),
.A2(n_1832),
.B1(n_1870),
.B2(n_1844),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1811),
.B(n_1765),
.Y(n_1955)
);

AO32x2_ASAP7_75t_L g1956 ( 
.A1(n_1790),
.A2(n_1820),
.A3(n_1801),
.B1(n_1843),
.B2(n_1841),
.Y(n_1956)
);

NAND4xp25_ASAP7_75t_L g1957 ( 
.A(n_1888),
.B(n_1802),
.C(n_1855),
.D(n_1808),
.Y(n_1957)
);

OA21x2_ASAP7_75t_L g1958 ( 
.A1(n_1818),
.A2(n_1812),
.B(n_1814),
.Y(n_1958)
);

HB1xp67_ASAP7_75t_L g1959 ( 
.A(n_1758),
.Y(n_1959)
);

AND2x2_ASAP7_75t_L g1960 ( 
.A(n_1840),
.B(n_1775),
.Y(n_1960)
);

NOR2xp33_ASAP7_75t_L g1961 ( 
.A(n_1850),
.B(n_1849),
.Y(n_1961)
);

AOI221xp5_ASAP7_75t_L g1962 ( 
.A1(n_1828),
.A2(n_1830),
.B1(n_1870),
.B2(n_1814),
.C(n_1812),
.Y(n_1962)
);

AND2x4_ASAP7_75t_L g1963 ( 
.A(n_1844),
.B(n_1759),
.Y(n_1963)
);

OA21x2_ASAP7_75t_L g1964 ( 
.A1(n_1828),
.A2(n_1830),
.B(n_1752),
.Y(n_1964)
);

CKINVDCx20_ASAP7_75t_R g1965 ( 
.A(n_1872),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1796),
.Y(n_1966)
);

AND2x4_ASAP7_75t_L g1967 ( 
.A(n_1759),
.B(n_1768),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1797),
.Y(n_1968)
);

HB1xp67_ASAP7_75t_L g1969 ( 
.A(n_1752),
.Y(n_1969)
);

AO32x2_ASAP7_75t_L g1970 ( 
.A1(n_1771),
.A2(n_1772),
.A3(n_1773),
.B1(n_1777),
.B2(n_1778),
.Y(n_1970)
);

OAI21x1_ASAP7_75t_L g1971 ( 
.A1(n_1852),
.A2(n_1861),
.B(n_1834),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1797),
.Y(n_1972)
);

NOR2x1_ASAP7_75t_SL g1973 ( 
.A(n_1850),
.B(n_1753),
.Y(n_1973)
);

OR2x6_ASAP7_75t_L g1974 ( 
.A(n_1792),
.B(n_1805),
.Y(n_1974)
);

INVx4_ASAP7_75t_L g1975 ( 
.A(n_1877),
.Y(n_1975)
);

AND2x6_ASAP7_75t_L g1976 ( 
.A(n_1792),
.B(n_1805),
.Y(n_1976)
);

NOR2xp33_ASAP7_75t_L g1977 ( 
.A(n_1888),
.B(n_1768),
.Y(n_1977)
);

AND2x2_ASAP7_75t_L g1978 ( 
.A(n_1794),
.B(n_1803),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_L g1979 ( 
.A(n_1811),
.B(n_1765),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_L g1980 ( 
.A(n_1811),
.B(n_1764),
.Y(n_1980)
);

NOR2x1_ASAP7_75t_SL g1981 ( 
.A(n_1753),
.B(n_1788),
.Y(n_1981)
);

AOI22xp5_ASAP7_75t_L g1982 ( 
.A1(n_1870),
.A2(n_1783),
.B1(n_1872),
.B2(n_1890),
.Y(n_1982)
);

NOR2xp33_ASAP7_75t_L g1983 ( 
.A(n_1768),
.B(n_1784),
.Y(n_1983)
);

OR2x6_ASAP7_75t_L g1984 ( 
.A(n_1792),
.B(n_1805),
.Y(n_1984)
);

OR2x2_ASAP7_75t_L g1985 ( 
.A(n_1803),
.B(n_1798),
.Y(n_1985)
);

CKINVDCx5p33_ASAP7_75t_R g1986 ( 
.A(n_1891),
.Y(n_1986)
);

NOR2xp33_ASAP7_75t_L g1987 ( 
.A(n_1784),
.B(n_1877),
.Y(n_1987)
);

NOR2xp33_ASAP7_75t_L g1988 ( 
.A(n_1877),
.B(n_1869),
.Y(n_1988)
);

OR2x6_ASAP7_75t_L g1989 ( 
.A(n_1805),
.B(n_1810),
.Y(n_1989)
);

AO32x2_ASAP7_75t_L g1990 ( 
.A1(n_1772),
.A2(n_1773),
.A3(n_1777),
.B1(n_1778),
.B2(n_1783),
.Y(n_1990)
);

INVx4_ASAP7_75t_L g1991 ( 
.A(n_1819),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_L g1992 ( 
.A(n_1798),
.B(n_1756),
.Y(n_1992)
);

AOI22xp33_ASAP7_75t_L g1993 ( 
.A1(n_1919),
.A2(n_1813),
.B1(n_1944),
.B2(n_1986),
.Y(n_1993)
);

AOI22xp33_ASAP7_75t_L g1994 ( 
.A1(n_1919),
.A2(n_1813),
.B1(n_1783),
.B2(n_1780),
.Y(n_1994)
);

HB1xp67_ASAP7_75t_L g1995 ( 
.A(n_1964),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1969),
.Y(n_1996)
);

AND2x4_ASAP7_75t_SL g1997 ( 
.A(n_1948),
.B(n_1829),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_L g1998 ( 
.A(n_1961),
.B(n_1744),
.Y(n_1998)
);

NOR2x1_ASAP7_75t_SL g1999 ( 
.A(n_1940),
.B(n_1762),
.Y(n_1999)
);

AOI22xp5_ASAP7_75t_L g2000 ( 
.A1(n_1944),
.A2(n_1783),
.B1(n_1780),
.B2(n_1760),
.Y(n_2000)
);

INVxp67_ASAP7_75t_SL g2001 ( 
.A(n_1901),
.Y(n_2001)
);

AND2x2_ASAP7_75t_L g2002 ( 
.A(n_1936),
.B(n_1990),
.Y(n_2002)
);

AND2x2_ASAP7_75t_L g2003 ( 
.A(n_1936),
.B(n_1760),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1901),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_L g2005 ( 
.A(n_1961),
.B(n_1744),
.Y(n_2005)
);

AOI22xp33_ASAP7_75t_SL g2006 ( 
.A1(n_1928),
.A2(n_1780),
.B1(n_1760),
.B2(n_1810),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1959),
.Y(n_2007)
);

OR2x2_ASAP7_75t_L g2008 ( 
.A(n_1980),
.B(n_1779),
.Y(n_2008)
);

HB1xp67_ASAP7_75t_L g2009 ( 
.A(n_1964),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1959),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_L g2011 ( 
.A(n_1952),
.B(n_1748),
.Y(n_2011)
);

OR2x2_ASAP7_75t_L g2012 ( 
.A(n_1980),
.B(n_1779),
.Y(n_2012)
);

AND2x2_ASAP7_75t_L g2013 ( 
.A(n_1990),
.B(n_1760),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_L g2014 ( 
.A(n_1958),
.B(n_1748),
.Y(n_2014)
);

INVx2_ASAP7_75t_L g2015 ( 
.A(n_1978),
.Y(n_2015)
);

AND2x2_ASAP7_75t_L g2016 ( 
.A(n_1990),
.B(n_1746),
.Y(n_2016)
);

HB1xp67_ASAP7_75t_L g2017 ( 
.A(n_1947),
.Y(n_2017)
);

AOI22xp33_ASAP7_75t_L g2018 ( 
.A1(n_1930),
.A2(n_1878),
.B1(n_1879),
.B2(n_1869),
.Y(n_2018)
);

BUFx3_ASAP7_75t_L g2019 ( 
.A(n_1976),
.Y(n_2019)
);

INVx2_ASAP7_75t_L g2020 ( 
.A(n_1966),
.Y(n_2020)
);

INVx2_ASAP7_75t_L g2021 ( 
.A(n_1968),
.Y(n_2021)
);

OR2x2_ASAP7_75t_L g2022 ( 
.A(n_1913),
.B(n_1938),
.Y(n_2022)
);

INVx2_ASAP7_75t_L g2023 ( 
.A(n_1972),
.Y(n_2023)
);

HB1xp67_ASAP7_75t_L g2024 ( 
.A(n_1947),
.Y(n_2024)
);

AOI22xp5_ASAP7_75t_L g2025 ( 
.A1(n_1897),
.A2(n_1896),
.B1(n_1933),
.B2(n_1930),
.Y(n_2025)
);

HB1xp67_ASAP7_75t_L g2026 ( 
.A(n_1958),
.Y(n_2026)
);

AND2x2_ASAP7_75t_L g2027 ( 
.A(n_1932),
.B(n_1949),
.Y(n_2027)
);

AND2x4_ASAP7_75t_L g2028 ( 
.A(n_1948),
.B(n_1781),
.Y(n_2028)
);

INVx2_ASAP7_75t_SL g2029 ( 
.A(n_1974),
.Y(n_2029)
);

INVx2_ASAP7_75t_SL g2030 ( 
.A(n_1974),
.Y(n_2030)
);

BUFx2_ASAP7_75t_SL g2031 ( 
.A(n_1965),
.Y(n_2031)
);

AND2x2_ASAP7_75t_L g2032 ( 
.A(n_1970),
.B(n_1747),
.Y(n_2032)
);

INVx8_ASAP7_75t_L g2033 ( 
.A(n_1906),
.Y(n_2033)
);

AND2x2_ASAP7_75t_L g2034 ( 
.A(n_1970),
.B(n_1750),
.Y(n_2034)
);

AND2x2_ASAP7_75t_L g2035 ( 
.A(n_1937),
.B(n_1781),
.Y(n_2035)
);

AND2x2_ASAP7_75t_L g2036 ( 
.A(n_1937),
.B(n_1762),
.Y(n_2036)
);

AND2x2_ASAP7_75t_L g2037 ( 
.A(n_1937),
.B(n_1762),
.Y(n_2037)
);

INVxp67_ASAP7_75t_L g2038 ( 
.A(n_1909),
.Y(n_2038)
);

NAND2xp5_ASAP7_75t_L g2039 ( 
.A(n_1950),
.B(n_1749),
.Y(n_2039)
);

AND2x2_ASAP7_75t_L g2040 ( 
.A(n_1941),
.B(n_1762),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1985),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_L g2042 ( 
.A(n_1950),
.B(n_1793),
.Y(n_2042)
);

AND2x2_ASAP7_75t_L g2043 ( 
.A(n_1914),
.B(n_1762),
.Y(n_2043)
);

OAI22xp5_ASAP7_75t_L g2044 ( 
.A1(n_1962),
.A2(n_1931),
.B1(n_1953),
.B2(n_1926),
.Y(n_2044)
);

NOR2xp33_ASAP7_75t_L g2045 ( 
.A(n_1912),
.B(n_1866),
.Y(n_2045)
);

HB1xp67_ASAP7_75t_L g2046 ( 
.A(n_1955),
.Y(n_2046)
);

INVx2_ASAP7_75t_L g2047 ( 
.A(n_1971),
.Y(n_2047)
);

BUFx6f_ASAP7_75t_L g2048 ( 
.A(n_1948),
.Y(n_2048)
);

OR2x2_ASAP7_75t_L g2049 ( 
.A(n_1955),
.B(n_1979),
.Y(n_2049)
);

AND2x2_ASAP7_75t_L g2050 ( 
.A(n_1929),
.B(n_1754),
.Y(n_2050)
);

AND2x2_ASAP7_75t_L g2051 ( 
.A(n_1956),
.B(n_1762),
.Y(n_2051)
);

OAI22xp5_ASAP7_75t_L g2052 ( 
.A1(n_1962),
.A2(n_1756),
.B1(n_1823),
.B2(n_1825),
.Y(n_2052)
);

AOI221xp5_ASAP7_75t_L g2053 ( 
.A1(n_2044),
.A2(n_1897),
.B1(n_2011),
.B2(n_2025),
.C(n_1896),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_2020),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_2020),
.Y(n_2055)
);

OR2x2_ASAP7_75t_L g2056 ( 
.A(n_2038),
.B(n_2022),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_2020),
.Y(n_2057)
);

OAI221xp5_ASAP7_75t_L g2058 ( 
.A1(n_2025),
.A2(n_1918),
.B1(n_1895),
.B2(n_1900),
.C(n_1926),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_2021),
.Y(n_2059)
);

OAI22xp5_ASAP7_75t_SL g2060 ( 
.A1(n_1993),
.A2(n_1923),
.B1(n_1895),
.B2(n_1906),
.Y(n_2060)
);

AOI221xp5_ASAP7_75t_L g2061 ( 
.A1(n_2044),
.A2(n_1957),
.B1(n_1951),
.B2(n_1935),
.C(n_1942),
.Y(n_2061)
);

AND2x2_ASAP7_75t_L g2062 ( 
.A(n_2036),
.B(n_1981),
.Y(n_2062)
);

INVx2_ASAP7_75t_SL g2063 ( 
.A(n_2033),
.Y(n_2063)
);

BUFx2_ASAP7_75t_L g2064 ( 
.A(n_2019),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_2021),
.Y(n_2065)
);

AOI21xp5_ASAP7_75t_L g2066 ( 
.A1(n_2042),
.A2(n_1894),
.B(n_1915),
.Y(n_2066)
);

AND2x4_ASAP7_75t_SL g2067 ( 
.A(n_2028),
.B(n_1991),
.Y(n_2067)
);

NOR2xp33_ASAP7_75t_L g2068 ( 
.A(n_2038),
.B(n_1957),
.Y(n_2068)
);

NAND5xp2_ASAP7_75t_L g2069 ( 
.A(n_1994),
.B(n_1982),
.C(n_1954),
.D(n_1929),
.E(n_1917),
.Y(n_2069)
);

HB1xp67_ASAP7_75t_L g2070 ( 
.A(n_2026),
.Y(n_2070)
);

AND2x2_ASAP7_75t_L g2071 ( 
.A(n_2036),
.B(n_1956),
.Y(n_2071)
);

INVx5_ASAP7_75t_SL g2072 ( 
.A(n_2048),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_2021),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_2023),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_2023),
.Y(n_2075)
);

AND2x4_ASAP7_75t_L g2076 ( 
.A(n_2019),
.B(n_1974),
.Y(n_2076)
);

INVx1_ASAP7_75t_SL g2077 ( 
.A(n_2031),
.Y(n_2077)
);

AOI22xp33_ASAP7_75t_SL g2078 ( 
.A1(n_2031),
.A2(n_1910),
.B1(n_1925),
.B2(n_1894),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_L g2079 ( 
.A(n_2022),
.B(n_1960),
.Y(n_2079)
);

NAND2xp5_ASAP7_75t_L g2080 ( 
.A(n_1998),
.B(n_1909),
.Y(n_2080)
);

AND2x2_ASAP7_75t_L g2081 ( 
.A(n_2037),
.B(n_1956),
.Y(n_2081)
);

AND2x4_ASAP7_75t_L g2082 ( 
.A(n_2019),
.B(n_1984),
.Y(n_2082)
);

OR2x6_ASAP7_75t_L g2083 ( 
.A(n_2048),
.B(n_1940),
.Y(n_2083)
);

AO21x2_ASAP7_75t_L g2084 ( 
.A1(n_2047),
.A2(n_1973),
.B(n_1917),
.Y(n_2084)
);

AND2x4_ASAP7_75t_L g2085 ( 
.A(n_2029),
.B(n_1984),
.Y(n_2085)
);

INVxp67_ASAP7_75t_SL g2086 ( 
.A(n_2017),
.Y(n_2086)
);

AND2x2_ASAP7_75t_L g2087 ( 
.A(n_2037),
.B(n_1946),
.Y(n_2087)
);

AND2x2_ASAP7_75t_L g2088 ( 
.A(n_2027),
.B(n_1984),
.Y(n_2088)
);

AOI22xp5_ASAP7_75t_L g2089 ( 
.A1(n_2029),
.A2(n_1940),
.B1(n_1983),
.B2(n_1977),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_2023),
.Y(n_2090)
);

INVx4_ASAP7_75t_L g2091 ( 
.A(n_2033),
.Y(n_2091)
);

NAND2x1_ASAP7_75t_L g2092 ( 
.A(n_2051),
.B(n_1976),
.Y(n_2092)
);

INVx5_ASAP7_75t_L g2093 ( 
.A(n_2048),
.Y(n_2093)
);

AOI22xp33_ASAP7_75t_L g2094 ( 
.A1(n_2048),
.A2(n_1921),
.B1(n_1977),
.B2(n_1963),
.Y(n_2094)
);

NOR3xp33_ASAP7_75t_L g2095 ( 
.A(n_2042),
.B(n_1908),
.C(n_1876),
.Y(n_2095)
);

NAND2x1p5_ASAP7_75t_L g2096 ( 
.A(n_2048),
.B(n_1991),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_2004),
.Y(n_2097)
);

OR2x2_ASAP7_75t_L g2098 ( 
.A(n_2008),
.B(n_1904),
.Y(n_2098)
);

AND2x2_ASAP7_75t_L g2099 ( 
.A(n_2027),
.B(n_1989),
.Y(n_2099)
);

BUFx3_ASAP7_75t_L g2100 ( 
.A(n_2033),
.Y(n_2100)
);

AND2x2_ASAP7_75t_L g2101 ( 
.A(n_2051),
.B(n_2040),
.Y(n_2101)
);

AO21x2_ASAP7_75t_L g2102 ( 
.A1(n_2047),
.A2(n_1786),
.B(n_1791),
.Y(n_2102)
);

HB1xp67_ASAP7_75t_L g2103 ( 
.A(n_2026),
.Y(n_2103)
);

OAI21xp33_ASAP7_75t_L g2104 ( 
.A1(n_2006),
.A2(n_1908),
.B(n_1988),
.Y(n_2104)
);

INVx2_ASAP7_75t_L g2105 ( 
.A(n_2032),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_2004),
.Y(n_2106)
);

INVxp67_ASAP7_75t_L g2107 ( 
.A(n_2041),
.Y(n_2107)
);

OAI33xp33_ASAP7_75t_L g2108 ( 
.A1(n_2011),
.A2(n_1905),
.A3(n_1992),
.B1(n_1903),
.B2(n_1821),
.B3(n_1827),
.Y(n_2108)
);

AND2x2_ASAP7_75t_L g2109 ( 
.A(n_2040),
.B(n_1989),
.Y(n_2109)
);

AO21x2_ASAP7_75t_L g2110 ( 
.A1(n_2047),
.A2(n_1786),
.B(n_1791),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_2007),
.Y(n_2111)
);

INVx3_ASAP7_75t_L g2112 ( 
.A(n_2048),
.Y(n_2112)
);

AND2x4_ASAP7_75t_L g2113 ( 
.A(n_2029),
.B(n_1989),
.Y(n_2113)
);

NOR2xp33_ASAP7_75t_L g2114 ( 
.A(n_2045),
.B(n_1920),
.Y(n_2114)
);

INVx2_ASAP7_75t_L g2115 ( 
.A(n_2032),
.Y(n_2115)
);

OAI33xp33_ASAP7_75t_L g2116 ( 
.A1(n_1998),
.A2(n_1992),
.A3(n_1827),
.B1(n_1824),
.B2(n_1821),
.B3(n_1825),
.Y(n_2116)
);

HB1xp67_ASAP7_75t_L g2117 ( 
.A(n_2046),
.Y(n_2117)
);

NAND2x1p5_ASAP7_75t_L g2118 ( 
.A(n_2048),
.B(n_1829),
.Y(n_2118)
);

OR2x2_ASAP7_75t_SL g2119 ( 
.A(n_2017),
.B(n_1939),
.Y(n_2119)
);

INVx1_ASAP7_75t_SL g2120 ( 
.A(n_2043),
.Y(n_2120)
);

INVx2_ASAP7_75t_SL g2121 ( 
.A(n_2033),
.Y(n_2121)
);

AND2x2_ASAP7_75t_L g2122 ( 
.A(n_2035),
.B(n_1943),
.Y(n_2122)
);

HB1xp67_ASAP7_75t_L g2123 ( 
.A(n_2046),
.Y(n_2123)
);

INVx2_ASAP7_75t_SL g2124 ( 
.A(n_2093),
.Y(n_2124)
);

AND2x4_ASAP7_75t_L g2125 ( 
.A(n_2093),
.B(n_1999),
.Y(n_2125)
);

OR2x2_ASAP7_75t_L g2126 ( 
.A(n_2056),
.B(n_2005),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_2097),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_L g2128 ( 
.A(n_2068),
.B(n_2005),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_2106),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_2111),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_2054),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_2055),
.Y(n_2132)
);

NAND2xp5_ASAP7_75t_L g2133 ( 
.A(n_2068),
.B(n_2041),
.Y(n_2133)
);

CKINVDCx20_ASAP7_75t_R g2134 ( 
.A(n_2077),
.Y(n_2134)
);

OR2x2_ASAP7_75t_L g2135 ( 
.A(n_2056),
.B(n_2024),
.Y(n_2135)
);

AND2x4_ASAP7_75t_L g2136 ( 
.A(n_2093),
.B(n_1999),
.Y(n_2136)
);

NOR3xp33_ASAP7_75t_SL g2137 ( 
.A(n_2058),
.B(n_2052),
.C(n_1987),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_2057),
.Y(n_2138)
);

NAND2xp5_ASAP7_75t_L g2139 ( 
.A(n_2080),
.B(n_2008),
.Y(n_2139)
);

INVx2_ASAP7_75t_L g2140 ( 
.A(n_2105),
.Y(n_2140)
);

AND2x2_ASAP7_75t_L g2141 ( 
.A(n_2071),
.B(n_2030),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_2059),
.Y(n_2142)
);

NOR4xp25_ASAP7_75t_SL g2143 ( 
.A(n_2053),
.B(n_1951),
.C(n_2001),
.D(n_1894),
.Y(n_2143)
);

INVx2_ASAP7_75t_L g2144 ( 
.A(n_2105),
.Y(n_2144)
);

AND2x2_ASAP7_75t_L g2145 ( 
.A(n_2071),
.B(n_2081),
.Y(n_2145)
);

NAND2xp5_ASAP7_75t_L g2146 ( 
.A(n_2095),
.B(n_2098),
.Y(n_2146)
);

AND2x2_ASAP7_75t_L g2147 ( 
.A(n_2081),
.B(n_2030),
.Y(n_2147)
);

INVx3_ASAP7_75t_SL g2148 ( 
.A(n_2119),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_2065),
.Y(n_2149)
);

AND2x2_ASAP7_75t_L g2150 ( 
.A(n_2062),
.B(n_2030),
.Y(n_2150)
);

AND2x2_ASAP7_75t_L g2151 ( 
.A(n_2062),
.B(n_2035),
.Y(n_2151)
);

HB1xp67_ASAP7_75t_L g2152 ( 
.A(n_2117),
.Y(n_2152)
);

INVx2_ASAP7_75t_L g2153 ( 
.A(n_2115),
.Y(n_2153)
);

AND2x2_ASAP7_75t_L g2154 ( 
.A(n_2101),
.B(n_2015),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_2073),
.Y(n_2155)
);

OAI21xp5_ASAP7_75t_L g2156 ( 
.A1(n_2061),
.A2(n_2052),
.B(n_2000),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_2074),
.Y(n_2157)
);

INVxp67_ASAP7_75t_SL g2158 ( 
.A(n_2070),
.Y(n_2158)
);

AND2x2_ASAP7_75t_L g2159 ( 
.A(n_2101),
.B(n_2015),
.Y(n_2159)
);

INVx2_ASAP7_75t_L g2160 ( 
.A(n_2115),
.Y(n_2160)
);

OR2x2_ASAP7_75t_L g2161 ( 
.A(n_2098),
.B(n_2024),
.Y(n_2161)
);

NAND2xp5_ASAP7_75t_L g2162 ( 
.A(n_2079),
.B(n_2012),
.Y(n_2162)
);

OAI33xp33_ASAP7_75t_L g2163 ( 
.A1(n_2060),
.A2(n_2039),
.A3(n_2014),
.B1(n_2007),
.B2(n_2010),
.B3(n_1996),
.Y(n_2163)
);

OR2x2_ASAP7_75t_L g2164 ( 
.A(n_2123),
.B(n_2012),
.Y(n_2164)
);

AND2x4_ASAP7_75t_L g2165 ( 
.A(n_2093),
.B(n_1997),
.Y(n_2165)
);

NAND2xp5_ASAP7_75t_L g2166 ( 
.A(n_2107),
.B(n_2016),
.Y(n_2166)
);

INVx2_ASAP7_75t_SL g2167 ( 
.A(n_2093),
.Y(n_2167)
);

AND2x2_ASAP7_75t_L g2168 ( 
.A(n_2072),
.B(n_2015),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_2075),
.Y(n_2169)
);

INVx2_ASAP7_75t_L g2170 ( 
.A(n_2102),
.Y(n_2170)
);

INVx3_ASAP7_75t_L g2171 ( 
.A(n_2092),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_2090),
.Y(n_2172)
);

BUFx2_ASAP7_75t_L g2173 ( 
.A(n_2083),
.Y(n_2173)
);

HB1xp67_ASAP7_75t_L g2174 ( 
.A(n_2103),
.Y(n_2174)
);

HB1xp67_ASAP7_75t_L g2175 ( 
.A(n_2087),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_2086),
.Y(n_2176)
);

NAND2xp5_ASAP7_75t_L g2177 ( 
.A(n_2066),
.B(n_2016),
.Y(n_2177)
);

OR2x2_ASAP7_75t_L g2178 ( 
.A(n_2112),
.B(n_2072),
.Y(n_2178)
);

INVx2_ASAP7_75t_L g2179 ( 
.A(n_2102),
.Y(n_2179)
);

NAND2x1p5_ASAP7_75t_L g2180 ( 
.A(n_2112),
.B(n_2000),
.Y(n_2180)
);

AND2x2_ASAP7_75t_L g2181 ( 
.A(n_2072),
.B(n_1997),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_2102),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_2127),
.Y(n_2183)
);

AND2x4_ASAP7_75t_L g2184 ( 
.A(n_2171),
.B(n_2076),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_2127),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_L g2186 ( 
.A(n_2128),
.B(n_2104),
.Y(n_2186)
);

INVx2_ASAP7_75t_L g2187 ( 
.A(n_2170),
.Y(n_2187)
);

NAND3xp33_ASAP7_75t_L g2188 ( 
.A(n_2156),
.B(n_2137),
.C(n_2143),
.Y(n_2188)
);

NOR2x1_ASAP7_75t_L g2189 ( 
.A(n_2134),
.B(n_1899),
.Y(n_2189)
);

INVx2_ASAP7_75t_L g2190 ( 
.A(n_2170),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_2129),
.Y(n_2191)
);

INVxp67_ASAP7_75t_SL g2192 ( 
.A(n_2180),
.Y(n_2192)
);

AND2x4_ASAP7_75t_L g2193 ( 
.A(n_2171),
.B(n_2076),
.Y(n_2193)
);

AND2x2_ASAP7_75t_L g2194 ( 
.A(n_2148),
.B(n_2112),
.Y(n_2194)
);

OAI21xp33_ASAP7_75t_L g2195 ( 
.A1(n_2156),
.A2(n_2069),
.B(n_2078),
.Y(n_2195)
);

NAND2xp5_ASAP7_75t_L g2196 ( 
.A(n_2133),
.B(n_2087),
.Y(n_2196)
);

HB1xp67_ASAP7_75t_L g2197 ( 
.A(n_2152),
.Y(n_2197)
);

OR2x2_ASAP7_75t_L g2198 ( 
.A(n_2177),
.B(n_2135),
.Y(n_2198)
);

OR2x2_ASAP7_75t_L g2199 ( 
.A(n_2177),
.B(n_2049),
.Y(n_2199)
);

OR2x2_ASAP7_75t_L g2200 ( 
.A(n_2135),
.B(n_2049),
.Y(n_2200)
);

NOR5xp2_ASAP7_75t_L g2201 ( 
.A(n_2174),
.B(n_1995),
.C(n_2009),
.D(n_2001),
.E(n_2010),
.Y(n_2201)
);

OR2x2_ASAP7_75t_L g2202 ( 
.A(n_2161),
.B(n_1995),
.Y(n_2202)
);

AND2x2_ASAP7_75t_L g2203 ( 
.A(n_2148),
.B(n_2072),
.Y(n_2203)
);

NAND2xp5_ASAP7_75t_L g2204 ( 
.A(n_2146),
.B(n_2094),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_2129),
.Y(n_2205)
);

NAND2xp5_ASAP7_75t_L g2206 ( 
.A(n_2139),
.B(n_2064),
.Y(n_2206)
);

INVx2_ASAP7_75t_L g2207 ( 
.A(n_2170),
.Y(n_2207)
);

INVx2_ASAP7_75t_SL g2208 ( 
.A(n_2165),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_2130),
.Y(n_2209)
);

OR2x2_ASAP7_75t_L g2210 ( 
.A(n_2161),
.B(n_2126),
.Y(n_2210)
);

AND2x2_ASAP7_75t_L g2211 ( 
.A(n_2148),
.B(n_2088),
.Y(n_2211)
);

NOR2x1_ASAP7_75t_L g2212 ( 
.A(n_2171),
.B(n_2173),
.Y(n_2212)
);

AND2x2_ASAP7_75t_L g2213 ( 
.A(n_2171),
.B(n_2088),
.Y(n_2213)
);

INVx2_ASAP7_75t_L g2214 ( 
.A(n_2179),
.Y(n_2214)
);

INVx2_ASAP7_75t_SL g2215 ( 
.A(n_2165),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_2130),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_2131),
.Y(n_2217)
);

INVx1_ASAP7_75t_SL g2218 ( 
.A(n_2173),
.Y(n_2218)
);

NAND2x1p5_ASAP7_75t_L g2219 ( 
.A(n_2125),
.B(n_2091),
.Y(n_2219)
);

INVxp67_ASAP7_75t_L g2220 ( 
.A(n_2163),
.Y(n_2220)
);

NAND2xp5_ASAP7_75t_L g2221 ( 
.A(n_2126),
.B(n_2120),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_2131),
.Y(n_2222)
);

AOI22xp5_ASAP7_75t_L g2223 ( 
.A1(n_2165),
.A2(n_2108),
.B1(n_2083),
.B2(n_2006),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_2132),
.Y(n_2224)
);

NOR2xp33_ASAP7_75t_SL g2225 ( 
.A(n_2165),
.B(n_2091),
.Y(n_2225)
);

INVx2_ASAP7_75t_L g2226 ( 
.A(n_2179),
.Y(n_2226)
);

OAI221xp5_ASAP7_75t_L g2227 ( 
.A1(n_2180),
.A2(n_2089),
.B1(n_2083),
.B2(n_2118),
.C(n_2096),
.Y(n_2227)
);

NAND3xp33_ASAP7_75t_L g2228 ( 
.A(n_2143),
.B(n_2018),
.C(n_1988),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_2132),
.Y(n_2229)
);

INVx2_ASAP7_75t_L g2230 ( 
.A(n_2179),
.Y(n_2230)
);

NAND2xp5_ASAP7_75t_L g2231 ( 
.A(n_2162),
.B(n_2099),
.Y(n_2231)
);

OR2x2_ASAP7_75t_L g2232 ( 
.A(n_2164),
.B(n_2175),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_2138),
.Y(n_2233)
);

BUFx3_ASAP7_75t_L g2234 ( 
.A(n_2124),
.Y(n_2234)
);

INVx1_ASAP7_75t_SL g2235 ( 
.A(n_2181),
.Y(n_2235)
);

AND2x2_ASAP7_75t_L g2236 ( 
.A(n_2145),
.B(n_2150),
.Y(n_2236)
);

OAI22xp5_ASAP7_75t_L g2237 ( 
.A1(n_2180),
.A2(n_2083),
.B1(n_2096),
.B2(n_2118),
.Y(n_2237)
);

OR2x2_ASAP7_75t_L g2238 ( 
.A(n_2166),
.B(n_2009),
.Y(n_2238)
);

INVx2_ASAP7_75t_SL g2239 ( 
.A(n_2124),
.Y(n_2239)
);

NAND2xp5_ASAP7_75t_L g2240 ( 
.A(n_2220),
.B(n_2141),
.Y(n_2240)
);

NAND2xp5_ASAP7_75t_L g2241 ( 
.A(n_2195),
.B(n_2141),
.Y(n_2241)
);

AND2x2_ASAP7_75t_L g2242 ( 
.A(n_2236),
.B(n_2145),
.Y(n_2242)
);

NOR2xp33_ASAP7_75t_SL g2243 ( 
.A(n_2189),
.B(n_2091),
.Y(n_2243)
);

OAI22xp33_ASAP7_75t_SL g2244 ( 
.A1(n_2186),
.A2(n_2167),
.B1(n_2178),
.B2(n_2136),
.Y(n_2244)
);

AOI22xp5_ASAP7_75t_L g2245 ( 
.A1(n_2188),
.A2(n_2235),
.B1(n_2211),
.B2(n_2225),
.Y(n_2245)
);

AND2x2_ASAP7_75t_L g2246 ( 
.A(n_2236),
.B(n_2150),
.Y(n_2246)
);

NOR2x1_ASAP7_75t_R g2247 ( 
.A(n_2203),
.B(n_1911),
.Y(n_2247)
);

NAND2xp5_ASAP7_75t_L g2248 ( 
.A(n_2218),
.B(n_2147),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_2183),
.Y(n_2249)
);

AND2x2_ASAP7_75t_SL g2250 ( 
.A(n_2201),
.B(n_1945),
.Y(n_2250)
);

AND2x2_ASAP7_75t_L g2251 ( 
.A(n_2211),
.B(n_2203),
.Y(n_2251)
);

NAND2xp5_ASAP7_75t_L g2252 ( 
.A(n_2204),
.B(n_2147),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_2185),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_2191),
.Y(n_2254)
);

NAND2xp5_ASAP7_75t_L g2255 ( 
.A(n_2197),
.B(n_2223),
.Y(n_2255)
);

NAND2x1p5_ASAP7_75t_L g2256 ( 
.A(n_2212),
.B(n_2125),
.Y(n_2256)
);

NAND2xp5_ASAP7_75t_L g2257 ( 
.A(n_2206),
.B(n_2154),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_2205),
.Y(n_2258)
);

NOR2x1_ASAP7_75t_L g2259 ( 
.A(n_2234),
.B(n_2178),
.Y(n_2259)
);

NAND2xp5_ASAP7_75t_L g2260 ( 
.A(n_2196),
.B(n_2154),
.Y(n_2260)
);

AOI211x1_ASAP7_75t_L g2261 ( 
.A1(n_2228),
.A2(n_2166),
.B(n_2151),
.C(n_2176),
.Y(n_2261)
);

OR2x2_ASAP7_75t_L g2262 ( 
.A(n_2198),
.B(n_2176),
.Y(n_2262)
);

NAND2xp5_ASAP7_75t_L g2263 ( 
.A(n_2231),
.B(n_2199),
.Y(n_2263)
);

INVx2_ASAP7_75t_L g2264 ( 
.A(n_2187),
.Y(n_2264)
);

AND2x2_ASAP7_75t_L g2265 ( 
.A(n_2194),
.B(n_2213),
.Y(n_2265)
);

NOR2xp33_ASAP7_75t_L g2266 ( 
.A(n_2227),
.B(n_1945),
.Y(n_2266)
);

AND2x2_ASAP7_75t_L g2267 ( 
.A(n_2194),
.B(n_2125),
.Y(n_2267)
);

AND2x2_ASAP7_75t_L g2268 ( 
.A(n_2213),
.B(n_2125),
.Y(n_2268)
);

OR2x2_ASAP7_75t_L g2269 ( 
.A(n_2198),
.B(n_2164),
.Y(n_2269)
);

INVxp67_ASAP7_75t_L g2270 ( 
.A(n_2234),
.Y(n_2270)
);

BUFx3_ASAP7_75t_L g2271 ( 
.A(n_2239),
.Y(n_2271)
);

AND2x2_ASAP7_75t_L g2272 ( 
.A(n_2184),
.B(n_2136),
.Y(n_2272)
);

NAND2xp5_ASAP7_75t_L g2273 ( 
.A(n_2199),
.B(n_2159),
.Y(n_2273)
);

OR2x2_ASAP7_75t_L g2274 ( 
.A(n_2232),
.B(n_2158),
.Y(n_2274)
);

AOI22xp33_ASAP7_75t_SL g2275 ( 
.A1(n_2192),
.A2(n_2136),
.B1(n_2033),
.B2(n_2013),
.Y(n_2275)
);

OAI21xp33_ASAP7_75t_L g2276 ( 
.A1(n_2208),
.A2(n_2013),
.B(n_2168),
.Y(n_2276)
);

OAI22xp5_ASAP7_75t_L g2277 ( 
.A1(n_2208),
.A2(n_2136),
.B1(n_2167),
.B2(n_2181),
.Y(n_2277)
);

HB1xp67_ASAP7_75t_L g2278 ( 
.A(n_2239),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_2209),
.Y(n_2279)
);

HB1xp67_ASAP7_75t_L g2280 ( 
.A(n_2210),
.Y(n_2280)
);

INVx2_ASAP7_75t_SL g2281 ( 
.A(n_2184),
.Y(n_2281)
);

AOI32xp33_ASAP7_75t_L g2282 ( 
.A1(n_2237),
.A2(n_2168),
.A3(n_2151),
.B1(n_2013),
.B2(n_2114),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_2280),
.Y(n_2283)
);

AOI21xp5_ASAP7_75t_L g2284 ( 
.A1(n_2255),
.A2(n_2215),
.B(n_2219),
.Y(n_2284)
);

NAND2xp5_ASAP7_75t_L g2285 ( 
.A(n_2240),
.B(n_2216),
.Y(n_2285)
);

NAND2xp5_ASAP7_75t_L g2286 ( 
.A(n_2270),
.B(n_2215),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_2249),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_2249),
.Y(n_2288)
);

NAND2x1_ASAP7_75t_L g2289 ( 
.A(n_2259),
.B(n_2184),
.Y(n_2289)
);

OAI22xp33_ASAP7_75t_L g2290 ( 
.A1(n_2245),
.A2(n_2219),
.B1(n_2221),
.B2(n_2210),
.Y(n_2290)
);

OR2x2_ASAP7_75t_L g2291 ( 
.A(n_2274),
.B(n_2200),
.Y(n_2291)
);

OAI21xp5_ASAP7_75t_L g2292 ( 
.A1(n_2250),
.A2(n_1916),
.B(n_2114),
.Y(n_2292)
);

AOI221xp5_ASAP7_75t_L g2293 ( 
.A1(n_2261),
.A2(n_2244),
.B1(n_2241),
.B2(n_2282),
.C(n_2252),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_2254),
.Y(n_2294)
);

A2O1A1Ixp33_ASAP7_75t_L g2295 ( 
.A1(n_2243),
.A2(n_2193),
.B(n_2002),
.C(n_2200),
.Y(n_2295)
);

INVx2_ASAP7_75t_SL g2296 ( 
.A(n_2271),
.Y(n_2296)
);

AOI322xp5_ASAP7_75t_L g2297 ( 
.A1(n_2250),
.A2(n_2002),
.A3(n_2193),
.B1(n_2159),
.B2(n_2003),
.C1(n_2229),
.C2(n_2224),
.Y(n_2297)
);

INVx1_ASAP7_75t_L g2298 ( 
.A(n_2254),
.Y(n_2298)
);

NAND2xp5_ASAP7_75t_L g2299 ( 
.A(n_2251),
.B(n_2193),
.Y(n_2299)
);

AOI221xp5_ASAP7_75t_L g2300 ( 
.A1(n_2276),
.A2(n_2233),
.B1(n_2217),
.B2(n_2222),
.C(n_2238),
.Y(n_2300)
);

NAND2xp5_ASAP7_75t_L g2301 ( 
.A(n_2242),
.B(n_2138),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_2258),
.Y(n_2302)
);

AND2x2_ASAP7_75t_L g2303 ( 
.A(n_2251),
.B(n_2109),
.Y(n_2303)
);

AOI22xp5_ASAP7_75t_L g2304 ( 
.A1(n_2266),
.A2(n_2116),
.B1(n_2076),
.B2(n_2082),
.Y(n_2304)
);

OAI22xp33_ASAP7_75t_SL g2305 ( 
.A1(n_2256),
.A2(n_2202),
.B1(n_2238),
.B2(n_2144),
.Y(n_2305)
);

NAND2xp5_ASAP7_75t_L g2306 ( 
.A(n_2265),
.B(n_2142),
.Y(n_2306)
);

NAND2xp5_ASAP7_75t_L g2307 ( 
.A(n_2265),
.B(n_2142),
.Y(n_2307)
);

AOI22xp5_ASAP7_75t_L g2308 ( 
.A1(n_2277),
.A2(n_2082),
.B1(n_2085),
.B2(n_2113),
.Y(n_2308)
);

INVx1_ASAP7_75t_L g2309 ( 
.A(n_2258),
.Y(n_2309)
);

OR2x2_ASAP7_75t_L g2310 ( 
.A(n_2274),
.B(n_2202),
.Y(n_2310)
);

NAND2xp5_ASAP7_75t_L g2311 ( 
.A(n_2242),
.B(n_2278),
.Y(n_2311)
);

OAI32xp33_ASAP7_75t_L g2312 ( 
.A1(n_2256),
.A2(n_2182),
.A3(n_2002),
.B1(n_2039),
.B2(n_2160),
.Y(n_2312)
);

INVx1_ASAP7_75t_SL g2313 ( 
.A(n_2289),
.Y(n_2313)
);

NAND2xp5_ASAP7_75t_L g2314 ( 
.A(n_2283),
.B(n_2253),
.Y(n_2314)
);

INVx1_ASAP7_75t_L g2315 ( 
.A(n_2287),
.Y(n_2315)
);

O2A1O1Ixp33_ASAP7_75t_L g2316 ( 
.A1(n_2292),
.A2(n_2256),
.B(n_2271),
.C(n_2281),
.Y(n_2316)
);

AND2x2_ASAP7_75t_L g2317 ( 
.A(n_2303),
.B(n_2272),
.Y(n_2317)
);

AOI221xp5_ASAP7_75t_L g2318 ( 
.A1(n_2293),
.A2(n_2281),
.B1(n_2279),
.B2(n_2263),
.C(n_2248),
.Y(n_2318)
);

OAI21xp33_ASAP7_75t_L g2319 ( 
.A1(n_2311),
.A2(n_2267),
.B(n_2275),
.Y(n_2319)
);

NAND4xp25_ASAP7_75t_L g2320 ( 
.A(n_2284),
.B(n_2267),
.C(n_2272),
.D(n_2268),
.Y(n_2320)
);

AOI21xp5_ASAP7_75t_L g2321 ( 
.A1(n_2292),
.A2(n_2247),
.B(n_2262),
.Y(n_2321)
);

AOI322xp5_ASAP7_75t_L g2322 ( 
.A1(n_2290),
.A2(n_2246),
.A3(n_2273),
.B1(n_2268),
.B2(n_2257),
.C1(n_2260),
.C2(n_2182),
.Y(n_2322)
);

OR2x2_ASAP7_75t_L g2323 ( 
.A(n_2291),
.B(n_2269),
.Y(n_2323)
);

AOI32xp33_ASAP7_75t_L g2324 ( 
.A1(n_2300),
.A2(n_2246),
.A3(n_2262),
.B1(n_2269),
.B2(n_2264),
.Y(n_2324)
);

NOR2xp67_ASAP7_75t_L g2325 ( 
.A(n_2296),
.B(n_2264),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_L g2326 ( 
.A(n_2286),
.B(n_2149),
.Y(n_2326)
);

NAND2xp5_ASAP7_75t_L g2327 ( 
.A(n_2285),
.B(n_2149),
.Y(n_2327)
);

NAND2xp5_ASAP7_75t_L g2328 ( 
.A(n_2285),
.B(n_2155),
.Y(n_2328)
);

OAI22xp5_ASAP7_75t_L g2329 ( 
.A1(n_2308),
.A2(n_2082),
.B1(n_2113),
.B2(n_2085),
.Y(n_2329)
);

INVxp67_ASAP7_75t_L g2330 ( 
.A(n_2299),
.Y(n_2330)
);

OAI31xp33_ASAP7_75t_L g2331 ( 
.A1(n_2305),
.A2(n_1907),
.A3(n_1911),
.B(n_2085),
.Y(n_2331)
);

AOI222xp33_ASAP7_75t_L g2332 ( 
.A1(n_2312),
.A2(n_2003),
.B1(n_2033),
.B2(n_2050),
.C1(n_2016),
.C2(n_2190),
.Y(n_2332)
);

OAI22xp5_ASAP7_75t_L g2333 ( 
.A1(n_2304),
.A2(n_2113),
.B1(n_2067),
.B2(n_2063),
.Y(n_2333)
);

AND2x2_ASAP7_75t_L g2334 ( 
.A(n_2310),
.B(n_2109),
.Y(n_2334)
);

NAND2xp5_ASAP7_75t_L g2335 ( 
.A(n_2288),
.B(n_2294),
.Y(n_2335)
);

NAND3xp33_ASAP7_75t_L g2336 ( 
.A(n_2297),
.B(n_2190),
.C(n_2187),
.Y(n_2336)
);

INVx1_ASAP7_75t_SL g2337 ( 
.A(n_2313),
.Y(n_2337)
);

INVxp33_ASAP7_75t_L g2338 ( 
.A(n_2323),
.Y(n_2338)
);

NOR2xp33_ASAP7_75t_L g2339 ( 
.A(n_2330),
.B(n_2306),
.Y(n_2339)
);

NAND2xp5_ASAP7_75t_L g2340 ( 
.A(n_2325),
.B(n_2298),
.Y(n_2340)
);

OAI21xp5_ASAP7_75t_L g2341 ( 
.A1(n_2316),
.A2(n_2295),
.B(n_2307),
.Y(n_2341)
);

INVx1_ASAP7_75t_SL g2342 ( 
.A(n_2317),
.Y(n_2342)
);

OAI21xp33_ASAP7_75t_L g2343 ( 
.A1(n_2319),
.A2(n_2301),
.B(n_2302),
.Y(n_2343)
);

NAND2x1p5_ASAP7_75t_L g2344 ( 
.A(n_2315),
.B(n_2309),
.Y(n_2344)
);

OAI22xp33_ASAP7_75t_L g2345 ( 
.A1(n_2321),
.A2(n_2301),
.B1(n_2121),
.B2(n_2063),
.Y(n_2345)
);

OAI21xp5_ASAP7_75t_L g2346 ( 
.A1(n_2322),
.A2(n_2214),
.B(n_2207),
.Y(n_2346)
);

AND2x2_ASAP7_75t_L g2347 ( 
.A(n_2334),
.B(n_2099),
.Y(n_2347)
);

AOI22xp5_ASAP7_75t_L g2348 ( 
.A1(n_2320),
.A2(n_2084),
.B1(n_1924),
.B2(n_2121),
.Y(n_2348)
);

INVx1_ASAP7_75t_L g2349 ( 
.A(n_2314),
.Y(n_2349)
);

NOR2xp33_ASAP7_75t_L g2350 ( 
.A(n_2314),
.B(n_2326),
.Y(n_2350)
);

NAND2xp5_ASAP7_75t_L g2351 ( 
.A(n_2318),
.B(n_2155),
.Y(n_2351)
);

NAND2xp5_ASAP7_75t_SL g2352 ( 
.A(n_2337),
.B(n_2331),
.Y(n_2352)
);

AOI31xp33_ASAP7_75t_L g2353 ( 
.A1(n_2338),
.A2(n_2335),
.A3(n_2329),
.B(n_2333),
.Y(n_2353)
);

NOR3xp33_ASAP7_75t_L g2354 ( 
.A(n_2343),
.B(n_2324),
.C(n_2336),
.Y(n_2354)
);

NAND2xp5_ASAP7_75t_L g2355 ( 
.A(n_2342),
.B(n_2328),
.Y(n_2355)
);

NAND3xp33_ASAP7_75t_L g2356 ( 
.A(n_2340),
.B(n_2332),
.C(n_2327),
.Y(n_2356)
);

INVx1_ASAP7_75t_L g2357 ( 
.A(n_2344),
.Y(n_2357)
);

NOR3xp33_ASAP7_75t_L g2358 ( 
.A(n_2345),
.B(n_2327),
.C(n_2214),
.Y(n_2358)
);

NAND4xp25_ASAP7_75t_L g2359 ( 
.A(n_2339),
.B(n_1924),
.C(n_2226),
.D(n_2207),
.Y(n_2359)
);

OAI21xp5_ASAP7_75t_L g2360 ( 
.A1(n_2351),
.A2(n_2230),
.B(n_2226),
.Y(n_2360)
);

NAND2xp5_ASAP7_75t_L g2361 ( 
.A(n_2350),
.B(n_2140),
.Y(n_2361)
);

NAND2xp5_ASAP7_75t_L g2362 ( 
.A(n_2349),
.B(n_2140),
.Y(n_2362)
);

NAND2xp5_ASAP7_75t_L g2363 ( 
.A(n_2344),
.B(n_2140),
.Y(n_2363)
);

O2A1O1Ixp33_ASAP7_75t_SL g2364 ( 
.A1(n_2341),
.A2(n_2230),
.B(n_2160),
.C(n_2144),
.Y(n_2364)
);

NAND3xp33_ASAP7_75t_L g2365 ( 
.A(n_2354),
.B(n_2346),
.C(n_2348),
.Y(n_2365)
);

NOR4xp25_ASAP7_75t_L g2366 ( 
.A(n_2357),
.B(n_2347),
.C(n_2172),
.D(n_2157),
.Y(n_2366)
);

OAI221xp5_ASAP7_75t_SL g2367 ( 
.A1(n_2356),
.A2(n_2100),
.B1(n_2144),
.B2(n_2153),
.C(n_2160),
.Y(n_2367)
);

AND2x2_ASAP7_75t_L g2368 ( 
.A(n_2352),
.B(n_2153),
.Y(n_2368)
);

OAI221xp5_ASAP7_75t_L g2369 ( 
.A1(n_2353),
.A2(n_2100),
.B1(n_2153),
.B2(n_2157),
.C(n_2169),
.Y(n_2369)
);

AOI221xp5_ASAP7_75t_L g2370 ( 
.A1(n_2364),
.A2(n_2172),
.B1(n_2169),
.B2(n_2003),
.C(n_2084),
.Y(n_2370)
);

XOR2xp5_ASAP7_75t_L g2371 ( 
.A(n_2355),
.B(n_1866),
.Y(n_2371)
);

NAND2xp5_ASAP7_75t_L g2372 ( 
.A(n_2358),
.B(n_2084),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_2361),
.Y(n_2373)
);

NOR3xp33_ASAP7_75t_L g2374 ( 
.A(n_2359),
.B(n_2362),
.C(n_2363),
.Y(n_2374)
);

OAI22xp33_ASAP7_75t_L g2375 ( 
.A1(n_2365),
.A2(n_2360),
.B1(n_1975),
.B2(n_1934),
.Y(n_2375)
);

INVx2_ASAP7_75t_L g2376 ( 
.A(n_2368),
.Y(n_2376)
);

NAND2xp5_ASAP7_75t_L g2377 ( 
.A(n_2366),
.B(n_2122),
.Y(n_2377)
);

OAI211xp5_ASAP7_75t_SL g2378 ( 
.A1(n_2369),
.A2(n_1893),
.B(n_1871),
.C(n_1873),
.Y(n_2378)
);

OAI211xp5_ASAP7_75t_L g2379 ( 
.A1(n_2367),
.A2(n_1887),
.B(n_1871),
.C(n_1873),
.Y(n_2379)
);

OAI211xp5_ASAP7_75t_SL g2380 ( 
.A1(n_2374),
.A2(n_1887),
.B(n_1884),
.C(n_1893),
.Y(n_2380)
);

O2A1O1Ixp33_ASAP7_75t_L g2381 ( 
.A1(n_2373),
.A2(n_1884),
.B(n_1876),
.C(n_1892),
.Y(n_2381)
);

AOI221xp5_ASAP7_75t_L g2382 ( 
.A1(n_2372),
.A2(n_1927),
.B1(n_1922),
.B2(n_1890),
.C(n_1892),
.Y(n_2382)
);

INVx1_ASAP7_75t_SL g2383 ( 
.A(n_2371),
.Y(n_2383)
);

NOR2x1p5_ASAP7_75t_L g2384 ( 
.A(n_2376),
.B(n_2370),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_2377),
.Y(n_2385)
);

HB1xp67_ASAP7_75t_L g2386 ( 
.A(n_2383),
.Y(n_2386)
);

AND2x2_ASAP7_75t_L g2387 ( 
.A(n_2382),
.B(n_2067),
.Y(n_2387)
);

AND3x4_ASAP7_75t_L g2388 ( 
.A(n_2380),
.B(n_1902),
.C(n_1875),
.Y(n_2388)
);

AOI22xp5_ASAP7_75t_L g2389 ( 
.A1(n_2375),
.A2(n_1983),
.B1(n_2122),
.B2(n_1902),
.Y(n_2389)
);

XNOR2xp5_ASAP7_75t_L g2390 ( 
.A(n_2379),
.B(n_1967),
.Y(n_2390)
);

NOR2x1p5_ASAP7_75t_L g2391 ( 
.A(n_2385),
.B(n_2378),
.Y(n_2391)
);

INVx1_ASAP7_75t_L g2392 ( 
.A(n_2386),
.Y(n_2392)
);

NAND4xp75_ASAP7_75t_L g2393 ( 
.A(n_2389),
.B(n_2381),
.C(n_1898),
.D(n_2034),
.Y(n_2393)
);

XNOR2x1_ASAP7_75t_L g2394 ( 
.A(n_2384),
.B(n_1875),
.Y(n_2394)
);

AOI21xp5_ASAP7_75t_L g2395 ( 
.A1(n_2392),
.A2(n_2390),
.B(n_2389),
.Y(n_2395)
);

INVx1_ASAP7_75t_L g2396 ( 
.A(n_2391),
.Y(n_2396)
);

INVx1_ASAP7_75t_L g2397 ( 
.A(n_2396),
.Y(n_2397)
);

AOI22xp5_ASAP7_75t_L g2398 ( 
.A1(n_2397),
.A2(n_2394),
.B1(n_2395),
.B2(n_2387),
.Y(n_2398)
);

OAI21x1_ASAP7_75t_SL g2399 ( 
.A1(n_2397),
.A2(n_2393),
.B(n_2388),
.Y(n_2399)
);

OAI22xp5_ASAP7_75t_L g2400 ( 
.A1(n_2398),
.A2(n_1875),
.B1(n_1889),
.B2(n_1885),
.Y(n_2400)
);

AOI21xp5_ASAP7_75t_L g2401 ( 
.A1(n_2399),
.A2(n_1875),
.B(n_1915),
.Y(n_2401)
);

OAI22xp5_ASAP7_75t_L g2402 ( 
.A1(n_2401),
.A2(n_1879),
.B1(n_1889),
.B2(n_1885),
.Y(n_2402)
);

INVx1_ASAP7_75t_L g2403 ( 
.A(n_2400),
.Y(n_2403)
);

OA21x2_ASAP7_75t_L g2404 ( 
.A1(n_2403),
.A2(n_1852),
.B(n_1861),
.Y(n_2404)
);

AOI22xp5_ASAP7_75t_L g2405 ( 
.A1(n_2404),
.A2(n_2402),
.B1(n_1987),
.B2(n_2110),
.Y(n_2405)
);

OAI22xp33_ASAP7_75t_L g2406 ( 
.A1(n_2405),
.A2(n_1860),
.B1(n_1845),
.B2(n_1858),
.Y(n_2406)
);

OAI221xp5_ASAP7_75t_R g2407 ( 
.A1(n_2406),
.A2(n_1915),
.B1(n_1819),
.B2(n_1864),
.C(n_2110),
.Y(n_2407)
);

AOI211xp5_ASAP7_75t_L g2408 ( 
.A1(n_2407),
.A2(n_1860),
.B(n_1845),
.C(n_1858),
.Y(n_2408)
);


endmodule