module fake_jpeg_25076_n_116 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_116);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_116;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_2),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_17),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_26),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_31),
.Y(n_48)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_0),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_51),
.B(n_40),
.Y(n_58)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_52),
.B(n_54),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

CKINVDCx6p67_ASAP7_75t_R g70 ( 
.A(n_53),
.Y(n_70)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_56),
.Y(n_64)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_46),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_39),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_58),
.B(n_59),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_51),
.B(n_37),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_50),
.B(n_37),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_66),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_57),
.A2(n_49),
.B1(n_43),
.B2(n_47),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_1),
.Y(n_74)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_51),
.B(n_48),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_56),
.A2(n_45),
.B1(n_42),
.B2(n_38),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_67),
.A2(n_69),
.B1(n_0),
.B2(n_1),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_51),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_68),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_56),
.A2(n_19),
.B1(n_36),
.B2(n_34),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_71),
.B(n_79),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_69),
.A2(n_16),
.B1(n_32),
.B2(n_30),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_72),
.A2(n_73),
.B1(n_78),
.B2(n_3),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_74),
.A2(n_5),
.B(n_6),
.Y(n_93)
);

A2O1A1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_67),
.A2(n_3),
.B(n_4),
.C(n_5),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_77),
.A2(n_74),
.B(n_83),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_70),
.A2(n_18),
.B1(n_29),
.B2(n_28),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

INVx3_ASAP7_75t_SL g80 ( 
.A(n_70),
.Y(n_80)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_80),
.Y(n_89)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_4),
.Y(n_91)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_82),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_87),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_93),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_90),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_91),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_94),
.B(n_84),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_86),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_95),
.B(n_100),
.Y(n_106)
);

OAI21xp33_ASAP7_75t_L g101 ( 
.A1(n_85),
.A2(n_6),
.B(n_7),
.Y(n_101)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_101),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_97),
.B(n_89),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_102),
.B(n_104),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_99),
.B(n_89),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_96),
.B(n_75),
.C(n_92),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_105),
.B(n_98),
.C(n_101),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_107),
.A2(n_103),
.B(n_106),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_109),
.B(n_108),
.Y(n_110)
);

AOI31xp33_ASAP7_75t_L g111 ( 
.A1(n_110),
.A2(n_8),
.A3(n_9),
.B(n_10),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_111),
.B(n_11),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_112),
.B(n_14),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_20),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_22),
.C(n_23),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_115),
.B(n_25),
.Y(n_116)
);


endmodule