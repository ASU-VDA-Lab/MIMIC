module real_jpeg_28365_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_215;
wire n_166;
wire n_176;
wire n_300;
wire n_292;
wire n_221;
wire n_286;
wire n_288;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_301;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_299;
wire n_243;
wire n_115;
wire n_255;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_275;
wire n_293;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_238;
wire n_76;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_302;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_298;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_297;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_167;
wire n_295;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_216;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_210;
wire n_53;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_0),
.A2(n_29),
.B1(n_30),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_0),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_0),
.A2(n_38),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_0),
.A2(n_33),
.B1(n_34),
.B2(n_38),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_0),
.A2(n_38),
.B1(n_47),
.B2(n_51),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_1),
.A2(n_33),
.B1(n_34),
.B2(n_44),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_1),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_1),
.A2(n_44),
.B1(n_47),
.B2(n_51),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_1),
.A2(n_44),
.B1(n_77),
.B2(n_78),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_44),
.Y(n_148)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_2),
.Y(n_92)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_2),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_3),
.A2(n_33),
.B1(n_34),
.B2(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_3),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_58),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_3),
.A2(n_58),
.B1(n_77),
.B2(n_78),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_3),
.A2(n_47),
.B1(n_51),
.B2(n_58),
.Y(n_115)
);

BUFx12_ASAP7_75t_L g75 ( 
.A(n_4),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_5),
.A2(n_29),
.B1(n_30),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_5),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_5),
.A2(n_33),
.B1(n_34),
.B2(n_40),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_5),
.A2(n_40),
.B1(n_47),
.B2(n_51),
.Y(n_142)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_7),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_8),
.A2(n_77),
.B1(n_78),
.B2(n_152),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_8),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_8),
.A2(n_29),
.B1(n_30),
.B2(n_152),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_8),
.A2(n_33),
.B1(n_34),
.B2(n_152),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_8),
.A2(n_47),
.B1(n_51),
.B2(n_152),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_9),
.A2(n_77),
.B1(n_78),
.B2(n_126),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_9),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_9),
.A2(n_29),
.B1(n_30),
.B2(n_126),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_9),
.A2(n_33),
.B1(n_34),
.B2(n_126),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_9),
.A2(n_47),
.B1(n_51),
.B2(n_126),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_10),
.A2(n_77),
.B1(n_78),
.B2(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_10),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_173),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_10),
.A2(n_33),
.B1(n_34),
.B2(n_173),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_10),
.A2(n_47),
.B1(n_51),
.B2(n_173),
.Y(n_259)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_12),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_12),
.B(n_73),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_12),
.B(n_29),
.Y(n_211)
);

AOI21xp33_ASAP7_75t_L g215 ( 
.A1(n_12),
.A2(n_29),
.B(n_211),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_12),
.A2(n_33),
.B1(n_34),
.B2(n_171),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_12),
.A2(n_47),
.B(n_52),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_12),
.B(n_120),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_12),
.A2(n_89),
.B1(n_93),
.B2(n_259),
.Y(n_261)
);

BUFx24_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx11_ASAP7_75t_SL g49 ( 
.A(n_15),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_130),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_128),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_103),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_19),
.B(n_103),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_86),
.B2(n_87),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_59),
.B2(n_60),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_23),
.A2(n_24),
.B(n_41),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_41),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_32),
.B1(n_36),
.B2(n_39),
.Y(n_24)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_25),
.B(n_70),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_25),
.A2(n_32),
.B1(n_167),
.B2(n_168),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_25),
.A2(n_32),
.B1(n_167),
.B2(n_196),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_25),
.A2(n_32),
.B1(n_196),
.B2(n_215),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_32),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_27),
.A2(n_28),
.B1(n_33),
.B2(n_34),
.Y(n_32)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_27),
.Y(n_210)
);

NAND2xp33_ASAP7_75t_SL g212 ( 
.A(n_27),
.B(n_34),
.Y(n_212)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_29),
.A2(n_30),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_29),
.B(n_74),
.Y(n_185)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_30),
.A2(n_81),
.B1(n_170),
.B2(n_185),
.Y(n_184)
);

AOI32xp33_ASAP7_75t_L g209 ( 
.A1(n_30),
.A2(n_33),
.A3(n_210),
.B1(n_211),
.B2(n_212),
.Y(n_209)
);

BUFx4f_ASAP7_75t_SL g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_32),
.B(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_32),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_32),
.B(n_148),
.Y(n_182)
);

OAI22xp33_ASAP7_75t_L g56 ( 
.A1(n_33),
.A2(n_34),
.B1(n_50),
.B2(n_52),
.Y(n_56)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

A2O1A1Ixp33_ASAP7_75t_L g237 ( 
.A1(n_34),
.A2(n_50),
.B(n_171),
.C(n_238),
.Y(n_237)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_37),
.A2(n_120),
.B(n_121),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_39),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_53),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_42),
.A2(n_55),
.B(n_219),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_43),
.B(n_45),
.Y(n_42)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_45),
.B(n_57),
.Y(n_99)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_56),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_46),
.A2(n_55),
.B(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_46),
.A2(n_55),
.B1(n_98),
.B2(n_118),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_46),
.A2(n_53),
.B(n_118),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_46),
.A2(n_55),
.B1(n_218),
.B2(n_219),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_46),
.A2(n_55),
.B1(n_235),
.B2(n_236),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_46),
.A2(n_55),
.B1(n_218),
.B2(n_236),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_46),
.B(n_171),
.Y(n_257)
);

OA22x2_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_46)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

BUFx4f_ASAP7_75t_SL g47 ( 
.A(n_48),
.Y(n_47)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_51),
.B(n_91),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_51),
.B(n_263),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_54),
.B(n_57),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_55),
.A2(n_98),
.B(n_99),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_55),
.A2(n_64),
.B(n_99),
.Y(n_164)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_71),
.B1(n_84),
.B2(n_85),
.Y(n_60)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_63),
.B1(n_65),
.B2(n_66),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_68),
.B(n_69),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_67),
.A2(n_69),
.B(n_147),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_67),
.A2(n_181),
.B(n_182),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_71),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_76),
.B(n_79),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_72),
.B(n_83),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_72),
.A2(n_124),
.B1(n_125),
.B2(n_151),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_72),
.A2(n_124),
.B1(n_151),
.B2(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

O2A1O1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_73),
.A2(n_74),
.B(n_78),
.C(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_73),
.B(n_101),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_73),
.A2(n_80),
.B1(n_170),
.B2(n_172),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_78),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_77),
.Y(n_78)
);

HAxp5_ASAP7_75t_SL g170 ( 
.A(n_78),
.B(n_171),
.CON(n_170),
.SN(n_170)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_80),
.B(n_82),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_80),
.A2(n_101),
.B(n_102),
.Y(n_100)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_80),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_96),
.B(n_100),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_88),
.B(n_97),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_88),
.A2(n_100),
.B1(n_106),
.B2(n_107),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_88),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_88),
.A2(n_97),
.B1(n_107),
.B2(n_138),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_93),
.B(n_94),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_89),
.A2(n_142),
.B(n_143),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_89),
.A2(n_92),
.B1(n_142),
.B2(n_187),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_89),
.A2(n_116),
.B(n_246),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_89),
.A2(n_200),
.B1(n_251),
.B2(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_90),
.B(n_114),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_90),
.A2(n_95),
.B(n_144),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_90),
.A2(n_91),
.B1(n_250),
.B2(n_252),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_91),
.B(n_95),
.Y(n_116)
);

INVx11_ASAP7_75t_L g200 ( 
.A(n_91),
.Y(n_200)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_93),
.B(n_115),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_93),
.B(n_171),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_96),
.B(n_105),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_97),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_100),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_108),
.C(n_109),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_104),
.B(n_108),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_109),
.A2(n_110),
.B1(n_154),
.B2(n_155),
.Y(n_153)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_119),
.C(n_122),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_111),
.B(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_117),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_112),
.B(n_117),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_116),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_113),
.A2(n_187),
.B(n_200),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_119),
.A2(n_122),
.B1(n_123),
.B2(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_119),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_125),
.B(n_127),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_156),
.B(n_302),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_153),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_132),
.B(n_153),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_137),
.C(n_139),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_133),
.A2(n_134),
.B1(n_137),
.B2(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_137),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_139),
.B(n_299),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_146),
.C(n_149),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_140),
.B(n_291),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_145),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_141),
.B(n_145),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_146),
.A2(n_149),
.B1(n_150),
.B2(n_292),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_146),
.Y(n_292)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_296),
.B(n_301),
.Y(n_156)
);

O2A1O1Ixp33_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_201),
.B(n_282),
.C(n_295),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_188),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_159),
.B(n_188),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_174),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_162),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_161),
.B(n_162),
.C(n_174),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_165),
.C(n_169),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_163),
.A2(n_164),
.B1(n_165),
.B2(n_166),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_168),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_169),
.B(n_191),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_172),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_175),
.B(n_183),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_177),
.B1(n_179),
.B2(n_180),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_176),
.B(n_180),
.C(n_183),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_186),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_184),
.B(n_186),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_192),
.C(n_194),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_189),
.A2(n_190),
.B1(n_277),
.B2(n_279),
.Y(n_276)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_192),
.A2(n_193),
.B1(n_194),
.B2(n_278),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_194),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_197),
.C(n_199),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_195),
.B(n_223),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_197),
.A2(n_198),
.B1(n_199),
.B2(n_224),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_198),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_199),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_281),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_274),
.B(n_280),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_229),
.B(n_273),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_220),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_205),
.B(n_220),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_213),
.C(n_216),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_206),
.A2(n_207),
.B1(n_270),
.B2(n_271),
.Y(n_269)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_208),
.B(n_209),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_213),
.A2(n_214),
.B1(n_216),
.B2(n_217),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_214),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_222),
.B1(n_225),
.B2(n_226),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_221),
.B(n_227),
.C(n_228),
.Y(n_275)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_267),
.B(n_272),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_247),
.B(n_266),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_239),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_232),
.B(n_239),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_233),
.B(n_237),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_233),
.A2(n_234),
.B1(n_237),
.B2(n_254),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_234),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_237),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_245),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_242),
.B1(n_243),
.B2(n_244),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_241),
.B(n_244),
.C(n_245),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_242),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_244),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_246),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_255),
.B(n_265),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_253),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_249),
.B(n_253),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_260),
.B(n_264),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_257),
.B(n_258),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_268),
.B(n_269),
.Y(n_272)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_275),
.B(n_276),
.Y(n_280)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_277),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_283),
.B(n_284),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_285),
.A2(n_286),
.B1(n_293),
.B2(n_294),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_288),
.B1(n_289),
.B2(n_290),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_287),
.B(n_290),
.C(n_294),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_293),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_297),
.B(n_298),
.Y(n_301)
);


endmodule