module real_aes_1217_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_841;
wire n_318;
wire n_718;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_815;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_292;
wire n_539;
wire n_400;
wire n_626;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_528;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_434;
wire n_502;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_749;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_L g587 ( .A(n_0), .B(n_242), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_1), .B(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g165 ( .A(n_2), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_3), .B(n_524), .Y(n_523) );
NAND2xp33_ASAP7_75t_SL g579 ( .A(n_4), .B(n_182), .Y(n_579) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_5), .B(n_226), .Y(n_234) );
INVx1_ASAP7_75t_L g572 ( .A(n_6), .Y(n_572) );
INVx1_ASAP7_75t_L g173 ( .A(n_7), .Y(n_173) );
CKINVDCx16_ASAP7_75t_R g113 ( .A(n_8), .Y(n_113) );
AOI22xp5_ASAP7_75t_SL g131 ( .A1(n_9), .A2(n_132), .B1(n_133), .B2(n_134), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_9), .Y(n_132) );
OAI22x1_ASAP7_75t_R g134 ( .A1(n_10), .A2(n_80), .B1(n_135), .B2(n_136), .Y(n_134) );
CKINVDCx20_ASAP7_75t_R g135 ( .A(n_10), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g199 ( .A(n_11), .Y(n_199) );
AND2x2_ASAP7_75t_L g521 ( .A(n_12), .B(n_214), .Y(n_521) );
INVx2_ASAP7_75t_L g155 ( .A(n_13), .Y(n_155) );
AND3x1_ASAP7_75t_L g110 ( .A(n_14), .B(n_39), .C(n_111), .Y(n_110) );
CKINVDCx16_ASAP7_75t_R g125 ( .A(n_14), .Y(n_125) );
INVx1_ASAP7_75t_L g243 ( .A(n_15), .Y(n_243) );
AOI221x1_ASAP7_75t_L g575 ( .A1(n_16), .A2(n_186), .B1(n_526), .B2(n_576), .C(n_578), .Y(n_575) );
NAND2xp5_ASAP7_75t_SL g559 ( .A(n_17), .B(n_524), .Y(n_559) );
INVx1_ASAP7_75t_L g109 ( .A(n_18), .Y(n_109) );
INVx1_ASAP7_75t_L g240 ( .A(n_19), .Y(n_240) );
INVx1_ASAP7_75t_SL g255 ( .A(n_20), .Y(n_255) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_21), .B(n_176), .Y(n_229) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_22), .Y(n_122) );
OAI22xp5_ASAP7_75t_L g839 ( .A1(n_23), .A2(n_30), .B1(n_512), .B2(n_840), .Y(n_839) );
INVx1_ASAP7_75t_L g840 ( .A(n_23), .Y(n_840) );
AOI33xp33_ASAP7_75t_L g280 ( .A1(n_24), .A2(n_54), .A3(n_160), .B1(n_168), .B2(n_281), .B3(n_282), .Y(n_280) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_25), .A2(n_526), .B(n_527), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_26), .B(n_242), .Y(n_528) );
AOI221xp5_ASAP7_75t_SL g551 ( .A1(n_27), .A2(n_44), .B1(n_524), .B2(n_526), .C(n_552), .Y(n_551) );
OAI21xp5_ASAP7_75t_L g826 ( .A1(n_28), .A2(n_827), .B(n_842), .Y(n_826) );
INVx1_ASAP7_75t_L g845 ( .A(n_28), .Y(n_845) );
INVx1_ASAP7_75t_L g191 ( .A(n_29), .Y(n_191) );
NOR3xp33_ASAP7_75t_L g144 ( .A(n_30), .B(n_145), .C(n_336), .Y(n_144) );
INVx1_ASAP7_75t_SL g512 ( .A(n_30), .Y(n_512) );
OA21x2_ASAP7_75t_L g154 ( .A1(n_31), .A2(n_92), .B(n_155), .Y(n_154) );
OR2x2_ASAP7_75t_L g215 ( .A(n_31), .B(n_92), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_32), .B(n_245), .Y(n_563) );
INVxp67_ASAP7_75t_L g574 ( .A(n_33), .Y(n_574) );
AND2x2_ASAP7_75t_L g547 ( .A(n_34), .B(n_213), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_35), .B(n_166), .Y(n_252) );
AOI21xp5_ASAP7_75t_L g585 ( .A1(n_36), .A2(n_526), .B(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_37), .B(n_245), .Y(n_553) );
INVx1_ASAP7_75t_L g159 ( .A(n_38), .Y(n_159) );
AND2x2_ASAP7_75t_L g171 ( .A(n_38), .B(n_162), .Y(n_171) );
AND2x2_ASAP7_75t_L g182 ( .A(n_38), .B(n_165), .Y(n_182) );
OR2x6_ASAP7_75t_L g127 ( .A(n_39), .B(n_128), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g194 ( .A(n_40), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_41), .B(n_166), .Y(n_207) );
AOI22xp5_ASAP7_75t_L g221 ( .A1(n_42), .A2(n_187), .B1(n_222), .B2(n_226), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_43), .B(n_231), .Y(n_230) );
AOI22xp5_ASAP7_75t_L g601 ( .A1(n_45), .A2(n_84), .B1(n_157), .B2(n_526), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_46), .B(n_176), .Y(n_256) );
CKINVDCx20_ASAP7_75t_R g847 ( .A(n_47), .Y(n_847) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_48), .B(n_242), .Y(n_545) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_49), .B(n_153), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_50), .B(n_176), .Y(n_175) );
CKINVDCx5p33_ASAP7_75t_R g225 ( .A(n_51), .Y(n_225) );
AND2x2_ASAP7_75t_L g590 ( .A(n_52), .B(n_213), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_53), .B(n_213), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_55), .B(n_176), .Y(n_211) );
INVx1_ASAP7_75t_L g164 ( .A(n_56), .Y(n_164) );
INVx1_ASAP7_75t_L g178 ( .A(n_56), .Y(n_178) );
AND2x2_ASAP7_75t_L g212 ( .A(n_57), .B(n_213), .Y(n_212) );
AOI221xp5_ASAP7_75t_L g156 ( .A1(n_58), .A2(n_76), .B1(n_157), .B2(n_166), .C(n_172), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_59), .B(n_166), .Y(n_268) );
NAND2xp5_ASAP7_75t_SL g546 ( .A(n_60), .B(n_524), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_61), .B(n_187), .Y(n_201) );
AOI21xp5_ASAP7_75t_SL g264 ( .A1(n_62), .A2(n_157), .B(n_265), .Y(n_264) );
AND2x2_ASAP7_75t_L g538 ( .A(n_63), .B(n_213), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_64), .B(n_245), .Y(n_588) );
INVx1_ASAP7_75t_L g237 ( .A(n_65), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_66), .B(n_242), .Y(n_536) );
AND2x2_ASAP7_75t_SL g564 ( .A(n_67), .B(n_214), .Y(n_564) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_68), .A2(n_526), .B(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g210 ( .A(n_69), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_70), .B(n_245), .Y(n_529) );
AND2x2_ASAP7_75t_SL g602 ( .A(n_71), .B(n_153), .Y(n_602) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_72), .A2(n_157), .B(n_209), .Y(n_208) );
AOI22xp5_ASAP7_75t_L g815 ( .A1(n_73), .A2(n_131), .B1(n_816), .B2(n_820), .Y(n_815) );
INVx1_ASAP7_75t_L g162 ( .A(n_74), .Y(n_162) );
INVx1_ASAP7_75t_L g180 ( .A(n_74), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_75), .B(n_166), .Y(n_283) );
AND2x2_ASAP7_75t_L g257 ( .A(n_77), .B(n_186), .Y(n_257) );
INVx1_ASAP7_75t_L g238 ( .A(n_78), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_79), .A2(n_157), .B(n_254), .Y(n_253) );
CKINVDCx20_ASAP7_75t_R g136 ( .A(n_80), .Y(n_136) );
A2O1A1Ixp33_ASAP7_75t_L g227 ( .A1(n_81), .A2(n_157), .B(n_228), .C(n_232), .Y(n_227) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_82), .B(n_524), .Y(n_537) );
AOI22xp5_ASAP7_75t_L g600 ( .A1(n_83), .A2(n_87), .B1(n_166), .B2(n_524), .Y(n_600) );
NOR2xp33_ASAP7_75t_L g108 ( .A(n_85), .B(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g129 ( .A(n_85), .Y(n_129) );
AND2x2_ASAP7_75t_SL g262 ( .A(n_86), .B(n_186), .Y(n_262) );
AOI22xp5_ASAP7_75t_L g277 ( .A1(n_88), .A2(n_157), .B1(n_278), .B2(n_279), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_89), .B(n_242), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_90), .B(n_242), .Y(n_554) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_91), .A2(n_526), .B(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g266 ( .A(n_93), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_94), .B(n_245), .Y(n_535) );
AND2x2_ASAP7_75t_L g284 ( .A(n_95), .B(n_186), .Y(n_284) );
A2O1A1Ixp33_ASAP7_75t_L g188 ( .A1(n_96), .A2(n_189), .B(n_190), .C(n_193), .Y(n_188) );
INVxp67_ASAP7_75t_L g577 ( .A(n_97), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_98), .B(n_524), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_99), .B(n_245), .Y(n_544) );
AOI21xp5_ASAP7_75t_L g560 ( .A1(n_100), .A2(n_526), .B(n_561), .Y(n_560) );
BUFx2_ASAP7_75t_L g119 ( .A(n_101), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_102), .B(n_176), .Y(n_267) );
OAI22xp5_ASAP7_75t_SL g837 ( .A1(n_103), .A2(n_838), .B1(n_839), .B2(n_841), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_103), .Y(n_838) );
AOI21xp33_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_114), .B(n_846), .Y(n_104) );
INVx2_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx2_ASAP7_75t_L g848 ( .A(n_106), .Y(n_848) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
AND2x2_ASAP7_75t_SL g107 ( .A(n_108), .B(n_110), .Y(n_107) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_109), .B(n_129), .Y(n_128) );
INVx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
OA22x2_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_130), .B1(n_824), .B2(n_826), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_116), .B(n_120), .Y(n_115) );
CKINVDCx11_ASAP7_75t_R g116 ( .A(n_117), .Y(n_116) );
BUFx3_ASAP7_75t_L g825 ( .A(n_117), .Y(n_825) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_118), .Y(n_117) );
HB1xp67_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVxp67_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
AOI21xp33_ASAP7_75t_L g842 ( .A1(n_121), .A2(n_843), .B(n_844), .Y(n_842) );
NOR2xp33_ASAP7_75t_L g121 ( .A(n_122), .B(n_123), .Y(n_121) );
BUFx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
BUFx3_ASAP7_75t_L g831 ( .A(n_124), .Y(n_831) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_125), .B(n_126), .Y(n_124) );
AND2x6_ASAP7_75t_SL g142 ( .A(n_125), .B(n_127), .Y(n_142) );
OR2x6_ASAP7_75t_SL g814 ( .A(n_125), .B(n_126), .Y(n_814) );
OR2x2_ASAP7_75t_L g823 ( .A(n_125), .B(n_127), .Y(n_823) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_127), .Y(n_126) );
OAI21xp5_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_137), .B(n_815), .Y(n_130) );
INVxp33_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
OAI22xp5_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_143), .B1(n_514), .B2(n_812), .Y(n_138) );
CKINVDCx6p67_ASAP7_75t_R g139 ( .A(n_140), .Y(n_139) );
CKINVDCx11_ASAP7_75t_R g819 ( .A(n_140), .Y(n_819) );
INVx3_ASAP7_75t_SL g140 ( .A(n_141), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_142), .Y(n_141) );
AOI211xp5_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_407), .B(n_510), .C(n_513), .Y(n_143) );
AOI21xp5_ASAP7_75t_L g817 ( .A1(n_144), .A2(n_407), .B(n_510), .Y(n_817) );
INVx1_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_146), .A2(n_408), .B(n_512), .Y(n_513) );
NAND2xp5_ASAP7_75t_SL g835 ( .A(n_146), .B(n_485), .Y(n_835) );
NOR2x1_ASAP7_75t_L g146 ( .A(n_147), .B(n_314), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_148), .B(n_297), .Y(n_147) );
AOI221xp5_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_216), .B1(n_258), .B2(n_272), .C(n_287), .Y(n_148) );
AND2x2_ASAP7_75t_L g149 ( .A(n_150), .B(n_203), .Y(n_149) );
NAND2x1_ASAP7_75t_SL g323 ( .A(n_150), .B(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g350 ( .A(n_150), .B(n_320), .Y(n_350) );
HB1xp67_ASAP7_75t_L g396 ( .A(n_150), .Y(n_396) );
AND2x2_ASAP7_75t_L g404 ( .A(n_150), .B(n_405), .Y(n_404) );
INVx3_ASAP7_75t_L g508 ( .A(n_150), .Y(n_508) );
AND2x4_ASAP7_75t_L g150 ( .A(n_151), .B(n_184), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
HB1xp67_ASAP7_75t_L g286 ( .A(n_152), .Y(n_286) );
INVx1_ASAP7_75t_L g302 ( .A(n_152), .Y(n_302) );
AND2x4_ASAP7_75t_L g309 ( .A(n_152), .B(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g319 ( .A(n_152), .B(n_184), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_152), .B(n_305), .Y(n_346) );
INVx1_ASAP7_75t_L g357 ( .A(n_152), .Y(n_357) );
INVxp67_ASAP7_75t_L g391 ( .A(n_152), .Y(n_391) );
OA21x2_ASAP7_75t_L g152 ( .A1(n_153), .A2(n_156), .B(n_183), .Y(n_152) );
INVx2_ASAP7_75t_SL g232 ( .A(n_153), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g558 ( .A1(n_153), .A2(n_559), .B(n_560), .Y(n_558) );
BUFx4f_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx3_ASAP7_75t_L g187 ( .A(n_154), .Y(n_187) );
AND2x2_ASAP7_75t_SL g214 ( .A(n_155), .B(n_215), .Y(n_214) );
AND2x4_ASAP7_75t_L g226 ( .A(n_155), .B(n_215), .Y(n_226) );
INVxp67_ASAP7_75t_L g200 ( .A(n_157), .Y(n_200) );
AOI22xp5_ASAP7_75t_L g570 ( .A1(n_157), .A2(n_166), .B1(n_571), .B2(n_573), .Y(n_570) );
AND2x4_ASAP7_75t_L g157 ( .A(n_158), .B(n_163), .Y(n_157) );
NOR2x1p5_ASAP7_75t_L g158 ( .A(n_159), .B(n_160), .Y(n_158) );
INVx1_ASAP7_75t_L g282 ( .A(n_160), .Y(n_282) );
INVx3_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
OR2x6_ASAP7_75t_L g174 ( .A(n_161), .B(n_168), .Y(n_174) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
AND2x6_ASAP7_75t_L g242 ( .A(n_162), .B(n_177), .Y(n_242) );
AND2x6_ASAP7_75t_L g526 ( .A(n_163), .B(n_171), .Y(n_526) );
AND2x2_ASAP7_75t_L g163 ( .A(n_164), .B(n_165), .Y(n_163) );
INVx2_ASAP7_75t_L g168 ( .A(n_164), .Y(n_168) );
AND2x4_ASAP7_75t_L g245 ( .A(n_164), .B(n_179), .Y(n_245) );
HB1xp67_ASAP7_75t_L g169 ( .A(n_165), .Y(n_169) );
INVx1_ASAP7_75t_L g202 ( .A(n_166), .Y(n_202) );
AND2x4_ASAP7_75t_L g166 ( .A(n_167), .B(n_170), .Y(n_166) );
INVx1_ASAP7_75t_L g223 ( .A(n_167), .Y(n_223) );
AND2x2_ASAP7_75t_L g167 ( .A(n_168), .B(n_169), .Y(n_167) );
INVxp33_ASAP7_75t_L g281 ( .A(n_168), .Y(n_281) );
INVx1_ASAP7_75t_L g224 ( .A(n_170), .Y(n_224) );
BUFx3_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
O2A1O1Ixp33_ASAP7_75t_SL g172 ( .A1(n_173), .A2(n_174), .B(n_175), .C(n_181), .Y(n_172) );
INVxp67_ASAP7_75t_L g189 ( .A(n_174), .Y(n_189) );
O2A1O1Ixp33_ASAP7_75t_L g209 ( .A1(n_174), .A2(n_181), .B(n_210), .C(n_211), .Y(n_209) );
INVx2_ASAP7_75t_L g231 ( .A(n_174), .Y(n_231) );
OAI22xp5_ASAP7_75t_L g236 ( .A1(n_174), .A2(n_192), .B1(n_237), .B2(n_238), .Y(n_236) );
O2A1O1Ixp33_ASAP7_75t_SL g254 ( .A1(n_174), .A2(n_181), .B(n_255), .C(n_256), .Y(n_254) );
O2A1O1Ixp33_ASAP7_75t_L g265 ( .A1(n_174), .A2(n_181), .B(n_266), .C(n_267), .Y(n_265) );
INVx1_ASAP7_75t_L g192 ( .A(n_176), .Y(n_192) );
AND2x4_ASAP7_75t_L g524 ( .A(n_176), .B(n_182), .Y(n_524) );
AND2x4_ASAP7_75t_L g176 ( .A(n_177), .B(n_179), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_181), .A2(n_229), .B(n_230), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_181), .B(n_226), .Y(n_246) );
INVx1_ASAP7_75t_L g278 ( .A(n_181), .Y(n_278) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_181), .A2(n_528), .B(n_529), .Y(n_527) );
AOI21xp5_ASAP7_75t_L g534 ( .A1(n_181), .A2(n_535), .B(n_536), .Y(n_534) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_181), .A2(n_544), .B(n_545), .Y(n_543) );
AOI21xp5_ASAP7_75t_L g552 ( .A1(n_181), .A2(n_553), .B(n_554), .Y(n_552) );
AOI21xp5_ASAP7_75t_L g561 ( .A1(n_181), .A2(n_562), .B(n_563), .Y(n_561) );
AOI21xp5_ASAP7_75t_L g586 ( .A1(n_181), .A2(n_587), .B(n_588), .Y(n_586) );
INVx5_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
HB1xp67_ASAP7_75t_L g193 ( .A(n_182), .Y(n_193) );
INVx2_ASAP7_75t_L g274 ( .A(n_184), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_184), .B(n_205), .Y(n_290) );
INVx1_ASAP7_75t_L g308 ( .A(n_184), .Y(n_308) );
INVx1_ASAP7_75t_L g355 ( .A(n_184), .Y(n_355) );
OR2x2_ASAP7_75t_L g184 ( .A(n_185), .B(n_196), .Y(n_184) );
OAI22xp5_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_188), .B1(n_194), .B2(n_195), .Y(n_185) );
INVx3_ASAP7_75t_L g195 ( .A(n_186), .Y(n_195) );
INVx4_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_187), .B(n_198), .Y(n_197) );
AOI21x1_ASAP7_75t_L g583 ( .A1(n_187), .A2(n_584), .B(n_590), .Y(n_583) );
NOR2xp33_ASAP7_75t_L g190 ( .A(n_191), .B(n_192), .Y(n_190) );
NOR3xp33_ASAP7_75t_L g578 ( .A(n_192), .B(n_226), .C(n_579), .Y(n_578) );
AO21x2_ASAP7_75t_L g205 ( .A1(n_195), .A2(n_206), .B(n_212), .Y(n_205) );
AO21x2_ASAP7_75t_L g322 ( .A1(n_195), .A2(n_206), .B(n_212), .Y(n_322) );
OAI22xp5_ASAP7_75t_L g196 ( .A1(n_197), .A2(n_200), .B1(n_201), .B2(n_202), .Y(n_196) );
INVx1_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_203), .B(n_327), .Y(n_332) );
AND2x2_ASAP7_75t_L g344 ( .A(n_203), .B(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g363 ( .A(n_203), .B(n_309), .Y(n_363) );
INVx1_ASAP7_75t_L g372 ( .A(n_203), .Y(n_372) );
AND2x2_ASAP7_75t_L g420 ( .A(n_203), .B(n_319), .Y(n_420) );
OR2x2_ASAP7_75t_L g463 ( .A(n_203), .B(n_464), .Y(n_463) );
INVx3_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
AND2x4_ASAP7_75t_L g303 ( .A(n_204), .B(n_304), .Y(n_303) );
NAND2x1p5_ASAP7_75t_L g428 ( .A(n_204), .B(n_429), .Y(n_428) );
INVx3_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
AND2x2_ASAP7_75t_L g285 ( .A(n_205), .B(n_286), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_205), .B(n_305), .Y(n_383) );
HB1xp67_ASAP7_75t_L g406 ( .A(n_205), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_207), .B(n_208), .Y(n_206) );
CKINVDCx5p33_ASAP7_75t_R g250 ( .A(n_213), .Y(n_250) );
OA21x2_ASAP7_75t_L g550 ( .A1(n_213), .A2(n_551), .B(n_555), .Y(n_550) );
BUFx6f_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
INVx1_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
OR2x2_ASAP7_75t_L g217 ( .A(n_218), .B(n_247), .Y(n_217) );
NOR2x1_ASAP7_75t_L g387 ( .A(n_218), .B(n_342), .Y(n_387) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
AND2x2_ASAP7_75t_L g349 ( .A(n_219), .B(n_340), .Y(n_349) );
AND2x2_ASAP7_75t_L g219 ( .A(n_220), .B(n_233), .Y(n_219) );
INVx1_ASAP7_75t_L g269 ( .A(n_220), .Y(n_269) );
AND2x4_ASAP7_75t_L g295 ( .A(n_220), .B(n_296), .Y(n_295) );
INVx2_ASAP7_75t_L g299 ( .A(n_220), .Y(n_299) );
HB1xp67_ASAP7_75t_L g335 ( .A(n_220), .Y(n_335) );
AND2x2_ASAP7_75t_L g505 ( .A(n_220), .B(n_261), .Y(n_505) );
AND2x2_ASAP7_75t_L g220 ( .A(n_221), .B(n_227), .Y(n_220) );
NOR3xp33_ASAP7_75t_L g222 ( .A(n_223), .B(n_224), .C(n_225), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g263 ( .A1(n_226), .A2(n_264), .B(n_268), .Y(n_263) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_226), .A2(n_523), .B(n_525), .Y(n_522) );
NOR2xp33_ASAP7_75t_L g571 ( .A(n_226), .B(n_572), .Y(n_571) );
NOR2xp33_ASAP7_75t_L g573 ( .A(n_226), .B(n_574), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g576 ( .A(n_226), .B(n_577), .Y(n_576) );
AO21x2_ASAP7_75t_L g275 ( .A1(n_232), .A2(n_276), .B(n_284), .Y(n_275) );
AO21x2_ASAP7_75t_L g305 ( .A1(n_232), .A2(n_276), .B(n_284), .Y(n_305) );
AOI21x1_ASAP7_75t_L g598 ( .A1(n_232), .A2(n_599), .B(n_602), .Y(n_598) );
INVx3_ASAP7_75t_L g296 ( .A(n_233), .Y(n_296) );
INVx2_ASAP7_75t_L g313 ( .A(n_233), .Y(n_313) );
NOR2x1_ASAP7_75t_SL g330 ( .A(n_233), .B(n_261), .Y(n_330) );
AND2x2_ASAP7_75t_L g368 ( .A(n_233), .B(n_249), .Y(n_368) );
AND2x4_ASAP7_75t_L g233 ( .A(n_234), .B(n_235), .Y(n_233) );
OAI21xp5_ASAP7_75t_L g235 ( .A1(n_236), .A2(n_239), .B(n_246), .Y(n_235) );
OAI22xp5_ASAP7_75t_L g239 ( .A1(n_240), .A2(n_241), .B1(n_243), .B2(n_244), .Y(n_239) );
INVxp67_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
INVxp67_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
INVx1_ASAP7_75t_L g442 ( .A(n_247), .Y(n_442) );
HB1xp67_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
INVx2_ASAP7_75t_L g271 ( .A(n_248), .Y(n_271) );
INVx2_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
HB1xp67_ASAP7_75t_L g327 ( .A(n_249), .Y(n_327) );
INVx1_ASAP7_75t_L g340 ( .A(n_249), .Y(n_340) );
INVx1_ASAP7_75t_L g400 ( .A(n_249), .Y(n_400) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_249), .Y(n_419) );
OR2x2_ASAP7_75t_L g425 ( .A(n_249), .B(n_261), .Y(n_425) );
AND2x2_ASAP7_75t_L g469 ( .A(n_249), .B(n_296), .Y(n_469) );
AO21x2_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_251), .B(n_257), .Y(n_249) );
AO21x2_ASAP7_75t_L g531 ( .A1(n_250), .A2(n_532), .B(n_538), .Y(n_531) );
AO21x2_ASAP7_75t_L g540 ( .A1(n_250), .A2(n_541), .B(n_547), .Y(n_540) );
AO21x2_ASAP7_75t_L g679 ( .A1(n_250), .A2(n_541), .B(n_547), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_252), .B(n_253), .Y(n_251) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_260), .B(n_270), .Y(n_259) );
AND2x2_ASAP7_75t_L g311 ( .A(n_260), .B(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g465 ( .A(n_260), .B(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g470 ( .A(n_260), .Y(n_470) );
AND2x2_ASAP7_75t_L g482 ( .A(n_260), .B(n_368), .Y(n_482) );
AND2x4_ASAP7_75t_L g260 ( .A(n_261), .B(n_269), .Y(n_260) );
INVx4_ASAP7_75t_L g293 ( .A(n_261), .Y(n_293) );
INVx2_ASAP7_75t_L g343 ( .A(n_261), .Y(n_343) );
BUFx6f_ASAP7_75t_L g375 ( .A(n_261), .Y(n_375) );
NAND2xp5_ASAP7_75t_SL g443 ( .A(n_261), .B(n_401), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_261), .B(n_271), .Y(n_474) );
AND2x2_ASAP7_75t_L g500 ( .A(n_261), .B(n_313), .Y(n_500) );
OR2x6_ASAP7_75t_L g261 ( .A(n_262), .B(n_263), .Y(n_261) );
AND2x4_ASAP7_75t_L g402 ( .A(n_269), .B(n_293), .Y(n_402) );
AND2x2_ASAP7_75t_L g329 ( .A(n_270), .B(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g347 ( .A(n_270), .B(n_334), .Y(n_347) );
INVx1_ASAP7_75t_L g381 ( .A(n_270), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_270), .B(n_295), .Y(n_437) );
INVx3_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
HB1xp67_ASAP7_75t_L g361 ( .A(n_271), .Y(n_361) );
AOI22xp5_ASAP7_75t_L g497 ( .A1(n_272), .A2(n_354), .B1(n_498), .B2(n_501), .Y(n_497) );
AND2x4_ASAP7_75t_L g272 ( .A(n_273), .B(n_285), .Y(n_272) );
INVx1_ASAP7_75t_L g427 ( .A(n_273), .Y(n_427) );
AND2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
AND2x2_ASAP7_75t_L g301 ( .A(n_274), .B(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g450 ( .A(n_274), .B(n_322), .Y(n_450) );
NOR2xp67_ASAP7_75t_L g459 ( .A(n_274), .B(n_322), .Y(n_459) );
INVx2_ASAP7_75t_L g310 ( .A(n_275), .Y(n_310) );
AND2x4_ASAP7_75t_L g320 ( .A(n_275), .B(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g324 ( .A(n_275), .Y(n_324) );
NAND2xp5_ASAP7_75t_SL g276 ( .A(n_277), .B(n_283), .Y(n_276) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_286), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g287 ( .A(n_288), .B(n_291), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
NAND2x1p5_ASAP7_75t_L g389 ( .A(n_289), .B(n_390), .Y(n_389) );
AND2x2_ASAP7_75t_L g394 ( .A(n_289), .B(n_309), .Y(n_394) );
INVx2_ASAP7_75t_SL g289 ( .A(n_290), .Y(n_289) );
OR2x2_ASAP7_75t_L g432 ( .A(n_290), .B(n_346), .Y(n_432) );
INVxp33_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
BUFx2_ASAP7_75t_L g413 ( .A(n_292), .Y(n_413) );
NOR2x1_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
AND2x4_ASAP7_75t_SL g334 ( .A(n_293), .B(n_335), .Y(n_334) );
HB1xp67_ASAP7_75t_L g359 ( .A(n_293), .Y(n_359) );
INVx2_ASAP7_75t_L g423 ( .A(n_294), .Y(n_423) );
NAND2xp33_ASAP7_75t_SL g498 ( .A(n_294), .B(n_499), .Y(n_498) );
INVx4_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g364 ( .A(n_295), .B(n_343), .Y(n_364) );
AND2x2_ASAP7_75t_L g298 ( .A(n_296), .B(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g401 ( .A(n_296), .Y(n_401) );
AOI22xp5_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_300), .B1(n_306), .B2(n_311), .Y(n_297) );
AND2x2_ASAP7_75t_L g326 ( .A(n_298), .B(n_327), .Y(n_326) );
INVx2_ASAP7_75t_L g431 ( .A(n_298), .Y(n_431) );
INVx1_ASAP7_75t_L g380 ( .A(n_299), .Y(n_380) );
AOI22xp33_ASAP7_75t_SL g338 ( .A1(n_300), .A2(n_339), .B1(n_344), .B2(n_347), .Y(n_338) );
AND2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_303), .Y(n_300) );
INVx2_ASAP7_75t_L g464 ( .A(n_301), .Y(n_464) );
BUFx3_ASAP7_75t_L g429 ( .A(n_302), .Y(n_429) );
INVx1_ASAP7_75t_L g452 ( .A(n_303), .Y(n_452) );
AND2x2_ASAP7_75t_L g390 ( .A(n_304), .B(n_391), .Y(n_390) );
AND2x2_ASAP7_75t_L g457 ( .A(n_304), .B(n_322), .Y(n_457) );
INVx1_ASAP7_75t_L g491 ( .A(n_304), .Y(n_491) );
INVx2_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
OAI21xp33_ASAP7_75t_L g328 ( .A1(n_306), .A2(n_329), .B(n_331), .Y(n_328) );
OA21x2_ASAP7_75t_L g362 ( .A1(n_306), .A2(n_363), .B(n_364), .Y(n_362) );
AND2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_309), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g439 ( .A(n_308), .Y(n_439) );
AND2x2_ASAP7_75t_L g456 ( .A(n_308), .B(n_457), .Y(n_456) );
AND2x2_ASAP7_75t_L g446 ( .A(n_309), .B(n_405), .Y(n_446) );
AND2x2_ASAP7_75t_L g449 ( .A(n_309), .B(n_450), .Y(n_449) );
AND2x4_ASAP7_75t_L g458 ( .A(n_309), .B(n_459), .Y(n_458) );
AND2x2_ASAP7_75t_L g403 ( .A(n_312), .B(n_402), .Y(n_403) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
NOR2x1_ASAP7_75t_L g341 ( .A(n_313), .B(n_342), .Y(n_341) );
NAND2x1_ASAP7_75t_L g417 ( .A(n_313), .B(n_418), .Y(n_417) );
OAI21xp5_ASAP7_75t_SL g314 ( .A1(n_315), .A2(n_325), .B(n_328), .Y(n_314) );
INVxp67_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_317), .B(n_323), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
AOI22xp5_ASAP7_75t_L g369 ( .A1(n_318), .A2(n_334), .B1(n_359), .B2(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
INVx2_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
NOR2x1_ASAP7_75t_L g356 ( .A(n_322), .B(n_357), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_324), .B(n_354), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_324), .B(n_472), .Y(n_471) );
INVx2_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
BUFx2_ASAP7_75t_L g466 ( .A(n_327), .Y(n_466) );
AND2x2_ASAP7_75t_L g453 ( .A(n_330), .B(n_454), .Y(n_453) );
NOR2xp33_ASAP7_75t_R g331 ( .A(n_332), .B(n_333), .Y(n_331) );
INVx2_ASAP7_75t_SL g333 ( .A(n_334), .Y(n_333) );
NOR2xp33_ASAP7_75t_L g509 ( .A(n_334), .B(n_417), .Y(n_509) );
INVx1_ASAP7_75t_L g511 ( .A(n_336), .Y(n_511) );
OR3x2_ASAP7_75t_L g834 ( .A(n_336), .B(n_409), .C(n_835), .Y(n_834) );
NAND3x1_ASAP7_75t_SL g336 ( .A(n_337), .B(n_351), .C(n_365), .Y(n_336) );
AND2x2_ASAP7_75t_L g337 ( .A(n_338), .B(n_348), .Y(n_337) );
AOI22xp33_ASAP7_75t_L g448 ( .A1(n_339), .A2(n_449), .B1(n_451), .B2(n_453), .Y(n_448) );
AND2x2_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
NAND2xp5_ASAP7_75t_SL g393 ( .A(n_340), .B(n_379), .Y(n_393) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_345), .B(n_372), .Y(n_371) );
AND2x2_ASAP7_75t_L g414 ( .A(n_345), .B(n_355), .Y(n_414) );
AND2x2_ASAP7_75t_L g438 ( .A(n_345), .B(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_349), .B(n_350), .Y(n_348) );
OAI21xp5_ASAP7_75t_L g444 ( .A1(n_349), .A2(n_445), .B(n_446), .Y(n_444) );
AND2x2_ASAP7_75t_L g496 ( .A(n_349), .B(n_375), .Y(n_496) );
AOI22xp5_ASAP7_75t_L g502 ( .A1(n_350), .A2(n_503), .B1(n_506), .B2(n_509), .Y(n_502) );
AOI21xp5_ASAP7_75t_SL g351 ( .A1(n_352), .A2(n_358), .B(n_362), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g354 ( .A(n_355), .B(n_356), .Y(n_354) );
BUFx2_ASAP7_75t_L g472 ( .A(n_355), .Y(n_472) );
INVx1_ASAP7_75t_SL g479 ( .A(n_355), .Y(n_479) );
HB1xp67_ASAP7_75t_L g440 ( .A(n_356), .Y(n_440) );
NOR2xp33_ASAP7_75t_L g358 ( .A(n_359), .B(n_360), .Y(n_358) );
HB1xp67_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
NOR2x1_ASAP7_75t_L g365 ( .A(n_366), .B(n_385), .Y(n_365) );
OAI21xp5_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_369), .B(n_373), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g374 ( .A(n_368), .B(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_SL g460 ( .A(n_368), .B(n_379), .Y(n_460) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
OAI21xp5_ASAP7_75t_SL g373 ( .A1(n_374), .A2(n_376), .B(n_382), .Y(n_373) );
OR2x6_ASAP7_75t_L g430 ( .A(n_375), .B(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_378), .B(n_381), .Y(n_377) );
INVx2_ASAP7_75t_SL g378 ( .A(n_379), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
NOR2xp33_ASAP7_75t_L g382 ( .A(n_383), .B(n_384), .Y(n_382) );
INVx1_ASAP7_75t_L g480 ( .A(n_383), .Y(n_480) );
OR2x2_ASAP7_75t_L g507 ( .A(n_383), .B(n_508), .Y(n_507) );
NOR2xp33_ASAP7_75t_L g451 ( .A(n_384), .B(n_452), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_386), .B(n_395), .Y(n_385) );
AOI22xp5_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_388), .B1(n_392), .B2(n_394), .Y(n_386) );
INVx3_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
HB1xp67_ASAP7_75t_L g487 ( .A(n_389), .Y(n_487) );
INVxp67_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
AOI22xp5_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_397), .B1(n_403), .B2(n_404), .Y(n_395) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_399), .B(n_402), .Y(n_398) );
AND2x4_ASAP7_75t_SL g399 ( .A(n_400), .B(n_401), .Y(n_399) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
AND2x2_ASAP7_75t_L g407 ( .A(n_408), .B(n_483), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
NAND3xp33_ASAP7_75t_L g409 ( .A(n_410), .B(n_433), .C(n_461), .Y(n_409) );
NOR2xp33_ASAP7_75t_L g410 ( .A(n_411), .B(n_421), .Y(n_410) );
NAND2xp5_ASAP7_75t_SL g411 ( .A(n_412), .B(n_415), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_413), .B(n_414), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_416), .B(n_420), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g454 ( .A(n_418), .Y(n_454) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
OAI22xp33_ASAP7_75t_SL g421 ( .A1(n_422), .A2(n_426), .B1(n_430), .B2(n_432), .Y(n_421) );
NAND2x1_ASAP7_75t_L g422 ( .A(n_423), .B(n_424), .Y(n_422) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_423), .B(n_505), .Y(n_504) );
INVx2_ASAP7_75t_SL g424 ( .A(n_425), .Y(n_424) );
NOR2x1_ASAP7_75t_L g501 ( .A(n_425), .B(n_431), .Y(n_501) );
OR2x2_ASAP7_75t_L g426 ( .A(n_427), .B(n_428), .Y(n_426) );
INVx3_ASAP7_75t_L g489 ( .A(n_429), .Y(n_489) );
INVx2_ASAP7_75t_L g493 ( .A(n_430), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g433 ( .A(n_434), .B(n_447), .Y(n_433) );
NAND2xp5_ASAP7_75t_SL g434 ( .A(n_435), .B(n_444), .Y(n_434) );
AOI22xp33_ASAP7_75t_SL g435 ( .A1(n_436), .A2(n_438), .B1(n_440), .B2(n_441), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
NOR2x1_ASAP7_75t_L g441 ( .A(n_442), .B(n_443), .Y(n_441) );
INVxp67_ASAP7_75t_SL g445 ( .A(n_443), .Y(n_445) );
NAND2xp5_ASAP7_75t_SL g447 ( .A(n_448), .B(n_455), .Y(n_447) );
NAND2x1p5_ASAP7_75t_L g490 ( .A(n_450), .B(n_491), .Y(n_490) );
OAI21xp5_ASAP7_75t_L g455 ( .A1(n_456), .A2(n_458), .B(n_460), .Y(n_455) );
INVx1_ASAP7_75t_L g475 ( .A(n_458), .Y(n_475) );
AOI211xp5_ASAP7_75t_L g461 ( .A1(n_462), .A2(n_465), .B(n_467), .C(n_476), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
OAI211xp5_ASAP7_75t_L g494 ( .A1(n_464), .A2(n_495), .B(n_497), .C(n_502), .Y(n_494) );
OAI22xp5_ASAP7_75t_L g467 ( .A1(n_468), .A2(n_471), .B1(n_473), .B2(n_475), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_469), .B(n_470), .Y(n_468) );
HB1xp67_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_477), .B(n_481), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_479), .B(n_480), .Y(n_478) );
INVxp67_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
AOI21xp5_ASAP7_75t_SL g510 ( .A1(n_483), .A2(n_511), .B(n_512), .Y(n_510) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
NOR2xp67_ASAP7_75t_L g485 ( .A(n_486), .B(n_494), .Y(n_485) );
AOI21xp33_ASAP7_75t_SL g486 ( .A1(n_487), .A2(n_488), .B(n_492), .Y(n_486) );
OR2x2_ASAP7_75t_L g488 ( .A(n_489), .B(n_490), .Y(n_488) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVxp33_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
NOR2xp33_ASAP7_75t_L g818 ( .A(n_513), .B(n_819), .Y(n_818) );
AO22x2_ASAP7_75t_L g816 ( .A1(n_514), .A2(n_813), .B1(n_817), .B2(n_818), .Y(n_816) );
INVx4_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
AND2x4_ASAP7_75t_L g515 ( .A(n_516), .B(n_723), .Y(n_515) );
NOR3xp33_ASAP7_75t_L g516 ( .A(n_517), .B(n_645), .C(n_695), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_518), .B(n_612), .Y(n_517) );
AOI221xp5_ASAP7_75t_L g518 ( .A1(n_519), .A2(n_548), .B1(n_565), .B2(n_595), .C(n_604), .Y(n_518) );
INVx1_ASAP7_75t_SL g694 ( .A(n_519), .Y(n_694) );
AND2x4_ASAP7_75t_SL g519 ( .A(n_520), .B(n_530), .Y(n_519) );
INVx2_ASAP7_75t_L g616 ( .A(n_520), .Y(n_616) );
OR2x2_ASAP7_75t_L g638 ( .A(n_520), .B(n_629), .Y(n_638) );
HB1xp67_ASAP7_75t_L g653 ( .A(n_520), .Y(n_653) );
INVx5_ASAP7_75t_L g660 ( .A(n_520), .Y(n_660) );
AND2x4_ASAP7_75t_L g666 ( .A(n_520), .B(n_540), .Y(n_666) );
AND2x2_ASAP7_75t_SL g669 ( .A(n_520), .B(n_597), .Y(n_669) );
OR2x2_ASAP7_75t_L g678 ( .A(n_520), .B(n_679), .Y(n_678) );
AND2x2_ASAP7_75t_L g685 ( .A(n_520), .B(n_531), .Y(n_685) );
AND2x2_ASAP7_75t_L g786 ( .A(n_520), .B(n_539), .Y(n_786) );
OR2x6_ASAP7_75t_L g520 ( .A(n_521), .B(n_522), .Y(n_520) );
INVx3_ASAP7_75t_SL g637 ( .A(n_530), .Y(n_637) );
AND2x2_ASAP7_75t_L g681 ( .A(n_530), .B(n_597), .Y(n_681) );
OAI21xp5_ASAP7_75t_L g684 ( .A1(n_530), .A2(n_685), .B(n_686), .Y(n_684) );
AND2x2_ASAP7_75t_L g722 ( .A(n_530), .B(n_660), .Y(n_722) );
AND2x4_ASAP7_75t_L g530 ( .A(n_531), .B(n_539), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_531), .B(n_540), .Y(n_603) );
OR2x2_ASAP7_75t_L g607 ( .A(n_531), .B(n_540), .Y(n_607) );
INVx1_ASAP7_75t_L g615 ( .A(n_531), .Y(n_615) );
HB1xp67_ASAP7_75t_L g627 ( .A(n_531), .Y(n_627) );
INVx2_ASAP7_75t_L g635 ( .A(n_531), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_531), .B(n_660), .Y(n_659) );
AND2x2_ASAP7_75t_L g744 ( .A(n_531), .B(n_629), .Y(n_744) );
AND2x2_ASAP7_75t_L g759 ( .A(n_531), .B(n_597), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_533), .B(n_537), .Y(n_532) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g628 ( .A(n_540), .B(n_629), .Y(n_628) );
HB1xp67_ASAP7_75t_L g699 ( .A(n_540), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_542), .B(n_546), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_548), .B(n_752), .Y(n_751) );
NOR2x1p5_ASAP7_75t_L g548 ( .A(n_549), .B(n_556), .Y(n_548) );
BUFx3_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g581 ( .A(n_550), .B(n_582), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_550), .B(n_557), .Y(n_610) );
INVx1_ASAP7_75t_L g620 ( .A(n_550), .Y(n_620) );
INVx2_ASAP7_75t_L g643 ( .A(n_550), .Y(n_643) );
INVx2_ASAP7_75t_L g649 ( .A(n_550), .Y(n_649) );
HB1xp67_ASAP7_75t_L g719 ( .A(n_550), .Y(n_719) );
OR2x2_ASAP7_75t_L g750 ( .A(n_550), .B(n_557), .Y(n_750) );
OR2x2_ASAP7_75t_L g766 ( .A(n_556), .B(n_767), .Y(n_766) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
AND2x4_ASAP7_75t_SL g568 ( .A(n_557), .B(n_569), .Y(n_568) );
AND2x4_ASAP7_75t_L g593 ( .A(n_557), .B(n_594), .Y(n_593) );
OR2x2_ASAP7_75t_L g630 ( .A(n_557), .B(n_631), .Y(n_630) );
OR2x2_ASAP7_75t_L g642 ( .A(n_557), .B(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g655 ( .A(n_557), .B(n_621), .Y(n_655) );
OR2x2_ASAP7_75t_L g663 ( .A(n_557), .B(n_569), .Y(n_663) );
INVx2_ASAP7_75t_L g690 ( .A(n_557), .Y(n_690) );
INVx1_ASAP7_75t_L g708 ( .A(n_557), .Y(n_708) );
NOR2xp33_ASAP7_75t_R g741 ( .A(n_557), .B(n_582), .Y(n_741) );
OR2x6_ASAP7_75t_L g557 ( .A(n_558), .B(n_564), .Y(n_557) );
NAND2xp5_ASAP7_75t_SL g565 ( .A(n_566), .B(n_591), .Y(n_565) );
OAI22xp5_ASAP7_75t_L g632 ( .A1(n_566), .A2(n_633), .B1(n_636), .B2(n_639), .Y(n_632) );
OR2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_580), .Y(n_566) );
INVx1_ASAP7_75t_SL g567 ( .A(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g647 ( .A(n_568), .B(n_648), .Y(n_647) );
AND2x2_ASAP7_75t_L g682 ( .A(n_568), .B(n_683), .Y(n_682) );
AND2x4_ASAP7_75t_L g761 ( .A(n_568), .B(n_739), .Y(n_761) );
INVx3_ASAP7_75t_L g594 ( .A(n_569), .Y(n_594) );
AND2x4_ASAP7_75t_L g621 ( .A(n_569), .B(n_622), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_569), .B(n_582), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_569), .B(n_643), .Y(n_688) );
AND2x2_ASAP7_75t_L g693 ( .A(n_569), .B(n_690), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_569), .B(n_581), .Y(n_730) );
INVx1_ASAP7_75t_L g800 ( .A(n_569), .Y(n_800) );
NAND2xp5_ASAP7_75t_L g811 ( .A(n_569), .B(n_718), .Y(n_811) );
AND2x4_ASAP7_75t_L g569 ( .A(n_570), .B(n_575), .Y(n_569) );
INVx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g592 ( .A(n_582), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_582), .B(n_594), .Y(n_611) );
INVx2_ASAP7_75t_L g622 ( .A(n_582), .Y(n_622) );
AND2x2_ASAP7_75t_L g648 ( .A(n_582), .B(n_649), .Y(n_648) );
OR2x2_ASAP7_75t_L g664 ( .A(n_582), .B(n_643), .Y(n_664) );
HB1xp67_ASAP7_75t_L g683 ( .A(n_582), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_582), .B(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g753 ( .A(n_582), .Y(n_753) );
INVx3_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_585), .B(n_589), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_592), .B(n_620), .Y(n_631) );
AOI221x1_ASAP7_75t_SL g725 ( .A1(n_593), .A2(n_726), .B1(n_729), .B2(n_731), .C(n_735), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_593), .B(n_774), .Y(n_773) );
AND2x2_ASAP7_75t_L g783 ( .A(n_593), .B(n_648), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g804 ( .A(n_593), .B(n_805), .Y(n_804) );
OR2x2_ASAP7_75t_L g714 ( .A(n_594), .B(n_642), .Y(n_714) );
AND2x2_ASAP7_75t_L g752 ( .A(n_594), .B(n_753), .Y(n_752) );
INVx1_ASAP7_75t_SL g595 ( .A(n_596), .Y(n_595) );
OR2x2_ASAP7_75t_L g596 ( .A(n_597), .B(n_603), .Y(n_596) );
AND2x2_ASAP7_75t_L g605 ( .A(n_597), .B(n_606), .Y(n_605) );
INVx2_ASAP7_75t_L g700 ( .A(n_597), .Y(n_700) );
NOR2xp33_ASAP7_75t_L g705 ( .A(n_597), .B(n_616), .Y(n_705) );
AND2x4_ASAP7_75t_L g734 ( .A(n_597), .B(n_635), .Y(n_734) );
NAND2xp5_ASAP7_75t_SL g770 ( .A(n_597), .B(n_666), .Y(n_770) );
OR2x2_ASAP7_75t_L g788 ( .A(n_597), .B(n_719), .Y(n_788) );
NOR2xp33_ASAP7_75t_L g798 ( .A(n_597), .B(n_679), .Y(n_798) );
BUFx6f_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx2_ASAP7_75t_L g629 ( .A(n_598), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_600), .B(n_601), .Y(n_599) );
INVx1_ASAP7_75t_L g654 ( .A(n_603), .Y(n_654) );
OAI22xp5_ASAP7_75t_L g661 ( .A1(n_603), .A2(n_662), .B1(n_665), .B2(n_667), .Y(n_661) );
AND2x2_ASAP7_75t_L g604 ( .A(n_605), .B(n_608), .Y(n_604) );
INVx2_ASAP7_75t_L g617 ( .A(n_605), .Y(n_617) );
AND2x2_ASAP7_75t_L g756 ( .A(n_606), .B(n_616), .Y(n_756) );
AND2x2_ASAP7_75t_L g802 ( .A(n_606), .B(n_669), .Y(n_802) );
AND2x2_ASAP7_75t_L g807 ( .A(n_606), .B(n_658), .Y(n_807) );
INVx2_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
AOI32xp33_ASAP7_75t_L g776 ( .A1(n_608), .A2(n_678), .A3(n_758), .B1(n_777), .B2(n_779), .Y(n_776) );
INVx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
OR2x2_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .Y(n_609) );
INVx1_ASAP7_75t_L g644 ( .A(n_611), .Y(n_644) );
AOI211xp5_ASAP7_75t_SL g612 ( .A1(n_613), .A2(n_618), .B(n_623), .C(n_632), .Y(n_612) );
OAI21xp5_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_616), .B(n_617), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_615), .B(n_666), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_616), .B(n_634), .Y(n_633) );
INVx2_ASAP7_75t_L g796 ( .A(n_616), .Y(n_796) );
AND2x2_ASAP7_75t_L g706 ( .A(n_618), .B(n_707), .Y(n_706) );
AND2x2_ASAP7_75t_SL g618 ( .A(n_619), .B(n_621), .Y(n_618) );
HB1xp67_ASAP7_75t_L g806 ( .A(n_619), .Y(n_806) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVxp67_ASAP7_75t_SL g675 ( .A(n_620), .Y(n_675) );
HB1xp67_ASAP7_75t_L g775 ( .A(n_620), .Y(n_775) );
INVx1_ASAP7_75t_L g672 ( .A(n_621), .Y(n_672) );
AND2x2_ASAP7_75t_L g738 ( .A(n_621), .B(n_739), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_621), .B(n_749), .Y(n_778) );
NOR2xp33_ASAP7_75t_L g623 ( .A(n_624), .B(n_630), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
OAI21xp33_ASAP7_75t_L g704 ( .A1(n_625), .A2(n_705), .B(n_706), .Y(n_704) );
AND2x2_ASAP7_75t_SL g625 ( .A(n_626), .B(n_628), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g634 ( .A(n_629), .B(n_635), .Y(n_634) );
BUFx2_ASAP7_75t_L g658 ( .A(n_629), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_634), .B(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g765 ( .A(n_634), .Y(n_765) );
AND2x2_ASAP7_75t_L g795 ( .A(n_634), .B(n_796), .Y(n_795) );
HB1xp67_ASAP7_75t_L g772 ( .A(n_635), .Y(n_772) );
OR2x2_ASAP7_75t_L g636 ( .A(n_637), .B(n_638), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_637), .B(n_785), .Y(n_784) );
INVx1_ASAP7_75t_SL g712 ( .A(n_638), .Y(n_712) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
AND2x4_ASAP7_75t_L g640 ( .A(n_641), .B(n_644), .Y(n_640) );
INVx2_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
OR2x2_ASAP7_75t_L g671 ( .A(n_642), .B(n_672), .Y(n_671) );
HB1xp67_ASAP7_75t_L g739 ( .A(n_643), .Y(n_739) );
AND2x2_ASAP7_75t_L g748 ( .A(n_644), .B(n_749), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_646), .B(n_668), .Y(n_645) );
AOI221xp5_ASAP7_75t_L g646 ( .A1(n_647), .A2(n_650), .B1(n_655), .B2(n_656), .C(n_661), .Y(n_646) );
INVx1_ASAP7_75t_L g767 ( .A(n_648), .Y(n_767) );
INVxp33_ASAP7_75t_SL g799 ( .A(n_648), .Y(n_799) );
AOI21xp5_ASAP7_75t_L g745 ( .A1(n_650), .A2(n_746), .B(n_754), .Y(n_745) );
INVx2_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
NAND2xp5_ASAP7_75t_SL g651 ( .A(n_652), .B(n_654), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_654), .B(n_712), .Y(n_711) );
INVx2_ASAP7_75t_L g667 ( .A(n_655), .Y(n_667) );
AND2x2_ASAP7_75t_L g702 ( .A(n_655), .B(n_703), .Y(n_702) );
AND2x2_ASAP7_75t_L g721 ( .A(n_655), .B(n_722), .Y(n_721) );
AOI22xp33_ASAP7_75t_SL g782 ( .A1(n_655), .A2(n_783), .B1(n_784), .B2(n_787), .Y(n_782) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
OR2x2_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .Y(n_657) );
OR2x2_ASAP7_75t_L g677 ( .A(n_658), .B(n_678), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_658), .B(n_666), .Y(n_716) );
AND2x4_ASAP7_75t_L g733 ( .A(n_660), .B(n_679), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_660), .B(n_734), .Y(n_780) );
AND2x2_ASAP7_75t_L g792 ( .A(n_660), .B(n_744), .Y(n_792) );
NAND2xp33_ASAP7_75t_L g777 ( .A(n_662), .B(n_778), .Y(n_777) );
OR2x2_ASAP7_75t_L g662 ( .A(n_663), .B(n_664), .Y(n_662) );
INVx1_ASAP7_75t_SL g720 ( .A(n_663), .Y(n_720) );
INVx1_ASAP7_75t_L g791 ( .A(n_664), .Y(n_791) );
INVx2_ASAP7_75t_SL g743 ( .A(n_666), .Y(n_743) );
AOI211xp5_ASAP7_75t_SL g668 ( .A1(n_669), .A2(n_670), .B(n_673), .C(n_691), .Y(n_668) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
OAI211xp5_ASAP7_75t_L g673 ( .A1(n_674), .A2(n_677), .B(n_680), .C(n_684), .Y(n_673) );
OR2x6_ASAP7_75t_SL g674 ( .A(n_675), .B(n_676), .Y(n_674) );
INVx1_ASAP7_75t_L g703 ( .A(n_675), .Y(n_703) );
INVx1_ASAP7_75t_SL g728 ( .A(n_678), .Y(n_728) );
NOR2xp33_ASAP7_75t_L g787 ( .A(n_678), .B(n_788), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_681), .B(n_682), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_683), .B(n_693), .Y(n_692) );
INVx2_ASAP7_75t_SL g686 ( .A(n_687), .Y(n_686) );
OAI22xp33_ASAP7_75t_L g769 ( .A1(n_687), .A2(n_770), .B1(n_771), .B2(n_773), .Y(n_769) );
OR2x2_ASAP7_75t_L g687 ( .A(n_688), .B(n_689), .Y(n_687) );
NOR2xp33_ASAP7_75t_L g691 ( .A(n_692), .B(n_694), .Y(n_691) );
OAI211xp5_ASAP7_75t_SL g695 ( .A1(n_696), .A2(n_701), .B(n_704), .C(n_709), .Y(n_695) );
INVxp67_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
NOR2xp33_ASAP7_75t_L g697 ( .A(n_698), .B(n_700), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
AOI221xp5_ASAP7_75t_L g709 ( .A1(n_710), .A2(n_713), .B1(n_715), .B2(n_717), .C(n_721), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_SL g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
AND2x2_ASAP7_75t_L g717 ( .A(n_718), .B(n_720), .Y(n_717) );
HB1xp67_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
AOI222xp33_ASAP7_75t_L g801 ( .A1(n_720), .A2(n_802), .B1(n_803), .B2(n_807), .C1(n_808), .C2(n_810), .Y(n_801) );
INVx2_ASAP7_75t_L g736 ( .A(n_722), .Y(n_736) );
NOR3xp33_ASAP7_75t_L g723 ( .A(n_724), .B(n_762), .C(n_781), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_725), .B(n_745), .Y(n_724) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVxp67_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_733), .B(n_734), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_733), .B(n_772), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_734), .B(n_796), .Y(n_809) );
OAI22xp33_ASAP7_75t_L g735 ( .A1(n_736), .A2(n_737), .B1(n_740), .B2(n_742), .Y(n_735) );
INVx1_ASAP7_75t_SL g737 ( .A(n_738), .Y(n_737) );
INVxp33_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_743), .B(n_744), .Y(n_742) );
NOR2xp33_ASAP7_75t_L g764 ( .A(n_743), .B(n_765), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_747), .B(n_751), .Y(n_746) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_SL g749 ( .A(n_750), .Y(n_749) );
OAI22xp5_ASAP7_75t_L g754 ( .A1(n_751), .A2(n_755), .B1(n_757), .B2(n_760), .Y(n_754) );
INVx2_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
BUFx2_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
CKINVDCx16_ASAP7_75t_R g760 ( .A(n_761), .Y(n_760) );
OAI211xp5_ASAP7_75t_SL g762 ( .A1(n_763), .A2(n_766), .B(n_768), .C(n_776), .Y(n_762) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
INVxp67_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
INVx1_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
NAND3xp33_ASAP7_75t_L g781 ( .A(n_782), .B(n_789), .C(n_801), .Y(n_781) );
INVx2_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
OAI21xp5_ASAP7_75t_L g789 ( .A1(n_790), .A2(n_793), .B(n_800), .Y(n_789) );
AND2x2_ASAP7_75t_L g790 ( .A(n_791), .B(n_792), .Y(n_790) );
AOI21xp5_ASAP7_75t_L g793 ( .A1(n_794), .A2(n_797), .B(n_799), .Y(n_793) );
INVx1_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
INVx1_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
INVx1_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
INVx1_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
INVx1_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
INVx1_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
CKINVDCx5p33_ASAP7_75t_R g812 ( .A(n_813), .Y(n_812) );
CKINVDCx11_ASAP7_75t_R g813 ( .A(n_814), .Y(n_813) );
CKINVDCx5p33_ASAP7_75t_R g820 ( .A(n_821), .Y(n_820) );
CKINVDCx5p33_ASAP7_75t_R g821 ( .A(n_822), .Y(n_821) );
INVx3_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
CKINVDCx5p33_ASAP7_75t_R g824 ( .A(n_825), .Y(n_824) );
NAND2xp5_ASAP7_75t_L g827 ( .A(n_828), .B(n_832), .Y(n_827) );
INVx1_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
NOR2xp33_ASAP7_75t_L g844 ( .A(n_829), .B(n_845), .Y(n_844) );
BUFx2_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
CKINVDCx20_ASAP7_75t_R g830 ( .A(n_831), .Y(n_830) );
INVxp67_ASAP7_75t_L g843 ( .A(n_832), .Y(n_843) );
AOI22x1_ASAP7_75t_L g832 ( .A1(n_833), .A2(n_834), .B1(n_836), .B2(n_837), .Y(n_832) );
INVx2_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
INVx1_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
INVx1_ASAP7_75t_L g841 ( .A(n_839), .Y(n_841) );
NOR2xp33_ASAP7_75t_L g846 ( .A(n_847), .B(n_848), .Y(n_846) );
endmodule