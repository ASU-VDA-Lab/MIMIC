module fake_jpeg_3961_n_91 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_91);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_91;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

CKINVDCx14_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

AND2x2_ASAP7_75t_L g16 ( 
.A(n_1),
.B(n_0),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_4),
.B(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_11),
.B(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_31),
.Y(n_34)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_25),
.B(n_31),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_19),
.A2(n_11),
.B1(n_10),
.B2(n_7),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_26),
.A2(n_27),
.B1(n_3),
.B2(n_4),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g27 ( 
.A1(n_16),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_16),
.B(n_21),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_28),
.B(n_29),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_18),
.Y(n_29)
);

CKINVDCx12_ASAP7_75t_R g30 ( 
.A(n_17),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_30),
.B(n_22),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

HB1xp67_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_33),
.B(n_6),
.Y(n_52)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_2),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_41),
.Y(n_59)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_40),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_24),
.B(n_2),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_29),
.A2(n_15),
.B1(n_20),
.B2(n_14),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_42),
.A2(n_40),
.B1(n_37),
.B2(n_51),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_3),
.Y(n_43)
);

XOR2xp5_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_47),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_32),
.A2(n_23),
.B1(n_13),
.B2(n_12),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_44),
.A2(n_6),
.B1(n_7),
.B2(n_42),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

O2A1O1Ixp33_ASAP7_75t_L g63 ( 
.A1(n_46),
.A2(n_35),
.B(n_41),
.C(n_47),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_3),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_30),
.B(n_14),
.C(n_23),
.Y(n_48)
);

XOR2xp5_ASAP7_75t_L g65 ( 
.A(n_48),
.B(n_51),
.Y(n_65)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_SL g64 ( 
.A(n_50),
.B(n_53),
.C(n_39),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_28),
.B(n_5),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_52),
.A2(n_45),
.B(n_43),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

CKINVDCx14_ASAP7_75t_R g71 ( 
.A(n_54),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_58),
.A2(n_62),
.B1(n_63),
.B2(n_49),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_35),
.A2(n_46),
.B1(n_36),
.B2(n_48),
.Y(n_62)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_67),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_34),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_50),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_68),
.B(n_70),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g69 ( 
.A(n_65),
.B(n_38),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_74),
.C(n_75),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_38),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_53),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_58),
.C(n_56),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_68),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_76),
.B(n_78),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_77),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_72),
.B(n_61),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_73),
.A2(n_60),
.B(n_57),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_76),
.B(n_67),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_84),
.B(n_80),
.Y(n_86)
);

AOI322xp5_ASAP7_75t_L g89 ( 
.A1(n_86),
.A2(n_87),
.A3(n_88),
.B1(n_74),
.B2(n_79),
.C1(n_84),
.C2(n_81),
.Y(n_89)
);

AOI322xp5_ASAP7_75t_L g87 ( 
.A1(n_83),
.A2(n_79),
.A3(n_81),
.B1(n_71),
.B2(n_69),
.C1(n_75),
.C2(n_80),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_85),
.B(n_82),
.Y(n_88)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_89),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_90),
.Y(n_91)
);


endmodule