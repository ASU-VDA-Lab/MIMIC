module fake_jpeg_5476_n_54 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_54);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_54;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_1),
.Y(n_7)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_0),
.B(n_5),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

INVx3_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx5_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g16 ( 
.A(n_7),
.B(n_1),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_16),
.B(n_17),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g17 ( 
.A(n_7),
.B(n_15),
.Y(n_17)
);

A2O1A1Ixp33_ASAP7_75t_L g18 ( 
.A1(n_11),
.A2(n_4),
.B(n_5),
.C(n_6),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_18),
.B(n_20),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g20 ( 
.A(n_15),
.B(n_4),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_23),
.Y(n_25)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_24),
.A2(n_11),
.B1(n_8),
.B2(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

OAI32xp33_ASAP7_75t_L g28 ( 
.A1(n_18),
.A2(n_8),
.A3(n_10),
.B1(n_12),
.B2(n_14),
.Y(n_28)
);

NAND3xp33_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_33),
.C(n_34),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_16),
.B(n_14),
.C(n_6),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_34),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_24),
.A2(n_23),
.B1(n_21),
.B2(n_17),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_26),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_35),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_37),
.A2(n_28),
.B1(n_33),
.B2(n_29),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_32),
.B(n_22),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_40),
.Y(n_48)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_20),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

NOR3xp33_ASAP7_75t_SL g44 ( 
.A(n_42),
.B(n_19),
.C(n_33),
.Y(n_44)
);

AOI322xp5_ASAP7_75t_L g49 ( 
.A1(n_43),
.A2(n_25),
.A3(n_39),
.B1(n_40),
.B2(n_44),
.C1(n_45),
.C2(n_46),
.Y(n_49)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_36),
.A2(n_39),
.B1(n_27),
.B2(n_42),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_47),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_49),
.A2(n_50),
.B(n_36),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_51),
.A2(n_48),
.B(n_47),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g54 ( 
.A(n_52),
.B(n_53),
.Y(n_54)
);


endmodule