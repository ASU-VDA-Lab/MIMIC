module fake_netlist_5_2155_n_1634 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1634);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1634;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_775;
wire n_219;
wire n_157;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_284;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_254;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_433;
wire n_314;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_233;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_833;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1419;
wire n_338;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_253;
wire n_1116;
wire n_1212;
wire n_1541;
wire n_172;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_768;
wire n_1475;
wire n_1302;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_462;
wire n_1193;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1540;
wire n_229;
wire n_437;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_97),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_130),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_59),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_151),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_31),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_147),
.Y(n_162)
);

BUFx10_ASAP7_75t_L g163 ( 
.A(n_77),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_113),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_19),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_120),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_36),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_1),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_132),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_44),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_68),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_118),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_110),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_105),
.Y(n_174)
);

INVx4_ASAP7_75t_R g175 ( 
.A(n_19),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_52),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_115),
.Y(n_177)
);

INVxp33_ASAP7_75t_SL g178 ( 
.A(n_91),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_64),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_22),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_1),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_52),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_87),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_143),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_156),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_140),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_79),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_83),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_116),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_20),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_102),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_107),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_128),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_119),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_71),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_137),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_98),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_114),
.Y(n_198)
);

BUFx10_ASAP7_75t_L g199 ( 
.A(n_126),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_89),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_95),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_149),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_134),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_58),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_33),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_55),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_100),
.Y(n_207)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_31),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_150),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_7),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_57),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_92),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_60),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_67),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_112),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_17),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_7),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_81),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_36),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_73),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_104),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_65),
.Y(n_222)
);

INVxp67_ASAP7_75t_SL g223 ( 
.A(n_123),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_78),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g225 ( 
.A(n_125),
.Y(n_225)
);

BUFx8_ASAP7_75t_SL g226 ( 
.A(n_93),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_135),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_133),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_41),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_136),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_35),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_46),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_145),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_48),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_57),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_90),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_124),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_75),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_11),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_61),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_131),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_33),
.Y(n_242)
);

INVx2_ASAP7_75t_SL g243 ( 
.A(n_86),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_30),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_106),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_38),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_17),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_0),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_6),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_141),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_22),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_138),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_88),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_8),
.Y(n_254)
);

BUFx10_ASAP7_75t_L g255 ( 
.A(n_85),
.Y(n_255)
);

BUFx10_ASAP7_75t_L g256 ( 
.A(n_23),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_96),
.Y(n_257)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_69),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_18),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_20),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_29),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_49),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_66),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_6),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_56),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_152),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_127),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_74),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_39),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_25),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_55),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_144),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_43),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_153),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_28),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_70),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_23),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g278 ( 
.A(n_82),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_16),
.Y(n_279)
);

BUFx8_ASAP7_75t_SL g280 ( 
.A(n_99),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_63),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_10),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_46),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_2),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_42),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_41),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_101),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_129),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_122),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_35),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_13),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_3),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_50),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_45),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_146),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_13),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_9),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_39),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_103),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_40),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_9),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_8),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_27),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_155),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_38),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_94),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_48),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_3),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_4),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_47),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_139),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_117),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_30),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_53),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_27),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_56),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_154),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_47),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_176),
.Y(n_319)
);

INVxp67_ASAP7_75t_SL g320 ( 
.A(n_258),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_176),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_176),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_176),
.Y(n_323)
);

NOR2xp67_ASAP7_75t_L g324 ( 
.A(n_208),
.B(n_2),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_226),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_176),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_180),
.Y(n_327)
);

NOR2xp67_ASAP7_75t_L g328 ( 
.A(n_208),
.B(n_4),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_309),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_158),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_280),
.Y(n_331)
);

INVxp67_ASAP7_75t_SL g332 ( 
.A(n_208),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_178),
.B(n_5),
.Y(n_333)
);

INVxp33_ASAP7_75t_SL g334 ( 
.A(n_297),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_180),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_161),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_157),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_173),
.Y(n_338)
);

INVxp67_ASAP7_75t_SL g339 ( 
.A(n_185),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_194),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_243),
.B(n_5),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_159),
.Y(n_342)
);

INVxp33_ASAP7_75t_SL g343 ( 
.A(n_182),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_212),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_214),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_180),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_180),
.Y(n_347)
);

BUFx3_ASAP7_75t_L g348 ( 
.A(n_185),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_160),
.Y(n_349)
);

BUFx3_ASAP7_75t_L g350 ( 
.A(n_191),
.Y(n_350)
);

CKINVDCx14_ASAP7_75t_R g351 ( 
.A(n_164),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_166),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_180),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_171),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_172),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_236),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_234),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_234),
.Y(n_358)
);

BUFx3_ASAP7_75t_L g359 ( 
.A(n_191),
.Y(n_359)
);

CKINVDCx16_ASAP7_75t_R g360 ( 
.A(n_309),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_234),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_234),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_177),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_234),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_183),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_186),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_187),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_243),
.B(n_10),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_287),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_165),
.Y(n_370)
);

BUFx2_ASAP7_75t_L g371 ( 
.A(n_190),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_165),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_188),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_189),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_169),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_167),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_167),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_162),
.B(n_174),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_268),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_219),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_219),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_318),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_197),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_318),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_190),
.B(n_161),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_205),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_168),
.Y(n_387)
);

NOR2xp67_ASAP7_75t_L g388 ( 
.A(n_259),
.B(n_11),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_198),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_200),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_268),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_201),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_168),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_210),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_210),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_229),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_202),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_203),
.Y(n_398)
);

HB1xp67_ASAP7_75t_L g399 ( 
.A(n_206),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_229),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_232),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_232),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_204),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_207),
.Y(n_404)
);

INVxp33_ASAP7_75t_SL g405 ( 
.A(n_211),
.Y(n_405)
);

HB1xp67_ASAP7_75t_L g406 ( 
.A(n_216),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_319),
.Y(n_407)
);

BUFx2_ASAP7_75t_L g408 ( 
.A(n_379),
.Y(n_408)
);

BUFx2_ASAP7_75t_L g409 ( 
.A(n_391),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_337),
.Y(n_410)
);

INVx3_ASAP7_75t_L g411 ( 
.A(n_375),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_375),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_375),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_342),
.Y(n_414)
);

AND2x4_ASAP7_75t_L g415 ( 
.A(n_324),
.B(n_195),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_330),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_349),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_319),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_321),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_352),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_322),
.Y(n_421)
);

NAND2xp33_ASAP7_75t_L g422 ( 
.A(n_341),
.B(n_217),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_322),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_338),
.Y(n_424)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_323),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_323),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_326),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_332),
.B(n_195),
.Y(n_428)
);

INVx3_ASAP7_75t_L g429 ( 
.A(n_326),
.Y(n_429)
);

OR2x2_ASAP7_75t_L g430 ( 
.A(n_371),
.B(n_269),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_327),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_378),
.B(n_209),
.Y(n_432)
);

OR2x2_ASAP7_75t_L g433 ( 
.A(n_371),
.B(n_249),
.Y(n_433)
);

BUFx2_ASAP7_75t_L g434 ( 
.A(n_329),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_354),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_385),
.B(n_225),
.Y(n_436)
);

AND2x4_ASAP7_75t_L g437 ( 
.A(n_324),
.B(n_328),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_385),
.B(n_225),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_355),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_360),
.B(n_199),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_335),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_363),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_335),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_346),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_346),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_365),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_340),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_347),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_347),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_366),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_R g451 ( 
.A(n_351),
.B(n_213),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_344),
.Y(n_452)
);

BUFx2_ASAP7_75t_L g453 ( 
.A(n_386),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_339),
.B(n_215),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_L g455 ( 
.A1(n_360),
.A2(n_181),
.B1(n_170),
.B2(n_242),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_353),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_367),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_353),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_373),
.Y(n_459)
);

XNOR2x1_ASAP7_75t_L g460 ( 
.A(n_388),
.B(n_231),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_357),
.Y(n_461)
);

OAI21x1_ASAP7_75t_L g462 ( 
.A1(n_368),
.A2(n_221),
.B(n_192),
.Y(n_462)
);

INVx3_ASAP7_75t_L g463 ( 
.A(n_357),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_358),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_358),
.B(n_361),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_361),
.B(n_218),
.Y(n_466)
);

AND2x4_ASAP7_75t_L g467 ( 
.A(n_328),
.B(n_267),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_362),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_362),
.Y(n_469)
);

HB1xp67_ASAP7_75t_L g470 ( 
.A(n_399),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_374),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_383),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_389),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_364),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_393),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_334),
.A2(n_292),
.B1(n_271),
.B2(n_273),
.Y(n_476)
);

AND2x2_ASAP7_75t_SL g477 ( 
.A(n_333),
.B(n_192),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_394),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_345),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_477),
.B(n_390),
.Y(n_480)
);

NOR2x1p5_ASAP7_75t_L g481 ( 
.A(n_410),
.B(n_325),
.Y(n_481)
);

OR2x2_ASAP7_75t_L g482 ( 
.A(n_430),
.B(n_406),
.Y(n_482)
);

AOI22xp33_ASAP7_75t_L g483 ( 
.A1(n_477),
.A2(n_320),
.B1(n_271),
.B2(n_273),
.Y(n_483)
);

AND2x4_ASAP7_75t_L g484 ( 
.A(n_437),
.B(n_267),
.Y(n_484)
);

BUFx2_ASAP7_75t_L g485 ( 
.A(n_434),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_L g486 ( 
.A1(n_477),
.A2(n_397),
.B1(n_398),
.B2(n_388),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_407),
.Y(n_487)
);

AND2x6_ASAP7_75t_L g488 ( 
.A(n_437),
.B(n_221),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_418),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_436),
.B(n_348),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_437),
.B(n_392),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_432),
.B(n_343),
.Y(n_492)
);

NOR2x1p5_ASAP7_75t_L g493 ( 
.A(n_414),
.B(n_331),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_417),
.B(n_403),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_475),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_420),
.B(n_404),
.Y(n_496)
);

INVx3_ASAP7_75t_L g497 ( 
.A(n_412),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_407),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_421),
.Y(n_499)
);

INVx1_ASAP7_75t_SL g500 ( 
.A(n_416),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_421),
.Y(n_501)
);

INVx4_ASAP7_75t_L g502 ( 
.A(n_419),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_423),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_432),
.B(n_405),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_460),
.A2(n_356),
.B1(n_369),
.B2(n_274),
.Y(n_505)
);

AOI22xp33_ASAP7_75t_L g506 ( 
.A1(n_437),
.A2(n_294),
.B1(n_296),
.B2(n_293),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_423),
.Y(n_507)
);

INVx5_ASAP7_75t_L g508 ( 
.A(n_412),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_475),
.Y(n_509)
);

INVx2_ASAP7_75t_SL g510 ( 
.A(n_436),
.Y(n_510)
);

BUFx10_ASAP7_75t_L g511 ( 
.A(n_435),
.Y(n_511)
);

INVx1_ASAP7_75t_SL g512 ( 
.A(n_424),
.Y(n_512)
);

INVx2_ASAP7_75t_SL g513 ( 
.A(n_438),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_439),
.B(n_199),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_418),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_426),
.Y(n_516)
);

OAI221xp5_ASAP7_75t_L g517 ( 
.A1(n_478),
.A2(n_336),
.B1(n_387),
.B2(n_395),
.C(n_303),
.Y(n_517)
);

INVx3_ASAP7_75t_L g518 ( 
.A(n_412),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_438),
.B(n_348),
.Y(n_519)
);

OR2x6_ASAP7_75t_L g520 ( 
.A(n_433),
.B(n_440),
.Y(n_520)
);

OR2x2_ASAP7_75t_L g521 ( 
.A(n_430),
.B(n_350),
.Y(n_521)
);

NAND2xp33_ASAP7_75t_L g522 ( 
.A(n_466),
.B(n_169),
.Y(n_522)
);

AOI22xp33_ASAP7_75t_L g523 ( 
.A1(n_428),
.A2(n_293),
.B1(n_294),
.B2(n_296),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_L g524 ( 
.A1(n_460),
.A2(n_453),
.B1(n_470),
.B2(n_422),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_454),
.B(n_350),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_438),
.B(n_428),
.Y(n_526)
);

INVx5_ASAP7_75t_L g527 ( 
.A(n_412),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_454),
.B(n_350),
.Y(n_528)
);

AOI22xp33_ASAP7_75t_L g529 ( 
.A1(n_428),
.A2(n_282),
.B1(n_277),
.B2(n_283),
.Y(n_529)
);

INVxp67_ASAP7_75t_SL g530 ( 
.A(n_466),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_443),
.Y(n_531)
);

INVx6_ASAP7_75t_L g532 ( 
.A(n_415),
.Y(n_532)
);

AOI22xp33_ASAP7_75t_L g533 ( 
.A1(n_415),
.A2(n_467),
.B1(n_460),
.B2(n_462),
.Y(n_533)
);

INVxp67_ASAP7_75t_SL g534 ( 
.A(n_412),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_415),
.B(n_359),
.Y(n_535)
);

OR2x2_ASAP7_75t_L g536 ( 
.A(n_434),
.B(n_359),
.Y(n_536)
);

INVx3_ASAP7_75t_L g537 ( 
.A(n_419),
.Y(n_537)
);

INVxp67_ASAP7_75t_SL g538 ( 
.A(n_465),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_426),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_442),
.B(n_199),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_446),
.B(n_450),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_L g542 ( 
.A1(n_433),
.A2(n_270),
.B1(n_261),
.B2(n_260),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_457),
.B(n_255),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_443),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_415),
.B(n_359),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_427),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_467),
.B(n_370),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_443),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_459),
.B(n_278),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_471),
.B(n_472),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_473),
.B(n_196),
.Y(n_551)
);

INVxp33_ASAP7_75t_SL g552 ( 
.A(n_455),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_448),
.Y(n_553)
);

AOI22xp33_ASAP7_75t_L g554 ( 
.A1(n_467),
.A2(n_284),
.B1(n_314),
.B2(n_277),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_431),
.B(n_227),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_431),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_470),
.B(n_453),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_SL g558 ( 
.A(n_455),
.B(n_163),
.Y(n_558)
);

NOR2x1p5_ASAP7_75t_L g559 ( 
.A(n_433),
.B(n_235),
.Y(n_559)
);

AOI22xp33_ASAP7_75t_L g560 ( 
.A1(n_462),
.A2(n_284),
.B1(n_283),
.B2(n_303),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_451),
.B(n_255),
.Y(n_561)
);

AND2x4_ASAP7_75t_L g562 ( 
.A(n_462),
.B(n_162),
.Y(n_562)
);

NAND2xp33_ASAP7_75t_SL g563 ( 
.A(n_476),
.B(n_239),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_444),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_419),
.Y(n_565)
);

NAND2xp33_ASAP7_75t_SL g566 ( 
.A(n_476),
.B(n_244),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_444),
.B(n_246),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g568 ( 
.A(n_419),
.Y(n_568)
);

OAI22xp33_ASAP7_75t_L g569 ( 
.A1(n_465),
.A2(n_251),
.B1(n_254),
.B2(n_316),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_445),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_448),
.Y(n_571)
);

AND2x6_ASAP7_75t_L g572 ( 
.A(n_445),
.B(n_230),
.Y(n_572)
);

HB1xp67_ASAP7_75t_L g573 ( 
.A(n_408),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_449),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_458),
.B(n_228),
.Y(n_575)
);

OAI22xp5_ASAP7_75t_L g576 ( 
.A1(n_458),
.A2(n_302),
.B1(n_301),
.B2(n_300),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_468),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_468),
.B(n_370),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_469),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_469),
.B(n_247),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_449),
.B(n_372),
.Y(n_581)
);

BUFx3_ASAP7_75t_L g582 ( 
.A(n_441),
.Y(n_582)
);

INVx3_ASAP7_75t_L g583 ( 
.A(n_441),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_449),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_456),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_425),
.Y(n_586)
);

BUFx3_ASAP7_75t_L g587 ( 
.A(n_441),
.Y(n_587)
);

INVx4_ASAP7_75t_L g588 ( 
.A(n_441),
.Y(n_588)
);

INVx1_ASAP7_75t_SL g589 ( 
.A(n_447),
.Y(n_589)
);

INVx1_ASAP7_75t_SL g590 ( 
.A(n_452),
.Y(n_590)
);

INVx2_ASAP7_75t_SL g591 ( 
.A(n_425),
.Y(n_591)
);

OR2x2_ASAP7_75t_L g592 ( 
.A(n_409),
.B(n_396),
.Y(n_592)
);

AOI22xp33_ASAP7_75t_L g593 ( 
.A1(n_429),
.A2(n_308),
.B1(n_310),
.B2(n_230),
.Y(n_593)
);

BUFx10_ASAP7_75t_L g594 ( 
.A(n_461),
.Y(n_594)
);

AOI22xp33_ASAP7_75t_L g595 ( 
.A1(n_429),
.A2(n_308),
.B1(n_310),
.B2(n_304),
.Y(n_595)
);

INVx2_ASAP7_75t_SL g596 ( 
.A(n_429),
.Y(n_596)
);

BUFx6f_ASAP7_75t_L g597 ( 
.A(n_461),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_463),
.B(n_248),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_463),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_409),
.B(n_163),
.Y(n_600)
);

INVx2_ASAP7_75t_SL g601 ( 
.A(n_463),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_463),
.B(n_238),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_461),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_461),
.B(n_262),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_456),
.Y(n_605)
);

AOI22xp33_ASAP7_75t_L g606 ( 
.A1(n_456),
.A2(n_304),
.B1(n_317),
.B2(n_233),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_533),
.B(n_169),
.Y(n_607)
);

INVx2_ASAP7_75t_SL g608 ( 
.A(n_536),
.Y(n_608)
);

INVxp67_ASAP7_75t_L g609 ( 
.A(n_557),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_530),
.B(n_461),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_547),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_538),
.B(n_174),
.Y(n_612)
);

NOR2x1p5_ASAP7_75t_L g613 ( 
.A(n_592),
.B(n_264),
.Y(n_613)
);

BUFx2_ASAP7_75t_L g614 ( 
.A(n_485),
.Y(n_614)
);

AOI22xp33_ASAP7_75t_L g615 ( 
.A1(n_562),
.A2(n_241),
.B1(n_257),
.B2(n_306),
.Y(n_615)
);

INVxp67_ASAP7_75t_L g616 ( 
.A(n_485),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_492),
.B(n_179),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_504),
.B(n_179),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_525),
.B(n_184),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_526),
.B(n_240),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_526),
.B(n_549),
.Y(n_621)
);

INVxp67_ASAP7_75t_L g622 ( 
.A(n_536),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_510),
.B(n_245),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_581),
.Y(n_624)
);

BUFx3_ASAP7_75t_L g625 ( 
.A(n_490),
.Y(n_625)
);

AOI22xp5_ASAP7_75t_L g626 ( 
.A1(n_480),
.A2(n_223),
.B1(n_263),
.B2(n_250),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_581),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_528),
.B(n_184),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_521),
.B(n_265),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_521),
.B(n_275),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_491),
.B(n_279),
.Y(n_631)
);

AND2x6_ASAP7_75t_SL g632 ( 
.A(n_550),
.B(n_551),
.Y(n_632)
);

HB1xp67_ASAP7_75t_L g633 ( 
.A(n_592),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_487),
.Y(n_634)
);

A2O1A1Ixp33_ASAP7_75t_L g635 ( 
.A1(n_510),
.A2(n_237),
.B(n_241),
.C(n_233),
.Y(n_635)
);

INVx5_ASAP7_75t_L g636 ( 
.A(n_488),
.Y(n_636)
);

OR2x6_ASAP7_75t_L g637 ( 
.A(n_573),
.B(n_193),
.Y(n_637)
);

BUFx3_ASAP7_75t_L g638 ( 
.A(n_490),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_513),
.B(n_252),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_486),
.B(n_253),
.Y(n_640)
);

BUFx8_ASAP7_75t_L g641 ( 
.A(n_482),
.Y(n_641)
);

AOI21xp5_ASAP7_75t_L g642 ( 
.A1(n_535),
.A2(n_545),
.B(n_534),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_598),
.B(n_193),
.Y(n_643)
);

OAI22xp5_ASAP7_75t_L g644 ( 
.A1(n_483),
.A2(n_237),
.B1(n_224),
.B2(n_222),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_562),
.B(n_169),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_482),
.B(n_285),
.Y(n_646)
);

A2O1A1Ixp33_ASAP7_75t_L g647 ( 
.A1(n_562),
.A2(n_224),
.B(n_222),
.C(n_220),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_487),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_558),
.B(n_524),
.Y(n_649)
);

BUFx3_ASAP7_75t_L g650 ( 
.A(n_519),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_519),
.B(n_266),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_569),
.B(n_272),
.Y(n_652)
);

OAI22xp33_ASAP7_75t_L g653 ( 
.A1(n_520),
.A2(n_295),
.B1(n_220),
.B2(n_257),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_498),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_498),
.Y(n_655)
);

OAI21xp5_ASAP7_75t_L g656 ( 
.A1(n_560),
.A2(n_596),
.B(n_591),
.Y(n_656)
);

INVx2_ASAP7_75t_SL g657 ( 
.A(n_484),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_484),
.B(n_281),
.Y(n_658)
);

NOR2x1p5_ASAP7_75t_L g659 ( 
.A(n_495),
.B(n_286),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_509),
.B(n_276),
.Y(n_660)
);

BUFx3_ASAP7_75t_L g661 ( 
.A(n_532),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_567),
.B(n_288),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_578),
.Y(n_663)
);

INVxp33_ASAP7_75t_SL g664 ( 
.A(n_505),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_511),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_591),
.B(n_169),
.Y(n_666)
);

OAI22xp33_ASAP7_75t_L g667 ( 
.A1(n_520),
.A2(n_295),
.B1(n_311),
.B2(n_317),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_596),
.B(n_306),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_601),
.B(n_311),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_601),
.B(n_411),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_546),
.B(n_556),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_499),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_520),
.B(n_290),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_578),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_499),
.Y(n_675)
);

OR2x2_ASAP7_75t_L g676 ( 
.A(n_520),
.B(n_396),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_494),
.B(n_291),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_586),
.B(n_312),
.Y(n_678)
);

AOI22xp5_ASAP7_75t_L g679 ( 
.A1(n_559),
.A2(n_488),
.B1(n_604),
.B2(n_555),
.Y(n_679)
);

AND2x6_ASAP7_75t_L g680 ( 
.A(n_586),
.B(n_312),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_501),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_501),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_503),
.B(n_411),
.Y(n_683)
);

AOI22xp5_ASAP7_75t_L g684 ( 
.A1(n_488),
.A2(n_289),
.B1(n_299),
.B2(n_163),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_503),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_511),
.B(n_256),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_507),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_516),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_539),
.Y(n_689)
);

NOR3xp33_ASAP7_75t_L g690 ( 
.A(n_600),
.B(n_313),
.C(n_298),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_539),
.B(n_474),
.Y(n_691)
);

AOI22xp5_ASAP7_75t_L g692 ( 
.A1(n_488),
.A2(n_312),
.B1(n_479),
.B2(n_315),
.Y(n_692)
);

INVx2_ASAP7_75t_SL g693 ( 
.A(n_575),
.Y(n_693)
);

AOI22xp33_ASAP7_75t_L g694 ( 
.A1(n_523),
.A2(n_312),
.B1(n_256),
.B2(n_402),
.Y(n_694)
);

OAI22xp5_ASAP7_75t_L g695 ( 
.A1(n_506),
.A2(n_312),
.B1(n_307),
.B2(n_305),
.Y(n_695)
);

AND2x6_ASAP7_75t_SL g696 ( 
.A(n_563),
.B(n_400),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_564),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_564),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_570),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_570),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_577),
.B(n_464),
.Y(n_701)
);

BUFx3_ASAP7_75t_L g702 ( 
.A(n_511),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_580),
.B(n_256),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_577),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_496),
.B(n_256),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_579),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_579),
.B(n_413),
.Y(n_707)
);

AOI22xp5_ASAP7_75t_L g708 ( 
.A1(n_488),
.A2(n_402),
.B1(n_401),
.B2(n_400),
.Y(n_708)
);

INVx2_ASAP7_75t_SL g709 ( 
.A(n_500),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_599),
.Y(n_710)
);

AOI22xp33_ASAP7_75t_SL g711 ( 
.A1(n_552),
.A2(n_175),
.B1(n_382),
.B2(n_381),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_602),
.B(n_384),
.Y(n_712)
);

AOI22xp5_ASAP7_75t_L g713 ( 
.A1(n_514),
.A2(n_384),
.B1(n_382),
.B2(n_381),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_529),
.B(n_380),
.Y(n_714)
);

NOR3xp33_ASAP7_75t_L g715 ( 
.A(n_563),
.B(n_566),
.C(n_540),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_554),
.B(n_377),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_489),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_543),
.B(n_12),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_542),
.B(n_377),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_561),
.B(n_12),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_552),
.B(n_376),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_537),
.B(n_372),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_515),
.Y(n_723)
);

AND2x6_ASAP7_75t_SL g724 ( 
.A(n_566),
.B(n_14),
.Y(n_724)
);

INVxp67_ASAP7_75t_L g725 ( 
.A(n_576),
.Y(n_725)
);

BUFx3_ASAP7_75t_L g726 ( 
.A(n_572),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_515),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_603),
.B(n_148),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_583),
.B(n_142),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_517),
.B(n_14),
.Y(n_730)
);

OR2x6_ASAP7_75t_L g731 ( 
.A(n_541),
.B(n_15),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_L g732 ( 
.A(n_582),
.B(n_16),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_497),
.B(n_121),
.Y(n_733)
);

AOI22xp5_ASAP7_75t_L g734 ( 
.A1(n_522),
.A2(n_111),
.B1(n_109),
.B2(n_108),
.Y(n_734)
);

AOI21xp5_ASAP7_75t_L g735 ( 
.A1(n_610),
.A2(n_588),
.B(n_502),
.Y(n_735)
);

OAI21xp5_ASAP7_75t_L g736 ( 
.A1(n_656),
.A2(n_522),
.B(n_605),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_609),
.B(n_590),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_636),
.B(n_497),
.Y(n_738)
);

BUFx2_ASAP7_75t_L g739 ( 
.A(n_614),
.Y(n_739)
);

BUFx6f_ASAP7_75t_L g740 ( 
.A(n_661),
.Y(n_740)
);

OAI22xp5_ASAP7_75t_L g741 ( 
.A1(n_725),
.A2(n_606),
.B1(n_593),
.B2(n_595),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_634),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_693),
.B(n_587),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_634),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_633),
.B(n_589),
.Y(n_745)
);

A2O1A1Ixp33_ASAP7_75t_L g746 ( 
.A1(n_730),
.A2(n_605),
.B(n_585),
.C(n_584),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_621),
.B(n_512),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_624),
.B(n_518),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_622),
.B(n_518),
.Y(n_749)
);

OAI22xp5_ASAP7_75t_L g750 ( 
.A1(n_615),
.A2(n_481),
.B1(n_493),
.B2(n_497),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_646),
.B(n_544),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_646),
.B(n_544),
.Y(n_752)
);

BUFx3_ASAP7_75t_L g753 ( 
.A(n_625),
.Y(n_753)
);

INVx3_ASAP7_75t_L g754 ( 
.A(n_661),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_679),
.B(n_518),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_648),
.Y(n_756)
);

O2A1O1Ixp33_ASAP7_75t_L g757 ( 
.A1(n_644),
.A2(n_531),
.B(n_548),
.C(n_553),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_627),
.B(n_574),
.Y(n_758)
);

BUFx8_ASAP7_75t_L g759 ( 
.A(n_709),
.Y(n_759)
);

OAI22xp5_ASAP7_75t_L g760 ( 
.A1(n_615),
.A2(n_574),
.B1(n_531),
.B2(n_585),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_654),
.Y(n_761)
);

OAI22xp5_ASAP7_75t_L g762 ( 
.A1(n_627),
.A2(n_571),
.B1(n_553),
.B2(n_584),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_654),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_608),
.B(n_629),
.Y(n_764)
);

BUFx4f_ASAP7_75t_L g765 ( 
.A(n_731),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_655),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_675),
.B(n_572),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_655),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_672),
.B(n_597),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_721),
.B(n_597),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_682),
.B(n_572),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_672),
.Y(n_772)
);

NOR2x1p5_ASAP7_75t_SL g773 ( 
.A(n_717),
.B(n_594),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_685),
.B(n_568),
.Y(n_774)
);

AOI21xp5_ASAP7_75t_L g775 ( 
.A1(n_657),
.A2(n_568),
.B(n_565),
.Y(n_775)
);

BUFx4f_ASAP7_75t_L g776 ( 
.A(n_731),
.Y(n_776)
);

NOR2xp67_ASAP7_75t_L g777 ( 
.A(n_665),
.B(n_84),
.Y(n_777)
);

INVx3_ASAP7_75t_L g778 ( 
.A(n_681),
.Y(n_778)
);

INVx2_ASAP7_75t_SL g779 ( 
.A(n_659),
.Y(n_779)
);

OAI22xp5_ASAP7_75t_L g780 ( 
.A1(n_612),
.A2(n_568),
.B1(n_565),
.B2(n_527),
.Y(n_780)
);

AOI22xp5_ASAP7_75t_L g781 ( 
.A1(n_649),
.A2(n_568),
.B1(n_565),
.B2(n_594),
.Y(n_781)
);

BUFx6f_ASAP7_75t_L g782 ( 
.A(n_726),
.Y(n_782)
);

AND2x2_ASAP7_75t_L g783 ( 
.A(n_630),
.B(n_18),
.Y(n_783)
);

BUFx6f_ASAP7_75t_L g784 ( 
.A(n_726),
.Y(n_784)
);

OAI21xp5_ASAP7_75t_L g785 ( 
.A1(n_611),
.A2(n_527),
.B(n_508),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_687),
.B(n_527),
.Y(n_786)
);

OAI21xp5_ASAP7_75t_L g787 ( 
.A1(n_688),
.A2(n_80),
.B(n_76),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_688),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_689),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_698),
.B(n_21),
.Y(n_790)
);

AOI21xp5_ASAP7_75t_L g791 ( 
.A1(n_671),
.A2(n_712),
.B(n_670),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_689),
.B(n_72),
.Y(n_792)
);

BUFx2_ASAP7_75t_L g793 ( 
.A(n_616),
.Y(n_793)
);

AO21x1_ASAP7_75t_L g794 ( 
.A1(n_653),
.A2(n_21),
.B(n_24),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_697),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_699),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_L g797 ( 
.A1(n_691),
.A2(n_62),
.B(n_26),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_699),
.Y(n_798)
);

HB1xp67_ASAP7_75t_L g799 ( 
.A(n_625),
.Y(n_799)
);

AOI22xp5_ASAP7_75t_L g800 ( 
.A1(n_631),
.A2(n_24),
.B1(n_26),
.B2(n_28),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_700),
.Y(n_801)
);

NOR2x1_ASAP7_75t_L g802 ( 
.A(n_702),
.B(n_638),
.Y(n_802)
);

AOI21xp5_ASAP7_75t_L g803 ( 
.A1(n_701),
.A2(n_29),
.B(n_32),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_707),
.A2(n_32),
.B(n_34),
.Y(n_804)
);

AND2x6_ASAP7_75t_SL g805 ( 
.A(n_731),
.B(n_34),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_L g806 ( 
.A(n_638),
.B(n_650),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_700),
.B(n_37),
.Y(n_807)
);

OAI21xp33_ASAP7_75t_L g808 ( 
.A1(n_705),
.A2(n_37),
.B(n_40),
.Y(n_808)
);

OAI21xp5_ASAP7_75t_L g809 ( 
.A1(n_704),
.A2(n_42),
.B(n_43),
.Y(n_809)
);

OAI21xp5_ASAP7_75t_L g810 ( 
.A1(n_704),
.A2(n_44),
.B(n_45),
.Y(n_810)
);

OAI22xp5_ASAP7_75t_L g811 ( 
.A1(n_650),
.A2(n_54),
.B1(n_50),
.B2(n_51),
.Y(n_811)
);

AND2x2_ASAP7_75t_SL g812 ( 
.A(n_715),
.B(n_49),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_706),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_683),
.A2(n_51),
.B(n_53),
.Y(n_814)
);

INVx3_ASAP7_75t_L g815 ( 
.A(n_706),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_631),
.B(n_54),
.Y(n_816)
);

AND2x2_ASAP7_75t_L g817 ( 
.A(n_630),
.B(n_686),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_663),
.B(n_674),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_619),
.B(n_628),
.Y(n_819)
);

OR2x2_ASAP7_75t_L g820 ( 
.A(n_676),
.B(n_620),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_719),
.B(n_710),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_651),
.A2(n_658),
.B(n_623),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_692),
.B(n_708),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_639),
.A2(n_729),
.B(n_733),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_717),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_722),
.Y(n_826)
);

AND2x4_ASAP7_75t_L g827 ( 
.A(n_702),
.B(n_613),
.Y(n_827)
);

OR2x2_ASAP7_75t_L g828 ( 
.A(n_637),
.B(n_673),
.Y(n_828)
);

AOI22xp5_ASAP7_75t_L g829 ( 
.A1(n_705),
.A2(n_677),
.B1(n_673),
.B2(n_640),
.Y(n_829)
);

AOI21x1_ASAP7_75t_L g830 ( 
.A1(n_668),
.A2(n_669),
.B(n_666),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_718),
.B(n_667),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_677),
.B(n_637),
.Y(n_832)
);

OAI21xp33_ASAP7_75t_L g833 ( 
.A1(n_718),
.A2(n_730),
.B(n_720),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_711),
.B(n_720),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_727),
.Y(n_835)
);

OAI22xp5_ASAP7_75t_L g836 ( 
.A1(n_626),
.A2(n_684),
.B1(n_664),
.B2(n_662),
.Y(n_836)
);

O2A1O1Ixp5_ASAP7_75t_SL g837 ( 
.A1(n_703),
.A2(n_652),
.B(n_678),
.C(n_728),
.Y(n_837)
);

AOI33xp33_ASAP7_75t_L g838 ( 
.A1(n_694),
.A2(n_713),
.A3(n_724),
.B1(n_734),
.B2(n_723),
.B3(n_696),
.Y(n_838)
);

AND2x2_ASAP7_75t_L g839 ( 
.A(n_637),
.B(n_690),
.Y(n_839)
);

INVxp67_ASAP7_75t_L g840 ( 
.A(n_732),
.Y(n_840)
);

NOR2x1_ASAP7_75t_L g841 ( 
.A(n_728),
.B(n_732),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_660),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_678),
.Y(n_843)
);

O2A1O1Ixp33_ASAP7_75t_L g844 ( 
.A1(n_647),
.A2(n_635),
.B(n_714),
.C(n_716),
.Y(n_844)
);

AOI21xp5_ASAP7_75t_L g845 ( 
.A1(n_694),
.A2(n_695),
.B(n_680),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_632),
.B(n_680),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_680),
.A2(n_610),
.B(n_642),
.Y(n_847)
);

BUFx8_ASAP7_75t_SL g848 ( 
.A(n_641),
.Y(n_848)
);

O2A1O1Ixp33_ASAP7_75t_L g849 ( 
.A1(n_680),
.A2(n_641),
.B(n_607),
.C(n_644),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_680),
.A2(n_610),
.B(n_642),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_610),
.A2(n_642),
.B(n_656),
.Y(n_851)
);

O2A1O1Ixp33_ASAP7_75t_SL g852 ( 
.A1(n_607),
.A2(n_647),
.B(n_645),
.C(n_618),
.Y(n_852)
);

AND2x4_ASAP7_75t_L g853 ( 
.A(n_625),
.B(n_638),
.Y(n_853)
);

NOR2x1_ASAP7_75t_L g854 ( 
.A(n_702),
.B(n_481),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_609),
.B(n_621),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_617),
.B(n_530),
.Y(n_856)
);

INVx3_ASAP7_75t_L g857 ( 
.A(n_661),
.Y(n_857)
);

AOI22xp5_ASAP7_75t_L g858 ( 
.A1(n_621),
.A2(n_504),
.B1(n_492),
.B2(n_530),
.Y(n_858)
);

OAI22xp5_ASAP7_75t_L g859 ( 
.A1(n_725),
.A2(n_617),
.B1(n_618),
.B2(n_615),
.Y(n_859)
);

OAI21xp33_ASAP7_75t_L g860 ( 
.A1(n_617),
.A2(n_618),
.B(n_558),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_636),
.B(n_679),
.Y(n_861)
);

INVx3_ASAP7_75t_L g862 ( 
.A(n_661),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_610),
.A2(n_642),
.B(n_656),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_634),
.Y(n_864)
);

AOI21xp5_ASAP7_75t_L g865 ( 
.A1(n_610),
.A2(n_642),
.B(n_656),
.Y(n_865)
);

A2O1A1Ixp33_ASAP7_75t_L g866 ( 
.A1(n_730),
.A2(n_718),
.B(n_720),
.C(n_617),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_609),
.B(n_621),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_617),
.B(n_530),
.Y(n_868)
);

AO21x1_ASAP7_75t_L g869 ( 
.A1(n_607),
.A2(n_643),
.B(n_618),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_617),
.B(n_530),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_617),
.B(n_530),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_617),
.B(n_530),
.Y(n_872)
);

BUFx6f_ASAP7_75t_L g873 ( 
.A(n_661),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_617),
.B(n_530),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_609),
.B(n_621),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_610),
.A2(n_642),
.B(n_656),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_617),
.B(n_530),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_634),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_617),
.B(n_530),
.Y(n_879)
);

NAND3xp33_ASAP7_75t_L g880 ( 
.A(n_609),
.B(n_558),
.C(n_504),
.Y(n_880)
);

BUFx2_ASAP7_75t_SL g881 ( 
.A(n_739),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_866),
.B(n_751),
.Y(n_882)
);

INVx3_ASAP7_75t_L g883 ( 
.A(n_782),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_866),
.B(n_752),
.Y(n_884)
);

AOI22xp33_ASAP7_75t_SL g885 ( 
.A1(n_765),
.A2(n_776),
.B1(n_812),
.B2(n_832),
.Y(n_885)
);

BUFx6f_ASAP7_75t_L g886 ( 
.A(n_740),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_819),
.B(n_842),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_817),
.B(n_764),
.Y(n_888)
);

OAI21x1_ASAP7_75t_L g889 ( 
.A1(n_847),
.A2(n_850),
.B(n_735),
.Y(n_889)
);

AOI21x1_ASAP7_75t_L g890 ( 
.A1(n_755),
.A2(n_861),
.B(n_769),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_851),
.A2(n_865),
.B(n_863),
.Y(n_891)
);

OR2x2_ASAP7_75t_L g892 ( 
.A(n_745),
.B(n_793),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_SL g893 ( 
.A1(n_787),
.A2(n_823),
.B(n_736),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_768),
.Y(n_894)
);

OAI22x1_ASAP7_75t_L g895 ( 
.A1(n_834),
.A2(n_831),
.B1(n_875),
.B2(n_867),
.Y(n_895)
);

AO31x2_ASAP7_75t_L g896 ( 
.A1(n_869),
.A2(n_746),
.A3(n_876),
.B(n_859),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_833),
.B(n_855),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_853),
.B(n_855),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_852),
.A2(n_868),
.B(n_856),
.Y(n_899)
);

BUFx6f_ASAP7_75t_L g900 ( 
.A(n_740),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_737),
.B(n_853),
.Y(n_901)
);

AOI22xp5_ASAP7_75t_L g902 ( 
.A1(n_836),
.A2(n_747),
.B1(n_875),
.B2(n_867),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_791),
.A2(n_824),
.B(n_870),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_871),
.B(n_872),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_778),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_874),
.B(n_877),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_742),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_879),
.B(n_840),
.Y(n_908)
);

OA22x2_ASAP7_75t_L g909 ( 
.A1(n_808),
.A2(n_831),
.B1(n_800),
.B2(n_860),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_840),
.B(n_826),
.Y(n_910)
);

OAI21x1_ASAP7_75t_L g911 ( 
.A1(n_769),
.A2(n_830),
.B(n_762),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_806),
.B(n_821),
.Y(n_912)
);

INVx1_ASAP7_75t_SL g913 ( 
.A(n_820),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_737),
.B(n_747),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_778),
.Y(n_915)
);

NOR2xp33_ASAP7_75t_L g916 ( 
.A(n_799),
.B(n_806),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_815),
.Y(n_917)
);

AOI21xp33_ASAP7_75t_L g918 ( 
.A1(n_783),
.A2(n_810),
.B(n_849),
.Y(n_918)
);

INVx3_ASAP7_75t_L g919 ( 
.A(n_782),
.Y(n_919)
);

BUFx3_ASAP7_75t_L g920 ( 
.A(n_759),
.Y(n_920)
);

CKINVDCx20_ASAP7_75t_R g921 ( 
.A(n_848),
.Y(n_921)
);

OAI22x1_ASAP7_75t_L g922 ( 
.A1(n_828),
.A2(n_839),
.B1(n_799),
.B2(n_827),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_753),
.B(n_818),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_SL g924 ( 
.A(n_753),
.B(n_765),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_744),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_776),
.B(n_838),
.Y(n_926)
);

NOR2x1_ASAP7_75t_L g927 ( 
.A(n_854),
.B(n_802),
.Y(n_927)
);

BUFx6f_ASAP7_75t_L g928 ( 
.A(n_740),
.Y(n_928)
);

AO31x2_ASAP7_75t_L g929 ( 
.A1(n_746),
.A2(n_760),
.A3(n_807),
.B(n_794),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_815),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_L g931 ( 
.A(n_743),
.B(n_846),
.Y(n_931)
);

AND2x4_ASAP7_75t_L g932 ( 
.A(n_779),
.B(n_827),
.Y(n_932)
);

INVx1_ASAP7_75t_SL g933 ( 
.A(n_790),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_766),
.Y(n_934)
);

BUFx6f_ASAP7_75t_L g935 ( 
.A(n_740),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_878),
.B(n_788),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_761),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_758),
.A2(n_767),
.B(n_771),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_785),
.A2(n_841),
.B(n_748),
.Y(n_939)
);

AND2x4_ASAP7_75t_L g940 ( 
.A(n_873),
.B(n_862),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_738),
.A2(n_822),
.B(n_774),
.Y(n_941)
);

BUFx2_ASAP7_75t_L g942 ( 
.A(n_759),
.Y(n_942)
);

OAI21xp5_ASAP7_75t_L g943 ( 
.A1(n_837),
.A2(n_845),
.B(n_757),
.Y(n_943)
);

INVx5_ASAP7_75t_L g944 ( 
.A(n_782),
.Y(n_944)
);

INVx1_ASAP7_75t_SL g945 ( 
.A(n_812),
.Y(n_945)
);

OAI21x1_ASAP7_75t_L g946 ( 
.A1(n_775),
.A2(n_757),
.B(n_786),
.Y(n_946)
);

OAI22xp5_ASAP7_75t_L g947 ( 
.A1(n_741),
.A2(n_784),
.B1(n_782),
.B2(n_801),
.Y(n_947)
);

OAI21x1_ASAP7_75t_L g948 ( 
.A1(n_772),
.A2(n_798),
.B(n_864),
.Y(n_948)
);

NOR2x1_ASAP7_75t_SL g949 ( 
.A(n_784),
.B(n_738),
.Y(n_949)
);

AOI21x1_ASAP7_75t_L g950 ( 
.A1(n_763),
.A2(n_789),
.B(n_813),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_795),
.B(n_796),
.Y(n_951)
);

BUFx2_ASAP7_75t_L g952 ( 
.A(n_805),
.Y(n_952)
);

NAND2x1_ASAP7_75t_L g953 ( 
.A(n_784),
.B(n_862),
.Y(n_953)
);

HB1xp67_ASAP7_75t_L g954 ( 
.A(n_749),
.Y(n_954)
);

A2O1A1Ixp33_ASAP7_75t_L g955 ( 
.A1(n_844),
.A2(n_838),
.B(n_770),
.C(n_750),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_873),
.B(n_777),
.Y(n_956)
);

A2O1A1Ixp33_ASAP7_75t_L g957 ( 
.A1(n_770),
.A2(n_749),
.B(n_843),
.C(n_803),
.Y(n_957)
);

BUFx6f_ASAP7_75t_L g958 ( 
.A(n_873),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_825),
.B(n_835),
.Y(n_959)
);

NAND2x1p5_ASAP7_75t_L g960 ( 
.A(n_754),
.B(n_857),
.Y(n_960)
);

OAI21xp5_ASAP7_75t_L g961 ( 
.A1(n_792),
.A2(n_781),
.B(n_780),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_754),
.B(n_857),
.Y(n_962)
);

AND2x4_ASAP7_75t_L g963 ( 
.A(n_773),
.B(n_814),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_804),
.B(n_811),
.Y(n_964)
);

O2A1O1Ixp5_ASAP7_75t_L g965 ( 
.A1(n_797),
.A2(n_617),
.B(n_618),
.C(n_866),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_848),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_851),
.A2(n_636),
.B(n_863),
.Y(n_967)
);

AOI21xp33_ASAP7_75t_L g968 ( 
.A1(n_833),
.A2(n_816),
.B(n_829),
.Y(n_968)
);

CKINVDCx20_ASAP7_75t_R g969 ( 
.A(n_848),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_866),
.B(n_751),
.Y(n_970)
);

AOI21xp33_ASAP7_75t_L g971 ( 
.A1(n_833),
.A2(n_816),
.B(n_829),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_866),
.B(n_751),
.Y(n_972)
);

BUFx2_ASAP7_75t_L g973 ( 
.A(n_739),
.Y(n_973)
);

A2O1A1Ixp33_ASAP7_75t_L g974 ( 
.A1(n_833),
.A2(n_866),
.B(n_829),
.C(n_858),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_756),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_851),
.A2(n_636),
.B(n_863),
.Y(n_976)
);

HB1xp67_ASAP7_75t_L g977 ( 
.A(n_739),
.Y(n_977)
);

INVx3_ASAP7_75t_L g978 ( 
.A(n_782),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_L g979 ( 
.A(n_737),
.B(n_609),
.Y(n_979)
);

AOI21xp33_ASAP7_75t_L g980 ( 
.A1(n_833),
.A2(n_816),
.B(n_829),
.Y(n_980)
);

CKINVDCx11_ASAP7_75t_R g981 ( 
.A(n_805),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_866),
.B(n_751),
.Y(n_982)
);

OR2x6_ASAP7_75t_L g983 ( 
.A(n_739),
.B(n_709),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_851),
.A2(n_636),
.B(n_863),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_756),
.Y(n_985)
);

INVx3_ASAP7_75t_L g986 ( 
.A(n_782),
.Y(n_986)
);

AND2x6_ASAP7_75t_L g987 ( 
.A(n_782),
.B(n_784),
.Y(n_987)
);

INVx8_ASAP7_75t_L g988 ( 
.A(n_740),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_756),
.Y(n_989)
);

AOI22xp5_ASAP7_75t_L g990 ( 
.A1(n_829),
.A2(n_492),
.B1(n_504),
.B2(n_817),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_817),
.B(n_609),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_866),
.B(n_751),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_866),
.B(n_751),
.Y(n_993)
);

A2O1A1Ixp33_ASAP7_75t_L g994 ( 
.A1(n_833),
.A2(n_866),
.B(n_829),
.C(n_858),
.Y(n_994)
);

AOI211x1_ASAP7_75t_L g995 ( 
.A1(n_833),
.A2(n_834),
.B(n_809),
.C(n_810),
.Y(n_995)
);

AND2x4_ASAP7_75t_L g996 ( 
.A(n_853),
.B(n_753),
.Y(n_996)
);

NOR2xp67_ASAP7_75t_L g997 ( 
.A(n_880),
.B(n_665),
.Y(n_997)
);

AND2x2_ASAP7_75t_L g998 ( 
.A(n_817),
.B(n_609),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_817),
.B(n_609),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_851),
.A2(n_865),
.B(n_863),
.Y(n_1000)
);

A2O1A1Ixp33_ASAP7_75t_L g1001 ( 
.A1(n_833),
.A2(n_866),
.B(n_829),
.C(n_858),
.Y(n_1001)
);

O2A1O1Ixp5_ASAP7_75t_L g1002 ( 
.A1(n_866),
.A2(n_617),
.B(n_618),
.C(n_831),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_756),
.Y(n_1003)
);

AND2x6_ASAP7_75t_L g1004 ( 
.A(n_782),
.B(n_784),
.Y(n_1004)
);

OAI22xp5_ASAP7_75t_L g1005 ( 
.A1(n_990),
.A2(n_902),
.B1(n_887),
.B2(n_994),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_887),
.B(n_908),
.Y(n_1006)
);

BUFx6f_ASAP7_75t_L g1007 ( 
.A(n_886),
.Y(n_1007)
);

CKINVDCx6p67_ASAP7_75t_R g1008 ( 
.A(n_920),
.Y(n_1008)
);

XNOR2xp5_ASAP7_75t_L g1009 ( 
.A(n_921),
.B(n_969),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_893),
.A2(n_903),
.B(n_899),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_907),
.Y(n_1011)
);

NOR2xp33_ASAP7_75t_SL g1012 ( 
.A(n_974),
.B(n_1001),
.Y(n_1012)
);

AOI22xp33_ASAP7_75t_L g1013 ( 
.A1(n_909),
.A2(n_968),
.B1(n_971),
.B2(n_980),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_894),
.Y(n_1014)
);

BUFx3_ASAP7_75t_L g1015 ( 
.A(n_973),
.Y(n_1015)
);

AND2x4_ASAP7_75t_L g1016 ( 
.A(n_996),
.B(n_932),
.Y(n_1016)
);

INVx3_ASAP7_75t_L g1017 ( 
.A(n_987),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_881),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_983),
.Y(n_1019)
);

OAI21xp33_ASAP7_75t_L g1020 ( 
.A1(n_979),
.A2(n_914),
.B(n_897),
.Y(n_1020)
);

CKINVDCx20_ASAP7_75t_R g1021 ( 
.A(n_977),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_901),
.B(n_991),
.Y(n_1022)
);

CKINVDCx6p67_ASAP7_75t_R g1023 ( 
.A(n_983),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_908),
.B(n_912),
.Y(n_1024)
);

AO21x1_ASAP7_75t_L g1025 ( 
.A1(n_968),
.A2(n_980),
.B(n_971),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_1000),
.A2(n_891),
.B(n_967),
.Y(n_1026)
);

AND2x2_ASAP7_75t_L g1027 ( 
.A(n_998),
.B(n_999),
.Y(n_1027)
);

NAND2xp33_ASAP7_75t_L g1028 ( 
.A(n_987),
.B(n_1004),
.Y(n_1028)
);

AND2x4_ASAP7_75t_L g1029 ( 
.A(n_996),
.B(n_932),
.Y(n_1029)
);

NOR2xp67_ASAP7_75t_L g1030 ( 
.A(n_944),
.B(n_895),
.Y(n_1030)
);

BUFx8_ASAP7_75t_L g1031 ( 
.A(n_942),
.Y(n_1031)
);

INVx2_ASAP7_75t_SL g1032 ( 
.A(n_983),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_925),
.Y(n_1033)
);

AOI22xp5_ASAP7_75t_L g1034 ( 
.A1(n_888),
.A2(n_909),
.B1(n_926),
.B2(n_945),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_1000),
.A2(n_984),
.B(n_976),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_912),
.B(n_897),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_923),
.B(n_913),
.Y(n_1037)
);

AND2x2_ASAP7_75t_L g1038 ( 
.A(n_913),
.B(n_916),
.Y(n_1038)
);

OAI22xp5_ASAP7_75t_L g1039 ( 
.A1(n_904),
.A2(n_906),
.B1(n_955),
.B2(n_995),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_904),
.B(n_906),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_L g1041 ( 
.A(n_898),
.B(n_945),
.Y(n_1041)
);

NAND2xp33_ASAP7_75t_L g1042 ( 
.A(n_1004),
.B(n_944),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_L g1043 ( 
.A(n_933),
.B(n_892),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_937),
.Y(n_1044)
);

BUFx4_ASAP7_75t_SL g1045 ( 
.A(n_966),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_981),
.Y(n_1046)
);

OR2x2_ASAP7_75t_L g1047 ( 
.A(n_910),
.B(n_933),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_910),
.B(n_931),
.Y(n_1048)
);

INVxp67_ASAP7_75t_SL g1049 ( 
.A(n_900),
.Y(n_1049)
);

INVx5_ASAP7_75t_L g1050 ( 
.A(n_1004),
.Y(n_1050)
);

BUFx12f_ASAP7_75t_L g1051 ( 
.A(n_952),
.Y(n_1051)
);

OAI22xp5_ASAP7_75t_SL g1052 ( 
.A1(n_885),
.A2(n_922),
.B1(n_882),
.B2(n_993),
.Y(n_1052)
);

INVx5_ASAP7_75t_L g1053 ( 
.A(n_988),
.Y(n_1053)
);

INVx2_ASAP7_75t_SL g1054 ( 
.A(n_988),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_954),
.B(n_882),
.Y(n_1055)
);

OAI22xp5_ASAP7_75t_L g1056 ( 
.A1(n_884),
.A2(n_982),
.B1(n_972),
.B2(n_970),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_884),
.B(n_970),
.Y(n_1057)
);

INVx3_ASAP7_75t_L g1058 ( 
.A(n_940),
.Y(n_1058)
);

CKINVDCx6p67_ASAP7_75t_R g1059 ( 
.A(n_988),
.Y(n_1059)
);

BUFx10_ASAP7_75t_L g1060 ( 
.A(n_940),
.Y(n_1060)
);

BUFx6f_ASAP7_75t_L g1061 ( 
.A(n_900),
.Y(n_1061)
);

BUFx2_ASAP7_75t_L g1062 ( 
.A(n_900),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_939),
.A2(n_941),
.B(n_943),
.Y(n_1063)
);

AOI21xp33_ASAP7_75t_L g1064 ( 
.A1(n_1002),
.A2(n_918),
.B(n_993),
.Y(n_1064)
);

INVx5_ASAP7_75t_L g1065 ( 
.A(n_928),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_972),
.B(n_982),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_924),
.B(n_927),
.Y(n_1067)
);

AND2x6_ASAP7_75t_L g1068 ( 
.A(n_883),
.B(n_919),
.Y(n_1068)
);

AND2x4_ASAP7_75t_L g1069 ( 
.A(n_997),
.B(n_986),
.Y(n_1069)
);

AND2x4_ASAP7_75t_L g1070 ( 
.A(n_978),
.B(n_986),
.Y(n_1070)
);

AND2x2_ASAP7_75t_L g1071 ( 
.A(n_934),
.B(n_905),
.Y(n_1071)
);

NOR2x1_ASAP7_75t_SL g1072 ( 
.A(n_956),
.B(n_947),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_935),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_939),
.A2(n_943),
.B(n_938),
.Y(n_1074)
);

AND2x2_ASAP7_75t_L g1075 ( 
.A(n_915),
.B(n_930),
.Y(n_1075)
);

HB1xp67_ASAP7_75t_L g1076 ( 
.A(n_958),
.Y(n_1076)
);

AND2x4_ASAP7_75t_L g1077 ( 
.A(n_978),
.B(n_958),
.Y(n_1077)
);

AOI22xp33_ASAP7_75t_L g1078 ( 
.A1(n_918),
.A2(n_964),
.B1(n_992),
.B2(n_917),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_L g1079 ( 
.A(n_992),
.B(n_947),
.Y(n_1079)
);

AOI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_936),
.A2(n_963),
.B1(n_989),
.B2(n_985),
.Y(n_1080)
);

BUFx10_ASAP7_75t_L g1081 ( 
.A(n_963),
.Y(n_1081)
);

OA21x2_ASAP7_75t_L g1082 ( 
.A1(n_911),
.A2(n_889),
.B(n_961),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_961),
.A2(n_957),
.B(n_965),
.Y(n_1083)
);

NOR2xp67_ASAP7_75t_L g1084 ( 
.A(n_962),
.B(n_951),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_936),
.B(n_951),
.Y(n_1085)
);

OR2x6_ASAP7_75t_L g1086 ( 
.A(n_953),
.B(n_960),
.Y(n_1086)
);

OR2x6_ASAP7_75t_L g1087 ( 
.A(n_960),
.B(n_962),
.Y(n_1087)
);

AND2x2_ASAP7_75t_L g1088 ( 
.A(n_1003),
.B(n_975),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_959),
.Y(n_1089)
);

NOR2x1_ASAP7_75t_L g1090 ( 
.A(n_959),
.B(n_949),
.Y(n_1090)
);

INVx1_ASAP7_75t_SL g1091 ( 
.A(n_948),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_950),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_890),
.Y(n_1093)
);

AND2x4_ASAP7_75t_L g1094 ( 
.A(n_946),
.B(n_896),
.Y(n_1094)
);

OR2x2_ASAP7_75t_L g1095 ( 
.A(n_929),
.B(n_896),
.Y(n_1095)
);

AOI22xp33_ASAP7_75t_SL g1096 ( 
.A1(n_929),
.A2(n_558),
.B1(n_552),
.B2(n_664),
.Y(n_1096)
);

INVx3_ASAP7_75t_L g1097 ( 
.A(n_929),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_SL g1098 ( 
.A(n_896),
.B(n_990),
.Y(n_1098)
);

AND2x4_ASAP7_75t_L g1099 ( 
.A(n_996),
.B(n_853),
.Y(n_1099)
);

BUFx2_ASAP7_75t_L g1100 ( 
.A(n_973),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_907),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_887),
.B(n_908),
.Y(n_1102)
);

OR2x2_ASAP7_75t_L g1103 ( 
.A(n_892),
.B(n_500),
.Y(n_1103)
);

BUFx6f_ASAP7_75t_L g1104 ( 
.A(n_886),
.Y(n_1104)
);

A2O1A1Ixp33_ASAP7_75t_L g1105 ( 
.A1(n_990),
.A2(n_833),
.B(n_829),
.C(n_866),
.Y(n_1105)
);

INVxp67_ASAP7_75t_SL g1106 ( 
.A(n_916),
.Y(n_1106)
);

OAI22xp5_ASAP7_75t_L g1107 ( 
.A1(n_990),
.A2(n_902),
.B1(n_887),
.B2(n_994),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_894),
.Y(n_1108)
);

AND2x2_ASAP7_75t_L g1109 ( 
.A(n_914),
.B(n_901),
.Y(n_1109)
);

AOI22xp5_ASAP7_75t_L g1110 ( 
.A1(n_990),
.A2(n_833),
.B1(n_902),
.B2(n_831),
.Y(n_1110)
);

AND2x2_ASAP7_75t_L g1111 ( 
.A(n_914),
.B(n_901),
.Y(n_1111)
);

NOR2xp67_ASAP7_75t_L g1112 ( 
.A(n_944),
.B(n_693),
.Y(n_1112)
);

INVx4_ASAP7_75t_L g1113 ( 
.A(n_944),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_SL g1114 ( 
.A(n_990),
.B(n_902),
.Y(n_1114)
);

OAI22xp5_ASAP7_75t_L g1115 ( 
.A1(n_990),
.A2(n_902),
.B1(n_887),
.B2(n_994),
.Y(n_1115)
);

OR2x2_ASAP7_75t_L g1116 ( 
.A(n_892),
.B(n_500),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_894),
.Y(n_1117)
);

BUFx3_ASAP7_75t_L g1118 ( 
.A(n_973),
.Y(n_1118)
);

OR2x2_ASAP7_75t_L g1119 ( 
.A(n_892),
.B(n_500),
.Y(n_1119)
);

AND2x2_ASAP7_75t_L g1120 ( 
.A(n_914),
.B(n_901),
.Y(n_1120)
);

AOI221x1_ASAP7_75t_L g1121 ( 
.A1(n_893),
.A2(n_918),
.B1(n_971),
.B2(n_980),
.C(n_968),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_887),
.B(n_908),
.Y(n_1122)
);

BUFx2_ASAP7_75t_L g1123 ( 
.A(n_973),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_921),
.Y(n_1124)
);

INVx2_ASAP7_75t_SL g1125 ( 
.A(n_983),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_893),
.A2(n_903),
.B(n_899),
.Y(n_1126)
);

INVx3_ASAP7_75t_L g1127 ( 
.A(n_987),
.Y(n_1127)
);

AND2x2_ASAP7_75t_L g1128 ( 
.A(n_914),
.B(n_901),
.Y(n_1128)
);

NOR2x1_ASAP7_75t_SL g1129 ( 
.A(n_944),
.B(n_956),
.Y(n_1129)
);

BUFx2_ASAP7_75t_L g1130 ( 
.A(n_973),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_893),
.A2(n_903),
.B(n_899),
.Y(n_1131)
);

NOR2xp67_ASAP7_75t_L g1132 ( 
.A(n_944),
.B(n_693),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_SL g1133 ( 
.A(n_990),
.B(n_902),
.Y(n_1133)
);

OR2x2_ASAP7_75t_L g1134 ( 
.A(n_892),
.B(n_500),
.Y(n_1134)
);

AND2x2_ASAP7_75t_L g1135 ( 
.A(n_914),
.B(n_901),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_894),
.Y(n_1136)
);

NOR2xp33_ASAP7_75t_L g1137 ( 
.A(n_1109),
.B(n_1111),
.Y(n_1137)
);

OAI22xp5_ASAP7_75t_L g1138 ( 
.A1(n_1048),
.A2(n_1040),
.B1(n_1106),
.B2(n_1096),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1006),
.B(n_1102),
.Y(n_1139)
);

OA21x2_ASAP7_75t_L g1140 ( 
.A1(n_1121),
.A2(n_1083),
.B(n_1074),
.Y(n_1140)
);

AOI22xp33_ASAP7_75t_L g1141 ( 
.A1(n_1052),
.A2(n_1012),
.B1(n_1115),
.B2(n_1107),
.Y(n_1141)
);

CKINVDCx20_ASAP7_75t_R g1142 ( 
.A(n_1009),
.Y(n_1142)
);

OAI22xp5_ASAP7_75t_L g1143 ( 
.A1(n_1122),
.A2(n_1110),
.B1(n_1034),
.B2(n_1024),
.Y(n_1143)
);

OA21x2_ASAP7_75t_L g1144 ( 
.A1(n_1063),
.A2(n_1026),
.B(n_1035),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1011),
.Y(n_1145)
);

AND2x2_ASAP7_75t_L g1146 ( 
.A(n_1110),
.B(n_1036),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_1108),
.Y(n_1147)
);

NAND2x1p5_ASAP7_75t_L g1148 ( 
.A(n_1030),
.B(n_1050),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_1117),
.Y(n_1149)
);

HB1xp67_ASAP7_75t_L g1150 ( 
.A(n_1037),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1033),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1092),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_1136),
.Y(n_1153)
);

NAND3xp33_ASAP7_75t_L g1154 ( 
.A(n_1105),
.B(n_1013),
.C(n_1012),
.Y(n_1154)
);

BUFx2_ASAP7_75t_R g1155 ( 
.A(n_1124),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_1088),
.Y(n_1156)
);

BUFx8_ASAP7_75t_L g1157 ( 
.A(n_1051),
.Y(n_1157)
);

BUFx2_ASAP7_75t_L g1158 ( 
.A(n_1038),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1097),
.Y(n_1159)
);

NAND2x1p5_ASAP7_75t_L g1160 ( 
.A(n_1030),
.B(n_1080),
.Y(n_1160)
);

BUFx3_ASAP7_75t_L g1161 ( 
.A(n_1015),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1120),
.B(n_1128),
.Y(n_1162)
);

CKINVDCx20_ASAP7_75t_R g1163 ( 
.A(n_1031),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1097),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1095),
.Y(n_1165)
);

AOI22xp33_ASAP7_75t_L g1166 ( 
.A1(n_1052),
.A2(n_1005),
.B1(n_1115),
.B2(n_1107),
.Y(n_1166)
);

CKINVDCx11_ASAP7_75t_R g1167 ( 
.A(n_1021),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_1089),
.Y(n_1168)
);

AND2x2_ASAP7_75t_L g1169 ( 
.A(n_1034),
.B(n_1020),
.Y(n_1169)
);

AOI22xp33_ASAP7_75t_SL g1170 ( 
.A1(n_1005),
.A2(n_1072),
.B1(n_1079),
.B2(n_1041),
.Y(n_1170)
);

BUFx3_ASAP7_75t_L g1171 ( 
.A(n_1118),
.Y(n_1171)
);

INVx8_ASAP7_75t_L g1172 ( 
.A(n_1053),
.Y(n_1172)
);

NAND2x1p5_ASAP7_75t_L g1173 ( 
.A(n_1080),
.B(n_1094),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1135),
.B(n_1027),
.Y(n_1174)
);

OAI22xp33_ASAP7_75t_L g1175 ( 
.A1(n_1047),
.A2(n_1134),
.B1(n_1116),
.B2(n_1103),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1044),
.Y(n_1176)
);

NOR2xp33_ASAP7_75t_L g1177 ( 
.A(n_1022),
.B(n_1020),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1101),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1071),
.Y(n_1179)
);

OA21x2_ASAP7_75t_L g1180 ( 
.A1(n_1010),
.A2(n_1131),
.B(n_1126),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1075),
.Y(n_1181)
);

AOI22xp33_ASAP7_75t_SL g1182 ( 
.A1(n_1067),
.A2(n_1043),
.B1(n_1039),
.B2(n_1019),
.Y(n_1182)
);

OR2x6_ASAP7_75t_L g1183 ( 
.A(n_1098),
.B(n_1087),
.Y(n_1183)
);

BUFx3_ASAP7_75t_L g1184 ( 
.A(n_1100),
.Y(n_1184)
);

AOI21x1_ASAP7_75t_L g1185 ( 
.A1(n_1025),
.A2(n_1039),
.B(n_1082),
.Y(n_1185)
);

AOI22xp33_ASAP7_75t_L g1186 ( 
.A1(n_1056),
.A2(n_1066),
.B1(n_1057),
.B2(n_1119),
.Y(n_1186)
);

CKINVDCx11_ASAP7_75t_R g1187 ( 
.A(n_1008),
.Y(n_1187)
);

AOI21x1_ASAP7_75t_L g1188 ( 
.A1(n_1057),
.A2(n_1084),
.B(n_1055),
.Y(n_1188)
);

AOI22xp33_ASAP7_75t_L g1189 ( 
.A1(n_1032),
.A2(n_1125),
.B1(n_1078),
.B2(n_1064),
.Y(n_1189)
);

OAI21x1_ASAP7_75t_L g1190 ( 
.A1(n_1090),
.A2(n_1084),
.B(n_1017),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1091),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1085),
.Y(n_1192)
);

HB1xp67_ASAP7_75t_L g1193 ( 
.A(n_1123),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1087),
.Y(n_1194)
);

AOI22xp33_ASAP7_75t_SL g1195 ( 
.A1(n_1069),
.A2(n_1129),
.B1(n_1018),
.B2(n_1031),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_1058),
.B(n_1087),
.Y(n_1196)
);

AOI22xp33_ASAP7_75t_L g1197 ( 
.A1(n_1064),
.A2(n_1130),
.B1(n_1099),
.B2(n_1029),
.Y(n_1197)
);

INVx1_ASAP7_75t_SL g1198 ( 
.A(n_1016),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1081),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1081),
.Y(n_1200)
);

INVxp67_ASAP7_75t_L g1201 ( 
.A(n_1076),
.Y(n_1201)
);

BUFx6f_ASAP7_75t_L g1202 ( 
.A(n_1065),
.Y(n_1202)
);

OAI22xp5_ASAP7_75t_L g1203 ( 
.A1(n_1023),
.A2(n_1132),
.B1(n_1112),
.B2(n_1016),
.Y(n_1203)
);

BUFx3_ASAP7_75t_L g1204 ( 
.A(n_1073),
.Y(n_1204)
);

AOI22xp33_ASAP7_75t_L g1205 ( 
.A1(n_1099),
.A2(n_1029),
.B1(n_1070),
.B2(n_1086),
.Y(n_1205)
);

OR2x2_ASAP7_75t_L g1206 ( 
.A(n_1086),
.B(n_1049),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1070),
.B(n_1077),
.Y(n_1207)
);

AND2x2_ASAP7_75t_L g1208 ( 
.A(n_1077),
.B(n_1086),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1062),
.B(n_1132),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1127),
.Y(n_1210)
);

AOI22xp33_ASAP7_75t_L g1211 ( 
.A1(n_1060),
.A2(n_1112),
.B1(n_1054),
.B2(n_1059),
.Y(n_1211)
);

AOI22xp33_ASAP7_75t_SL g1212 ( 
.A1(n_1042),
.A2(n_1028),
.B1(n_1053),
.B2(n_1113),
.Y(n_1212)
);

BUFx2_ASAP7_75t_L g1213 ( 
.A(n_1068),
.Y(n_1213)
);

BUFx3_ASAP7_75t_L g1214 ( 
.A(n_1053),
.Y(n_1214)
);

HB1xp67_ASAP7_75t_L g1215 ( 
.A(n_1065),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1065),
.B(n_1007),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1061),
.Y(n_1217)
);

NOR2xp33_ASAP7_75t_L g1218 ( 
.A(n_1046),
.B(n_1104),
.Y(n_1218)
);

INVx1_ASAP7_75t_SL g1219 ( 
.A(n_1045),
.Y(n_1219)
);

NOR2xp33_ASAP7_75t_L g1220 ( 
.A(n_1109),
.B(n_330),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_1014),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1011),
.Y(n_1222)
);

CKINVDCx11_ASAP7_75t_R g1223 ( 
.A(n_1051),
.Y(n_1223)
);

AND2x2_ASAP7_75t_L g1224 ( 
.A(n_1110),
.B(n_895),
.Y(n_1224)
);

INVx2_ASAP7_75t_L g1225 ( 
.A(n_1014),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_1014),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1093),
.Y(n_1227)
);

AND2x2_ASAP7_75t_L g1228 ( 
.A(n_1110),
.B(n_895),
.Y(n_1228)
);

BUFx3_ASAP7_75t_L g1229 ( 
.A(n_1015),
.Y(n_1229)
);

OAI22xp5_ASAP7_75t_SL g1230 ( 
.A1(n_1096),
.A2(n_552),
.B1(n_885),
.B2(n_812),
.Y(n_1230)
);

AND2x2_ASAP7_75t_L g1231 ( 
.A(n_1110),
.B(n_895),
.Y(n_1231)
);

OR2x2_ASAP7_75t_L g1232 ( 
.A(n_1057),
.B(n_1066),
.Y(n_1232)
);

HB1xp67_ASAP7_75t_L g1233 ( 
.A(n_1037),
.Y(n_1233)
);

AND2x2_ASAP7_75t_L g1234 ( 
.A(n_1110),
.B(n_895),
.Y(n_1234)
);

AOI22xp33_ASAP7_75t_L g1235 ( 
.A1(n_1114),
.A2(n_1133),
.B1(n_649),
.B2(n_1096),
.Y(n_1235)
);

AOI22xp33_ASAP7_75t_L g1236 ( 
.A1(n_1114),
.A2(n_1133),
.B1(n_649),
.B2(n_1096),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1093),
.Y(n_1237)
);

AOI22xp33_ASAP7_75t_L g1238 ( 
.A1(n_1114),
.A2(n_1133),
.B1(n_649),
.B2(n_1096),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_1152),
.Y(n_1239)
);

HB1xp67_ASAP7_75t_L g1240 ( 
.A(n_1158),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1232),
.B(n_1146),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1232),
.B(n_1146),
.Y(n_1242)
);

HB1xp67_ASAP7_75t_L g1243 ( 
.A(n_1158),
.Y(n_1243)
);

NOR2xp33_ASAP7_75t_L g1244 ( 
.A(n_1220),
.B(n_1162),
.Y(n_1244)
);

AND2x2_ASAP7_75t_L g1245 ( 
.A(n_1224),
.B(n_1228),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1192),
.B(n_1186),
.Y(n_1246)
);

AND2x2_ASAP7_75t_L g1247 ( 
.A(n_1224),
.B(n_1228),
.Y(n_1247)
);

OAI22xp5_ASAP7_75t_SL g1248 ( 
.A1(n_1230),
.A2(n_1182),
.B1(n_1141),
.B2(n_1166),
.Y(n_1248)
);

NOR2xp33_ASAP7_75t_L g1249 ( 
.A(n_1174),
.B(n_1137),
.Y(n_1249)
);

AND2x2_ASAP7_75t_L g1250 ( 
.A(n_1231),
.B(n_1234),
.Y(n_1250)
);

OR2x6_ASAP7_75t_L g1251 ( 
.A(n_1173),
.B(n_1183),
.Y(n_1251)
);

BUFx3_ASAP7_75t_L g1252 ( 
.A(n_1213),
.Y(n_1252)
);

AND2x2_ASAP7_75t_L g1253 ( 
.A(n_1231),
.B(n_1234),
.Y(n_1253)
);

CKINVDCx20_ASAP7_75t_R g1254 ( 
.A(n_1167),
.Y(n_1254)
);

HB1xp67_ASAP7_75t_L g1255 ( 
.A(n_1150),
.Y(n_1255)
);

NOR2x1_ASAP7_75t_R g1256 ( 
.A(n_1187),
.B(n_1223),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_1227),
.Y(n_1257)
);

OR2x2_ASAP7_75t_L g1258 ( 
.A(n_1165),
.B(n_1191),
.Y(n_1258)
);

BUFx2_ASAP7_75t_L g1259 ( 
.A(n_1183),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_1169),
.B(n_1165),
.Y(n_1260)
);

AND2x2_ASAP7_75t_L g1261 ( 
.A(n_1169),
.B(n_1237),
.Y(n_1261)
);

BUFx2_ASAP7_75t_L g1262 ( 
.A(n_1183),
.Y(n_1262)
);

AND2x2_ASAP7_75t_L g1263 ( 
.A(n_1156),
.B(n_1170),
.Y(n_1263)
);

BUFx3_ASAP7_75t_L g1264 ( 
.A(n_1213),
.Y(n_1264)
);

INVx4_ASAP7_75t_L g1265 ( 
.A(n_1172),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_1159),
.Y(n_1266)
);

NOR2xp33_ASAP7_75t_L g1267 ( 
.A(n_1198),
.B(n_1175),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1192),
.B(n_1143),
.Y(n_1268)
);

BUFx2_ASAP7_75t_L g1269 ( 
.A(n_1183),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_1159),
.Y(n_1270)
);

BUFx3_ASAP7_75t_L g1271 ( 
.A(n_1148),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1164),
.Y(n_1272)
);

AND2x2_ASAP7_75t_L g1273 ( 
.A(n_1156),
.B(n_1177),
.Y(n_1273)
);

BUFx2_ASAP7_75t_L g1274 ( 
.A(n_1194),
.Y(n_1274)
);

CKINVDCx9p33_ASAP7_75t_R g1275 ( 
.A(n_1218),
.Y(n_1275)
);

OAI21x1_ASAP7_75t_L g1276 ( 
.A1(n_1185),
.A2(n_1180),
.B(n_1190),
.Y(n_1276)
);

HB1xp67_ASAP7_75t_L g1277 ( 
.A(n_1233),
.Y(n_1277)
);

HB1xp67_ASAP7_75t_L g1278 ( 
.A(n_1193),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1191),
.Y(n_1279)
);

OAI21x1_ASAP7_75t_L g1280 ( 
.A1(n_1180),
.A2(n_1144),
.B(n_1188),
.Y(n_1280)
);

AND2x4_ASAP7_75t_L g1281 ( 
.A(n_1196),
.B(n_1208),
.Y(n_1281)
);

HB1xp67_ASAP7_75t_L g1282 ( 
.A(n_1168),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1188),
.Y(n_1283)
);

BUFx6f_ASAP7_75t_L g1284 ( 
.A(n_1148),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1173),
.Y(n_1285)
);

OR2x2_ASAP7_75t_L g1286 ( 
.A(n_1140),
.B(n_1154),
.Y(n_1286)
);

HB1xp67_ASAP7_75t_L g1287 ( 
.A(n_1168),
.Y(n_1287)
);

OR2x2_ASAP7_75t_L g1288 ( 
.A(n_1140),
.B(n_1138),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1173),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1140),
.Y(n_1290)
);

NOR2xp33_ASAP7_75t_L g1291 ( 
.A(n_1207),
.B(n_1184),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_1140),
.Y(n_1292)
);

AO21x2_ASAP7_75t_L g1293 ( 
.A1(n_1145),
.A2(n_1178),
.B(n_1151),
.Y(n_1293)
);

BUFx2_ASAP7_75t_L g1294 ( 
.A(n_1160),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1176),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1222),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1160),
.Y(n_1297)
);

BUFx3_ASAP7_75t_L g1298 ( 
.A(n_1148),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1160),
.Y(n_1299)
);

INVx3_ASAP7_75t_L g1300 ( 
.A(n_1196),
.Y(n_1300)
);

INVx2_ASAP7_75t_SL g1301 ( 
.A(n_1206),
.Y(n_1301)
);

NOR2xp33_ASAP7_75t_L g1302 ( 
.A(n_1184),
.B(n_1142),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1139),
.B(n_1238),
.Y(n_1303)
);

HB1xp67_ASAP7_75t_L g1304 ( 
.A(n_1179),
.Y(n_1304)
);

NOR2xp33_ASAP7_75t_L g1305 ( 
.A(n_1142),
.B(n_1155),
.Y(n_1305)
);

BUFx3_ASAP7_75t_L g1306 ( 
.A(n_1172),
.Y(n_1306)
);

NOR2x1_ASAP7_75t_R g1307 ( 
.A(n_1204),
.B(n_1229),
.Y(n_1307)
);

NAND2x1p5_ASAP7_75t_L g1308 ( 
.A(n_1199),
.B(n_1200),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1239),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1268),
.B(n_1236),
.Y(n_1310)
);

AND2x2_ASAP7_75t_L g1311 ( 
.A(n_1290),
.B(n_1235),
.Y(n_1311)
);

AND2x4_ASAP7_75t_L g1312 ( 
.A(n_1300),
.B(n_1208),
.Y(n_1312)
);

INVx4_ASAP7_75t_SL g1313 ( 
.A(n_1284),
.Y(n_1313)
);

INVxp67_ASAP7_75t_L g1314 ( 
.A(n_1240),
.Y(n_1314)
);

BUFx6f_ASAP7_75t_L g1315 ( 
.A(n_1290),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1292),
.B(n_1189),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1292),
.B(n_1197),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1260),
.B(n_1210),
.Y(n_1318)
);

BUFx3_ASAP7_75t_L g1319 ( 
.A(n_1308),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1268),
.B(n_1181),
.Y(n_1320)
);

OR2x2_ASAP7_75t_L g1321 ( 
.A(n_1286),
.B(n_1288),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1260),
.B(n_1266),
.Y(n_1322)
);

OAI221xp5_ASAP7_75t_SL g1323 ( 
.A1(n_1288),
.A2(n_1195),
.B1(n_1219),
.B2(n_1205),
.C(n_1211),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1241),
.B(n_1226),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1241),
.B(n_1226),
.Y(n_1325)
);

HB1xp67_ASAP7_75t_L g1326 ( 
.A(n_1243),
.Y(n_1326)
);

HB1xp67_ASAP7_75t_L g1327 ( 
.A(n_1255),
.Y(n_1327)
);

OAI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1303),
.A2(n_1206),
.B1(n_1204),
.B2(n_1163),
.Y(n_1328)
);

HB1xp67_ASAP7_75t_L g1329 ( 
.A(n_1277),
.Y(n_1329)
);

INVx2_ASAP7_75t_SL g1330 ( 
.A(n_1257),
.Y(n_1330)
);

OR2x2_ASAP7_75t_L g1331 ( 
.A(n_1286),
.B(n_1201),
.Y(n_1331)
);

AOI221xp5_ASAP7_75t_L g1332 ( 
.A1(n_1248),
.A2(n_1203),
.B1(n_1147),
.B2(n_1149),
.C(n_1153),
.Y(n_1332)
);

INVxp67_ASAP7_75t_SL g1333 ( 
.A(n_1283),
.Y(n_1333)
);

NOR2x1_ASAP7_75t_L g1334 ( 
.A(n_1283),
.B(n_1214),
.Y(n_1334)
);

NOR3xp33_ASAP7_75t_SL g1335 ( 
.A(n_1248),
.B(n_1209),
.C(n_1216),
.Y(n_1335)
);

BUFx3_ASAP7_75t_L g1336 ( 
.A(n_1271),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1270),
.B(n_1272),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1242),
.B(n_1221),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1242),
.B(n_1221),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1261),
.B(n_1225),
.Y(n_1340)
);

INVxp67_ASAP7_75t_L g1341 ( 
.A(n_1293),
.Y(n_1341)
);

INVx2_ASAP7_75t_SL g1342 ( 
.A(n_1251),
.Y(n_1342)
);

OAI22xp33_ASAP7_75t_L g1343 ( 
.A1(n_1303),
.A2(n_1163),
.B1(n_1171),
.B2(n_1229),
.Y(n_1343)
);

CKINVDCx12_ASAP7_75t_R g1344 ( 
.A(n_1256),
.Y(n_1344)
);

OR2x2_ASAP7_75t_L g1345 ( 
.A(n_1258),
.B(n_1217),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1327),
.B(n_1245),
.Y(n_1346)
);

NAND3xp33_ASAP7_75t_L g1347 ( 
.A(n_1335),
.B(n_1267),
.C(n_1244),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1329),
.B(n_1245),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1322),
.B(n_1247),
.Y(n_1349)
);

NAND3xp33_ASAP7_75t_L g1350 ( 
.A(n_1335),
.B(n_1246),
.C(n_1249),
.Y(n_1350)
);

AOI22xp33_ASAP7_75t_L g1351 ( 
.A1(n_1328),
.A2(n_1251),
.B1(n_1263),
.B2(n_1294),
.Y(n_1351)
);

AOI221xp5_ASAP7_75t_L g1352 ( 
.A1(n_1332),
.A2(n_1278),
.B1(n_1253),
.B2(n_1247),
.C(n_1250),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1326),
.B(n_1250),
.Y(n_1353)
);

AOI22xp33_ASAP7_75t_L g1354 ( 
.A1(n_1332),
.A2(n_1251),
.B1(n_1263),
.B2(n_1259),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1324),
.B(n_1253),
.Y(n_1355)
);

NAND3xp33_ASAP7_75t_L g1356 ( 
.A(n_1310),
.B(n_1246),
.C(n_1304),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1324),
.B(n_1301),
.Y(n_1357)
);

NAND4xp25_ASAP7_75t_SL g1358 ( 
.A(n_1334),
.B(n_1254),
.C(n_1321),
.D(n_1320),
.Y(n_1358)
);

AOI22xp33_ASAP7_75t_L g1359 ( 
.A1(n_1343),
.A2(n_1251),
.B1(n_1262),
.B2(n_1269),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1325),
.B(n_1273),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1309),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1338),
.B(n_1273),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1337),
.B(n_1285),
.Y(n_1363)
);

OA21x2_ASAP7_75t_L g1364 ( 
.A1(n_1341),
.A2(n_1280),
.B(n_1276),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1339),
.B(n_1293),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1317),
.B(n_1289),
.Y(n_1366)
);

OAI22xp5_ASAP7_75t_L g1367 ( 
.A1(n_1323),
.A2(n_1252),
.B1(n_1264),
.B2(n_1212),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_SL g1368 ( 
.A(n_1319),
.B(n_1284),
.Y(n_1368)
);

NAND3xp33_ASAP7_75t_L g1369 ( 
.A(n_1323),
.B(n_1291),
.C(n_1295),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1314),
.B(n_1293),
.Y(n_1370)
);

NAND3xp33_ASAP7_75t_L g1371 ( 
.A(n_1320),
.B(n_1331),
.C(n_1296),
.Y(n_1371)
);

NAND3xp33_ASAP7_75t_L g1372 ( 
.A(n_1331),
.B(n_1295),
.C(n_1296),
.Y(n_1372)
);

OAI221xp5_ASAP7_75t_L g1373 ( 
.A1(n_1342),
.A2(n_1302),
.B1(n_1297),
.B2(n_1299),
.C(n_1305),
.Y(n_1373)
);

OAI22xp5_ASAP7_75t_L g1374 ( 
.A1(n_1340),
.A2(n_1264),
.B1(n_1252),
.B2(n_1345),
.Y(n_1374)
);

OAI221xp5_ASAP7_75t_L g1375 ( 
.A1(n_1342),
.A2(n_1298),
.B1(n_1271),
.B2(n_1161),
.C(n_1171),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1317),
.B(n_1274),
.Y(n_1376)
);

AOI21xp5_ASAP7_75t_SL g1377 ( 
.A1(n_1319),
.A2(n_1307),
.B(n_1306),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1318),
.B(n_1282),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1317),
.B(n_1274),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1318),
.B(n_1287),
.Y(n_1380)
);

NAND3xp33_ASAP7_75t_L g1381 ( 
.A(n_1334),
.B(n_1284),
.C(n_1279),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1312),
.B(n_1281),
.Y(n_1382)
);

NAND3xp33_ASAP7_75t_L g1383 ( 
.A(n_1341),
.B(n_1284),
.C(n_1279),
.Y(n_1383)
);

OR2x2_ASAP7_75t_L g1384 ( 
.A(n_1370),
.B(n_1321),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1361),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1361),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1365),
.B(n_1333),
.Y(n_1387)
);

INVx4_ASAP7_75t_L g1388 ( 
.A(n_1364),
.Y(n_1388)
);

AOI22xp33_ASAP7_75t_L g1389 ( 
.A1(n_1347),
.A2(n_1358),
.B1(n_1350),
.B2(n_1367),
.Y(n_1389)
);

HB1xp67_ASAP7_75t_L g1390 ( 
.A(n_1376),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1372),
.Y(n_1391)
);

BUFx3_ASAP7_75t_L g1392 ( 
.A(n_1375),
.Y(n_1392)
);

INVx5_ASAP7_75t_L g1393 ( 
.A(n_1377),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1349),
.B(n_1363),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1349),
.B(n_1315),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1372),
.Y(n_1396)
);

INVx1_ASAP7_75t_SL g1397 ( 
.A(n_1376),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1371),
.B(n_1333),
.Y(n_1398)
);

OR2x2_ASAP7_75t_L g1399 ( 
.A(n_1371),
.B(n_1330),
.Y(n_1399)
);

BUFx2_ASAP7_75t_L g1400 ( 
.A(n_1379),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1378),
.Y(n_1401)
);

BUFx2_ASAP7_75t_L g1402 ( 
.A(n_1379),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1366),
.B(n_1342),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1356),
.B(n_1330),
.Y(n_1404)
);

BUFx2_ASAP7_75t_L g1405 ( 
.A(n_1366),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1356),
.B(n_1316),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1382),
.B(n_1311),
.Y(n_1407)
);

OR2x2_ASAP7_75t_L g1408 ( 
.A(n_1353),
.B(n_1309),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1364),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1380),
.Y(n_1410)
);

AND2x4_ASAP7_75t_L g1411 ( 
.A(n_1368),
.B(n_1313),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1357),
.B(n_1316),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1355),
.B(n_1311),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1405),
.B(n_1312),
.Y(n_1414)
);

NOR2xp33_ASAP7_75t_L g1415 ( 
.A(n_1392),
.B(n_1344),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1386),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1386),
.Y(n_1417)
);

OR2x2_ASAP7_75t_L g1418 ( 
.A(n_1384),
.B(n_1391),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1399),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1405),
.B(n_1312),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1407),
.B(n_1312),
.Y(n_1421)
);

AOI22xp33_ASAP7_75t_L g1422 ( 
.A1(n_1389),
.A2(n_1392),
.B1(n_1347),
.B2(n_1350),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1385),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1407),
.B(n_1412),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1385),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1407),
.B(n_1346),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1385),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1400),
.B(n_1348),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_SL g1429 ( 
.A(n_1392),
.B(n_1369),
.Y(n_1429)
);

OR2x2_ASAP7_75t_L g1430 ( 
.A(n_1384),
.B(n_1360),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1399),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1399),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1400),
.B(n_1336),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1402),
.B(n_1336),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1408),
.Y(n_1435)
);

OR2x2_ASAP7_75t_L g1436 ( 
.A(n_1391),
.B(n_1362),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1409),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1402),
.B(n_1395),
.Y(n_1438)
);

OAI21xp33_ASAP7_75t_SL g1439 ( 
.A1(n_1396),
.A2(n_1377),
.B(n_1352),
.Y(n_1439)
);

INVx2_ASAP7_75t_SL g1440 ( 
.A(n_1403),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1408),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1408),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1395),
.B(n_1390),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1409),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1398),
.Y(n_1445)
);

OR2x2_ASAP7_75t_L g1446 ( 
.A(n_1396),
.B(n_1374),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1398),
.Y(n_1447)
);

OR2x2_ASAP7_75t_L g1448 ( 
.A(n_1387),
.B(n_1374),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1412),
.B(n_1311),
.Y(n_1449)
);

HB1xp67_ASAP7_75t_L g1450 ( 
.A(n_1404),
.Y(n_1450)
);

OR2x2_ASAP7_75t_L g1451 ( 
.A(n_1387),
.B(n_1383),
.Y(n_1451)
);

INVx1_ASAP7_75t_SL g1452 ( 
.A(n_1404),
.Y(n_1452)
);

OR2x2_ASAP7_75t_L g1453 ( 
.A(n_1446),
.B(n_1406),
.Y(n_1453)
);

AND2x4_ASAP7_75t_L g1454 ( 
.A(n_1438),
.B(n_1393),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1416),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1438),
.B(n_1390),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1422),
.B(n_1429),
.Y(n_1457)
);

AND2x4_ASAP7_75t_L g1458 ( 
.A(n_1443),
.B(n_1393),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1437),
.Y(n_1459)
);

AOI32xp33_ASAP7_75t_L g1460 ( 
.A1(n_1439),
.A2(n_1406),
.A3(n_1367),
.B1(n_1411),
.B2(n_1397),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1443),
.B(n_1394),
.Y(n_1461)
);

OR2x6_ASAP7_75t_L g1462 ( 
.A(n_1419),
.B(n_1284),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1437),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1421),
.B(n_1394),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1450),
.B(n_1401),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1416),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1452),
.B(n_1401),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1421),
.B(n_1394),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1417),
.Y(n_1469)
);

NOR2xp33_ASAP7_75t_L g1470 ( 
.A(n_1415),
.B(n_1256),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1414),
.B(n_1420),
.Y(n_1471)
);

INVxp67_ASAP7_75t_L g1472 ( 
.A(n_1436),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1414),
.B(n_1393),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1420),
.B(n_1440),
.Y(n_1474)
);

AND2x4_ASAP7_75t_L g1475 ( 
.A(n_1431),
.B(n_1432),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1452),
.B(n_1410),
.Y(n_1476)
);

AND2x2_ASAP7_75t_SL g1477 ( 
.A(n_1446),
.B(n_1351),
.Y(n_1477)
);

AOI32xp33_ASAP7_75t_L g1478 ( 
.A1(n_1439),
.A2(n_1447),
.A3(n_1445),
.B1(n_1434),
.B2(n_1433),
.Y(n_1478)
);

OAI22xp5_ASAP7_75t_L g1479 ( 
.A1(n_1448),
.A2(n_1354),
.B1(n_1369),
.B2(n_1393),
.Y(n_1479)
);

NOR2xp67_ASAP7_75t_L g1480 ( 
.A(n_1440),
.B(n_1393),
.Y(n_1480)
);

NOR2x1_ASAP7_75t_L g1481 ( 
.A(n_1418),
.B(n_1381),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1433),
.B(n_1393),
.Y(n_1482)
);

INVx2_ASAP7_75t_SL g1483 ( 
.A(n_1434),
.Y(n_1483)
);

NOR2xp33_ASAP7_75t_L g1484 ( 
.A(n_1426),
.B(n_1157),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1417),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1428),
.B(n_1393),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1436),
.B(n_1410),
.Y(n_1487)
);

NOR2x1_ASAP7_75t_L g1488 ( 
.A(n_1418),
.B(n_1381),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1431),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1428),
.B(n_1393),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1424),
.B(n_1395),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1445),
.B(n_1413),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_SL g1493 ( 
.A(n_1430),
.B(n_1411),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1432),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1419),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1455),
.Y(n_1496)
);

NAND2xp33_ASAP7_75t_SL g1497 ( 
.A(n_1457),
.B(n_1448),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1459),
.Y(n_1498)
);

INVx1_ASAP7_75t_SL g1499 ( 
.A(n_1482),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1482),
.B(n_1419),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1455),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1466),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1466),
.Y(n_1503)
);

OAI22xp5_ASAP7_75t_L g1504 ( 
.A1(n_1460),
.A2(n_1373),
.B1(n_1359),
.B2(n_1411),
.Y(n_1504)
);

AND2x4_ASAP7_75t_L g1505 ( 
.A(n_1480),
.B(n_1447),
.Y(n_1505)
);

BUFx2_ASAP7_75t_L g1506 ( 
.A(n_1483),
.Y(n_1506)
);

INVx1_ASAP7_75t_SL g1507 ( 
.A(n_1453),
.Y(n_1507)
);

AND2x4_ASAP7_75t_L g1508 ( 
.A(n_1454),
.B(n_1435),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1469),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1469),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1477),
.B(n_1449),
.Y(n_1511)
);

HB1xp67_ASAP7_75t_L g1512 ( 
.A(n_1483),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1459),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1477),
.B(n_1451),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1456),
.B(n_1435),
.Y(n_1515)
);

OR2x2_ASAP7_75t_L g1516 ( 
.A(n_1453),
.B(n_1451),
.Y(n_1516)
);

OR2x2_ASAP7_75t_L g1517 ( 
.A(n_1487),
.B(n_1441),
.Y(n_1517)
);

OR2x2_ASAP7_75t_L g1518 ( 
.A(n_1472),
.B(n_1441),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_SL g1519 ( 
.A(n_1478),
.B(n_1411),
.Y(n_1519)
);

INVx1_ASAP7_75t_SL g1520 ( 
.A(n_1470),
.Y(n_1520)
);

INVx3_ASAP7_75t_L g1521 ( 
.A(n_1454),
.Y(n_1521)
);

OR2x2_ASAP7_75t_L g1522 ( 
.A(n_1465),
.B(n_1492),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1485),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1462),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1485),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1462),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1456),
.B(n_1442),
.Y(n_1527)
);

HB1xp67_ASAP7_75t_L g1528 ( 
.A(n_1481),
.Y(n_1528)
);

OR2x6_ASAP7_75t_L g1529 ( 
.A(n_1488),
.B(n_1265),
.Y(n_1529)
);

INVx1_ASAP7_75t_SL g1530 ( 
.A(n_1486),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1461),
.B(n_1442),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1496),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1506),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1520),
.B(n_1461),
.Y(n_1534)
);

XOR2x2_ASAP7_75t_L g1535 ( 
.A(n_1514),
.B(n_1484),
.Y(n_1535)
);

AOI222xp33_ASAP7_75t_L g1536 ( 
.A1(n_1497),
.A2(n_1479),
.B1(n_1467),
.B2(n_1476),
.C1(n_1494),
.C2(n_1489),
.Y(n_1536)
);

OAI22xp5_ASAP7_75t_L g1537 ( 
.A1(n_1528),
.A2(n_1493),
.B1(n_1383),
.B2(n_1454),
.Y(n_1537)
);

INVxp67_ASAP7_75t_L g1538 ( 
.A(n_1512),
.Y(n_1538)
);

AOI22xp33_ASAP7_75t_L g1539 ( 
.A1(n_1519),
.A2(n_1511),
.B1(n_1504),
.B2(n_1530),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1496),
.Y(n_1540)
);

NAND2x1_ASAP7_75t_L g1541 ( 
.A(n_1529),
.B(n_1458),
.Y(n_1541)
);

NOR2xp33_ASAP7_75t_L g1542 ( 
.A(n_1507),
.B(n_1157),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1501),
.Y(n_1543)
);

AOI22xp5_ASAP7_75t_L g1544 ( 
.A1(n_1499),
.A2(n_1458),
.B1(n_1486),
.B2(n_1490),
.Y(n_1544)
);

OAI33xp33_ASAP7_75t_L g1545 ( 
.A1(n_1501),
.A2(n_1494),
.A3(n_1489),
.B1(n_1495),
.B2(n_1463),
.B3(n_1425),
.Y(n_1545)
);

OR2x2_ASAP7_75t_L g1546 ( 
.A(n_1516),
.B(n_1491),
.Y(n_1546)
);

OAI22xp5_ASAP7_75t_L g1547 ( 
.A1(n_1529),
.A2(n_1490),
.B1(n_1458),
.B2(n_1474),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1502),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1506),
.Y(n_1549)
);

AND2x4_ASAP7_75t_L g1550 ( 
.A(n_1521),
.B(n_1475),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1521),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1502),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1503),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1503),
.Y(n_1554)
);

OAI21xp33_ASAP7_75t_L g1555 ( 
.A1(n_1522),
.A2(n_1475),
.B(n_1473),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1509),
.Y(n_1556)
);

AOI221xp5_ASAP7_75t_L g1557 ( 
.A1(n_1509),
.A2(n_1475),
.B1(n_1495),
.B2(n_1463),
.C(n_1388),
.Y(n_1557)
);

NOR2xp33_ASAP7_75t_L g1558 ( 
.A(n_1542),
.B(n_1534),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1533),
.B(n_1515),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_SL g1560 ( 
.A(n_1536),
.B(n_1521),
.Y(n_1560)
);

NOR2xp33_ASAP7_75t_L g1561 ( 
.A(n_1538),
.B(n_1522),
.Y(n_1561)
);

OAI22xp5_ASAP7_75t_L g1562 ( 
.A1(n_1539),
.A2(n_1529),
.B1(n_1516),
.B2(n_1521),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1549),
.B(n_1515),
.Y(n_1563)
);

INVx1_ASAP7_75t_SL g1564 ( 
.A(n_1550),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1555),
.B(n_1527),
.Y(n_1565)
);

HB1xp67_ASAP7_75t_L g1566 ( 
.A(n_1550),
.Y(n_1566)
);

INVxp67_ASAP7_75t_L g1567 ( 
.A(n_1535),
.Y(n_1567)
);

INVx1_ASAP7_75t_SL g1568 ( 
.A(n_1546),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1536),
.B(n_1551),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1532),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1544),
.B(n_1527),
.Y(n_1571)
);

AOI22xp33_ASAP7_75t_L g1572 ( 
.A1(n_1537),
.A2(n_1529),
.B1(n_1508),
.B2(n_1547),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1541),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1540),
.Y(n_1574)
);

OR2x6_ASAP7_75t_L g1575 ( 
.A(n_1543),
.B(n_1529),
.Y(n_1575)
);

HB1xp67_ASAP7_75t_L g1576 ( 
.A(n_1548),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1547),
.B(n_1500),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1566),
.Y(n_1578)
);

AOI21xp5_ASAP7_75t_L g1579 ( 
.A1(n_1560),
.A2(n_1537),
.B(n_1545),
.Y(n_1579)
);

OAI211xp5_ASAP7_75t_L g1580 ( 
.A1(n_1560),
.A2(n_1572),
.B(n_1569),
.C(n_1567),
.Y(n_1580)
);

OAI22xp33_ASAP7_75t_L g1581 ( 
.A1(n_1562),
.A2(n_1557),
.B1(n_1518),
.B2(n_1517),
.Y(n_1581)
);

OAI211xp5_ASAP7_75t_SL g1582 ( 
.A1(n_1558),
.A2(n_1568),
.B(n_1561),
.C(n_1564),
.Y(n_1582)
);

NAND4xp25_ASAP7_75t_L g1583 ( 
.A(n_1565),
.B(n_1557),
.C(n_1553),
.D(n_1554),
.Y(n_1583)
);

OAI22xp5_ASAP7_75t_L g1584 ( 
.A1(n_1559),
.A2(n_1518),
.B1(n_1473),
.B2(n_1505),
.Y(n_1584)
);

AOI21xp5_ASAP7_75t_L g1585 ( 
.A1(n_1573),
.A2(n_1545),
.B(n_1552),
.Y(n_1585)
);

OAI21xp33_ASAP7_75t_L g1586 ( 
.A1(n_1571),
.A2(n_1500),
.B(n_1508),
.Y(n_1586)
);

AOI221xp5_ASAP7_75t_L g1587 ( 
.A1(n_1571),
.A2(n_1563),
.B1(n_1576),
.B2(n_1577),
.C(n_1570),
.Y(n_1587)
);

OAI211xp5_ASAP7_75t_SL g1588 ( 
.A1(n_1573),
.A2(n_1556),
.B(n_1510),
.C(n_1523),
.Y(n_1588)
);

OAI21xp33_ASAP7_75t_SL g1589 ( 
.A1(n_1577),
.A2(n_1523),
.B(n_1510),
.Y(n_1589)
);

CKINVDCx20_ASAP7_75t_R g1590 ( 
.A(n_1574),
.Y(n_1590)
);

NAND4xp75_ASAP7_75t_L g1591 ( 
.A(n_1579),
.B(n_1578),
.C(n_1587),
.D(n_1585),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1580),
.B(n_1574),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1586),
.B(n_1508),
.Y(n_1593)
);

INVxp67_ASAP7_75t_L g1594 ( 
.A(n_1583),
.Y(n_1594)
);

NAND4xp75_ASAP7_75t_L g1595 ( 
.A(n_1589),
.B(n_1582),
.C(n_1581),
.D(n_1590),
.Y(n_1595)
);

BUFx2_ASAP7_75t_L g1596 ( 
.A(n_1584),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1588),
.Y(n_1597)
);

OAI22xp33_ASAP7_75t_L g1598 ( 
.A1(n_1579),
.A2(n_1575),
.B1(n_1517),
.B2(n_1462),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1578),
.B(n_1531),
.Y(n_1599)
);

NAND4xp75_ASAP7_75t_L g1600 ( 
.A(n_1579),
.B(n_1525),
.C(n_1498),
.D(n_1513),
.Y(n_1600)
);

AOI211xp5_ASAP7_75t_L g1601 ( 
.A1(n_1580),
.A2(n_1307),
.B(n_1505),
.C(n_1525),
.Y(n_1601)
);

NAND4xp25_ASAP7_75t_L g1602 ( 
.A(n_1601),
.B(n_1508),
.C(n_1505),
.D(n_1498),
.Y(n_1602)
);

OAI21xp33_ASAP7_75t_L g1603 ( 
.A1(n_1594),
.A2(n_1575),
.B(n_1526),
.Y(n_1603)
);

AOI22xp33_ASAP7_75t_L g1604 ( 
.A1(n_1596),
.A2(n_1575),
.B1(n_1505),
.B2(n_1526),
.Y(n_1604)
);

NOR2x1_ASAP7_75t_L g1605 ( 
.A(n_1595),
.B(n_1575),
.Y(n_1605)
);

NOR2xp67_ASAP7_75t_L g1606 ( 
.A(n_1599),
.B(n_1498),
.Y(n_1606)
);

AOI211xp5_ASAP7_75t_L g1607 ( 
.A1(n_1598),
.A2(n_1524),
.B(n_1513),
.C(n_1531),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1606),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1603),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1607),
.Y(n_1610)
);

OAI22xp5_ASAP7_75t_L g1611 ( 
.A1(n_1604),
.A2(n_1591),
.B1(n_1592),
.B2(n_1600),
.Y(n_1611)
);

NOR2x1_ASAP7_75t_L g1612 ( 
.A(n_1605),
.B(n_1597),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_1602),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1604),
.B(n_1601),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_1608),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1609),
.B(n_1593),
.Y(n_1616)
);

NOR2xp33_ASAP7_75t_R g1617 ( 
.A(n_1610),
.B(n_1157),
.Y(n_1617)
);

NAND3x1_ASAP7_75t_L g1618 ( 
.A(n_1612),
.B(n_1474),
.C(n_1471),
.Y(n_1618)
);

NAND4xp75_ASAP7_75t_L g1619 ( 
.A(n_1614),
.B(n_1513),
.C(n_1524),
.D(n_1471),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1618),
.Y(n_1620)
);

NOR2xp33_ASAP7_75t_L g1621 ( 
.A(n_1619),
.B(n_1611),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1616),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1620),
.Y(n_1623)
);

OR4x2_ASAP7_75t_L g1624 ( 
.A(n_1623),
.B(n_1617),
.C(n_1621),
.D(n_1622),
.Y(n_1624)
);

AOI21xp5_ASAP7_75t_L g1625 ( 
.A1(n_1624),
.A2(n_1615),
.B(n_1613),
.Y(n_1625)
);

OAI22x1_ASAP7_75t_L g1626 ( 
.A1(n_1624),
.A2(n_1444),
.B1(n_1437),
.B2(n_1215),
.Y(n_1626)
);

AOI21x1_ASAP7_75t_L g1627 ( 
.A1(n_1625),
.A2(n_1462),
.B(n_1444),
.Y(n_1627)
);

NOR2x1p5_ASAP7_75t_L g1628 ( 
.A(n_1626),
.B(n_1161),
.Y(n_1628)
);

OAI22x1_ASAP7_75t_L g1629 ( 
.A1(n_1627),
.A2(n_1444),
.B1(n_1491),
.B2(n_1388),
.Y(n_1629)
);

OR2x2_ASAP7_75t_L g1630 ( 
.A(n_1628),
.B(n_1464),
.Y(n_1630)
);

OAI21xp5_ASAP7_75t_L g1631 ( 
.A1(n_1630),
.A2(n_1468),
.B(n_1464),
.Y(n_1631)
);

AOI322xp5_ASAP7_75t_L g1632 ( 
.A1(n_1631),
.A2(n_1629),
.A3(n_1468),
.B1(n_1411),
.B2(n_1427),
.C1(n_1423),
.C2(n_1425),
.Y(n_1632)
);

AOI221xp5_ASAP7_75t_L g1633 ( 
.A1(n_1632),
.A2(n_1423),
.B1(n_1427),
.B2(n_1214),
.C(n_1388),
.Y(n_1633)
);

AOI211xp5_ASAP7_75t_L g1634 ( 
.A1(n_1633),
.A2(n_1202),
.B(n_1275),
.C(n_1306),
.Y(n_1634)
);


endmodule