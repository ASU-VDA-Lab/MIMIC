module fake_netlist_6_750_n_738 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_738);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_738;

wire n_591;
wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_578;
wire n_703;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_725;
wire n_358;
wire n_160;
wire n_449;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_255;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_222;
wire n_179;
wire n_248;
wire n_300;
wire n_517;
wire n_718;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_532;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_506;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_344;
wire n_581;
wire n_428;
wire n_609;
wire n_432;
wire n_641;
wire n_693;
wire n_167;
wire n_631;
wire n_174;
wire n_516;
wire n_153;
wire n_720;
wire n_525;
wire n_611;
wire n_156;
wire n_491;
wire n_656;
wire n_666;
wire n_371;
wire n_567;
wire n_189;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_155;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_163;
wire n_717;
wire n_330;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_699;
wire n_154;
wire n_551;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_252;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_152;
wire n_623;
wire n_599;
wire n_513;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_527;
wire n_474;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_325;
wire n_329;
wire n_464;
wire n_600;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_505;
wire n_240;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_556;
wire n_159;
wire n_157;
wire n_162;
wire n_692;
wire n_733;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_652;
wire n_553;
wire n_560;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_426;
wire n_317;
wire n_149;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_728;
wire n_681;
wire n_729;
wire n_151;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_410;
wire n_398;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_83),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_7),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_78),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_102),
.Y(n_152)
);

INVx1_ASAP7_75t_SL g153 ( 
.A(n_134),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_54),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_63),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_72),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_136),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_120),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g159 ( 
.A(n_118),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_46),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_6),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_96),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_141),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_16),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_99),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_52),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_127),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_71),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_143),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_115),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_20),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_77),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_135),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_23),
.Y(n_174)
);

BUFx2_ASAP7_75t_L g175 ( 
.A(n_15),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_25),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_111),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_79),
.B(n_104),
.Y(n_178)
);

BUFx2_ASAP7_75t_L g179 ( 
.A(n_125),
.Y(n_179)
);

INVx4_ASAP7_75t_R g180 ( 
.A(n_139),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_41),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_44),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_112),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_76),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_74),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_107),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_17),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_100),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_4),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_106),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_5),
.Y(n_191)
);

BUFx10_ASAP7_75t_L g192 ( 
.A(n_14),
.Y(n_192)
);

NOR2xp67_ASAP7_75t_L g193 ( 
.A(n_39),
.B(n_58),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_105),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_114),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_48),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_57),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_94),
.Y(n_198)
);

AND2x4_ASAP7_75t_L g199 ( 
.A(n_156),
.B(n_18),
.Y(n_199)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_156),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_179),
.B(n_0),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_159),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_170),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_191),
.Y(n_204)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_190),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_170),
.Y(n_206)
);

BUFx8_ASAP7_75t_SL g207 ( 
.A(n_175),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_190),
.Y(n_208)
);

OAI21x1_ASAP7_75t_L g209 ( 
.A1(n_155),
.A2(n_1),
.B(n_2),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_155),
.B(n_3),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_152),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_170),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_187),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_157),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_150),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_187),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_163),
.B(n_3),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_163),
.B(n_5),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_192),
.B(n_6),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_159),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_170),
.Y(n_221)
);

AND2x4_ASAP7_75t_L g222 ( 
.A(n_160),
.B(n_19),
.Y(n_222)
);

BUFx8_ASAP7_75t_SL g223 ( 
.A(n_186),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_162),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_192),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_225)
);

AND2x4_ASAP7_75t_L g226 ( 
.A(n_169),
.B(n_21),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_176),
.Y(n_227)
);

CKINVDCx11_ASAP7_75t_R g228 ( 
.A(n_192),
.Y(n_228)
);

OA21x2_ASAP7_75t_L g229 ( 
.A1(n_183),
.A2(n_10),
.B(n_11),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_186),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_161),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_184),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_195),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_196),
.B(n_11),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_197),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_198),
.Y(n_236)
);

INVx5_ASAP7_75t_L g237 ( 
.A(n_193),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_213),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_203),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_203),
.Y(n_240)
);

AND3x2_ASAP7_75t_L g241 ( 
.A(n_199),
.B(n_178),
.C(n_180),
.Y(n_241)
);

AND3x2_ASAP7_75t_L g242 ( 
.A(n_199),
.B(n_189),
.C(n_164),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_203),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_237),
.B(n_153),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_208),
.B(n_151),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_213),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_237),
.B(n_201),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_203),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_216),
.Y(n_249)
);

OR2x6_ASAP7_75t_L g250 ( 
.A(n_219),
.B(n_149),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_216),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_223),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_199),
.B(n_194),
.Y(n_253)
);

AND3x2_ASAP7_75t_L g254 ( 
.A(n_215),
.B(n_12),
.C(n_13),
.Y(n_254)
);

BUFx3_ASAP7_75t_L g255 ( 
.A(n_200),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_206),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_206),
.Y(n_257)
);

AO21x2_ASAP7_75t_L g258 ( 
.A1(n_210),
.A2(n_218),
.B(n_217),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_206),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_237),
.B(n_154),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_206),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_200),
.B(n_188),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_221),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_221),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_221),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_221),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_237),
.B(n_230),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_212),
.Y(n_268)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_212),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_235),
.Y(n_270)
);

AO21x2_ASAP7_75t_L g271 ( 
.A1(n_209),
.A2(n_234),
.B(n_219),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_237),
.B(n_158),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_212),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_212),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_212),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_223),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_204),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_236),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_233),
.Y(n_279)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_222),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_233),
.Y(n_281)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_222),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_282),
.B(n_280),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_239),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_282),
.B(n_222),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_282),
.B(n_226),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_239),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_R g288 ( 
.A(n_252),
.B(n_231),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_280),
.B(n_226),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_267),
.B(n_231),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_280),
.B(n_262),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_250),
.A2(n_166),
.B1(n_167),
.B2(n_168),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_253),
.B(n_220),
.Y(n_293)
);

INVx2_ASAP7_75t_SL g294 ( 
.A(n_245),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_250),
.B(n_207),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_245),
.B(n_165),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_279),
.Y(n_297)
);

OR2x6_ASAP7_75t_L g298 ( 
.A(n_250),
.B(n_202),
.Y(n_298)
);

NAND2xp33_ASAP7_75t_L g299 ( 
.A(n_247),
.B(n_171),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_255),
.B(n_228),
.Y(n_300)
);

NAND2xp33_ASAP7_75t_L g301 ( 
.A(n_277),
.B(n_172),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_255),
.B(n_205),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_258),
.B(n_205),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_258),
.B(n_211),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_250),
.A2(n_225),
.B1(n_174),
.B2(n_177),
.Y(n_305)
);

BUFx8_ASAP7_75t_L g306 ( 
.A(n_277),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_279),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_263),
.Y(n_308)
);

INVx8_ASAP7_75t_L g309 ( 
.A(n_252),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_240),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_258),
.B(n_214),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_244),
.B(n_228),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_L g313 ( 
.A1(n_271),
.A2(n_229),
.B1(n_232),
.B2(n_224),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_263),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_266),
.B(n_240),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_242),
.B(n_207),
.Y(n_316)
);

NAND2x1_ASAP7_75t_L g317 ( 
.A(n_269),
.B(n_229),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_260),
.B(n_173),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_266),
.B(n_233),
.Y(n_319)
);

NAND3xp33_ASAP7_75t_L g320 ( 
.A(n_270),
.B(n_229),
.C(n_235),
.Y(n_320)
);

BUFx5_ASAP7_75t_L g321 ( 
.A(n_273),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_272),
.B(n_181),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_278),
.B(n_182),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_243),
.Y(n_324)
);

INVx2_ASAP7_75t_SL g325 ( 
.A(n_241),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_243),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_248),
.B(n_233),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_248),
.Y(n_328)
);

INVx1_ASAP7_75t_SL g329 ( 
.A(n_276),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_271),
.B(n_227),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_256),
.B(n_236),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_256),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_271),
.B(n_227),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_278),
.B(n_185),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_257),
.B(n_259),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_257),
.B(n_209),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_259),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_261),
.Y(n_338)
);

INVx8_ASAP7_75t_L g339 ( 
.A(n_281),
.Y(n_339)
);

NAND2xp33_ASAP7_75t_L g340 ( 
.A(n_261),
.B(n_12),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_238),
.B(n_13),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_264),
.B(n_22),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_264),
.B(n_24),
.Y(n_343)
);

INVx1_ASAP7_75t_SL g344 ( 
.A(n_329),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_330),
.B(n_333),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_283),
.A2(n_291),
.B(n_286),
.Y(n_346)
);

INVx3_ASAP7_75t_L g347 ( 
.A(n_284),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_285),
.A2(n_281),
.B(n_275),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_289),
.A2(n_281),
.B(n_275),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_331),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_342),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_315),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_294),
.B(n_238),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_L g354 ( 
.A1(n_303),
.A2(n_274),
.B(n_273),
.Y(n_354)
);

A2O1A1Ixp33_ASAP7_75t_L g355 ( 
.A1(n_304),
.A2(n_246),
.B(n_249),
.C(n_251),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_311),
.B(n_265),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_302),
.B(n_265),
.Y(n_357)
);

INVx4_ASAP7_75t_L g358 ( 
.A(n_339),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_305),
.B(n_281),
.Y(n_359)
);

INVx4_ASAP7_75t_L g360 ( 
.A(n_339),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_339),
.A2(n_281),
.B(n_268),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_293),
.B(n_246),
.Y(n_362)
);

AND2x4_ASAP7_75t_L g363 ( 
.A(n_325),
.B(n_297),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_307),
.B(n_269),
.Y(n_364)
);

AOI221x1_ASAP7_75t_L g365 ( 
.A1(n_320),
.A2(n_274),
.B1(n_269),
.B2(n_268),
.C(n_251),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_335),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_334),
.B(n_249),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_312),
.B(n_254),
.Y(n_368)
);

BUFx12f_ASAP7_75t_L g369 ( 
.A(n_306),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_336),
.A2(n_81),
.B(n_147),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_317),
.A2(n_80),
.B(n_146),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_326),
.Y(n_372)
);

INVx3_ASAP7_75t_L g373 ( 
.A(n_287),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_313),
.B(n_308),
.Y(n_374)
);

BUFx12f_ASAP7_75t_L g375 ( 
.A(n_306),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_314),
.B(n_26),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_319),
.A2(n_82),
.B(n_145),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_300),
.B(n_14),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_296),
.B(n_292),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_321),
.B(n_27),
.Y(n_380)
);

AND2x4_ASAP7_75t_L g381 ( 
.A(n_323),
.B(n_28),
.Y(n_381)
);

A2O1A1Ixp33_ASAP7_75t_L g382 ( 
.A1(n_320),
.A2(n_15),
.B(n_16),
.C(n_17),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_290),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_327),
.A2(n_29),
.B(n_30),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_321),
.B(n_31),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_321),
.B(n_310),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_321),
.B(n_32),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_298),
.B(n_33),
.Y(n_388)
);

AOI21xp33_ASAP7_75t_L g389 ( 
.A1(n_298),
.A2(n_148),
.B(n_35),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_318),
.B(n_34),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_332),
.Y(n_391)
);

BUFx2_ASAP7_75t_L g392 ( 
.A(n_298),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_L g393 ( 
.A1(n_324),
.A2(n_36),
.B(n_37),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_343),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_338),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_340),
.A2(n_38),
.B1(n_40),
.B2(n_42),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_328),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_337),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_L g399 ( 
.A1(n_301),
.A2(n_43),
.B(n_45),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_295),
.Y(n_400)
);

INVx4_ASAP7_75t_L g401 ( 
.A(n_321),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_341),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_322),
.A2(n_47),
.B(n_49),
.Y(n_403)
);

OAI21xp33_ASAP7_75t_L g404 ( 
.A1(n_299),
.A2(n_50),
.B(n_51),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_316),
.A2(n_53),
.B(n_55),
.Y(n_405)
);

NOR2x1_ASAP7_75t_R g406 ( 
.A(n_288),
.B(n_56),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_309),
.B(n_59),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_309),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_309),
.B(n_60),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_330),
.B(n_61),
.Y(n_410)
);

INVx3_ASAP7_75t_L g411 ( 
.A(n_347),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_346),
.A2(n_62),
.B(n_64),
.Y(n_412)
);

NAND2xp33_ASAP7_75t_L g413 ( 
.A(n_345),
.B(n_65),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_397),
.Y(n_414)
);

BUFx3_ASAP7_75t_L g415 ( 
.A(n_344),
.Y(n_415)
);

AO31x2_ASAP7_75t_L g416 ( 
.A1(n_365),
.A2(n_66),
.A3(n_67),
.B(n_68),
.Y(n_416)
);

OAI21xp33_ASAP7_75t_L g417 ( 
.A1(n_402),
.A2(n_69),
.B(n_70),
.Y(n_417)
);

BUFx3_ASAP7_75t_L g418 ( 
.A(n_344),
.Y(n_418)
);

INVx8_ASAP7_75t_L g419 ( 
.A(n_363),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_352),
.B(n_73),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_350),
.B(n_75),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_366),
.B(n_84),
.Y(n_422)
);

OAI21x1_ASAP7_75t_L g423 ( 
.A1(n_348),
.A2(n_349),
.B(n_386),
.Y(n_423)
);

AOI21x1_ASAP7_75t_SL g424 ( 
.A1(n_410),
.A2(n_85),
.B(n_86),
.Y(n_424)
);

OAI21x1_ASAP7_75t_L g425 ( 
.A1(n_357),
.A2(n_144),
.B(n_88),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_353),
.B(n_383),
.Y(n_426)
);

OAI21x1_ASAP7_75t_L g427 ( 
.A1(n_364),
.A2(n_142),
.B(n_89),
.Y(n_427)
);

NAND3xp33_ASAP7_75t_SL g428 ( 
.A(n_379),
.B(n_87),
.C(n_90),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_398),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_367),
.B(n_91),
.Y(n_430)
);

A2O1A1Ixp33_ASAP7_75t_L g431 ( 
.A1(n_354),
.A2(n_92),
.B(n_93),
.C(n_95),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_378),
.B(n_97),
.Y(n_432)
);

AO21x1_ASAP7_75t_L g433 ( 
.A1(n_359),
.A2(n_389),
.B(n_356),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_362),
.B(n_98),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_372),
.Y(n_435)
);

OAI21x1_ASAP7_75t_L g436 ( 
.A1(n_371),
.A2(n_387),
.B(n_385),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_374),
.B(n_101),
.Y(n_437)
);

INVx2_ASAP7_75t_SL g438 ( 
.A(n_363),
.Y(n_438)
);

OR2x2_ASAP7_75t_L g439 ( 
.A(n_392),
.B(n_103),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_408),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_401),
.A2(n_108),
.B(n_109),
.Y(n_441)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_401),
.A2(n_110),
.B(n_113),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_L g443 ( 
.A1(n_355),
.A2(n_116),
.B(n_117),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_391),
.B(n_119),
.Y(n_444)
);

AO31x2_ASAP7_75t_L g445 ( 
.A1(n_382),
.A2(n_121),
.A3(n_122),
.B(n_123),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_395),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_381),
.B(n_124),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_373),
.Y(n_448)
);

AOI21xp5_ASAP7_75t_L g449 ( 
.A1(n_358),
.A2(n_126),
.B(n_128),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_400),
.B(n_129),
.Y(n_450)
);

BUFx10_ASAP7_75t_L g451 ( 
.A(n_409),
.Y(n_451)
);

AOI21x1_ASAP7_75t_L g452 ( 
.A1(n_361),
.A2(n_130),
.B(n_131),
.Y(n_452)
);

AND2x4_ASAP7_75t_L g453 ( 
.A(n_407),
.B(n_132),
.Y(n_453)
);

OAI22x1_ASAP7_75t_L g454 ( 
.A1(n_368),
.A2(n_133),
.B1(n_137),
.B2(n_138),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_381),
.B(n_140),
.Y(n_455)
);

OAI21xp33_ASAP7_75t_L g456 ( 
.A1(n_388),
.A2(n_404),
.B(n_390),
.Y(n_456)
);

AOI21x1_ASAP7_75t_L g457 ( 
.A1(n_376),
.A2(n_380),
.B(n_370),
.Y(n_457)
);

OAI21x1_ASAP7_75t_L g458 ( 
.A1(n_373),
.A2(n_399),
.B(n_403),
.Y(n_458)
);

OAI21x1_ASAP7_75t_L g459 ( 
.A1(n_393),
.A2(n_377),
.B(n_384),
.Y(n_459)
);

OAI22x1_ASAP7_75t_L g460 ( 
.A1(n_396),
.A2(n_375),
.B1(n_369),
.B2(n_406),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_351),
.B(n_394),
.Y(n_461)
);

A2O1A1Ixp33_ASAP7_75t_L g462 ( 
.A1(n_404),
.A2(n_396),
.B(n_405),
.C(n_394),
.Y(n_462)
);

OAI21x1_ASAP7_75t_L g463 ( 
.A1(n_351),
.A2(n_394),
.B(n_358),
.Y(n_463)
);

AOI21x1_ASAP7_75t_SL g464 ( 
.A1(n_351),
.A2(n_410),
.B(n_381),
.Y(n_464)
);

AO21x1_ASAP7_75t_L g465 ( 
.A1(n_443),
.A2(n_360),
.B(n_437),
.Y(n_465)
);

OAI21x1_ASAP7_75t_L g466 ( 
.A1(n_464),
.A2(n_458),
.B(n_459),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_461),
.A2(n_360),
.B(n_462),
.Y(n_467)
);

OA21x2_ASAP7_75t_L g468 ( 
.A1(n_433),
.A2(n_436),
.B(n_423),
.Y(n_468)
);

OR2x2_ASAP7_75t_L g469 ( 
.A(n_415),
.B(n_418),
.Y(n_469)
);

BUFx3_ASAP7_75t_L g470 ( 
.A(n_419),
.Y(n_470)
);

HB1xp67_ASAP7_75t_L g471 ( 
.A(n_426),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_446),
.Y(n_472)
);

INVx4_ASAP7_75t_L g473 ( 
.A(n_453),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_L g474 ( 
.A1(n_420),
.A2(n_430),
.B(n_422),
.Y(n_474)
);

BUFx3_ASAP7_75t_L g475 ( 
.A(n_419),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_448),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_440),
.Y(n_477)
);

A2O1A1Ixp33_ASAP7_75t_L g478 ( 
.A1(n_456),
.A2(n_447),
.B(n_455),
.C(n_432),
.Y(n_478)
);

OAI21x1_ASAP7_75t_L g479 ( 
.A1(n_463),
.A2(n_457),
.B(n_424),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_446),
.B(n_453),
.Y(n_480)
);

BUFx3_ASAP7_75t_L g481 ( 
.A(n_440),
.Y(n_481)
);

AO21x2_ASAP7_75t_L g482 ( 
.A1(n_428),
.A2(n_421),
.B(n_431),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_435),
.Y(n_483)
);

OAI21x1_ASAP7_75t_L g484 ( 
.A1(n_425),
.A2(n_427),
.B(n_452),
.Y(n_484)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_413),
.A2(n_434),
.B(n_444),
.Y(n_485)
);

AO21x2_ASAP7_75t_L g486 ( 
.A1(n_412),
.A2(n_417),
.B(n_449),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_451),
.Y(n_487)
);

BUFx2_ASAP7_75t_R g488 ( 
.A(n_439),
.Y(n_488)
);

OR3x4_ASAP7_75t_SL g489 ( 
.A(n_460),
.B(n_454),
.C(n_438),
.Y(n_489)
);

OA21x2_ASAP7_75t_L g490 ( 
.A1(n_414),
.A2(n_429),
.B(n_442),
.Y(n_490)
);

BUFx3_ASAP7_75t_L g491 ( 
.A(n_440),
.Y(n_491)
);

OAI21x1_ASAP7_75t_L g492 ( 
.A1(n_441),
.A2(n_411),
.B(n_414),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_411),
.B(n_450),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_429),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_451),
.Y(n_495)
);

BUFx12f_ASAP7_75t_L g496 ( 
.A(n_445),
.Y(n_496)
);

INVxp67_ASAP7_75t_SL g497 ( 
.A(n_445),
.Y(n_497)
);

AOI21xp5_ASAP7_75t_L g498 ( 
.A1(n_416),
.A2(n_401),
.B(n_345),
.Y(n_498)
);

OAI21x1_ASAP7_75t_L g499 ( 
.A1(n_416),
.A2(n_464),
.B(n_458),
.Y(n_499)
);

NAND2x1p5_ASAP7_75t_L g500 ( 
.A(n_445),
.B(n_463),
.Y(n_500)
);

OAI21x1_ASAP7_75t_L g501 ( 
.A1(n_464),
.A2(n_458),
.B(n_459),
.Y(n_501)
);

BUFx12f_ASAP7_75t_L g502 ( 
.A(n_415),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_448),
.Y(n_503)
);

NAND2x1p5_ASAP7_75t_L g504 ( 
.A(n_463),
.B(n_453),
.Y(n_504)
);

OAI21xp5_ASAP7_75t_L g505 ( 
.A1(n_437),
.A2(n_345),
.B(n_333),
.Y(n_505)
);

AND2x4_ASAP7_75t_L g506 ( 
.A(n_453),
.B(n_435),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_446),
.Y(n_507)
);

NAND2x1p5_ASAP7_75t_L g508 ( 
.A(n_473),
.B(n_492),
.Y(n_508)
);

OR2x2_ASAP7_75t_L g509 ( 
.A(n_471),
.B(n_507),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_472),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_494),
.Y(n_511)
);

BUFx2_ASAP7_75t_L g512 ( 
.A(n_469),
.Y(n_512)
);

AOI21xp33_ASAP7_75t_L g513 ( 
.A1(n_478),
.A2(n_505),
.B(n_480),
.Y(n_513)
);

BUFx3_ASAP7_75t_L g514 ( 
.A(n_502),
.Y(n_514)
);

HB1xp67_ASAP7_75t_L g515 ( 
.A(n_469),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_476),
.Y(n_516)
);

HB1xp67_ASAP7_75t_L g517 ( 
.A(n_502),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_480),
.B(n_506),
.Y(n_518)
);

AOI22xp33_ASAP7_75t_L g519 ( 
.A1(n_506),
.A2(n_473),
.B1(n_483),
.B2(n_465),
.Y(n_519)
);

BUFx2_ASAP7_75t_L g520 ( 
.A(n_506),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_476),
.Y(n_521)
);

BUFx2_ASAP7_75t_L g522 ( 
.A(n_481),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_477),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_477),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_503),
.Y(n_525)
);

INVx1_ASAP7_75t_SL g526 ( 
.A(n_487),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_503),
.Y(n_527)
);

NAND2x1p5_ASAP7_75t_L g528 ( 
.A(n_473),
.B(n_492),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_490),
.Y(n_529)
);

HB1xp67_ASAP7_75t_L g530 ( 
.A(n_481),
.Y(n_530)
);

OA21x2_ASAP7_75t_L g531 ( 
.A1(n_498),
.A2(n_499),
.B(n_466),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_491),
.Y(n_532)
);

OAI21x1_ASAP7_75t_L g533 ( 
.A1(n_466),
.A2(n_501),
.B(n_479),
.Y(n_533)
);

HB1xp67_ASAP7_75t_L g534 ( 
.A(n_491),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_477),
.Y(n_535)
);

INVx2_ASAP7_75t_SL g536 ( 
.A(n_477),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_504),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_490),
.Y(n_538)
);

INVx4_ASAP7_75t_SL g539 ( 
.A(n_496),
.Y(n_539)
);

HB1xp67_ASAP7_75t_L g540 ( 
.A(n_470),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_490),
.Y(n_541)
);

OR2x2_ASAP7_75t_L g542 ( 
.A(n_493),
.B(n_478),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_500),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_497),
.Y(n_544)
);

BUFx2_ASAP7_75t_SL g545 ( 
.A(n_470),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_516),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_518),
.B(n_487),
.Y(n_547)
);

BUFx2_ASAP7_75t_L g548 ( 
.A(n_512),
.Y(n_548)
);

OR2x2_ASAP7_75t_L g549 ( 
.A(n_542),
.B(n_468),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_518),
.B(n_495),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_525),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_525),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_527),
.Y(n_553)
);

BUFx3_ASAP7_75t_L g554 ( 
.A(n_512),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_516),
.Y(n_555)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_523),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_515),
.B(n_495),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_521),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_509),
.B(n_495),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_509),
.B(n_495),
.Y(n_560)
);

BUFx2_ASAP7_75t_L g561 ( 
.A(n_520),
.Y(n_561)
);

OAI22xp5_ASAP7_75t_L g562 ( 
.A1(n_510),
.A2(n_488),
.B1(n_496),
.B2(n_467),
.Y(n_562)
);

OR2x2_ASAP7_75t_L g563 ( 
.A(n_542),
.B(n_468),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_526),
.B(n_475),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_538),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g566 ( 
.A(n_520),
.B(n_482),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_511),
.B(n_475),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_529),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_541),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_514),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_529),
.Y(n_571)
);

BUFx2_ASAP7_75t_L g572 ( 
.A(n_522),
.Y(n_572)
);

AOI22xp33_ASAP7_75t_SL g573 ( 
.A1(n_545),
.A2(n_474),
.B1(n_482),
.B2(n_489),
.Y(n_573)
);

INVx5_ASAP7_75t_SL g574 ( 
.A(n_523),
.Y(n_574)
);

INVx3_ASAP7_75t_L g575 ( 
.A(n_537),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_523),
.Y(n_576)
);

OR2x2_ASAP7_75t_L g577 ( 
.A(n_544),
.B(n_468),
.Y(n_577)
);

BUFx3_ASAP7_75t_L g578 ( 
.A(n_522),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_543),
.Y(n_579)
);

BUFx3_ASAP7_75t_L g580 ( 
.A(n_514),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_543),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_535),
.B(n_513),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_519),
.B(n_482),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_533),
.Y(n_584)
);

AND2x4_ASAP7_75t_L g585 ( 
.A(n_575),
.B(n_539),
.Y(n_585)
);

AND2x4_ASAP7_75t_L g586 ( 
.A(n_575),
.B(n_539),
.Y(n_586)
);

OR2x2_ASAP7_75t_L g587 ( 
.A(n_548),
.B(n_530),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_565),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_565),
.Y(n_589)
);

AOI22xp33_ASAP7_75t_L g590 ( 
.A1(n_562),
.A2(n_465),
.B1(n_486),
.B2(n_545),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_568),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_550),
.B(n_532),
.Y(n_592)
);

OR2x2_ASAP7_75t_L g593 ( 
.A(n_548),
.B(n_534),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_554),
.B(n_536),
.Y(n_594)
);

AOI22xp33_ASAP7_75t_L g595 ( 
.A1(n_562),
.A2(n_486),
.B1(n_517),
.B2(n_540),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_568),
.Y(n_596)
);

AOI221xp5_ASAP7_75t_L g597 ( 
.A1(n_573),
.A2(n_485),
.B1(n_486),
.B2(n_489),
.C(n_537),
.Y(n_597)
);

BUFx3_ASAP7_75t_L g598 ( 
.A(n_578),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_569),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_569),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_546),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_571),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_546),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_555),
.Y(n_604)
);

AND2x4_ASAP7_75t_L g605 ( 
.A(n_575),
.B(n_539),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_555),
.Y(n_606)
);

HB1xp67_ASAP7_75t_L g607 ( 
.A(n_577),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_558),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_554),
.B(n_561),
.Y(n_609)
);

OR2x2_ASAP7_75t_L g610 ( 
.A(n_572),
.B(n_537),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_558),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_571),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_561),
.B(n_536),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_559),
.B(n_537),
.Y(n_614)
);

OR2x2_ASAP7_75t_L g615 ( 
.A(n_572),
.B(n_537),
.Y(n_615)
);

AOI21xp5_ASAP7_75t_SL g616 ( 
.A1(n_583),
.A2(n_528),
.B(n_508),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_560),
.B(n_524),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_579),
.Y(n_618)
);

BUFx3_ASAP7_75t_L g619 ( 
.A(n_578),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_570),
.Y(n_620)
);

NAND2x1p5_ASAP7_75t_L g621 ( 
.A(n_582),
.B(n_531),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_588),
.Y(n_622)
);

INVxp67_ASAP7_75t_SL g623 ( 
.A(n_607),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_621),
.B(n_566),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_589),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_614),
.B(n_582),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_599),
.Y(n_627)
);

BUFx2_ASAP7_75t_SL g628 ( 
.A(n_598),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_600),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_621),
.B(n_566),
.Y(n_630)
);

HB1xp67_ASAP7_75t_L g631 ( 
.A(n_607),
.Y(n_631)
);

INVx3_ASAP7_75t_L g632 ( 
.A(n_585),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_601),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_614),
.B(n_557),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_603),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_604),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_609),
.B(n_581),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_606),
.B(n_583),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_612),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_592),
.B(n_619),
.Y(n_640)
);

NAND3xp33_ASAP7_75t_L g641 ( 
.A(n_595),
.B(n_567),
.C(n_547),
.Y(n_641)
);

AND2x4_ASAP7_75t_L g642 ( 
.A(n_585),
.B(n_539),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_602),
.B(n_549),
.Y(n_643)
);

AND2x4_ASAP7_75t_SL g644 ( 
.A(n_585),
.B(n_556),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_602),
.B(n_549),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_608),
.Y(n_646)
);

OR2x2_ASAP7_75t_L g647 ( 
.A(n_587),
.B(n_563),
.Y(n_647)
);

OR2x6_ASAP7_75t_L g648 ( 
.A(n_616),
.B(n_563),
.Y(n_648)
);

HB1xp67_ASAP7_75t_L g649 ( 
.A(n_631),
.Y(n_649)
);

INVxp67_ASAP7_75t_SL g650 ( 
.A(n_631),
.Y(n_650)
);

NOR2xp67_ASAP7_75t_L g651 ( 
.A(n_632),
.B(n_620),
.Y(n_651)
);

AND2x4_ASAP7_75t_L g652 ( 
.A(n_632),
.B(n_598),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_629),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_629),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_640),
.B(n_619),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_622),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_625),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_627),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_624),
.B(n_616),
.Y(n_659)
);

NAND4xp75_ASAP7_75t_L g660 ( 
.A(n_626),
.B(n_597),
.C(n_564),
.D(n_594),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_637),
.B(n_611),
.Y(n_661)
);

OR2x2_ASAP7_75t_L g662 ( 
.A(n_647),
.B(n_593),
.Y(n_662)
);

NAND2x1p5_ASAP7_75t_L g663 ( 
.A(n_632),
.B(n_610),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_624),
.B(n_584),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_659),
.B(n_655),
.Y(n_665)
);

AOI22xp33_ASAP7_75t_L g666 ( 
.A1(n_659),
.A2(n_595),
.B1(n_641),
.B2(n_590),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_649),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_649),
.Y(n_668)
);

INVx3_ASAP7_75t_SL g669 ( 
.A(n_652),
.Y(n_669)
);

NAND4xp25_ASAP7_75t_L g670 ( 
.A(n_660),
.B(n_590),
.C(n_634),
.D(n_580),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_662),
.B(n_630),
.Y(n_671)
);

AOI22xp33_ASAP7_75t_L g672 ( 
.A1(n_652),
.A2(n_648),
.B1(n_642),
.B2(n_630),
.Y(n_672)
);

HB1xp67_ASAP7_75t_L g673 ( 
.A(n_650),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_661),
.B(n_638),
.Y(n_674)
);

OA21x2_ASAP7_75t_L g675 ( 
.A1(n_667),
.A2(n_650),
.B(n_654),
.Y(n_675)
);

AOI22xp5_ASAP7_75t_L g676 ( 
.A1(n_670),
.A2(n_642),
.B1(n_648),
.B2(n_651),
.Y(n_676)
);

OAI21xp33_ASAP7_75t_L g677 ( 
.A1(n_670),
.A2(n_656),
.B(n_658),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_669),
.B(n_652),
.Y(n_678)
);

OA21x2_ASAP7_75t_L g679 ( 
.A1(n_668),
.A2(n_673),
.B(n_653),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_671),
.Y(n_680)
);

AOI211xp5_ASAP7_75t_L g681 ( 
.A1(n_677),
.A2(n_657),
.B(n_570),
.C(n_580),
.Y(n_681)
);

AOI21xp33_ASAP7_75t_SL g682 ( 
.A1(n_676),
.A2(n_620),
.B(n_666),
.Y(n_682)
);

NAND3xp33_ASAP7_75t_L g683 ( 
.A(n_676),
.B(n_672),
.C(n_646),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_680),
.B(n_665),
.Y(n_684)
);

OAI221xp5_ASAP7_75t_SL g685 ( 
.A1(n_678),
.A2(n_648),
.B1(n_674),
.B2(n_664),
.C(n_615),
.Y(n_685)
);

NAND3x1_ASAP7_75t_L g686 ( 
.A(n_684),
.B(n_617),
.C(n_679),
.Y(n_686)
);

NAND3xp33_ASAP7_75t_L g687 ( 
.A(n_682),
.B(n_679),
.C(n_675),
.Y(n_687)
);

NOR2xp67_ASAP7_75t_SL g688 ( 
.A(n_683),
.B(n_628),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_681),
.Y(n_689)
);

NAND4xp75_ASAP7_75t_L g690 ( 
.A(n_689),
.B(n_675),
.C(n_685),
.D(n_613),
.Y(n_690)
);

NOR2x1_ASAP7_75t_L g691 ( 
.A(n_687),
.B(n_642),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_688),
.Y(n_692)
);

OAI322xp33_ASAP7_75t_L g693 ( 
.A1(n_686),
.A2(n_639),
.A3(n_633),
.B1(n_636),
.B2(n_635),
.C1(n_663),
.C2(n_623),
.Y(n_693)
);

NAND3xp33_ASAP7_75t_SL g694 ( 
.A(n_692),
.B(n_663),
.C(n_664),
.Y(n_694)
);

NAND4xp75_ASAP7_75t_L g695 ( 
.A(n_691),
.B(n_690),
.C(n_693),
.D(n_638),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_692),
.B(n_605),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_692),
.B(n_645),
.Y(n_697)
);

NOR3xp33_ASAP7_75t_L g698 ( 
.A(n_692),
.B(n_586),
.C(n_605),
.Y(n_698)
);

OAI221xp5_ASAP7_75t_L g699 ( 
.A1(n_698),
.A2(n_648),
.B1(n_618),
.B2(n_508),
.C(n_528),
.Y(n_699)
);

NOR2x1_ASAP7_75t_L g700 ( 
.A(n_695),
.B(n_524),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_697),
.Y(n_701)
);

HB1xp67_ASAP7_75t_L g702 ( 
.A(n_696),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_694),
.Y(n_703)
);

NOR2x1_ASAP7_75t_L g704 ( 
.A(n_695),
.B(n_524),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_697),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_702),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_703),
.Y(n_707)
);

AOI22xp5_ASAP7_75t_L g708 ( 
.A1(n_700),
.A2(n_605),
.B1(n_586),
.B2(n_644),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_701),
.B(n_705),
.Y(n_709)
);

NOR2x1_ASAP7_75t_SL g710 ( 
.A(n_704),
.B(n_524),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_699),
.Y(n_711)
);

AND2x4_ASAP7_75t_L g712 ( 
.A(n_706),
.B(n_586),
.Y(n_712)
);

OAI22xp33_ASAP7_75t_L g713 ( 
.A1(n_707),
.A2(n_576),
.B1(n_556),
.B2(n_524),
.Y(n_713)
);

HB1xp67_ASAP7_75t_L g714 ( 
.A(n_709),
.Y(n_714)
);

NOR3xp33_ASAP7_75t_L g715 ( 
.A(n_711),
.B(n_484),
.C(n_479),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_710),
.Y(n_716)
);

AND3x1_ASAP7_75t_L g717 ( 
.A(n_708),
.B(n_579),
.C(n_581),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_706),
.Y(n_718)
);

AOI22xp5_ASAP7_75t_L g719 ( 
.A1(n_707),
.A2(n_644),
.B1(n_645),
.B2(n_643),
.Y(n_719)
);

OA22x2_ASAP7_75t_L g720 ( 
.A1(n_707),
.A2(n_643),
.B1(n_596),
.B2(n_591),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_718),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_716),
.Y(n_722)
);

OAI22x1_ASAP7_75t_L g723 ( 
.A1(n_714),
.A2(n_551),
.B1(n_553),
.B2(n_552),
.Y(n_723)
);

AOI22xp5_ASAP7_75t_L g724 ( 
.A1(n_712),
.A2(n_576),
.B1(n_556),
.B2(n_574),
.Y(n_724)
);

INVx4_ASAP7_75t_L g725 ( 
.A(n_720),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_715),
.Y(n_726)
);

OAI22xp5_ASAP7_75t_L g727 ( 
.A1(n_719),
.A2(n_574),
.B1(n_556),
.B2(n_576),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_717),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_722),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_721),
.Y(n_730)
);

XOR2xp5_ASAP7_75t_L g731 ( 
.A(n_728),
.B(n_713),
.Y(n_731)
);

AO22x2_ASAP7_75t_L g732 ( 
.A1(n_725),
.A2(n_551),
.B1(n_553),
.B2(n_552),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_729),
.B(n_726),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_730),
.Y(n_734)
);

AOI21xp5_ASAP7_75t_L g735 ( 
.A1(n_733),
.A2(n_731),
.B(n_732),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_735),
.B(n_734),
.Y(n_736)
);

OR2x2_ASAP7_75t_L g737 ( 
.A(n_736),
.B(n_727),
.Y(n_737)
);

AOI22xp33_ASAP7_75t_SL g738 ( 
.A1(n_737),
.A2(n_723),
.B1(n_724),
.B2(n_523),
.Y(n_738)
);


endmodule