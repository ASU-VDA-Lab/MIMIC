module fake_jpeg_12873_n_387 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_387);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_387;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_13),
.B(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_8),
.B(n_10),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_7),
.B(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx4f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_1),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_10),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_6),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

BUFx10_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_5),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g131 ( 
.A(n_55),
.Y(n_131)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_56),
.Y(n_143)
);

AOI21xp33_ASAP7_75t_L g57 ( 
.A1(n_22),
.A2(n_2),
.B(n_6),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_57),
.B(n_99),
.C(n_35),
.Y(n_151)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx11_ASAP7_75t_L g176 ( 
.A(n_58),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_59),
.Y(n_172)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_60),
.Y(n_119)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_61),
.Y(n_120)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_62),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_27),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_63),
.B(n_66),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_64),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_65),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_31),
.Y(n_66)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g153 ( 
.A(n_67),
.Y(n_153)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_68),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_21),
.B(n_14),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_69),
.B(n_79),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_70),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_30),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_71),
.Y(n_129)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_19),
.Y(n_72)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_72),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_73),
.Y(n_135)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_74),
.Y(n_149)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_20),
.Y(n_75)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_75),
.Y(n_121)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_76),
.Y(n_152)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_77),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_52),
.B(n_11),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_78),
.B(n_81),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_21),
.B(n_11),
.Y(n_79)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_19),
.Y(n_80)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_80),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_39),
.B(n_11),
.Y(n_81)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_82),
.Y(n_169)
);

BUFx16f_ASAP7_75t_L g83 ( 
.A(n_19),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_83),
.B(n_84),
.Y(n_141)
);

INVx6_ASAP7_75t_SL g84 ( 
.A(n_50),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_19),
.Y(n_85)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_85),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_33),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_86),
.B(n_91),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_87),
.Y(n_160)
);

BUFx24_ASAP7_75t_L g88 ( 
.A(n_18),
.Y(n_88)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_88),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_89),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_45),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_90),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_33),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_39),
.B(n_12),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_92),
.B(n_93),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_42),
.B(n_12),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_37),
.Y(n_94)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_94),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_33),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_95),
.B(n_98),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_37),
.Y(n_96)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_96),
.Y(n_132)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_43),
.Y(n_97)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_97),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_42),
.B(n_12),
.Y(n_98)
);

AOI21xp33_ASAP7_75t_L g99 ( 
.A1(n_48),
.A2(n_40),
.B(n_23),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_48),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_100),
.B(n_104),
.Y(n_112)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_45),
.Y(n_101)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_101),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_44),
.Y(n_102)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_102),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_44),
.Y(n_103)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_103),
.Y(n_165)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_23),
.B(n_41),
.Y(n_104)
);

INVx11_ASAP7_75t_L g105 ( 
.A(n_18),
.Y(n_105)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_105),
.Y(n_167)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_45),
.Y(n_106)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_106),
.Y(n_168)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_44),
.Y(n_107)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_107),
.Y(n_147)
);

BUFx24_ASAP7_75t_L g108 ( 
.A(n_18),
.Y(n_108)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_108),
.Y(n_156)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_54),
.Y(n_109)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_109),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_49),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_110),
.B(n_111),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_24),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_104),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_114),
.B(n_118),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_78),
.B(n_24),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_115),
.B(n_126),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_59),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_65),
.A2(n_49),
.B1(n_53),
.B2(n_28),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_125),
.A2(n_138),
.B1(n_140),
.B2(n_159),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_80),
.B(n_40),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_101),
.B(n_41),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_133),
.B(n_144),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_88),
.A2(n_53),
.B1(n_28),
.B2(n_49),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_134),
.A2(n_173),
.B(n_175),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_88),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_136),
.B(n_139),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_110),
.A2(n_25),
.B1(n_26),
.B2(n_32),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_108),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_70),
.A2(n_25),
.B1(n_26),
.B2(n_32),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_107),
.B(n_35),
.Y(n_144)
);

NOR2x1_ASAP7_75t_L g203 ( 
.A(n_151),
.B(n_25),
.Y(n_203)
);

AO22x1_ASAP7_75t_SL g159 ( 
.A1(n_108),
.A2(n_38),
.B1(n_46),
.B2(n_47),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_67),
.B(n_51),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_161),
.B(n_135),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_85),
.A2(n_38),
.B1(n_46),
.B2(n_47),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_163),
.B(n_83),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_105),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_171),
.B(n_167),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_76),
.A2(n_97),
.B1(n_56),
.B2(n_64),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_56),
.A2(n_89),
.B1(n_97),
.B2(n_64),
.Y(n_175)
);

OR2x2_ASAP7_75t_L g177 ( 
.A(n_112),
.B(n_51),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_177),
.B(n_210),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_128),
.A2(n_90),
.B1(n_87),
.B2(n_89),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_178),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_146),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_179),
.B(n_186),
.Y(n_240)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_165),
.Y(n_180)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_180),
.Y(n_233)
);

NOR2x1_ASAP7_75t_L g261 ( 
.A(n_181),
.B(n_208),
.Y(n_261)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_128),
.Y(n_182)
);

BUFx2_ASAP7_75t_L g242 ( 
.A(n_182),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_125),
.A2(n_103),
.B1(n_71),
.B2(n_73),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_183),
.A2(n_185),
.B1(n_228),
.B2(n_223),
.Y(n_248)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_119),
.Y(n_184)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_184),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_113),
.A2(n_94),
.B1(n_96),
.B2(n_102),
.Y(n_185)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_141),
.Y(n_186)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_137),
.Y(n_187)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_187),
.Y(n_245)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_120),
.Y(n_188)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_188),
.Y(n_247)
);

INVx8_ASAP7_75t_L g189 ( 
.A(n_152),
.Y(n_189)
);

INVx3_ASAP7_75t_SL g251 ( 
.A(n_189),
.Y(n_251)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_121),
.Y(n_190)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_190),
.Y(n_255)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_137),
.Y(n_191)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_191),
.Y(n_258)
);

BUFx12f_ASAP7_75t_L g192 ( 
.A(n_143),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_192),
.B(n_193),
.Y(n_241)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_142),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_159),
.A2(n_172),
.B1(n_130),
.B2(n_149),
.Y(n_194)
);

OA22x2_ASAP7_75t_L g270 ( 
.A1(n_194),
.A2(n_207),
.B1(n_108),
.B2(n_88),
.Y(n_270)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_155),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_195),
.B(n_201),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_156),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_196),
.Y(n_257)
);

INVx6_ASAP7_75t_SL g198 ( 
.A(n_148),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_198),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_158),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_SL g269 ( 
.A(n_203),
.B(n_151),
.C(n_78),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_127),
.B(n_150),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_204),
.B(n_211),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_157),
.B(n_122),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_205),
.B(n_206),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_168),
.B(n_147),
.Y(n_206)
);

NAND2x1p5_ASAP7_75t_L g207 ( 
.A(n_148),
.B(n_169),
.Y(n_207)
);

A2O1A1Ixp33_ASAP7_75t_L g208 ( 
.A1(n_117),
.A2(n_134),
.B(n_175),
.C(n_173),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_166),
.B(n_145),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_153),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_212),
.B(n_213),
.Y(n_246)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_153),
.Y(n_213)
);

OAI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_116),
.A2(n_123),
.B1(n_135),
.B2(n_129),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_214),
.A2(n_227),
.B1(n_228),
.B2(n_185),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_162),
.B(n_152),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_215),
.B(n_226),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_176),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_216),
.B(n_217),
.Y(n_250)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_124),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_160),
.B(n_170),
.C(n_164),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_218),
.B(n_221),
.C(n_228),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_143),
.A2(n_154),
.B1(n_170),
.B2(n_160),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_219),
.A2(n_183),
.B1(n_222),
.B2(n_208),
.Y(n_235)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_124),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_220),
.B(n_222),
.Y(n_265)
);

MAJx2_ASAP7_75t_L g221 ( 
.A(n_154),
.B(n_131),
.C(n_164),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_131),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_132),
.B(n_174),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_223),
.B(n_230),
.Y(n_238)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_132),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_224),
.B(n_229),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_174),
.B(n_131),
.Y(n_226)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_116),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_123),
.B(n_129),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_146),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_197),
.A2(n_225),
.B1(n_200),
.B2(n_202),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_234),
.A2(n_259),
.B1(n_266),
.B2(n_267),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_235),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_239),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_248),
.B(n_270),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_206),
.B(n_205),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_252),
.B(n_253),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_209),
.B(n_181),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_203),
.B(n_196),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_254),
.B(n_264),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_197),
.A2(n_218),
.B1(n_177),
.B2(n_188),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_180),
.A2(n_207),
.B1(n_189),
.B2(n_195),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_263),
.A2(n_239),
.B1(n_248),
.B2(n_257),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_207),
.B(n_199),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_221),
.A2(n_191),
.B1(n_187),
.B2(n_198),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_216),
.A2(n_194),
.B1(n_197),
.B2(n_225),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_182),
.B(n_192),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_268),
.B(n_262),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_269),
.A2(n_253),
.B(n_261),
.Y(n_273)
);

AND2x6_ASAP7_75t_L g271 ( 
.A(n_269),
.B(n_192),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_271),
.B(n_279),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_232),
.B(n_252),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_272),
.B(n_287),
.C(n_245),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_273),
.Y(n_304)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_247),
.Y(n_274)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_274),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_231),
.B(n_260),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_275),
.Y(n_320)
);

NAND2x1_ASAP7_75t_SL g276 ( 
.A(n_256),
.B(n_264),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_276),
.A2(n_266),
.B(n_267),
.Y(n_301)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_247),
.Y(n_277)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_277),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_246),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_278),
.Y(n_315)
);

AND2x6_ASAP7_75t_L g279 ( 
.A(n_254),
.B(n_261),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_236),
.Y(n_280)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_280),
.Y(n_313)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_236),
.Y(n_281)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_281),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_240),
.B(n_232),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_282),
.B(n_289),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_268),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_285),
.Y(n_322)
);

MAJx2_ASAP7_75t_L g287 ( 
.A(n_238),
.B(n_256),
.C(n_234),
.Y(n_287)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_255),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_241),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_291),
.B(n_292),
.Y(n_309)
);

NOR3xp33_ASAP7_75t_SL g292 ( 
.A(n_237),
.B(n_238),
.C(n_243),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_293),
.B(n_294),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_244),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_233),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_295),
.B(n_296),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_255),
.B(n_265),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_259),
.B(n_250),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_297),
.B(n_300),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_299),
.A2(n_251),
.B1(n_258),
.B2(n_245),
.Y(n_316)
);

INVx13_ASAP7_75t_L g300 ( 
.A(n_242),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_301),
.Y(n_338)
);

NOR2x1_ASAP7_75t_L g303 ( 
.A(n_288),
.B(n_263),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_303),
.B(n_314),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_272),
.B(n_270),
.Y(n_306)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_306),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_290),
.A2(n_249),
.B1(n_270),
.B2(n_251),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_307),
.A2(n_298),
.B1(n_299),
.B2(n_284),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_286),
.A2(n_249),
.B(n_270),
.Y(n_308)
);

AOI211xp5_ASAP7_75t_L g329 ( 
.A1(n_308),
.A2(n_286),
.B(n_298),
.C(n_288),
.Y(n_329)
);

NOR2x1_ASAP7_75t_L g314 ( 
.A(n_288),
.B(n_258),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_316),
.A2(n_293),
.B1(n_289),
.B2(n_281),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_321),
.B(n_284),
.Y(n_326)
);

NAND3xp33_ASAP7_75t_L g323 ( 
.A(n_309),
.B(n_273),
.C(n_283),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_323),
.B(n_324),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_315),
.B(n_283),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_325),
.B(n_328),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_326),
.B(n_337),
.C(n_321),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_320),
.B(n_292),
.Y(n_328)
);

OA21x2_ASAP7_75t_L g348 ( 
.A1(n_329),
.A2(n_306),
.B(n_307),
.Y(n_348)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_313),
.Y(n_330)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_330),
.Y(n_342)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_313),
.Y(n_331)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_331),
.Y(n_344)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_317),
.Y(n_332)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_332),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_310),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_333),
.B(n_336),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_335),
.A2(n_339),
.B1(n_301),
.B2(n_308),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_315),
.B(n_280),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_321),
.B(n_287),
.C(n_276),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_307),
.A2(n_290),
.B1(n_276),
.B2(n_271),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_340),
.B(n_346),
.C(n_351),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_341),
.A2(n_329),
.B1(n_327),
.B2(n_308),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_337),
.B(n_304),
.C(n_306),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_SL g347 ( 
.A(n_326),
.B(n_327),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_347),
.B(n_349),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_SL g357 ( 
.A1(n_348),
.A2(n_303),
.B(n_314),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_339),
.B(n_302),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_335),
.B(n_301),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_343),
.B(n_310),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_L g364 ( 
.A1(n_353),
.A2(n_355),
.B(n_305),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_352),
.A2(n_338),
.B1(n_334),
.B2(n_302),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_354),
.A2(n_341),
.B1(n_309),
.B2(n_348),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_345),
.B(n_322),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_351),
.A2(n_338),
.B(n_314),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_SL g369 ( 
.A1(n_356),
.A2(n_361),
.B(n_319),
.Y(n_369)
);

NAND3xp33_ASAP7_75t_SL g370 ( 
.A(n_357),
.B(n_279),
.C(n_316),
.Y(n_370)
);

INVx11_ASAP7_75t_L g359 ( 
.A(n_342),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_359),
.B(n_360),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_349),
.A2(n_303),
.B(n_322),
.Y(n_361)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_364),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_358),
.B(n_340),
.C(n_346),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_365),
.B(n_367),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_L g374 ( 
.A1(n_366),
.A2(n_370),
.B(n_361),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_354),
.A2(n_319),
.B1(n_348),
.B2(n_305),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_353),
.B(n_355),
.Y(n_368)
);

OAI21x1_ASAP7_75t_L g376 ( 
.A1(n_368),
.A2(n_318),
.B(n_356),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_369),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_374),
.B(n_376),
.Y(n_377)
);

AOI322xp5_ASAP7_75t_L g375 ( 
.A1(n_363),
.A2(n_357),
.A3(n_359),
.B1(n_360),
.B2(n_350),
.C1(n_344),
.C2(n_330),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_375),
.B(n_318),
.Y(n_380)
);

OR2x6_ASAP7_75t_L g378 ( 
.A(n_373),
.B(n_362),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_378),
.A2(n_379),
.B1(n_380),
.B2(n_371),
.Y(n_381)
);

HB1xp67_ASAP7_75t_L g379 ( 
.A(n_372),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_SL g385 ( 
.A1(n_381),
.A2(n_382),
.B(n_383),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_SL g382 ( 
.A(n_377),
.B(n_372),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_379),
.B(n_365),
.C(n_358),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_383),
.A2(n_370),
.B1(n_316),
.B2(n_331),
.Y(n_384)
);

AOI322xp5_ASAP7_75t_L g386 ( 
.A1(n_384),
.A2(n_332),
.A3(n_347),
.B1(n_362),
.B2(n_317),
.C1(n_312),
.C2(n_311),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_386),
.B(n_385),
.Y(n_387)
);


endmodule