module real_jpeg_4669_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_470;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_475;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

AND2x2_ASAP7_75t_SL g55 ( 
.A(n_0),
.B(n_56),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_0),
.B(n_102),
.Y(n_101)
);

AND2x2_ASAP7_75t_SL g132 ( 
.A(n_0),
.B(n_133),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_0),
.B(n_146),
.Y(n_145)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

AND2x2_ASAP7_75t_SL g139 ( 
.A(n_2),
.B(n_39),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_2),
.B(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_2),
.B(n_229),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_2),
.B(n_256),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_2),
.B(n_282),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_2),
.B(n_369),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_2),
.B(n_374),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_2),
.B(n_403),
.Y(n_402)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_3),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_3),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_3),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_4),
.B(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_4),
.B(n_87),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_4),
.B(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_4),
.B(n_173),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g214 ( 
.A(n_4),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_4),
.B(n_240),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_4),
.B(n_27),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_4),
.B(n_337),
.Y(n_336)
);

AND2x2_ASAP7_75t_SL g30 ( 
.A(n_5),
.B(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_5),
.B(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_5),
.B(n_70),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_5),
.B(n_85),
.Y(n_84)
);

AND2x2_ASAP7_75t_SL g120 ( 
.A(n_5),
.B(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_5),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_5),
.B(n_189),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_5),
.B(n_201),
.Y(n_200)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_7),
.B(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_7),
.B(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_7),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_7),
.B(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_7),
.B(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_7),
.B(n_209),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_7),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_7),
.B(n_267),
.Y(n_266)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_8),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_8),
.Y(n_437)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_9),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_9),
.Y(n_89)
);

BUFx5_ASAP7_75t_L g146 ( 
.A(n_9),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_9),
.Y(n_221)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_10),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_11),
.B(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_11),
.B(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_11),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_11),
.B(n_269),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_11),
.B(n_385),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_11),
.B(n_398),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_11),
.B(n_428),
.Y(n_427)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_12),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_12),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_12),
.Y(n_204)
);

BUFx5_ASAP7_75t_L g269 ( 
.A(n_12),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_13),
.B(n_194),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_13),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_13),
.B(n_298),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_13),
.B(n_229),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_13),
.B(n_411),
.Y(n_410)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_14),
.Y(n_138)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_14),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_14),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_15),
.B(n_204),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_15),
.B(n_61),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_15),
.B(n_243),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_15),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_15),
.B(n_417),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_15),
.B(n_422),
.Y(n_421)
);

XNOR2x2_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_158),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_157),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_94),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_20),
.B(n_94),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_76),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_45),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_38),
.C(n_40),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_23),
.B(n_78),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_30),
.C(n_33),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_24),
.B(n_49),
.C(n_68),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_24),
.A2(n_49),
.B1(n_50),
.B2(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_24),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_24),
.A2(n_93),
.B1(n_150),
.B2(n_151),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_24),
.A2(n_93),
.B1(n_168),
.B2(n_171),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_24),
.B(n_168),
.C(n_172),
.Y(n_257)
);

OR2x2_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_26),
.Y(n_24)
);

OR2x2_ASAP7_75t_SL g34 ( 
.A(n_25),
.B(n_35),
.Y(n_34)
);

OR2x2_ASAP7_75t_SL g50 ( 
.A(n_25),
.B(n_51),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_25),
.B(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_28),
.B(n_218),
.Y(n_301)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx11_ASAP7_75t_L g114 ( 
.A(n_29),
.Y(n_114)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_29),
.Y(n_380)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_29),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_30),
.A2(n_33),
.B1(n_34),
.B2(n_152),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_30),
.Y(n_152)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_31),
.Y(n_226)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_33),
.A2(n_34),
.B1(n_98),
.B2(n_99),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_33),
.A2(n_34),
.B1(n_181),
.B2(n_294),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_34),
.B(n_101),
.C(n_105),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_34),
.B(n_179),
.C(n_181),
.Y(n_178)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_37),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_38),
.A2(n_40),
.B1(n_41),
.B2(n_79),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_38),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_44),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_64),
.B1(n_65),
.B2(n_75),
.Y(n_45)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_47),
.A2(n_48),
.B1(n_60),
.B2(n_63),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_50),
.B1(n_55),
.B2(n_59),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_49),
.A2(n_50),
.B1(n_197),
.B2(n_198),
.Y(n_196)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_50),
.B(n_199),
.C(n_203),
.Y(n_284)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_54),
.Y(n_119)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_54),
.Y(n_185)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_54),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_55),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_55),
.B(n_265),
.Y(n_264)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_57),
.Y(n_170)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_58),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_58),
.Y(n_244)
);

BUFx5_ASAP7_75t_L g300 ( 
.A(n_58),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_59),
.B(n_266),
.C(n_268),
.Y(n_320)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_60),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_60),
.A2(n_63),
.B1(n_116),
.B2(n_125),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_60),
.B(n_117),
.C(n_124),
.Y(n_153)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_62),
.Y(n_282)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_66),
.A2(n_67),
.B1(n_72),
.B2(n_73),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_68),
.A2(n_69),
.B1(n_91),
.B2(n_92),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_68),
.B(n_101),
.C(n_110),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_68),
.A2(n_69),
.B1(n_110),
.B2(n_111),
.Y(n_323)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_69),
.Y(n_68)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_80),
.C(n_90),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_77),
.B(n_156),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_80),
.B(n_90),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_83),
.C(n_86),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_81),
.A2(n_83),
.B1(n_84),
.B2(n_128),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_81),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_83),
.A2(n_84),
.B1(n_271),
.B2(n_272),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_84),
.B(n_132),
.C(n_188),
.Y(n_340)
);

INVx6_ASAP7_75t_L g230 ( 
.A(n_85),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_86),
.B(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_147),
.C(n_155),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_95),
.B(n_485),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_126),
.C(n_129),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_SL g478 ( 
.A(n_96),
.B(n_479),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_109),
.C(n_115),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_97),
.B(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_101),
.B1(n_105),
.B2(n_108),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_100),
.A2(n_101),
.B1(n_322),
.B2(n_323),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_101),
.B(n_200),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_101),
.B(n_200),
.Y(n_375)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_104),
.Y(n_400)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_105),
.Y(n_108)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_109),
.B(n_115),
.Y(n_349)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_114),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_114),
.Y(n_180)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_116),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_120),
.B1(n_123),
.B2(n_124),
.Y(n_116)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_117),
.Y(n_123)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_120),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_120),
.B(n_255),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_120),
.B(n_249),
.C(n_255),
.Y(n_263)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_126),
.B(n_129),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_140),
.C(n_144),
.Y(n_129)
);

AO22x1_ASAP7_75t_SL g356 ( 
.A1(n_130),
.A2(n_131),
.B1(n_357),
.B2(n_358),
.Y(n_356)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_135),
.C(n_139),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_132),
.A2(n_188),
.B1(n_273),
.B2(n_274),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_132),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_132),
.A2(n_139),
.B1(n_273),
.B2(n_326),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_132),
.B(n_367),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_132),
.A2(n_273),
.B1(n_367),
.B2(n_368),
.Y(n_404)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_134),
.Y(n_201)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_134),
.Y(n_211)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_134),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_134),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_135),
.A2(n_228),
.B1(n_231),
.B2(n_232),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_135),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_135),
.B(n_224),
.C(n_228),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_135),
.A2(n_231),
.B1(n_325),
.B2(n_327),
.Y(n_324)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_137),
.Y(n_135)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_137),
.Y(n_267)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_137),
.Y(n_374)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_138),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_139),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_140),
.A2(n_141),
.B1(n_144),
.B2(n_145),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g334 ( 
.A1(n_144),
.A2(n_145),
.B1(n_335),
.B2(n_336),
.Y(n_334)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_145),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_145),
.B(n_336),
.C(n_340),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_147),
.B(n_155),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_153),
.C(n_154),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_148),
.A2(n_149),
.B1(n_481),
.B2(n_482),
.Y(n_480)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_153),
.B(n_154),
.Y(n_482)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_475),
.B(n_489),
.Y(n_158)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_359),
.Y(n_159)
);

O2A1O1Ixp33_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_314),
.B(n_342),
.C(n_343),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_285),
.B(n_313),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_162),
.B(n_473),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_258),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_163),
.B(n_258),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_222),
.C(n_245),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_164),
.B(n_312),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_195),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_165),
.B(n_196),
.C(n_205),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_178),
.C(n_186),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_166),
.B(n_309),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_172),
.Y(n_166)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_168),
.Y(n_171)
);

BUFx12f_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

BUFx8_ASAP7_75t_L g371 ( 
.A(n_177),
.Y(n_371)
);

BUFx5_ASAP7_75t_L g434 ( 
.A(n_177),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_178),
.A2(n_186),
.B1(n_187),
.B2(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_178),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_SL g292 ( 
.A(n_179),
.B(n_293),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_181),
.Y(n_294)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx5_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx4_ASAP7_75t_L g306 ( 
.A(n_185),
.Y(n_306)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_192),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_188),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_188),
.A2(n_192),
.B1(n_193),
.B2(n_274),
.Y(n_307)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_191),
.Y(n_253)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_191),
.Y(n_425)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_205),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_199),
.A2(n_200),
.B1(n_202),
.B2(n_203),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_200),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_203),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_212),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_206),
.A2(n_207),
.B(n_208),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_206),
.B(n_213),
.C(n_217),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_210),
.Y(n_240)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_217),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

INVx8_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_222),
.B(n_245),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_233),
.C(n_235),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_223),
.A2(n_233),
.B1(n_234),
.B2(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_223),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_227),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_225),
.B(n_433),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_225),
.B(n_440),
.Y(n_439)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_228),
.Y(n_232)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g288 ( 
.A(n_235),
.B(n_289),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_238),
.C(n_241),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_236),
.A2(n_237),
.B1(n_462),
.B2(n_463),
.Y(n_461)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_238),
.A2(n_239),
.B1(n_241),
.B2(n_242),
.Y(n_463)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_244),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_257),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_247),
.B(n_248),
.C(n_257),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_249),
.B(n_254),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_259),
.B(n_261),
.C(n_275),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_275),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_270),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_263),
.B(n_264),
.C(n_270),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_268),
.Y(n_265)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_276),
.B(n_278),
.C(n_279),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_284),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_283),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_281),
.B(n_283),
.C(n_332),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_284),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_311),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_286),
.B(n_311),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_291),
.C(n_308),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_287),
.A2(n_288),
.B1(n_467),
.B2(n_468),
.Y(n_466)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_SL g467 ( 
.A(n_291),
.B(n_308),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_295),
.C(n_307),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_SL g456 ( 
.A(n_292),
.B(n_457),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_295),
.B(n_307),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_301),
.C(n_302),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_296),
.A2(n_297),
.B1(n_302),
.B2(n_390),
.Y(n_389)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

BUFx2_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx6_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_301),
.B(n_389),
.Y(n_388)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_302),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_304),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_303),
.B(n_379),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_303),
.B(n_436),
.Y(n_435)
);

INVx4_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx8_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_315),
.B(n_344),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

OR2x2_ASAP7_75t_L g342 ( 
.A(n_316),
.B(n_317),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_317),
.B(n_345),
.Y(n_344)
);

OR2x2_ASAP7_75t_L g474 ( 
.A(n_317),
.B(n_345),
.Y(n_474)
);

FAx1_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_328),
.CI(n_341),
.CON(n_317),
.SN(n_317)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_324),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_321),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_320),
.B(n_321),
.C(n_324),
.Y(n_352)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_325),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_SL g328 ( 
.A(n_329),
.B(n_330),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_329),
.B(n_331),
.C(n_333),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_333),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_340),
.Y(n_333)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_347),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_346),
.B(n_348),
.C(n_350),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_350),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_351),
.A2(n_352),
.B1(n_353),
.B2(n_354),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_351),
.B(n_355),
.C(n_356),
.Y(n_483)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_356),
.Y(n_354)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

OAI31xp33_ASAP7_75t_L g359 ( 
.A1(n_360),
.A2(n_471),
.A3(n_472),
.B(n_474),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_361),
.A2(n_465),
.B(n_470),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_SL g361 ( 
.A1(n_362),
.A2(n_452),
.B(n_464),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_L g362 ( 
.A1(n_363),
.A2(n_405),
.B(n_451),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_364),
.B(n_391),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_364),
.B(n_391),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_376),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_365),
.B(n_377),
.C(n_388),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_SL g365 ( 
.A(n_366),
.B(n_372),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_366),
.B(n_373),
.C(n_375),
.Y(n_460)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx8_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_375),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_388),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_381),
.C(n_383),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_SL g392 ( 
.A(n_378),
.B(n_393),
.Y(n_392)
);

INVx4_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_381),
.A2(n_382),
.B1(n_383),
.B2(n_384),
.Y(n_393)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx8_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

BUFx5_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_394),
.C(n_404),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_392),
.B(n_448),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_394),
.A2(n_395),
.B1(n_404),
.B2(n_449),
.Y(n_448)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_401),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_396),
.A2(n_397),
.B1(n_401),
.B2(n_402),
.Y(n_418)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx5_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_404),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_L g405 ( 
.A1(n_406),
.A2(n_445),
.B(n_450),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_L g406 ( 
.A1(n_407),
.A2(n_430),
.B(n_444),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_408),
.B(n_419),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_408),
.B(n_419),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_418),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_416),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_410),
.B(n_416),
.C(n_418),
.Y(n_446)
);

INVx3_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx5_ASAP7_75t_SL g412 ( 
.A(n_413),
.Y(n_412)
);

INVx4_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx4_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_420),
.B(n_426),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g442 ( 
.A1(n_420),
.A2(n_421),
.B1(n_426),
.B2(n_427),
.Y(n_442)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx6_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

INVx8_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_L g430 ( 
.A1(n_431),
.A2(n_438),
.B(n_443),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_435),
.Y(n_431)
);

INVx3_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx4_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_439),
.B(n_442),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_439),
.B(n_442),
.Y(n_443)
);

INVx4_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_447),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_446),
.B(n_447),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_454),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_453),
.B(n_454),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_455),
.A2(n_456),
.B1(n_458),
.B2(n_459),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_455),
.B(n_460),
.C(n_461),
.Y(n_469)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_460),
.B(n_461),
.Y(n_459)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_466),
.B(n_469),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_466),
.B(n_469),
.Y(n_470)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_467),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_486),
.Y(n_475)
);

OAI21xp33_ASAP7_75t_L g489 ( 
.A1(n_476),
.A2(n_490),
.B(n_491),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_477),
.B(n_484),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_477),
.B(n_484),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_478),
.B(n_480),
.C(n_483),
.Y(n_477)
);

FAx1_ASAP7_75t_SL g488 ( 
.A(n_478),
.B(n_480),
.CI(n_483),
.CON(n_488),
.SN(n_488)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_487),
.B(n_488),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_487),
.B(n_488),
.Y(n_490)
);

BUFx24_ASAP7_75t_SL g493 ( 
.A(n_488),
.Y(n_493)
);


endmodule