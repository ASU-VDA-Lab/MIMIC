module fake_jpeg_6634_n_340 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_340);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_340;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx13_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx11_ASAP7_75t_SL g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_35),
.B(n_36),
.Y(n_61)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_31),
.A2(n_15),
.B1(n_14),
.B2(n_12),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_37),
.A2(n_21),
.B1(n_28),
.B2(n_31),
.Y(n_62)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_25),
.B(n_0),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_21),
.Y(n_50)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_42),
.B(n_17),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_48),
.Y(n_75)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_50),
.B(n_62),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_23),
.C(n_29),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_51),
.B(n_17),
.Y(n_82)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_52),
.B(n_53),
.Y(n_80)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_43),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_55),
.Y(n_88)
);

NOR3xp33_ASAP7_75t_SL g57 ( 
.A(n_43),
.B(n_21),
.C(n_30),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_57),
.B(n_58),
.Y(n_97)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_59),
.Y(n_94)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_60),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_38),
.A2(n_30),
.B1(n_16),
.B2(n_31),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_63),
.A2(n_31),
.B1(n_30),
.B2(n_16),
.Y(n_77)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_66),
.Y(n_84)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_67),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_40),
.B(n_25),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_69),
.B(n_17),
.Y(n_91)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_70),
.Y(n_93)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_71),
.Y(n_95)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_77),
.A2(n_68),
.B1(n_65),
.B2(n_64),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_57),
.B(n_25),
.Y(n_78)
);

FAx1_ASAP7_75t_SL g106 ( 
.A(n_78),
.B(n_51),
.CI(n_69),
.CON(n_106),
.SN(n_106)
);

INVx2_ASAP7_75t_SL g79 ( 
.A(n_56),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_79),
.B(n_82),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_86),
.Y(n_105)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_89),
.B(n_90),
.Y(n_109)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_48),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_91),
.B(n_50),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_61),
.A2(n_16),
.B(n_32),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_96),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_81),
.A2(n_97),
.B1(n_80),
.B2(n_77),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_99),
.A2(n_100),
.B1(n_123),
.B2(n_117),
.Y(n_141)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_76),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_101),
.B(n_102),
.Y(n_134)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_76),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_103),
.B(n_106),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_91),
.Y(n_127)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_75),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_108),
.B(n_110),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_76),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_81),
.B(n_50),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_111),
.B(n_24),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_69),
.Y(n_112)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_112),
.Y(n_130)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_75),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_113),
.B(n_114),
.Y(n_144)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_85),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_87),
.B(n_58),
.Y(n_115)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_115),
.Y(n_137)
);

MAJx2_ASAP7_75t_L g116 ( 
.A(n_82),
.B(n_43),
.C(n_67),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_116),
.B(n_92),
.C(n_84),
.Y(n_145)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_80),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_117),
.B(n_119),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_96),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_79),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_120),
.B(n_121),
.Y(n_151)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_90),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_97),
.Y(n_122)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_122),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_81),
.A2(n_66),
.B1(n_35),
.B2(n_72),
.Y(n_123)
);

AOI22x1_ASAP7_75t_SL g124 ( 
.A1(n_91),
.A2(n_35),
.B1(n_44),
.B2(n_43),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_124),
.A2(n_68),
.B1(n_65),
.B2(n_73),
.Y(n_136)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_79),
.Y(n_125)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_125),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_127),
.B(n_128),
.Y(n_181)
);

OAI32xp33_ASAP7_75t_L g128 ( 
.A1(n_111),
.A2(n_91),
.A3(n_87),
.B1(n_78),
.B2(n_84),
.Y(n_128)
);

NOR2x1_ASAP7_75t_R g131 ( 
.A(n_124),
.B(n_116),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_131),
.A2(n_33),
.B(n_19),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_104),
.B(n_78),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_132),
.B(n_140),
.Y(n_172)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_101),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_133),
.B(n_141),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_136),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_118),
.A2(n_88),
.B1(n_59),
.B2(n_52),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_138),
.A2(n_146),
.B1(n_125),
.B2(n_120),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_99),
.B(n_73),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_108),
.A2(n_89),
.B1(n_86),
.B2(n_90),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_142),
.B(n_148),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_113),
.A2(n_83),
.B1(n_19),
.B2(n_26),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_143),
.A2(n_149),
.B1(n_154),
.B2(n_121),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_145),
.B(n_93),
.C(n_98),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_118),
.A2(n_92),
.B1(n_94),
.B2(n_26),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_147),
.B(n_18),
.Y(n_156)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_109),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_123),
.A2(n_119),
.B1(n_122),
.B2(n_106),
.Y(n_149)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_105),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_152),
.B(n_153),
.Y(n_177)
);

BUFx2_ASAP7_75t_L g153 ( 
.A(n_103),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_106),
.A2(n_26),
.B1(n_94),
.B2(n_95),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_155),
.A2(n_129),
.B1(n_133),
.B2(n_102),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_156),
.B(n_161),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_158),
.A2(n_159),
.B1(n_180),
.B2(n_126),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_140),
.B(n_95),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_131),
.A2(n_29),
.B(n_23),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_160),
.B(n_183),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_147),
.B(n_93),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_139),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_162),
.B(n_163),
.Y(n_199)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_151),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_144),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_164),
.B(n_167),
.Y(n_202)
);

XNOR2x1_ASAP7_75t_L g165 ( 
.A(n_145),
.B(n_114),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_165),
.B(n_173),
.C(n_136),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_134),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_166),
.Y(n_190)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_146),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_138),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_168),
.B(n_170),
.Y(n_185)
);

OA21x2_ASAP7_75t_L g170 ( 
.A1(n_150),
.A2(n_44),
.B(n_83),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_141),
.A2(n_98),
.B1(n_29),
.B2(n_23),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_174),
.A2(n_179),
.B1(n_137),
.B2(n_167),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_137),
.B(n_28),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_175),
.B(n_176),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_135),
.Y(n_176)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_154),
.Y(n_178)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_178),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_149),
.A2(n_28),
.B1(n_47),
.B2(n_49),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_126),
.A2(n_47),
.B1(n_49),
.B2(n_83),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_182),
.B(n_130),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_128),
.A2(n_18),
.B(n_19),
.Y(n_183)
);

NAND3xp33_ASAP7_75t_L g184 ( 
.A(n_165),
.B(n_127),
.C(n_132),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_184),
.B(n_187),
.Y(n_227)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_177),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_191),
.A2(n_27),
.B1(n_22),
.B2(n_18),
.Y(n_230)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_161),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_192),
.B(n_198),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_193),
.B(n_194),
.C(n_200),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_171),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_196),
.B(n_203),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_166),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_197),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_172),
.B(n_173),
.C(n_182),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_172),
.B(n_130),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_201),
.B(n_204),
.C(n_208),
.Y(n_229)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_155),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_181),
.B(n_152),
.C(n_148),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_205),
.A2(n_197),
.B1(n_190),
.B2(n_208),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_180),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_206),
.B(n_210),
.Y(n_232)
);

A2O1A1Ixp33_ASAP7_75t_L g207 ( 
.A1(n_181),
.A2(n_33),
.B(n_17),
.C(n_18),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_207),
.B(n_160),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_178),
.B(n_129),
.C(n_153),
.Y(n_208)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_163),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_209),
.A2(n_170),
.B1(n_22),
.B2(n_27),
.Y(n_223)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_174),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_164),
.B(n_110),
.Y(n_211)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_211),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_203),
.A2(n_169),
.B1(n_168),
.B2(n_176),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_212),
.A2(n_216),
.B1(n_221),
.B2(n_196),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_213),
.A2(n_218),
.B(n_234),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_214),
.A2(n_207),
.B1(n_189),
.B2(n_210),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_209),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_215),
.B(n_226),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_186),
.A2(n_157),
.B1(n_158),
.B2(n_183),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_200),
.B(n_159),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_217),
.B(n_222),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_186),
.A2(n_169),
.B(n_159),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_192),
.A2(n_179),
.B1(n_156),
.B2(n_162),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_201),
.B(n_170),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_223),
.Y(n_255)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_195),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_224),
.B(n_228),
.Y(n_239)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_188),
.Y(n_226)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_195),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_230),
.A2(n_235),
.B1(n_27),
.B2(n_18),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_191),
.A2(n_18),
.B(n_1),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_185),
.A2(n_27),
.B1(n_18),
.B2(n_33),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_189),
.B(n_204),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_236),
.B(n_2),
.Y(n_259)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_199),
.Y(n_237)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_237),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_225),
.B(n_193),
.C(n_194),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_240),
.B(n_252),
.C(n_257),
.Y(n_265)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_242),
.Y(n_267)
);

XNOR2x2_ASAP7_75t_L g243 ( 
.A(n_218),
.B(n_202),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_243),
.A2(n_247),
.B(n_248),
.Y(n_270)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_244),
.Y(n_272)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_214),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_245),
.B(n_250),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_213),
.A2(n_198),
.B(n_187),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_219),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_233),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_249),
.B(n_253),
.Y(n_271)
);

INVxp33_ASAP7_75t_L g250 ( 
.A(n_235),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_251),
.A2(n_260),
.B1(n_224),
.B2(n_234),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_225),
.B(n_33),
.C(n_32),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_232),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_236),
.B(n_33),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_256),
.B(n_259),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_229),
.B(n_0),
.C(n_1),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_237),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_258),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_216),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_238),
.B(n_217),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_261),
.B(n_264),
.Y(n_294)
);

AOI322xp5_ASAP7_75t_SL g263 ( 
.A1(n_243),
.A2(n_227),
.A3(n_229),
.B1(n_222),
.B2(n_220),
.C1(n_212),
.C2(n_221),
.Y(n_263)
);

NAND2xp33_ASAP7_75t_SL g282 ( 
.A(n_263),
.B(n_246),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_238),
.B(n_231),
.Y(n_264)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_266),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_256),
.B(n_14),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_268),
.B(n_269),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_240),
.B(n_14),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_247),
.B(n_12),
.Y(n_273)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_273),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_259),
.B(n_2),
.C(n_4),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_274),
.B(n_275),
.C(n_276),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_246),
.B(n_12),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_252),
.B(n_2),
.C(n_5),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_245),
.A2(n_11),
.B1(n_6),
.B2(n_7),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_277),
.A2(n_255),
.B1(n_241),
.B2(n_244),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_278),
.B(n_239),
.Y(n_281)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_281),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_282),
.A2(n_283),
.B(n_290),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_271),
.Y(n_283)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_284),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_264),
.B(n_239),
.C(n_257),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_286),
.B(n_295),
.C(n_274),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_279),
.A2(n_255),
.B1(n_258),
.B2(n_250),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_287),
.B(n_293),
.C(n_6),
.Y(n_307)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_278),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_270),
.B(n_254),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_291),
.B(n_285),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_272),
.A2(n_251),
.B(n_6),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_292),
.A2(n_291),
.B(n_280),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_267),
.A2(n_275),
.B(n_265),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_265),
.B(n_5),
.C(n_6),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_296),
.A2(n_298),
.B(n_299),
.Y(n_314)
);

INVxp33_ASAP7_75t_SL g297 ( 
.A(n_281),
.Y(n_297)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_297),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_286),
.B(n_262),
.C(n_261),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_294),
.B(n_262),
.C(n_269),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_294),
.B(n_268),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_301),
.B(n_305),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_289),
.B(n_276),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_303),
.B(n_304),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_293),
.B(n_5),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_307),
.A2(n_7),
.B(n_8),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_308),
.B(n_309),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_288),
.B(n_287),
.Y(n_309)
);

AO21x1_ASAP7_75t_L g310 ( 
.A1(n_297),
.A2(n_284),
.B(n_292),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_310),
.B(n_319),
.Y(n_321)
);

AOI21x1_ASAP7_75t_L g312 ( 
.A1(n_308),
.A2(n_285),
.B(n_295),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_312),
.A2(n_299),
.B(n_298),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_315),
.B(n_9),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_302),
.B(n_288),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_317),
.B(n_318),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_306),
.B(n_7),
.Y(n_318)
);

OAI21x1_ASAP7_75t_L g319 ( 
.A1(n_296),
.A2(n_7),
.B(n_8),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_317),
.B(n_300),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_322),
.B(n_323),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_313),
.B(n_8),
.Y(n_324)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_324),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_316),
.A2(n_8),
.B(n_9),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g334 ( 
.A(n_325),
.B(n_326),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_314),
.B(n_9),
.Y(n_328)
);

INVxp33_ASAP7_75t_L g333 ( 
.A(n_328),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g330 ( 
.A(n_321),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_330),
.A2(n_331),
.B(n_311),
.Y(n_335)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_327),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_335),
.A2(n_336),
.B1(n_329),
.B2(n_320),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_332),
.B(n_327),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_318),
.B(n_334),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_10),
.B1(n_333),
.B2(n_316),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_339),
.A2(n_10),
.B(n_270),
.Y(n_340)
);


endmodule