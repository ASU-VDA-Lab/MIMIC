module fake_jpeg_19066_n_172 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_172);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_172;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVxp33_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_28),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_31),
.A2(n_15),
.B1(n_26),
.B2(n_25),
.Y(n_52)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_17),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_36),
.Y(n_42)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_38),
.Y(n_48)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_40),
.Y(n_58)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_0),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_39),
.A2(n_15),
.B1(n_26),
.B2(n_14),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_45),
.A2(n_23),
.B1(n_20),
.B2(n_2),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_35),
.B(n_14),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_46),
.B(n_47),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_31),
.B(n_19),
.Y(n_47)
);

BUFx8_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_52),
.A2(n_53),
.B1(n_62),
.B2(n_23),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_33),
.A2(n_29),
.B1(n_25),
.B2(n_22),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_19),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_54),
.B(n_0),
.Y(n_74)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_17),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_61),
.B(n_18),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_37),
.A2(n_22),
.B1(n_18),
.B2(n_24),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_51),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_63),
.A2(n_66),
.B1(n_68),
.B2(n_70),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_64),
.B(n_73),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_24),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_65),
.B(n_84),
.Y(n_91)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_74),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_55),
.A2(n_20),
.B1(n_1),
.B2(n_3),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_42),
.B(n_20),
.Y(n_72)
);

OAI32xp33_ASAP7_75t_L g93 ( 
.A1(n_72),
.A2(n_60),
.A3(n_48),
.B1(n_43),
.B2(n_56),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_46),
.B(n_13),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_13),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_75),
.B(n_12),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_58),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_77)
);

A2O1A1Ixp33_ASAP7_75t_SL g92 ( 
.A1(n_77),
.A2(n_79),
.B(n_86),
.C(n_50),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_58),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_79)
);

INVx13_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

BUFx8_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_81),
.Y(n_103)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_43),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_52),
.A2(n_7),
.B1(n_8),
.B2(n_11),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_58),
.A2(n_49),
.B1(n_44),
.B2(n_59),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_48),
.B(n_7),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_87),
.B(n_57),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_92),
.A2(n_94),
.B(n_99),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_70),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_57),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_66),
.B(n_49),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_95),
.B(n_78),
.Y(n_118)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_96),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_81),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_98),
.B(n_104),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_71),
.B(n_56),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_64),
.B(n_65),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_102),
.B(n_107),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_88),
.B(n_87),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_105),
.B(n_108),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_84),
.B(n_76),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_76),
.B(n_80),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_67),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_109),
.B(n_78),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_94),
.B(n_63),
.C(n_85),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_110),
.B(n_111),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_106),
.A2(n_82),
.B1(n_69),
.B2(n_83),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_112),
.B(n_116),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_85),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_113),
.B(n_92),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_101),
.Y(n_114)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_114),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_118),
.A2(n_99),
.B(n_96),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_95),
.A2(n_81),
.B1(n_107),
.B2(n_91),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_120),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_121),
.B(n_126),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_90),
.B(n_91),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_123),
.B(n_124),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_98),
.A2(n_94),
.B1(n_102),
.B2(n_109),
.Y(n_124)
);

OA21x2_ASAP7_75t_SL g126 ( 
.A1(n_89),
.A2(n_99),
.B(n_92),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_128),
.B(n_134),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_131),
.B(n_135),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_122),
.Y(n_134)
);

MAJx2_ASAP7_75t_L g135 ( 
.A(n_117),
.B(n_92),
.C(n_100),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_117),
.A2(n_103),
.B(n_118),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_137),
.B(n_138),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_115),
.A2(n_103),
.B(n_113),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_129),
.B(n_119),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_140),
.B(n_148),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_127),
.B(n_124),
.C(n_111),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_141),
.B(n_127),
.Y(n_149)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_130),
.Y(n_142)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_142),
.Y(n_152)
);

BUFx2_ASAP7_75t_L g143 ( 
.A(n_132),
.Y(n_143)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_143),
.Y(n_155)
);

AO221x1_ASAP7_75t_L g144 ( 
.A1(n_128),
.A2(n_125),
.B1(n_116),
.B2(n_122),
.C(n_110),
.Y(n_144)
);

INVxp33_ASAP7_75t_SL g151 ( 
.A(n_144),
.Y(n_151)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_136),
.Y(n_146)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_146),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_138),
.B(n_115),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_149),
.B(n_150),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_141),
.B(n_137),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_139),
.A2(n_145),
.B(n_148),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_154),
.A2(n_145),
.B(n_151),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_120),
.Y(n_157)
);

OA21x2_ASAP7_75t_L g162 ( 
.A1(n_157),
.A2(n_158),
.B(n_133),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_153),
.B(n_143),
.Y(n_158)
);

OA21x2_ASAP7_75t_SL g159 ( 
.A1(n_151),
.A2(n_154),
.B(n_147),
.Y(n_159)
);

OAI31xp33_ASAP7_75t_L g164 ( 
.A1(n_159),
.A2(n_160),
.A3(n_147),
.B(n_135),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_162),
.B(n_163),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_160),
.A2(n_152),
.B(n_155),
.Y(n_163)
);

NOR2xp67_ASAP7_75t_L g167 ( 
.A(n_164),
.B(n_165),
.Y(n_167)
);

XOR2x1_ASAP7_75t_L g165 ( 
.A(n_161),
.B(n_131),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_162),
.B(n_112),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_168),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_166),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_170),
.B(n_167),
.Y(n_171)
);

NAND2xp33_ASAP7_75t_R g172 ( 
.A(n_171),
.B(n_169),
.Y(n_172)
);


endmodule