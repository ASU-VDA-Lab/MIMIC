module fake_jpeg_7916_n_269 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_269);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_269;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_223;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx4f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_34),
.B(n_39),
.Y(n_62)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_22),
.B(n_15),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_43),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_27),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_50),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_40),
.A2(n_18),
.B1(n_22),
.B2(n_25),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_47),
.A2(n_48),
.B1(n_63),
.B2(n_28),
.Y(n_75)
);

AO22x2_ASAP7_75t_L g48 ( 
.A1(n_39),
.A2(n_20),
.B1(n_32),
.B2(n_26),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_33),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_51),
.B(n_21),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_34),
.A2(n_18),
.B1(n_30),
.B2(n_25),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_52),
.A2(n_17),
.B1(n_30),
.B2(n_24),
.Y(n_69)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_33),
.Y(n_55)
);

OR2x2_ASAP7_75t_SL g86 ( 
.A(n_55),
.B(n_32),
.Y(n_86)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_60),
.Y(n_72)
);

NAND3xp33_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_15),
.C(n_14),
.Y(n_59)
);

INVx2_ASAP7_75t_R g78 ( 
.A(n_59),
.Y(n_78)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_38),
.A2(n_18),
.B1(n_16),
.B2(n_24),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_67),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_0),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_68),
.A2(n_69),
.B(n_71),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_48),
.B(n_55),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_73),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_48),
.A2(n_17),
.B1(n_28),
.B2(n_16),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_74),
.A2(n_79),
.B1(n_81),
.B2(n_64),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_75),
.B(n_88),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_55),
.B(n_1),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_32),
.C(n_26),
.Y(n_93)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_83),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_53),
.A2(n_20),
.B1(n_31),
.B2(n_29),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_53),
.A2(n_31),
.B1(n_29),
.B2(n_21),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_82),
.B(n_85),
.Y(n_91)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_63),
.B(n_11),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_86),
.B(n_89),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_61),
.A2(n_31),
.B1(n_29),
.B2(n_21),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_87),
.A2(n_54),
.B1(n_64),
.B2(n_57),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_65),
.B(n_19),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_72),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g128 ( 
.A(n_90),
.B(n_78),
.Y(n_128)
);

FAx1_ASAP7_75t_SL g120 ( 
.A(n_93),
.B(n_108),
.CI(n_78),
.CON(n_120),
.SN(n_120)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_96),
.A2(n_105),
.B1(n_83),
.B2(n_80),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_77),
.B(n_46),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_88),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_98),
.A2(n_101),
.B1(n_83),
.B2(n_80),
.Y(n_127)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_70),
.Y(n_99)
);

INVx5_ASAP7_75t_SL g117 ( 
.A(n_99),
.Y(n_117)
);

NAND2xp33_ASAP7_75t_SL g100 ( 
.A(n_71),
.B(n_65),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_100),
.A2(n_87),
.B(n_76),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_71),
.A2(n_85),
.B1(n_68),
.B2(n_75),
.Y(n_101)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_66),
.Y(n_103)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_103),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_71),
.A2(n_57),
.B1(n_44),
.B2(n_45),
.Y(n_105)
);

INVx13_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_106),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_84),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_107),
.Y(n_138)
);

FAx1_ASAP7_75t_SL g108 ( 
.A(n_86),
.B(n_44),
.CI(n_26),
.CON(n_108),
.SN(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_66),
.Y(n_109)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_109),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_82),
.B(n_1),
.Y(n_110)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_110),
.Y(n_123)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_72),
.Y(n_111)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_111),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_86),
.B(n_1),
.Y(n_112)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_112),
.Y(n_135)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_70),
.Y(n_114)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_114),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_113),
.A2(n_76),
.B(n_68),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_115),
.A2(n_120),
.B(n_122),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_116),
.B(n_129),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_111),
.B(n_78),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_125),
.B(n_128),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_126),
.A2(n_134),
.B1(n_98),
.B2(n_110),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_127),
.A2(n_130),
.B1(n_131),
.B2(n_133),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_95),
.B(n_76),
.Y(n_129)
);

OAI21xp33_ASAP7_75t_SL g130 ( 
.A1(n_102),
.A2(n_68),
.B(n_19),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_101),
.A2(n_89),
.B1(n_70),
.B2(n_79),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_95),
.A2(n_81),
.B1(n_19),
.B2(n_1),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_96),
.A2(n_8),
.B1(n_3),
.B2(n_4),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_113),
.A2(n_8),
.B(n_4),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_136),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_91),
.B(n_2),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_137),
.B(n_94),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_102),
.A2(n_2),
.B(n_5),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_139),
.B(n_140),
.C(n_112),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_105),
.B(n_6),
.C(n_7),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_138),
.B(n_90),
.Y(n_143)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_143),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_144),
.B(n_145),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_116),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_135),
.B(n_100),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_146),
.A2(n_118),
.B(n_114),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_138),
.B(n_94),
.Y(n_148)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_148),
.Y(n_180)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_131),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_149),
.B(n_150),
.Y(n_169)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_127),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_151),
.A2(n_152),
.B1(n_161),
.B2(n_135),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_133),
.A2(n_91),
.B1(n_109),
.B2(n_103),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_153),
.B(n_160),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_137),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_154),
.B(n_164),
.Y(n_178)
);

NAND2x1_ASAP7_75t_L g155 ( 
.A(n_115),
.B(n_136),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_155),
.A2(n_166),
.B(n_7),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_119),
.B(n_107),
.Y(n_157)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_157),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_129),
.B(n_93),
.C(n_97),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_158),
.B(n_128),
.C(n_124),
.Y(n_183)
);

OAI32xp33_ASAP7_75t_L g159 ( 
.A1(n_122),
.A2(n_108),
.A3(n_104),
.B1(n_92),
.B2(n_106),
.Y(n_159)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_159),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_119),
.B(n_108),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_126),
.A2(n_104),
.B1(n_108),
.B2(n_106),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_121),
.B(n_107),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_163),
.B(n_167),
.Y(n_187)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_117),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_132),
.B(n_104),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_165),
.Y(n_175)
);

NOR4xp25_ASAP7_75t_L g166 ( 
.A(n_120),
.B(n_6),
.C(n_7),
.D(n_8),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_117),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_156),
.B(n_120),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_168),
.B(n_182),
.C(n_183),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_171),
.B(n_189),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_163),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_172),
.B(n_184),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_150),
.A2(n_121),
.B1(n_132),
.B2(n_123),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_174),
.A2(n_185),
.B1(n_147),
.B2(n_166),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_155),
.B(n_140),
.Y(n_176)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_176),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_149),
.A2(n_134),
.B1(n_123),
.B2(n_124),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_177),
.A2(n_151),
.B1(n_147),
.B2(n_145),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_156),
.B(n_139),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_161),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_155),
.A2(n_107),
.B(n_10),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_186),
.B(n_188),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_153),
.Y(n_189)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_187),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_192),
.B(n_195),
.Y(n_212)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_187),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_183),
.B(n_158),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_197),
.B(n_204),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_178),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_198),
.B(n_201),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_199),
.B(n_177),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_182),
.B(n_162),
.Y(n_200)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_200),
.Y(n_222)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_169),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_168),
.B(n_141),
.C(n_160),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_202),
.B(n_204),
.C(n_207),
.Y(n_224)
);

XNOR2x1_ASAP7_75t_L g203 ( 
.A(n_176),
.B(n_159),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_203),
.B(n_188),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_173),
.B(n_141),
.C(n_142),
.Y(n_204)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_169),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_206),
.B(n_208),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_179),
.B(n_142),
.C(n_146),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_174),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_179),
.B(n_146),
.C(n_152),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_209),
.B(n_207),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_210),
.A2(n_186),
.B(n_184),
.Y(n_213)
);

INVx13_ASAP7_75t_L g211 ( 
.A(n_198),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_211),
.B(n_223),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_213),
.A2(n_144),
.B(n_154),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_203),
.A2(n_190),
.B1(n_170),
.B2(n_175),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_215),
.B(n_221),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_205),
.A2(n_180),
.B1(n_189),
.B2(n_171),
.Y(n_216)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_216),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_217),
.B(n_218),
.C(n_219),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_194),
.B(n_209),
.Y(n_219)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_220),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_191),
.A2(n_193),
.B1(n_200),
.B2(n_196),
.Y(n_223)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_202),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_226),
.B(n_176),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_219),
.B(n_194),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_228),
.B(n_224),
.C(n_218),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_230),
.Y(n_243)
);

NOR2xp67_ASAP7_75t_SL g231 ( 
.A(n_222),
.B(n_181),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_231),
.B(n_9),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_217),
.B(n_185),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_233),
.B(n_238),
.Y(n_246)
);

OAI321xp33_ASAP7_75t_L g240 ( 
.A1(n_236),
.A2(n_221),
.A3(n_215),
.B1(n_213),
.B2(n_225),
.C(n_224),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_211),
.B(n_164),
.Y(n_237)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_237),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_214),
.B(n_167),
.Y(n_238)
);

FAx1_ASAP7_75t_SL g239 ( 
.A(n_233),
.B(n_223),
.CI(n_212),
.CON(n_239),
.SN(n_239)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_239),
.B(n_241),
.Y(n_251)
);

OR2x2_ASAP7_75t_L g249 ( 
.A(n_240),
.B(n_244),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_229),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_242),
.B(n_227),
.C(n_99),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_232),
.B(n_234),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_247),
.B(n_9),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_246),
.A2(n_235),
.B(n_228),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_248),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_246),
.B(n_235),
.Y(n_250)
);

XNOR2x1_ASAP7_75t_L g256 ( 
.A(n_250),
.B(n_239),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_245),
.B(n_118),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_252),
.B(n_253),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_254),
.B(n_255),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_243),
.B(n_227),
.Y(n_255)
);

AOI322xp5_ASAP7_75t_L g264 ( 
.A1(n_256),
.A2(n_260),
.A3(n_9),
.B1(n_13),
.B2(n_14),
.C1(n_247),
.C2(n_246),
.Y(n_264)
);

FAx1_ASAP7_75t_SL g260 ( 
.A(n_255),
.B(n_15),
.CI(n_10),
.CON(n_260),
.SN(n_260)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_258),
.Y(n_261)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_261),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_259),
.B(n_249),
.Y(n_262)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_262),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_257),
.B(n_251),
.C(n_13),
.Y(n_263)
);

MAJx2_ASAP7_75t_L g267 ( 
.A(n_265),
.B(n_257),
.C(n_263),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_267),
.B(n_264),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_268),
.B(n_266),
.Y(n_269)
);


endmodule