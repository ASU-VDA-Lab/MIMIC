module real_jpeg_7583_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_525;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_531;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_534;
wire n_181;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp33_ASAP7_75t_L g276 ( 
.A1(n_0),
.A2(n_192),
.B1(n_210),
.B2(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_0),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g357 ( 
.A1(n_0),
.A2(n_119),
.B1(n_277),
.B2(n_358),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_0),
.A2(n_112),
.B1(n_277),
.B2(n_392),
.Y(n_391)
);

OAI22xp33_ASAP7_75t_L g454 ( 
.A1(n_0),
.A2(n_47),
.B1(n_277),
.B2(n_455),
.Y(n_454)
);

INVx8_ASAP7_75t_L g199 ( 
.A(n_1),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_1),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_1),
.Y(n_243)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_1),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_1),
.Y(n_417)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_2),
.Y(n_59)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_2),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g328 ( 
.A(n_2),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_2),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_2),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_2),
.Y(n_457)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_3),
.A2(n_58),
.B1(n_60),
.B2(n_64),
.Y(n_57)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_3),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_3),
.A2(n_64),
.B1(n_107),
.B2(n_109),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_SL g367 ( 
.A1(n_3),
.A2(n_64),
.B1(n_189),
.B2(n_368),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_3),
.A2(n_64),
.B1(n_402),
.B2(n_405),
.Y(n_401)
);

OAI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_4),
.A2(n_187),
.B1(n_191),
.B2(n_192),
.Y(n_186)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_4),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_4),
.A2(n_161),
.B1(n_191),
.B2(n_255),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_L g352 ( 
.A1(n_4),
.A2(n_191),
.B1(n_353),
.B2(n_355),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_4),
.A2(n_191),
.B1(n_347),
.B2(n_348),
.Y(n_397)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_5),
.A2(n_161),
.B1(n_162),
.B2(n_166),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_5),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_5),
.B(n_176),
.C(n_179),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_5),
.B(n_98),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_5),
.B(n_205),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_5),
.B(n_141),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_5),
.B(n_261),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_6),
.A2(n_40),
.B1(n_63),
.B2(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_6),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_6),
.A2(n_74),
.B1(n_305),
.B2(n_306),
.Y(n_304)
);

OAI22xp33_ASAP7_75t_SL g377 ( 
.A1(n_6),
.A2(n_74),
.B1(n_378),
.B2(n_382),
.Y(n_377)
);

AOI22xp33_ASAP7_75t_SL g394 ( 
.A1(n_6),
.A2(n_74),
.B1(n_96),
.B2(n_395),
.Y(n_394)
);

AOI22xp33_ASAP7_75t_L g214 ( 
.A1(n_7),
.A2(n_161),
.B1(n_215),
.B2(n_216),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_7),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_7),
.A2(n_187),
.B1(n_207),
.B2(n_215),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_7),
.A2(n_215),
.B1(n_294),
.B2(n_296),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_7),
.A2(n_51),
.B1(n_215),
.B2(n_421),
.Y(n_420)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

INVx3_ASAP7_75t_L g533 ( 
.A(n_9),
.Y(n_533)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_10),
.Y(n_123)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_10),
.Y(n_127)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_10),
.Y(n_132)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_11),
.Y(n_101)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_12),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_12),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_12),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_13),
.A2(n_47),
.B1(n_48),
.B2(n_54),
.Y(n_46)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_13),
.A2(n_54),
.B1(n_112),
.B2(n_113),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_13),
.A2(n_54),
.B1(n_100),
.B2(n_143),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_13),
.A2(n_54),
.B1(n_188),
.B2(n_373),
.Y(n_372)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_14),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_15),
.A2(n_76),
.B1(n_79),
.B2(n_81),
.Y(n_75)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_15),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g333 ( 
.A1(n_15),
.A2(n_81),
.B1(n_207),
.B2(n_334),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_15),
.A2(n_81),
.B1(n_217),
.B2(n_386),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_15),
.A2(n_81),
.B1(n_434),
.B2(n_439),
.Y(n_433)
);

INVxp33_ASAP7_75t_L g537 ( 
.A(n_16),
.Y(n_537)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_18),
.A2(n_144),
.B1(n_169),
.B2(n_172),
.Y(n_168)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_18),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_18),
.A2(n_172),
.B1(n_207),
.B2(n_210),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_18),
.A2(n_172),
.B1(n_267),
.B2(n_270),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_18),
.A2(n_61),
.B1(n_172),
.B2(n_347),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_532),
.B(n_534),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_67),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_66),
.Y(n_21)
);

OR2x2_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_55),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_23),
.B(n_55),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_35),
.B(n_45),
.Y(n_23)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_24),
.B(n_346),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_24),
.B(n_454),
.Y(n_453)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_25),
.B(n_166),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_25),
.A2(n_56),
.B1(n_397),
.B2(n_420),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_31),
.B2(n_33),
.Y(n_25)
);

INVx6_ASAP7_75t_L g354 ( 
.A(n_27),
.Y(n_354)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_28),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_29),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_29),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_29),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_29),
.Y(n_438)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_30),
.Y(n_97)
);

BUFx5_ASAP7_75t_L g264 ( 
.A(n_30),
.Y(n_264)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_30),
.Y(n_272)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx6_ASAP7_75t_SL g280 ( 
.A(n_32),
.Y(n_280)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_35),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_35),
.A2(n_342),
.B(n_344),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_35),
.B(n_346),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_40),
.B1(n_42),
.B2(n_43),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

OAI32xp33_ASAP7_75t_L g320 ( 
.A1(n_40),
.A2(n_321),
.A3(n_322),
.B1(n_323),
.B2(n_325),
.Y(n_320)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_43),
.Y(n_322)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_44),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_46),
.A2(n_56),
.B1(n_57),
.B2(n_65),
.Y(n_55)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_55),
.B(n_69),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_55),
.B(n_69),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_56),
.A2(n_65),
.B1(n_73),
.B2(n_75),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_56),
.A2(n_57),
.B1(n_65),
.B2(n_75),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g396 ( 
.A1(n_56),
.A2(n_345),
.B(n_397),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g503 ( 
.A1(n_56),
.A2(n_65),
.B1(n_73),
.B2(n_504),
.Y(n_503)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx3_ASAP7_75t_L g422 ( 
.A(n_63),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_L g468 ( 
.A1(n_65),
.A2(n_420),
.B(n_458),
.Y(n_468)
);

AO21x1_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_150),
.B(n_531),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_146),
.C(n_147),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g526 ( 
.A1(n_70),
.A2(n_71),
.B1(n_527),
.B2(n_528),
.Y(n_526)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_82),
.C(n_114),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_SL g518 ( 
.A(n_72),
.B(n_519),
.Y(n_518)
);

INVx2_ASAP7_75t_SL g76 ( 
.A(n_77),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_82),
.A2(n_114),
.B1(n_115),
.B2(n_520),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_82),
.Y(n_520)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_106),
.B1(n_110),
.B2(n_111),
.Y(n_82)
);

INVx3_ASAP7_75t_SL g148 ( 
.A(n_83),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_83),
.A2(n_110),
.B1(n_293),
.B2(n_352),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_83),
.A2(n_110),
.B1(n_391),
.B2(n_394),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g507 ( 
.A1(n_83),
.A2(n_106),
.B1(n_110),
.B2(n_508),
.Y(n_507)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_98),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_90),
.B1(n_91),
.B2(n_95),
.Y(n_84)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_89),
.Y(n_94)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_94),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_95),
.B(n_324),
.Y(n_323)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

OAI21xp33_ASAP7_75t_SL g258 ( 
.A1(n_96),
.A2(n_166),
.B(n_259),
.Y(n_258)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_97),
.Y(n_113)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_97),
.Y(n_295)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_98),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_98),
.A2(n_148),
.B(n_149),
.Y(n_147)
);

AOI22x1_ASAP7_75t_L g423 ( 
.A1(n_98),
.A2(n_148),
.B1(n_300),
.B2(n_424),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_98),
.A2(n_148),
.B1(n_432),
.B2(n_433),
.Y(n_431)
);

AO22x2_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_100),
.B1(n_102),
.B2(n_104),
.Y(n_98)
);

INVx5_ASAP7_75t_L g388 ( 
.A(n_100),
.Y(n_388)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx11_ASAP7_75t_L g103 ( 
.A(n_101),
.Y(n_103)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_101),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_101),
.Y(n_161)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_101),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g381 ( 
.A(n_101),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_103),
.Y(n_129)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_103),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_103),
.Y(n_358)
);

INVx6_ASAP7_75t_L g384 ( 
.A(n_103),
.Y(n_384)
);

AOI32xp33_ASAP7_75t_L g279 ( 
.A1(n_104),
.A2(n_161),
.A3(n_260),
.B1(n_280),
.B2(n_281),
.Y(n_279)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx2_ASAP7_75t_L g282 ( 
.A(n_105),
.Y(n_282)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_110),
.B(n_266),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_110),
.A2(n_293),
.B(n_299),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_111),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_114),
.A2(n_115),
.B1(n_506),
.B2(n_507),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_114),
.B(n_503),
.C(n_506),
.Y(n_514)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_140),
.B(n_142),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_116),
.A2(n_160),
.B(n_167),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_116),
.A2(n_140),
.B1(n_214),
.B2(n_254),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_116),
.A2(n_167),
.B(n_254),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_116),
.A2(n_140),
.B1(n_357),
.B2(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_SL g116 ( 
.A(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_117),
.B(n_168),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_117),
.A2(n_141),
.B1(n_377),
.B2(n_385),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_117),
.A2(n_141),
.B1(n_385),
.B2(n_401),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_117),
.A2(n_141),
.B1(n_401),
.B2(n_445),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_130),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_121),
.B1(n_124),
.B2(n_128),
.Y(n_118)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx5_ASAP7_75t_L g139 ( 
.A(n_127),
.Y(n_139)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx5_ASAP7_75t_L g406 ( 
.A(n_129),
.Y(n_406)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_130),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_130),
.A2(n_214),
.B(n_218),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_133),
.B1(n_137),
.B2(n_139),
.Y(n_130)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_132),
.Y(n_178)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_135),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_136),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_136),
.Y(n_183)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx8_ASAP7_75t_L g308 ( 
.A(n_138),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_140),
.A2(n_218),
.B(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_141),
.B(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_142),
.Y(n_445)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_143),
.Y(n_217)
);

INVx4_ASAP7_75t_SL g143 ( 
.A(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g528 ( 
.A(n_146),
.B(n_147),
.Y(n_528)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_148),
.A2(n_258),
.B(n_265),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_148),
.B(n_300),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_148),
.A2(n_265),
.B(n_471),
.Y(n_470)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_151),
.A2(n_525),
.B(n_530),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_152),
.A2(n_497),
.B(n_522),
.Y(n_151)
);

OAI311xp33_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_361),
.A3(n_473),
.B1(n_491),
.C1(n_492),
.Y(n_152)
);

AOI21x1_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_314),
.B(n_360),
.Y(n_153)
);

AO21x1_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_284),
.B(n_313),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_156),
.A2(n_248),
.B(n_283),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_221),
.B(n_247),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_184),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_158),
.B(n_184),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_173),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_159),
.A2(n_173),
.B1(n_174),
.B2(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_159),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_162),
.B(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx6_ASAP7_75t_L g404 ( 
.A(n_165),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_166),
.A2(n_196),
.B(n_203),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_166),
.B(n_326),
.Y(n_325)
);

OAI21xp33_ASAP7_75t_SL g342 ( 
.A1(n_166),
.A2(n_325),
.B(n_343),
.Y(n_342)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_170),
.Y(n_255)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_182),
.Y(n_210)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_183),
.Y(n_190)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_183),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_211),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_185),
.B(n_212),
.C(n_220),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_196),
.B(n_203),
.Y(n_185)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_186),
.Y(n_241)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx4_ASAP7_75t_SL g193 ( 
.A(n_194),
.Y(n_193)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_196),
.A2(n_278),
.B1(n_331),
.B2(n_332),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_196),
.A2(n_367),
.B1(n_370),
.B2(n_372),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_SL g407 ( 
.A1(n_196),
.A2(n_372),
.B(n_408),
.Y(n_407)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_197),
.B(n_206),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_197),
.A2(n_240),
.B1(n_241),
.B2(n_242),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_197),
.A2(n_276),
.B1(n_304),
.B2(n_309),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_197),
.A2(n_333),
.B1(n_415),
.B2(n_416),
.Y(n_414)
);

OR2x2_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_200),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_199),
.Y(n_408)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

BUFx5_ASAP7_75t_L g369 ( 
.A(n_202),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_206),
.Y(n_203)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_204),
.Y(n_234)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_205),
.Y(n_371)
);

INVx8_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

BUFx8_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_209),
.Y(n_335)
);

BUFx5_ASAP7_75t_L g375 ( 
.A(n_209),
.Y(n_375)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_210),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_212),
.A2(n_213),
.B1(n_219),
.B2(n_220),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

NAND2xp33_ASAP7_75t_SL g281 ( 
.A(n_216),
.B(n_282),
.Y(n_281)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_238),
.B(n_246),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_231),
.B(n_237),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_230),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_229),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx6_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_232),
.B(n_236),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_232),
.B(n_236),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_234),
.B(n_235),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_233),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_235),
.A2(n_275),
.B(n_278),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_244),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_239),
.B(n_244),
.Y(n_246)
);

INVx4_ASAP7_75t_L g278 ( 
.A(n_242),
.Y(n_278)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_249),
.B(n_250),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_273),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_253),
.B1(n_256),
.B2(n_257),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_253),
.B(n_256),
.C(n_273),
.Y(n_285)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVxp33_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

BUFx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx6_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_264),
.Y(n_298)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_264),
.Y(n_442)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_266),
.Y(n_300)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

BUFx12f_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_269),
.Y(n_393)
);

INVx8_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx4_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx4_ASAP7_75t_L g395 ( 
.A(n_272),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_279),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_274),
.B(n_279),
.Y(n_290)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_285),
.B(n_286),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_288),
.B1(n_291),
.B2(n_312),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_SL g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_289),
.B(n_290),
.C(n_312),
.Y(n_315)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_291),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_301),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_292),
.B(n_302),
.C(n_303),
.Y(n_336)
);

INVx5_ASAP7_75t_L g355 ( 
.A(n_294),
.Y(n_355)
);

INVx4_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_303),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_304),
.Y(n_331)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx4_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx5_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g360 ( 
.A(n_315),
.B(n_316),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_339),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_318),
.A2(n_336),
.B1(n_337),
.B2(n_338),
.Y(n_317)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_318),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_319),
.A2(n_320),
.B1(n_329),
.B2(n_330),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_320),
.B(n_329),
.Y(n_469)
);

INVx4_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_336),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_336),
.B(n_337),
.C(n_339),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_340),
.A2(n_341),
.B1(n_350),
.B2(n_359),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_340),
.B(n_351),
.C(n_356),
.Y(n_482)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx3_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx4_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_350),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_SL g350 ( 
.A(n_351),
.B(n_356),
.Y(n_350)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_352),
.Y(n_471)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

NAND2xp33_ASAP7_75t_SL g361 ( 
.A(n_362),
.B(n_459),
.Y(n_361)
);

A2O1A1Ixp33_ASAP7_75t_SL g492 ( 
.A1(n_362),
.A2(n_459),
.B(n_493),
.C(n_496),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_425),
.Y(n_362)
);

OR2x2_ASAP7_75t_L g491 ( 
.A(n_363),
.B(n_425),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_398),
.C(n_410),
.Y(n_363)
);

FAx1_ASAP7_75t_SL g472 ( 
.A(n_364),
.B(n_398),
.CI(n_410),
.CON(n_472),
.SN(n_472)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_389),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_365),
.B(n_390),
.C(n_396),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_376),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_366),
.B(n_376),
.Y(n_465)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_367),
.Y(n_415)
);

INVx5_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

BUFx3_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

CKINVDCx14_ASAP7_75t_R g373 ( 
.A(n_374),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_377),
.Y(n_413)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx3_ASAP7_75t_SL g382 ( 
.A(n_383),
.Y(n_382)
);

INVx8_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_396),
.Y(n_389)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_391),
.Y(n_424)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_394),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_399),
.A2(n_400),
.B1(n_407),
.B2(n_409),
.Y(n_398)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_400),
.B(n_407),
.Y(n_449)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_407),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_407),
.A2(n_409),
.B1(n_451),
.B2(n_452),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_L g500 ( 
.A1(n_407),
.A2(n_449),
.B(n_452),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_418),
.C(n_423),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_411),
.B(n_463),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_412),
.B(n_414),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_412),
.B(n_414),
.Y(n_481)
);

INVx3_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_418),
.A2(n_419),
.B1(n_423),
.B2(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_423),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_427),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_426),
.B(n_429),
.C(n_447),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_428),
.A2(n_429),
.B1(n_447),
.B2(n_448),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_430),
.A2(n_443),
.B(n_446),
.Y(n_429)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_431),
.B(n_444),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g508 ( 
.A(n_433),
.Y(n_508)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx4_ASAP7_75t_SL g436 ( 
.A(n_437),
.Y(n_436)
);

INVx5_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

FAx1_ASAP7_75t_SL g499 ( 
.A(n_446),
.B(n_500),
.CI(n_501),
.CON(n_499),
.SN(n_499)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_446),
.B(n_500),
.C(n_501),
.Y(n_521)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_450),
.Y(n_448)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_458),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g504 ( 
.A(n_454),
.Y(n_504)
);

INVx3_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

INVx8_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_460),
.B(n_472),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_460),
.B(n_472),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_465),
.C(n_466),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_461),
.A2(n_462),
.B1(n_465),
.B2(n_485),
.Y(n_484)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_465),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_466),
.B(n_484),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_469),
.C(n_470),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_467),
.A2(n_468),
.B1(n_470),
.B2(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_469),
.B(n_478),
.Y(n_477)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_470),
.Y(n_479)
);

BUFx24_ASAP7_75t_SL g539 ( 
.A(n_472),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_474),
.B(n_486),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

OAI21xp5_ASAP7_75t_L g493 ( 
.A1(n_475),
.A2(n_494),
.B(n_495),
.Y(n_493)
);

NOR2x1_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_483),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_476),
.B(n_483),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_477),
.B(n_480),
.C(n_482),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_477),
.B(n_489),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_480),
.A2(n_481),
.B1(n_482),
.B2(n_490),
.Y(n_489)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_482),
.Y(n_490)
);

OR2x2_ASAP7_75t_L g486 ( 
.A(n_487),
.B(n_488),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_487),
.B(n_488),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_498),
.B(n_511),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_SL g498 ( 
.A(n_499),
.B(n_510),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_499),
.B(n_510),
.Y(n_523)
);

BUFx24_ASAP7_75t_SL g538 ( 
.A(n_499),
.Y(n_538)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_502),
.A2(n_503),
.B1(n_505),
.B2(n_509),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_502),
.A2(n_503),
.B1(n_517),
.B2(n_518),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_502),
.B(n_513),
.C(n_517),
.Y(n_529)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_505),
.Y(n_509)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

OAI21xp5_ASAP7_75t_L g522 ( 
.A1(n_511),
.A2(n_523),
.B(n_524),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_SL g511 ( 
.A(n_512),
.B(n_521),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_512),
.B(n_521),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_L g512 ( 
.A1(n_513),
.A2(n_514),
.B1(n_515),
.B2(n_516),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_526),
.B(n_529),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_526),
.B(n_529),
.Y(n_530)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_528),
.Y(n_527)
);

INVx8_ASAP7_75t_L g532 ( 
.A(n_533),
.Y(n_532)
);

INVx13_ASAP7_75t_L g536 ( 
.A(n_533),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_535),
.B(n_537),
.Y(n_534)
);

BUFx12f_ASAP7_75t_L g535 ( 
.A(n_536),
.Y(n_535)
);


endmodule