module fake_jpeg_17719_n_19 (n_3, n_2, n_1, n_0, n_4, n_19);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;

output n_19;

wire n_13;
wire n_10;
wire n_6;
wire n_14;
wire n_18;
wire n_16;
wire n_9;
wire n_5;
wire n_11;
wire n_17;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

INVx1_ASAP7_75t_L g5 ( 
.A(n_4),
.Y(n_5)
);

INVx4_ASAP7_75t_L g6 ( 
.A(n_4),
.Y(n_6)
);

INVx1_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);

INVx8_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

MAJx2_ASAP7_75t_L g9 ( 
.A(n_6),
.B(n_0),
.C(n_1),
.Y(n_9)
);

MAJIxp5_ASAP7_75t_L g14 ( 
.A(n_9),
.B(n_7),
.C(n_2),
.Y(n_14)
);

AND2x2_ASAP7_75t_L g10 ( 
.A(n_5),
.B(n_0),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_10),
.B(n_11),
.Y(n_13)
);

OR2x2_ASAP7_75t_L g11 ( 
.A(n_5),
.B(n_0),
.Y(n_11)
);

MAJIxp5_ASAP7_75t_L g12 ( 
.A(n_10),
.B(n_5),
.C(n_7),
.Y(n_12)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_12),
.B(n_14),
.C(n_7),
.Y(n_15)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_15),
.B(n_16),
.C(n_6),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_13),
.A2(n_6),
.B1(n_8),
.B2(n_11),
.Y(n_16)
);

AOI332xp33_ASAP7_75t_L g18 ( 
.A1(n_17),
.A2(n_1),
.A3(n_2),
.B1(n_3),
.B2(n_8),
.B3(n_9),
.C1(n_15),
.C2(n_16),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_18),
.B(n_3),
.Y(n_19)
);


endmodule