module fake_netlist_1_6_n_789 (n_117, n_44, n_133, n_149, n_81, n_69, n_185, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_125, n_9, n_161, n_10, n_177, n_130, n_103, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_154, n_7, n_29, n_165, n_146, n_45, n_85, n_181, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_139, n_16, n_13, n_169, n_152, n_113, n_95, n_124, n_156, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_24, n_78, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_38, n_64, n_142, n_184, n_46, n_31, n_58, n_122, n_138, n_126, n_178, n_118, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_12, n_86, n_143, n_182, n_166, n_162, n_186, n_75, n_163, n_105, n_159, n_174, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_67, n_77, n_20, n_2, n_147, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_150, n_168, n_3, n_18, n_110, n_66, n_134, n_1, n_164, n_82, n_106, n_175, n_15, n_173, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_96, n_39, n_789);
input n_117;
input n_44;
input n_133;
input n_149;
input n_81;
input n_69;
input n_185;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_125;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_103;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_154;
input n_7;
input n_29;
input n_165;
input n_146;
input n_45;
input n_85;
input n_181;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_139;
input n_16;
input n_13;
input n_169;
input n_152;
input n_113;
input n_95;
input n_124;
input n_156;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_38;
input n_64;
input n_142;
input n_184;
input n_46;
input n_31;
input n_58;
input n_122;
input n_138;
input n_126;
input n_178;
input n_118;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_12;
input n_86;
input n_143;
input n_182;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_105;
input n_159;
input n_174;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_67;
input n_77;
input n_20;
input n_2;
input n_147;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_150;
input n_168;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_1;
input n_164;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_96;
input n_39;
output n_789;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_755;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_607;
wire n_431;
wire n_484;
wire n_496;
wire n_667;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_637;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_383;
wire n_288;
wire n_661;
wire n_762;
wire n_672;
wire n_627;
wire n_532;
wire n_758;
wire n_544;
wire n_400;
wire n_787;
wire n_296;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_476;
wire n_434;
wire n_384;
wire n_227;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_489;
wire n_777;
wire n_752;
wire n_732;
wire n_199;
wire n_351;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_517;
wire n_560;
wire n_479;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_608;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_767;
wire n_293;
wire n_506;
wire n_533;
wire n_393;
wire n_490;
wire n_247;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_322;
wire n_310;
wire n_708;
wire n_307;
wire n_191;
wire n_634;
wire n_610;
wire n_730;
wire n_771;
wire n_696;
wire n_735;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_415;
wire n_235;
wire n_243;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_760;
wire n_751;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_207;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_578;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_776;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_285;
wire n_195;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_673;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_409;
wire n_363;
wire n_315;
wire n_733;
wire n_295;
wire n_654;
wire n_263;
wire n_495;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_749;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_449;
wire n_300;
wire n_734;
wire n_524;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_766;
wire n_602;
wire n_198;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_410;
wire n_774;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_675;
wire n_291;
wire n_504;
wire n_581;
wire n_458;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_187;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_713;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_736;
wire n_194;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_781;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g187 ( .A(n_148), .Y(n_187) );
BUFx6f_ASAP7_75t_L g188 ( .A(n_63), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_105), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_175), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_135), .Y(n_191) );
CKINVDCx5p33_ASAP7_75t_R g192 ( .A(n_44), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_142), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_131), .Y(n_194) );
CKINVDCx14_ASAP7_75t_R g195 ( .A(n_93), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_61), .Y(n_196) );
CKINVDCx5p33_ASAP7_75t_R g197 ( .A(n_67), .Y(n_197) );
CKINVDCx20_ASAP7_75t_R g198 ( .A(n_181), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_112), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_64), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_74), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_119), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_143), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_57), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_11), .Y(n_205) );
BUFx3_ASAP7_75t_L g206 ( .A(n_52), .Y(n_206) );
INVx3_ASAP7_75t_L g207 ( .A(n_125), .Y(n_207) );
CKINVDCx14_ASAP7_75t_R g208 ( .A(n_100), .Y(n_208) );
CKINVDCx20_ASAP7_75t_R g209 ( .A(n_43), .Y(n_209) );
CKINVDCx5p33_ASAP7_75t_R g210 ( .A(n_48), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_133), .Y(n_211) );
CKINVDCx5p33_ASAP7_75t_R g212 ( .A(n_85), .Y(n_212) );
HB1xp67_ASAP7_75t_L g213 ( .A(n_164), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_81), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_165), .Y(n_215) );
CKINVDCx5p33_ASAP7_75t_R g216 ( .A(n_160), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_128), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_151), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_80), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_158), .Y(n_220) );
INVxp33_ASAP7_75t_SL g221 ( .A(n_41), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_55), .Y(n_222) );
CKINVDCx5p33_ASAP7_75t_R g223 ( .A(n_145), .Y(n_223) );
CKINVDCx5p33_ASAP7_75t_R g224 ( .A(n_153), .Y(n_224) );
INVx3_ASAP7_75t_L g225 ( .A(n_53), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_48), .Y(n_226) );
CKINVDCx5p33_ASAP7_75t_R g227 ( .A(n_174), .Y(n_227) );
HB1xp67_ASAP7_75t_L g228 ( .A(n_176), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_130), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_186), .Y(n_230) );
HB1xp67_ASAP7_75t_L g231 ( .A(n_113), .Y(n_231) );
BUFx3_ASAP7_75t_L g232 ( .A(n_132), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_184), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_58), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_139), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_177), .Y(n_236) );
BUFx2_ASAP7_75t_L g237 ( .A(n_109), .Y(n_237) );
HB1xp67_ASAP7_75t_L g238 ( .A(n_26), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_183), .Y(n_239) );
CKINVDCx20_ASAP7_75t_R g240 ( .A(n_185), .Y(n_240) );
NOR2xp67_ASAP7_75t_L g241 ( .A(n_20), .B(n_138), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_72), .Y(n_242) );
INVx2_ASAP7_75t_L g243 ( .A(n_180), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_116), .Y(n_244) );
BUFx2_ASAP7_75t_SL g245 ( .A(n_146), .Y(n_245) );
BUFx3_ASAP7_75t_L g246 ( .A(n_59), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_114), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_118), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_140), .Y(n_249) );
INVx2_ASAP7_75t_L g250 ( .A(n_120), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_124), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_94), .Y(n_252) );
INVx3_ASAP7_75t_L g253 ( .A(n_26), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_152), .Y(n_254) );
HB1xp67_ASAP7_75t_L g255 ( .A(n_53), .Y(n_255) );
CKINVDCx5p33_ASAP7_75t_R g256 ( .A(n_10), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_178), .Y(n_257) );
INVxp67_ASAP7_75t_SL g258 ( .A(n_126), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_76), .Y(n_259) );
CKINVDCx5p33_ASAP7_75t_R g260 ( .A(n_123), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_19), .Y(n_261) );
CKINVDCx20_ASAP7_75t_R g262 ( .A(n_122), .Y(n_262) );
CKINVDCx5p33_ASAP7_75t_R g263 ( .A(n_179), .Y(n_263) );
BUFx5_ASAP7_75t_L g264 ( .A(n_150), .Y(n_264) );
CKINVDCx5p33_ASAP7_75t_R g265 ( .A(n_17), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_7), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_172), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_137), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_51), .Y(n_269) );
CKINVDCx5p33_ASAP7_75t_R g270 ( .A(n_35), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_65), .Y(n_271) );
CKINVDCx5p33_ASAP7_75t_R g272 ( .A(n_117), .Y(n_272) );
CKINVDCx20_ASAP7_75t_R g273 ( .A(n_121), .Y(n_273) );
CKINVDCx5p33_ASAP7_75t_R g274 ( .A(n_66), .Y(n_274) );
CKINVDCx5p33_ASAP7_75t_R g275 ( .A(n_60), .Y(n_275) );
BUFx6f_ASAP7_75t_L g276 ( .A(n_11), .Y(n_276) );
CKINVDCx14_ASAP7_75t_R g277 ( .A(n_36), .Y(n_277) );
CKINVDCx20_ASAP7_75t_R g278 ( .A(n_14), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_78), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_149), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_115), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_141), .Y(n_282) );
INVxp67_ASAP7_75t_L g283 ( .A(n_134), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_12), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_24), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_108), .Y(n_286) );
BUFx6f_ASAP7_75t_L g287 ( .A(n_167), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_54), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_157), .Y(n_289) );
CKINVDCx20_ASAP7_75t_R g290 ( .A(n_110), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_102), .Y(n_291) );
BUFx6f_ASAP7_75t_L g292 ( .A(n_188), .Y(n_292) );
INVx3_ASAP7_75t_L g293 ( .A(n_225), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_207), .Y(n_294) );
CKINVDCx5p33_ASAP7_75t_R g295 ( .A(n_277), .Y(n_295) );
AND2x4_ASAP7_75t_L g296 ( .A(n_225), .B(n_0), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_225), .Y(n_297) );
AND2x4_ASAP7_75t_L g298 ( .A(n_253), .B(n_0), .Y(n_298) );
INVx3_ASAP7_75t_L g299 ( .A(n_253), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_207), .Y(n_300) );
NOR2x1_ASAP7_75t_L g301 ( .A(n_253), .B(n_1), .Y(n_301) );
BUFx6f_ASAP7_75t_L g302 ( .A(n_188), .Y(n_302) );
CKINVDCx5p33_ASAP7_75t_R g303 ( .A(n_277), .Y(n_303) );
BUFx6f_ASAP7_75t_L g304 ( .A(n_188), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_237), .B(n_1), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_205), .Y(n_306) );
AND2x2_ASAP7_75t_L g307 ( .A(n_195), .B(n_2), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_207), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_264), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_264), .Y(n_310) );
BUFx6f_ASAP7_75t_L g311 ( .A(n_188), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_205), .Y(n_312) );
AND2x2_ASAP7_75t_L g313 ( .A(n_195), .B(n_2), .Y(n_313) );
INVx3_ASAP7_75t_L g314 ( .A(n_206), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_222), .Y(n_315) );
BUFx6f_ASAP7_75t_L g316 ( .A(n_287), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_264), .Y(n_317) );
BUFx6f_ASAP7_75t_L g318 ( .A(n_287), .Y(n_318) );
INVxp67_ASAP7_75t_L g319 ( .A(n_213), .Y(n_319) );
INVx3_ASAP7_75t_L g320 ( .A(n_206), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_264), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_264), .Y(n_322) );
AND2x4_ASAP7_75t_L g323 ( .A(n_222), .B(n_3), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_264), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_226), .Y(n_325) );
BUFx6f_ASAP7_75t_L g326 ( .A(n_287), .Y(n_326) );
AOI22xp5_ASAP7_75t_L g327 ( .A1(n_221), .A2(n_5), .B1(n_3), .B2(n_4), .Y(n_327) );
AND2x4_ASAP7_75t_L g328 ( .A(n_293), .B(n_226), .Y(n_328) );
INVx3_ASAP7_75t_L g329 ( .A(n_296), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_309), .Y(n_330) );
BUFx12f_ASAP7_75t_L g331 ( .A(n_295), .Y(n_331) );
OAI22xp5_ASAP7_75t_L g332 ( .A1(n_327), .A2(n_209), .B1(n_278), .B2(n_221), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_309), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_309), .Y(n_334) );
NAND2x1p5_ASAP7_75t_L g335 ( .A(n_307), .B(n_187), .Y(n_335) );
NAND2x1p5_ASAP7_75t_L g336 ( .A(n_307), .B(n_189), .Y(n_336) );
AND2x2_ASAP7_75t_L g337 ( .A(n_319), .B(n_208), .Y(n_337) );
BUFx6f_ASAP7_75t_L g338 ( .A(n_292), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_310), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_292), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_310), .Y(n_341) );
AND2x2_ASAP7_75t_SL g342 ( .A(n_296), .B(n_228), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_307), .B(n_208), .Y(n_343) );
INVx4_ASAP7_75t_L g344 ( .A(n_296), .Y(n_344) );
INVx4_ASAP7_75t_L g345 ( .A(n_296), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_293), .B(n_231), .Y(n_346) );
OR2x2_ASAP7_75t_L g347 ( .A(n_305), .B(n_238), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_293), .B(n_190), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_310), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_317), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_293), .B(n_190), .Y(n_351) );
BUFx3_ASAP7_75t_L g352 ( .A(n_296), .Y(n_352) );
INVx5_ASAP7_75t_L g353 ( .A(n_299), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_317), .Y(n_354) );
AND2x2_ASAP7_75t_SL g355 ( .A(n_298), .B(n_313), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_292), .Y(n_356) );
BUFx10_ASAP7_75t_L g357 ( .A(n_303), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_292), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_321), .Y(n_359) );
INVx5_ASAP7_75t_L g360 ( .A(n_299), .Y(n_360) );
INVx3_ASAP7_75t_L g361 ( .A(n_298), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_299), .B(n_203), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_299), .B(n_255), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_321), .Y(n_364) );
INVx3_ASAP7_75t_L g365 ( .A(n_298), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_322), .Y(n_366) );
INVx2_ASAP7_75t_L g367 ( .A(n_344), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_344), .Y(n_368) );
INVx3_ASAP7_75t_L g369 ( .A(n_344), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_328), .Y(n_370) );
AND2x6_ASAP7_75t_L g371 ( .A(n_352), .B(n_298), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_355), .B(n_298), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_355), .B(n_323), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_355), .B(n_323), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_345), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_343), .B(n_320), .Y(n_376) );
AOI22xp5_ASAP7_75t_L g377 ( .A1(n_342), .A2(n_198), .B1(n_262), .B2(n_240), .Y(n_377) );
INVx3_ASAP7_75t_L g378 ( .A(n_345), .Y(n_378) );
NAND2xp5_ASAP7_75t_SL g379 ( .A(n_342), .B(n_197), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_328), .Y(n_380) );
AOI22xp5_ASAP7_75t_L g381 ( .A1(n_343), .A2(n_262), .B1(n_273), .B2(n_240), .Y(n_381) );
AND2x4_ASAP7_75t_L g382 ( .A(n_337), .B(n_327), .Y(n_382) );
BUFx6f_ASAP7_75t_L g383 ( .A(n_352), .Y(n_383) );
AOI22xp33_ASAP7_75t_L g384 ( .A1(n_352), .A2(n_300), .B1(n_308), .B2(n_294), .Y(n_384) );
INVxp67_ASAP7_75t_SL g385 ( .A(n_335), .Y(n_385) );
INVx5_ASAP7_75t_L g386 ( .A(n_345), .Y(n_386) );
BUFx3_ASAP7_75t_L g387 ( .A(n_331), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_363), .Y(n_388) );
AOI22xp33_ASAP7_75t_L g389 ( .A1(n_329), .A2(n_300), .B1(n_308), .B2(n_294), .Y(n_389) );
INVx3_ASAP7_75t_L g390 ( .A(n_329), .Y(n_390) );
BUFx3_ASAP7_75t_L g391 ( .A(n_331), .Y(n_391) );
OR2x2_ASAP7_75t_L g392 ( .A(n_347), .B(n_332), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_363), .B(n_320), .Y(n_393) );
NOR2xp33_ASAP7_75t_L g394 ( .A(n_346), .B(n_297), .Y(n_394) );
OAI22xp5_ASAP7_75t_SL g395 ( .A1(n_332), .A2(n_278), .B1(n_209), .B2(n_290), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_336), .Y(n_396) );
INVx2_ASAP7_75t_SL g397 ( .A(n_336), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_353), .Y(n_398) );
A2O1A1Ixp33_ASAP7_75t_L g399 ( .A1(n_329), .A2(n_300), .B(n_308), .C(n_294), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_353), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_329), .B(n_320), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_353), .Y(n_402) );
NAND2xp5_ASAP7_75t_SL g403 ( .A(n_336), .B(n_216), .Y(n_403) );
BUFx6f_ASAP7_75t_L g404 ( .A(n_353), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_361), .B(n_314), .Y(n_405) );
OR2x6_ASAP7_75t_L g406 ( .A(n_331), .B(n_301), .Y(n_406) );
INVx3_ASAP7_75t_L g407 ( .A(n_365), .Y(n_407) );
OR2x2_ASAP7_75t_L g408 ( .A(n_348), .B(n_256), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_330), .B(n_314), .Y(n_409) );
NAND2x1p5_ASAP7_75t_L g410 ( .A(n_353), .B(n_301), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_330), .B(n_322), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_351), .Y(n_412) );
BUFx6f_ASAP7_75t_L g413 ( .A(n_360), .Y(n_413) );
BUFx12f_ASAP7_75t_L g414 ( .A(n_357), .Y(n_414) );
NOR2xp33_ASAP7_75t_L g415 ( .A(n_357), .B(n_283), .Y(n_415) );
NAND2xp5_ASAP7_75t_SL g416 ( .A(n_360), .B(n_223), .Y(n_416) );
HB1xp67_ASAP7_75t_L g417 ( .A(n_362), .Y(n_417) );
BUFx8_ASAP7_75t_L g418 ( .A(n_333), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_362), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_360), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_360), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_333), .B(n_322), .Y(n_422) );
NAND2xp5_ASAP7_75t_SL g423 ( .A(n_360), .B(n_223), .Y(n_423) );
BUFx4f_ASAP7_75t_L g424 ( .A(n_334), .Y(n_424) );
BUFx6f_ASAP7_75t_L g425 ( .A(n_360), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_339), .Y(n_426) );
NAND2xp33_ASAP7_75t_L g427 ( .A(n_339), .B(n_264), .Y(n_427) );
NAND2x1p5_ASAP7_75t_L g428 ( .A(n_397), .B(n_306), .Y(n_428) );
NOR2xp33_ASAP7_75t_L g429 ( .A(n_388), .B(n_265), .Y(n_429) );
BUFx12f_ASAP7_75t_L g430 ( .A(n_418), .Y(n_430) );
OR2x2_ASAP7_75t_L g431 ( .A(n_392), .B(n_270), .Y(n_431) );
BUFx2_ASAP7_75t_L g432 ( .A(n_385), .Y(n_432) );
AOI21xp5_ASAP7_75t_L g433 ( .A1(n_401), .A2(n_349), .B(n_341), .Y(n_433) );
OAI21xp5_ASAP7_75t_L g434 ( .A1(n_372), .A2(n_349), .B(n_341), .Y(n_434) );
INVx3_ASAP7_75t_L g435 ( .A(n_386), .Y(n_435) );
AOI21x1_ASAP7_75t_L g436 ( .A1(n_405), .A2(n_354), .B(n_350), .Y(n_436) );
NOR2xp67_ASAP7_75t_L g437 ( .A(n_386), .B(n_56), .Y(n_437) );
O2A1O1Ixp33_ASAP7_75t_L g438 ( .A1(n_373), .A2(n_364), .B(n_366), .C(n_359), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_412), .B(n_364), .Y(n_439) );
NOR2xp33_ASAP7_75t_L g440 ( .A(n_382), .B(n_192), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_419), .B(n_366), .Y(n_441) );
OAI22xp5_ASAP7_75t_L g442 ( .A1(n_374), .A2(n_266), .B1(n_269), .B2(n_261), .Y(n_442) );
INVx2_ASAP7_75t_SL g443 ( .A(n_414), .Y(n_443) );
INVx3_ASAP7_75t_L g444 ( .A(n_386), .Y(n_444) );
BUFx6f_ASAP7_75t_L g445 ( .A(n_424), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_394), .B(n_324), .Y(n_446) );
INVx4_ASAP7_75t_L g447 ( .A(n_424), .Y(n_447) );
BUFx2_ASAP7_75t_L g448 ( .A(n_391), .Y(n_448) );
BUFx2_ASAP7_75t_L g449 ( .A(n_381), .Y(n_449) );
INVx3_ASAP7_75t_L g450 ( .A(n_383), .Y(n_450) );
BUFx2_ASAP7_75t_SL g451 ( .A(n_371), .Y(n_451) );
INVx4_ASAP7_75t_L g452 ( .A(n_371), .Y(n_452) );
INVx6_ASAP7_75t_L g453 ( .A(n_406), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_368), .Y(n_454) );
AOI21xp5_ASAP7_75t_L g455 ( .A1(n_376), .A2(n_258), .B(n_340), .Y(n_455) );
BUFx12f_ASAP7_75t_L g456 ( .A(n_406), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_393), .Y(n_457) );
BUFx6f_ASAP7_75t_L g458 ( .A(n_383), .Y(n_458) );
OAI22xp5_ASAP7_75t_L g459 ( .A1(n_377), .A2(n_284), .B1(n_288), .B2(n_285), .Y(n_459) );
AOI222xp33_ASAP7_75t_L g460 ( .A1(n_395), .A2(n_325), .B1(n_306), .B2(n_315), .C1(n_312), .C2(n_210), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_408), .B(n_260), .Y(n_461) );
AOI21x1_ASAP7_75t_L g462 ( .A1(n_411), .A2(n_356), .B(n_340), .Y(n_462) );
AND2x4_ASAP7_75t_L g463 ( .A(n_370), .B(n_241), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_393), .Y(n_464) );
OAI22xp5_ASAP7_75t_L g465 ( .A1(n_389), .A2(n_193), .B1(n_194), .B2(n_191), .Y(n_465) );
BUFx6f_ASAP7_75t_L g466 ( .A(n_404), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_375), .Y(n_467) );
INVx1_ASAP7_75t_SL g468 ( .A(n_371), .Y(n_468) );
BUFx6f_ASAP7_75t_L g469 ( .A(n_404), .Y(n_469) );
INVx3_ASAP7_75t_L g470 ( .A(n_369), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_390), .Y(n_471) );
INVx3_ASAP7_75t_L g472 ( .A(n_378), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_390), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_407), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_407), .Y(n_475) );
AOI21xp5_ASAP7_75t_L g476 ( .A1(n_411), .A2(n_358), .B(n_356), .Y(n_476) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_379), .A2(n_276), .B1(n_245), .B2(n_199), .Y(n_477) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_422), .A2(n_358), .B(n_200), .Y(n_478) );
A2O1A1Ixp33_ASAP7_75t_L g479 ( .A1(n_399), .A2(n_201), .B(n_202), .C(n_196), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_426), .Y(n_480) );
AO32x2_ASAP7_75t_L g481 ( .A1(n_427), .A2(n_292), .A3(n_311), .B1(n_304), .B2(n_302), .Y(n_481) );
BUFx6f_ASAP7_75t_L g482 ( .A(n_413), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_380), .Y(n_483) );
BUFx2_ASAP7_75t_L g484 ( .A(n_410), .Y(n_484) );
NAND3xp33_ASAP7_75t_L g485 ( .A(n_384), .B(n_276), .C(n_211), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_415), .B(n_263), .Y(n_486) );
CKINVDCx5p33_ASAP7_75t_R g487 ( .A(n_403), .Y(n_487) );
O2A1O1Ixp5_ASAP7_75t_L g488 ( .A1(n_416), .A2(n_204), .B(n_217), .C(n_203), .Y(n_488) );
A2O1A1Ixp33_ASAP7_75t_L g489 ( .A1(n_389), .A2(n_214), .B(n_219), .C(n_215), .Y(n_489) );
OR2x6_ASAP7_75t_L g490 ( .A(n_413), .B(n_276), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_422), .B(n_272), .Y(n_491) );
A2O1A1Ixp33_ASAP7_75t_SL g492 ( .A1(n_384), .A2(n_358), .B(n_217), .C(n_218), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_409), .B(n_274), .Y(n_493) );
NOR2x1_ASAP7_75t_SL g494 ( .A(n_425), .B(n_232), .Y(n_494) );
A2O1A1Ixp33_ASAP7_75t_L g495 ( .A1(n_409), .A2(n_229), .B(n_230), .C(n_220), .Y(n_495) );
OAI21xp33_ASAP7_75t_L g496 ( .A1(n_423), .A2(n_234), .B(n_233), .Y(n_496) );
A2O1A1Ixp33_ASAP7_75t_L g497 ( .A1(n_420), .A2(n_236), .B(n_239), .C(n_235), .Y(n_497) );
BUFx6f_ASAP7_75t_L g498 ( .A(n_425), .Y(n_498) );
INVx1_ASAP7_75t_SL g499 ( .A(n_425), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_421), .B(n_274), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_398), .Y(n_501) );
INVx3_ASAP7_75t_L g502 ( .A(n_400), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_402), .B(n_275), .Y(n_503) );
OR2x4_ASAP7_75t_L g504 ( .A(n_392), .B(n_276), .Y(n_504) );
AO22x1_ASAP7_75t_L g505 ( .A1(n_418), .A2(n_212), .B1(n_227), .B2(n_224), .Y(n_505) );
AOI21x1_ASAP7_75t_L g506 ( .A1(n_405), .A2(n_244), .B(n_242), .Y(n_506) );
INVx1_ASAP7_75t_SL g507 ( .A(n_417), .Y(n_507) );
AND2x6_ASAP7_75t_L g508 ( .A(n_396), .B(n_246), .Y(n_508) );
INVx2_ASAP7_75t_L g509 ( .A(n_367), .Y(n_509) );
BUFx6f_ASAP7_75t_SL g510 ( .A(n_387), .Y(n_510) );
AO32x2_ASAP7_75t_L g511 ( .A1(n_465), .A2(n_302), .A3(n_318), .B1(n_316), .B2(n_311), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_507), .Y(n_512) );
BUFx6f_ASAP7_75t_L g513 ( .A(n_466), .Y(n_513) );
AOI21x1_ASAP7_75t_L g514 ( .A1(n_506), .A2(n_247), .B(n_243), .Y(n_514) );
AO32x2_ASAP7_75t_L g515 ( .A1(n_465), .A2(n_302), .A3(n_318), .B1(n_316), .B2(n_311), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_449), .A2(n_249), .B1(n_251), .B2(n_248), .Y(n_516) );
OAI21x1_ASAP7_75t_L g517 ( .A1(n_462), .A2(n_247), .B(n_243), .Y(n_517) );
AOI21x1_ASAP7_75t_L g518 ( .A1(n_436), .A2(n_254), .B(n_250), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_428), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_478), .A2(n_268), .B(n_257), .Y(n_520) );
AO21x2_ASAP7_75t_L g521 ( .A1(n_492), .A2(n_259), .B(n_252), .Y(n_521) );
INVx1_ASAP7_75t_SL g522 ( .A(n_432), .Y(n_522) );
OA21x2_ASAP7_75t_L g523 ( .A1(n_476), .A2(n_268), .B(n_257), .Y(n_523) );
INVx6_ASAP7_75t_L g524 ( .A(n_430), .Y(n_524) );
OAI21xp5_ASAP7_75t_L g525 ( .A1(n_433), .A2(n_271), .B(n_267), .Y(n_525) );
OAI21x1_ASAP7_75t_L g526 ( .A1(n_437), .A2(n_280), .B(n_279), .Y(n_526) );
OR2x6_ASAP7_75t_L g527 ( .A(n_451), .B(n_281), .Y(n_527) );
OA21x2_ASAP7_75t_L g528 ( .A1(n_488), .A2(n_286), .B(n_282), .Y(n_528) );
OA21x2_ASAP7_75t_L g529 ( .A1(n_479), .A2(n_291), .B(n_289), .Y(n_529) );
BUFx8_ASAP7_75t_L g530 ( .A(n_510), .Y(n_530) );
INVx2_ASAP7_75t_L g531 ( .A(n_480), .Y(n_531) );
AO21x2_ASAP7_75t_L g532 ( .A1(n_485), .A2(n_302), .B(n_292), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_440), .A2(n_292), .B1(n_304), .B2(n_302), .Y(n_533) );
INVx3_ASAP7_75t_L g534 ( .A(n_452), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_457), .B(n_6), .Y(n_535) );
OAI21x1_ASAP7_75t_L g536 ( .A1(n_437), .A2(n_304), .B(n_302), .Y(n_536) );
OA21x2_ASAP7_75t_L g537 ( .A1(n_496), .A2(n_455), .B(n_489), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_460), .B(n_8), .Y(n_538) );
NAND3xp33_ASAP7_75t_L g539 ( .A(n_495), .B(n_311), .C(n_304), .Y(n_539) );
NAND2xp33_ASAP7_75t_SL g540 ( .A(n_445), .B(n_8), .Y(n_540) );
AOI22xp5_ASAP7_75t_L g541 ( .A1(n_429), .A2(n_311), .B1(n_316), .B2(n_304), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g542 ( .A1(n_459), .A2(n_311), .B1(n_316), .B2(n_304), .Y(n_542) );
OAI22xp5_ASAP7_75t_L g543 ( .A1(n_504), .A2(n_441), .B1(n_439), .B2(n_464), .Y(n_543) );
INVx4_ASAP7_75t_L g544 ( .A(n_445), .Y(n_544) );
BUFx6f_ASAP7_75t_L g545 ( .A(n_466), .Y(n_545) );
AO21x2_ASAP7_75t_L g546 ( .A1(n_494), .A2(n_326), .B(n_318), .Y(n_546) );
NAND3xp33_ASAP7_75t_L g547 ( .A(n_497), .B(n_326), .C(n_318), .Y(n_547) );
OAI21xp5_ASAP7_75t_L g548 ( .A1(n_438), .A2(n_326), .B(n_318), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_483), .Y(n_549) );
OA21x2_ASAP7_75t_L g550 ( .A1(n_496), .A2(n_326), .B(n_338), .Y(n_550) );
OAI21x1_ASAP7_75t_L g551 ( .A1(n_450), .A2(n_326), .B(n_338), .Y(n_551) );
INVx6_ASAP7_75t_L g552 ( .A(n_456), .Y(n_552) );
BUFx2_ASAP7_75t_SL g553 ( .A(n_443), .Y(n_553) );
NAND2x1p5_ASAP7_75t_L g554 ( .A(n_447), .B(n_9), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_431), .B(n_10), .Y(n_555) );
INVx2_ASAP7_75t_L g556 ( .A(n_454), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_463), .Y(n_557) );
BUFx8_ASAP7_75t_L g558 ( .A(n_448), .Y(n_558) );
INVx2_ASAP7_75t_L g559 ( .A(n_467), .Y(n_559) );
AO21x2_ASAP7_75t_L g560 ( .A1(n_446), .A2(n_338), .B(n_62), .Y(n_560) );
OAI22xp5_ASAP7_75t_L g561 ( .A1(n_434), .A2(n_12), .B1(n_13), .B2(n_15), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_491), .B(n_16), .Y(n_562) );
INVx2_ASAP7_75t_L g563 ( .A(n_509), .Y(n_563) );
NAND2xp33_ASAP7_75t_SL g564 ( .A(n_445), .B(n_18), .Y(n_564) );
OA21x2_ASAP7_75t_L g565 ( .A1(n_500), .A2(n_69), .B(n_68), .Y(n_565) );
OAI21x1_ASAP7_75t_L g566 ( .A1(n_502), .A2(n_71), .B(n_70), .Y(n_566) );
OAI21x1_ASAP7_75t_SL g567 ( .A1(n_447), .A2(n_18), .B(n_19), .Y(n_567) );
BUFx6f_ASAP7_75t_L g568 ( .A(n_466), .Y(n_568) );
OAI21x1_ASAP7_75t_L g569 ( .A1(n_435), .A2(n_75), .B(n_73), .Y(n_569) );
OAI21x1_ASAP7_75t_L g570 ( .A1(n_444), .A2(n_79), .B(n_77), .Y(n_570) );
NOR2xp33_ASAP7_75t_SL g571 ( .A(n_468), .B(n_82), .Y(n_571) );
OAI21x1_ASAP7_75t_L g572 ( .A1(n_444), .A2(n_84), .B(n_83), .Y(n_572) );
AOI21xp5_ASAP7_75t_L g573 ( .A1(n_493), .A2(n_87), .B(n_86), .Y(n_573) );
INVxp67_ASAP7_75t_SL g574 ( .A(n_458), .Y(n_574) );
INVx1_ASAP7_75t_SL g575 ( .A(n_499), .Y(n_575) );
BUFx10_ASAP7_75t_L g576 ( .A(n_453), .Y(n_576) );
OAI21x1_ASAP7_75t_L g577 ( .A1(n_471), .A2(n_89), .B(n_88), .Y(n_577) );
OR2x6_ASAP7_75t_L g578 ( .A(n_505), .B(n_21), .Y(n_578) );
OAI21x1_ASAP7_75t_L g579 ( .A1(n_501), .A2(n_91), .B(n_90), .Y(n_579) );
OAI22xp33_ASAP7_75t_L g580 ( .A1(n_461), .A2(n_22), .B1(n_23), .B2(n_24), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_442), .Y(n_581) );
OAI22xp5_ASAP7_75t_L g582 ( .A1(n_490), .A2(n_25), .B1(n_27), .B2(n_28), .Y(n_582) );
OA21x2_ASAP7_75t_L g583 ( .A1(n_477), .A2(n_95), .B(n_92), .Y(n_583) );
BUFx3_ASAP7_75t_L g584 ( .A(n_484), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_503), .Y(n_585) );
OAI21x1_ASAP7_75t_L g586 ( .A1(n_473), .A2(n_97), .B(n_96), .Y(n_586) );
HB1xp67_ASAP7_75t_L g587 ( .A(n_490), .Y(n_587) );
INVx2_ASAP7_75t_SL g588 ( .A(n_487), .Y(n_588) );
OAI21x1_ASAP7_75t_L g589 ( .A1(n_474), .A2(n_99), .B(n_98), .Y(n_589) );
AO31x2_ASAP7_75t_L g590 ( .A1(n_475), .A2(n_29), .A3(n_30), .B(n_31), .Y(n_590) );
OAI22xp5_ASAP7_75t_L g591 ( .A1(n_490), .A2(n_31), .B1(n_32), .B2(n_33), .Y(n_591) );
OR2x2_ASAP7_75t_L g592 ( .A(n_486), .B(n_32), .Y(n_592) );
OAI21x1_ASAP7_75t_L g593 ( .A1(n_536), .A2(n_472), .B(n_470), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_538), .B(n_508), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_512), .B(n_33), .Y(n_595) );
OAI22xp5_ASAP7_75t_L g596 ( .A1(n_543), .A2(n_498), .B1(n_482), .B2(n_469), .Y(n_596) );
OA21x2_ASAP7_75t_L g597 ( .A1(n_517), .A2(n_481), .B(n_129), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_581), .B(n_34), .Y(n_598) );
BUFx3_ASAP7_75t_L g599 ( .A(n_558), .Y(n_599) );
HB1xp67_ASAP7_75t_L g600 ( .A(n_522), .Y(n_600) );
OAI22xp5_ASAP7_75t_L g601 ( .A1(n_527), .A2(n_37), .B1(n_38), .B2(n_39), .Y(n_601) );
AND2x2_ASAP7_75t_L g602 ( .A(n_555), .B(n_38), .Y(n_602) );
INVx2_ASAP7_75t_L g603 ( .A(n_531), .Y(n_603) );
AOI22xp33_ASAP7_75t_SL g604 ( .A1(n_578), .A2(n_39), .B1(n_40), .B2(n_41), .Y(n_604) );
OAI211xp5_ASAP7_75t_SL g605 ( .A1(n_516), .A2(n_42), .B(n_45), .C(n_46), .Y(n_605) );
OAI211xp5_ASAP7_75t_SL g606 ( .A1(n_557), .A2(n_47), .B(n_49), .C(n_50), .Y(n_606) );
AO21x2_ASAP7_75t_L g607 ( .A1(n_548), .A2(n_144), .B(n_182), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_535), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_535), .Y(n_609) );
AOI21x1_ASAP7_75t_L g610 ( .A1(n_518), .A2(n_101), .B(n_103), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_585), .B(n_104), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_554), .Y(n_612) );
AOI22xp33_ASAP7_75t_SL g613 ( .A1(n_578), .A2(n_106), .B1(n_107), .B2(n_111), .Y(n_613) );
BUFx10_ASAP7_75t_L g614 ( .A(n_524), .Y(n_614) );
AOI211xp5_ASAP7_75t_L g615 ( .A1(n_561), .A2(n_591), .B(n_582), .C(n_580), .Y(n_615) );
BUFx2_ASAP7_75t_L g616 ( .A(n_584), .Y(n_616) );
INVx3_ASAP7_75t_L g617 ( .A(n_519), .Y(n_617) );
OR2x2_ASAP7_75t_L g618 ( .A(n_592), .B(n_127), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_549), .B(n_136), .Y(n_619) );
AND2x2_ASAP7_75t_L g620 ( .A(n_578), .B(n_147), .Y(n_620) );
OR2x2_ASAP7_75t_L g621 ( .A(n_553), .B(n_154), .Y(n_621) );
AOI22xp33_ASAP7_75t_SL g622 ( .A1(n_582), .A2(n_155), .B1(n_156), .B2(n_159), .Y(n_622) );
OR2x2_ASAP7_75t_L g623 ( .A(n_588), .B(n_161), .Y(n_623) );
AO21x2_ASAP7_75t_L g624 ( .A1(n_514), .A2(n_162), .B(n_163), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_561), .Y(n_625) );
AOI22xp5_ASAP7_75t_L g626 ( .A1(n_562), .A2(n_166), .B1(n_168), .B2(n_169), .Y(n_626) );
OR2x6_ASAP7_75t_L g627 ( .A(n_524), .B(n_170), .Y(n_627) );
OAI21x1_ASAP7_75t_L g628 ( .A1(n_551), .A2(n_171), .B(n_173), .Y(n_628) );
INVx2_ASAP7_75t_SL g629 ( .A(n_530), .Y(n_629) );
HB1xp67_ASAP7_75t_L g630 ( .A(n_575), .Y(n_630) );
INVx1_ASAP7_75t_SL g631 ( .A(n_587), .Y(n_631) );
INVx2_ASAP7_75t_L g632 ( .A(n_556), .Y(n_632) );
AOI22xp5_ASAP7_75t_L g633 ( .A1(n_552), .A2(n_591), .B1(n_540), .B2(n_564), .Y(n_633) );
AOI21xp5_ASAP7_75t_L g634 ( .A1(n_573), .A2(n_525), .B(n_523), .Y(n_634) );
OR2x6_ASAP7_75t_L g635 ( .A(n_552), .B(n_544), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_590), .Y(n_636) );
AOI21xp5_ASAP7_75t_L g637 ( .A1(n_523), .A2(n_520), .B(n_550), .Y(n_637) );
OAI22xp5_ASAP7_75t_L g638 ( .A1(n_539), .A2(n_547), .B1(n_529), .B2(n_541), .Y(n_638) );
OAI22xp33_ASAP7_75t_L g639 ( .A1(n_571), .A2(n_534), .B1(n_544), .B2(n_559), .Y(n_639) );
AOI22xp33_ASAP7_75t_SL g640 ( .A1(n_567), .A2(n_571), .B1(n_565), .B2(n_583), .Y(n_640) );
HB1xp67_ASAP7_75t_L g641 ( .A(n_563), .Y(n_641) );
AOI22xp33_ASAP7_75t_L g642 ( .A1(n_533), .A2(n_537), .B1(n_542), .B2(n_576), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_537), .B(n_520), .Y(n_643) );
OAI22xp33_ASAP7_75t_L g644 ( .A1(n_565), .A2(n_583), .B1(n_574), .B2(n_545), .Y(n_644) );
OAI22xp33_ASAP7_75t_L g645 ( .A1(n_574), .A2(n_568), .B1(n_513), .B2(n_545), .Y(n_645) );
OA21x2_ASAP7_75t_L g646 ( .A1(n_526), .A2(n_586), .B(n_589), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_513), .B(n_568), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_590), .Y(n_648) );
AND2x2_ASAP7_75t_L g649 ( .A(n_603), .B(n_511), .Y(n_649) );
A2O1A1Ixp33_ASAP7_75t_L g650 ( .A1(n_615), .A2(n_572), .B(n_570), .C(n_569), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_636), .Y(n_651) );
AND2x2_ASAP7_75t_L g652 ( .A(n_632), .B(n_515), .Y(n_652) );
OR2x2_ASAP7_75t_L g653 ( .A(n_600), .B(n_521), .Y(n_653) );
NOR2x1_ASAP7_75t_L g654 ( .A(n_627), .B(n_546), .Y(n_654) );
AND2x4_ASAP7_75t_L g655 ( .A(n_612), .B(n_566), .Y(n_655) );
AND2x2_ASAP7_75t_L g656 ( .A(n_608), .B(n_528), .Y(n_656) );
BUFx2_ASAP7_75t_L g657 ( .A(n_596), .Y(n_657) );
AND2x2_ASAP7_75t_L g658 ( .A(n_609), .B(n_577), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_648), .Y(n_659) );
AND2x2_ASAP7_75t_L g660 ( .A(n_641), .B(n_579), .Y(n_660) );
BUFx3_ASAP7_75t_L g661 ( .A(n_616), .Y(n_661) );
INVx2_ASAP7_75t_L g662 ( .A(n_643), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_625), .Y(n_663) );
INVx2_ASAP7_75t_L g664 ( .A(n_643), .Y(n_664) );
AND2x4_ASAP7_75t_L g665 ( .A(n_617), .B(n_560), .Y(n_665) );
AND2x2_ASAP7_75t_L g666 ( .A(n_617), .B(n_532), .Y(n_666) );
INVxp67_ASAP7_75t_L g667 ( .A(n_630), .Y(n_667) );
INVx2_ASAP7_75t_L g668 ( .A(n_593), .Y(n_668) );
AND2x2_ASAP7_75t_L g669 ( .A(n_594), .B(n_620), .Y(n_669) );
AND2x2_ASAP7_75t_L g670 ( .A(n_595), .B(n_598), .Y(n_670) );
INVx2_ASAP7_75t_SL g671 ( .A(n_635), .Y(n_671) );
OR2x2_ASAP7_75t_L g672 ( .A(n_631), .B(n_618), .Y(n_672) );
BUFx3_ASAP7_75t_L g673 ( .A(n_635), .Y(n_673) );
AND2x2_ASAP7_75t_L g674 ( .A(n_601), .B(n_627), .Y(n_674) );
INVx2_ASAP7_75t_L g675 ( .A(n_597), .Y(n_675) );
AND2x2_ASAP7_75t_L g676 ( .A(n_602), .B(n_604), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_623), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_621), .Y(n_678) );
INVx1_ASAP7_75t_SL g679 ( .A(n_599), .Y(n_679) );
BUFx3_ASAP7_75t_L g680 ( .A(n_614), .Y(n_680) );
INVx2_ASAP7_75t_L g681 ( .A(n_597), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_619), .Y(n_682) );
NOR2xp33_ASAP7_75t_L g683 ( .A(n_633), .B(n_629), .Y(n_683) );
AO21x2_ASAP7_75t_L g684 ( .A1(n_637), .A2(n_644), .B(n_634), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_619), .Y(n_685) );
INVx3_ASAP7_75t_L g686 ( .A(n_647), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_611), .Y(n_687) );
INVx2_ASAP7_75t_L g688 ( .A(n_628), .Y(n_688) );
BUFx6f_ASAP7_75t_L g689 ( .A(n_646), .Y(n_689) );
INVx3_ASAP7_75t_L g690 ( .A(n_607), .Y(n_690) );
INVx2_ASAP7_75t_L g691 ( .A(n_646), .Y(n_691) );
INVx2_ASAP7_75t_L g692 ( .A(n_624), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_606), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_605), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_607), .Y(n_695) );
AND2x4_ASAP7_75t_L g696 ( .A(n_663), .B(n_624), .Y(n_696) );
INVx3_ASAP7_75t_L g697 ( .A(n_655), .Y(n_697) );
NAND3xp33_ASAP7_75t_L g698 ( .A(n_683), .B(n_613), .C(n_622), .Y(n_698) );
INVx2_ASAP7_75t_SL g699 ( .A(n_661), .Y(n_699) );
INVx4_ASAP7_75t_L g700 ( .A(n_673), .Y(n_700) );
AOI21xp5_ASAP7_75t_L g701 ( .A1(n_650), .A2(n_639), .B(n_640), .Y(n_701) );
BUFx3_ASAP7_75t_L g702 ( .A(n_680), .Y(n_702) );
AND2x2_ASAP7_75t_L g703 ( .A(n_663), .B(n_638), .Y(n_703) );
INVx2_ASAP7_75t_L g704 ( .A(n_691), .Y(n_704) );
INVx2_ASAP7_75t_L g705 ( .A(n_691), .Y(n_705) );
AND2x2_ASAP7_75t_L g706 ( .A(n_669), .B(n_642), .Y(n_706) );
OR2x2_ASAP7_75t_L g707 ( .A(n_672), .B(n_638), .Y(n_707) );
INVx3_ASAP7_75t_L g708 ( .A(n_655), .Y(n_708) );
INVx3_ASAP7_75t_L g709 ( .A(n_655), .Y(n_709) );
INVx2_ASAP7_75t_L g710 ( .A(n_662), .Y(n_710) );
AND2x4_ASAP7_75t_L g711 ( .A(n_651), .B(n_626), .Y(n_711) );
AOI33xp33_ASAP7_75t_L g712 ( .A1(n_679), .A2(n_677), .A3(n_674), .B1(n_678), .B2(n_676), .B3(n_670), .Y(n_712) );
INVxp67_ASAP7_75t_SL g713 ( .A(n_654), .Y(n_713) );
OR2x2_ASAP7_75t_L g714 ( .A(n_667), .B(n_645), .Y(n_714) );
HB1xp67_ASAP7_75t_L g715 ( .A(n_662), .Y(n_715) );
HB1xp67_ASAP7_75t_L g716 ( .A(n_664), .Y(n_716) );
OAI21xp5_ASAP7_75t_L g717 ( .A1(n_693), .A2(n_610), .B(n_694), .Y(n_717) );
HB1xp67_ASAP7_75t_L g718 ( .A(n_664), .Y(n_718) );
NOR2x1_ASAP7_75t_SL g719 ( .A(n_671), .B(n_680), .Y(n_719) );
INVx3_ASAP7_75t_L g720 ( .A(n_665), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_659), .Y(n_721) );
INVx1_ASAP7_75t_L g722 ( .A(n_653), .Y(n_722) );
AND2x4_ASAP7_75t_L g723 ( .A(n_666), .B(n_686), .Y(n_723) );
AND2x2_ASAP7_75t_L g724 ( .A(n_686), .B(n_656), .Y(n_724) );
AO221x2_ASAP7_75t_L g725 ( .A1(n_695), .A2(n_675), .B1(n_681), .B2(n_687), .C(n_682), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_721), .Y(n_726) );
AO21x2_ASAP7_75t_L g727 ( .A1(n_717), .A2(n_692), .B(n_695), .Y(n_727) );
AND2x2_ASAP7_75t_L g728 ( .A(n_724), .B(n_657), .Y(n_728) );
INVx2_ASAP7_75t_SL g729 ( .A(n_699), .Y(n_729) );
INVx2_ASAP7_75t_L g730 ( .A(n_704), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_710), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_710), .Y(n_732) );
INVx1_ASAP7_75t_L g733 ( .A(n_715), .Y(n_733) );
AND2x4_ASAP7_75t_L g734 ( .A(n_697), .B(n_665), .Y(n_734) );
AND2x4_ASAP7_75t_L g735 ( .A(n_697), .B(n_665), .Y(n_735) );
INVx2_ASAP7_75t_L g736 ( .A(n_704), .Y(n_736) );
AOI211x1_ASAP7_75t_L g737 ( .A1(n_698), .A2(n_658), .B(n_660), .C(n_685), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_716), .Y(n_738) );
AND2x2_ASAP7_75t_L g739 ( .A(n_703), .B(n_649), .Y(n_739) );
AND2x2_ASAP7_75t_L g740 ( .A(n_703), .B(n_652), .Y(n_740) );
INVx6_ASAP7_75t_L g741 ( .A(n_702), .Y(n_741) );
INVx3_ASAP7_75t_L g742 ( .A(n_725), .Y(n_742) );
AND2x2_ASAP7_75t_L g743 ( .A(n_723), .B(n_684), .Y(n_743) );
INVx1_ASAP7_75t_L g744 ( .A(n_718), .Y(n_744) );
AND2x2_ASAP7_75t_L g745 ( .A(n_723), .B(n_684), .Y(n_745) );
OR2x2_ASAP7_75t_L g746 ( .A(n_707), .B(n_689), .Y(n_746) );
AND2x2_ASAP7_75t_L g747 ( .A(n_706), .B(n_689), .Y(n_747) );
AND3x1_ASAP7_75t_L g748 ( .A(n_712), .B(n_690), .C(n_681), .Y(n_748) );
OR2x2_ASAP7_75t_L g749 ( .A(n_722), .B(n_689), .Y(n_749) );
INVx2_ASAP7_75t_L g750 ( .A(n_705), .Y(n_750) );
AND2x4_ASAP7_75t_L g751 ( .A(n_697), .B(n_668), .Y(n_751) );
INVx1_ASAP7_75t_SL g752 ( .A(n_699), .Y(n_752) );
OR2x6_ASAP7_75t_L g753 ( .A(n_742), .B(n_708), .Y(n_753) );
AND2x2_ASAP7_75t_L g754 ( .A(n_739), .B(n_720), .Y(n_754) );
INVx2_ASAP7_75t_L g755 ( .A(n_730), .Y(n_755) );
NAND2x1_ASAP7_75t_L g756 ( .A(n_741), .B(n_742), .Y(n_756) );
AND2x2_ASAP7_75t_L g757 ( .A(n_740), .B(n_720), .Y(n_757) );
OR2x2_ASAP7_75t_L g758 ( .A(n_733), .B(n_709), .Y(n_758) );
AND2x2_ASAP7_75t_L g759 ( .A(n_747), .B(n_709), .Y(n_759) );
AND2x2_ASAP7_75t_L g760 ( .A(n_747), .B(n_709), .Y(n_760) );
OR2x6_ASAP7_75t_L g761 ( .A(n_742), .B(n_737), .Y(n_761) );
AND2x4_ASAP7_75t_L g762 ( .A(n_743), .B(n_713), .Y(n_762) );
CKINVDCx20_ASAP7_75t_R g763 ( .A(n_741), .Y(n_763) );
NAND2x1p5_ASAP7_75t_L g764 ( .A(n_748), .B(n_700), .Y(n_764) );
INVx2_ASAP7_75t_L g765 ( .A(n_730), .Y(n_765) );
INVx1_ASAP7_75t_L g766 ( .A(n_726), .Y(n_766) );
INVx2_ASAP7_75t_SL g767 ( .A(n_763), .Y(n_767) );
OAI222xp33_ASAP7_75t_L g768 ( .A1(n_761), .A2(n_752), .B1(n_729), .B2(n_745), .C1(n_743), .C2(n_728), .Y(n_768) );
INVx1_ASAP7_75t_L g769 ( .A(n_766), .Y(n_769) );
AOI31xp33_ASAP7_75t_L g770 ( .A1(n_764), .A2(n_719), .A3(n_714), .B(n_701), .Y(n_770) );
AND2x4_ASAP7_75t_L g771 ( .A(n_767), .B(n_753), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_769), .Y(n_772) );
O2A1O1Ixp33_ASAP7_75t_L g773 ( .A1(n_770), .A2(n_761), .B(n_756), .C(n_753), .Y(n_773) );
INVx1_ASAP7_75t_L g774 ( .A(n_772), .Y(n_774) );
AOI21xp5_ASAP7_75t_L g775 ( .A1(n_773), .A2(n_768), .B(n_756), .Y(n_775) );
AOI22xp33_ASAP7_75t_SL g776 ( .A1(n_771), .A2(n_762), .B1(n_757), .B2(n_754), .Y(n_776) );
AOI221xp5_ASAP7_75t_L g777 ( .A1(n_775), .A2(n_759), .B1(n_760), .B2(n_738), .C(n_744), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_774), .B(n_758), .Y(n_778) );
INVx1_ASAP7_75t_L g779 ( .A(n_778), .Y(n_779) );
OAI31xp33_ASAP7_75t_L g780 ( .A1(n_777), .A2(n_711), .A3(n_776), .B(n_696), .Y(n_780) );
INVx2_ASAP7_75t_L g781 ( .A(n_779), .Y(n_781) );
NAND3xp33_ASAP7_75t_SL g782 ( .A(n_780), .B(n_746), .C(n_749), .Y(n_782) );
BUFx8_ASAP7_75t_L g783 ( .A(n_781), .Y(n_783) );
OAI22xp5_ASAP7_75t_L g784 ( .A1(n_782), .A2(n_746), .B1(n_734), .B2(n_735), .Y(n_784) );
AOI21xp5_ASAP7_75t_L g785 ( .A1(n_783), .A2(n_711), .B(n_692), .Y(n_785) );
AOI222xp33_ASAP7_75t_SL g786 ( .A1(n_785), .A2(n_784), .B1(n_765), .B2(n_755), .C1(n_731), .C2(n_732), .Y(n_786) );
AOI22xp33_ASAP7_75t_L g787 ( .A1(n_786), .A2(n_751), .B1(n_727), .B2(n_732), .Y(n_787) );
OAI22xp33_ASAP7_75t_L g788 ( .A1(n_787), .A2(n_688), .B1(n_736), .B2(n_750), .Y(n_788) );
AOI21xp5_ASAP7_75t_L g789 ( .A1(n_788), .A2(n_688), .B(n_668), .Y(n_789) );
endmodule