module fake_netlist_6_3887_n_1748 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1748);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1748;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_297;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1736;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_535;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_82),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_24),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_25),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_40),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_28),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_142),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_106),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_134),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_120),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_23),
.Y(n_164)
);

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_91),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_87),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_74),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_78),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_124),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_98),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_131),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_24),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_153),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_39),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_84),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_99),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_34),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_83),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_39),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_17),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_19),
.Y(n_181)
);

INVx2_ASAP7_75t_SL g182 ( 
.A(n_72),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_107),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_13),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_123),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_69),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_19),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_148),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_15),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_108),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_49),
.Y(n_191)
);

BUFx5_ASAP7_75t_L g192 ( 
.A(n_96),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_56),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_73),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_16),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_130),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_152),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_117),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_149),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_147),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_125),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_64),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_71),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_55),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_128),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_5),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_150),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_30),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_41),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_16),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_65),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_100),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_101),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_89),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_68),
.Y(n_215)
);

INVx2_ASAP7_75t_SL g216 ( 
.A(n_22),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_94),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_42),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_116),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_132),
.Y(n_220)
);

INVx4_ASAP7_75t_R g221 ( 
.A(n_53),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_6),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_102),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_14),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_10),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_32),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_6),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_112),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_85),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_141),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_9),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_97),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_38),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_66),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_46),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_145),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_77),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_45),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_86),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_103),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_17),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_45),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_59),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_51),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_88),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_140),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_21),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_137),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_151),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_51),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_34),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_43),
.Y(n_252)
);

INVxp33_ASAP7_75t_SL g253 ( 
.A(n_15),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_75),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_129),
.Y(n_255)
);

CKINVDCx14_ASAP7_75t_R g256 ( 
.A(n_58),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_18),
.Y(n_257)
);

BUFx10_ASAP7_75t_L g258 ( 
.A(n_63),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_115),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_13),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_76),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_146),
.Y(n_262)
);

BUFx10_ASAP7_75t_L g263 ( 
.A(n_18),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_44),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_122),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_11),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_23),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_144),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_2),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_40),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_5),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_95),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_105),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_143),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_20),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_20),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_53),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_119),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_7),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_25),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_11),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_118),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_48),
.Y(n_283)
);

BUFx10_ASAP7_75t_L g284 ( 
.A(n_37),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_121),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_8),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g287 ( 
.A(n_33),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_139),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_50),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_60),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_28),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_4),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_32),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_9),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_67),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_7),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_10),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_4),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_0),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_104),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_57),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_50),
.Y(n_302)
);

INVx1_ASAP7_75t_SL g303 ( 
.A(n_70),
.Y(n_303)
);

BUFx10_ASAP7_75t_L g304 ( 
.A(n_127),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_54),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_79),
.Y(n_306)
);

INVx1_ASAP7_75t_SL g307 ( 
.A(n_113),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_257),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_203),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_246),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_190),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_206),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_193),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_194),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_165),
.B(n_0),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_257),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_257),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_263),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_257),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_199),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_257),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_184),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_201),
.Y(n_323)
);

BUFx2_ASAP7_75t_L g324 ( 
.A(n_157),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_207),
.Y(n_325)
);

NOR2xp67_ASAP7_75t_L g326 ( 
.A(n_216),
.B(n_1),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_184),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_192),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_244),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_249),
.Y(n_330)
);

INVx1_ASAP7_75t_SL g331 ( 
.A(n_189),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_157),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_211),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_288),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_301),
.Y(n_335)
);

INVxp67_ASAP7_75t_SL g336 ( 
.A(n_161),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_244),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_156),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_182),
.B(n_1),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_159),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_263),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_182),
.B(n_2),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_306),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_202),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_214),
.Y(n_345)
);

INVxp67_ASAP7_75t_SL g346 ( 
.A(n_162),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_164),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_205),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_219),
.Y(n_349)
);

NOR2xp67_ASAP7_75t_L g350 ( 
.A(n_216),
.B(n_3),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_180),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_263),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_220),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_228),
.Y(n_354)
);

BUFx2_ASAP7_75t_L g355 ( 
.A(n_172),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_234),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_208),
.Y(n_357)
);

INVxp33_ASAP7_75t_SL g358 ( 
.A(n_172),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_215),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_200),
.B(n_3),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_200),
.B(n_8),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_236),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_209),
.Y(n_363)
);

NOR2xp67_ASAP7_75t_L g364 ( 
.A(n_279),
.B(n_12),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_239),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_232),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_284),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_245),
.Y(n_368)
);

BUFx3_ASAP7_75t_L g369 ( 
.A(n_168),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_253),
.B(n_12),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_254),
.Y(n_371)
);

INVxp67_ASAP7_75t_SL g372 ( 
.A(n_176),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_222),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_225),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_255),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_226),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_256),
.Y(n_377)
);

INVxp67_ASAP7_75t_SL g378 ( 
.A(n_186),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_261),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_284),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_265),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_233),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_238),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_308),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_328),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_328),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_331),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_308),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_328),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_316),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_SL g391 ( 
.A(n_331),
.B(n_284),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_316),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_317),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_317),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_319),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_319),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_336),
.B(n_212),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_321),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_346),
.B(n_155),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_321),
.Y(n_400)
);

AND2x4_ASAP7_75t_L g401 ( 
.A(n_369),
.B(n_212),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_322),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_322),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_309),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_372),
.B(n_155),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_327),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_369),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_327),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_329),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_369),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_329),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_378),
.B(n_160),
.Y(n_412)
);

AND2x4_ASAP7_75t_L g413 ( 
.A(n_360),
.B(n_223),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_337),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_337),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g416 ( 
.A(n_332),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_361),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_338),
.Y(n_418)
);

AND2x2_ASAP7_75t_SL g419 ( 
.A(n_342),
.B(n_223),
.Y(n_419)
);

AND2x4_ASAP7_75t_L g420 ( 
.A(n_326),
.B(n_240),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_338),
.B(n_240),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_340),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_383),
.B(n_272),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_340),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_347),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_347),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_342),
.B(n_204),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_339),
.B(n_160),
.Y(n_428)
);

INVx3_ASAP7_75t_L g429 ( 
.A(n_351),
.Y(n_429)
);

INVx3_ASAP7_75t_L g430 ( 
.A(n_351),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_357),
.Y(n_431)
);

BUFx2_ASAP7_75t_L g432 ( 
.A(n_318),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_357),
.Y(n_433)
);

INVx5_ASAP7_75t_L g434 ( 
.A(n_324),
.Y(n_434)
);

INVx3_ASAP7_75t_L g435 ( 
.A(n_363),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_363),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_373),
.Y(n_437)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_373),
.Y(n_438)
);

BUFx3_ASAP7_75t_L g439 ( 
.A(n_374),
.Y(n_439)
);

BUFx2_ASAP7_75t_L g440 ( 
.A(n_341),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_374),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_376),
.Y(n_442)
);

BUFx2_ASAP7_75t_L g443 ( 
.A(n_352),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_376),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_382),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_382),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_383),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_326),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_350),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_350),
.Y(n_450)
);

INVx3_ASAP7_75t_L g451 ( 
.A(n_311),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_364),
.Y(n_452)
);

BUFx2_ASAP7_75t_L g453 ( 
.A(n_387),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_387),
.B(n_313),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_439),
.Y(n_455)
);

NAND3xp33_ASAP7_75t_L g456 ( 
.A(n_419),
.B(n_315),
.C(n_370),
.Y(n_456)
);

INVxp67_ASAP7_75t_L g457 ( 
.A(n_391),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_439),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_417),
.B(n_324),
.Y(n_459)
);

BUFx8_ASAP7_75t_SL g460 ( 
.A(n_404),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_439),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_434),
.B(n_314),
.Y(n_462)
);

INVx2_ASAP7_75t_SL g463 ( 
.A(n_434),
.Y(n_463)
);

BUFx3_ASAP7_75t_L g464 ( 
.A(n_407),
.Y(n_464)
);

AND3x2_ASAP7_75t_L g465 ( 
.A(n_391),
.B(n_272),
.C(n_367),
.Y(n_465)
);

AND2x4_ASAP7_75t_L g466 ( 
.A(n_401),
.B(n_196),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_385),
.Y(n_467)
);

BUFx3_ASAP7_75t_L g468 ( 
.A(n_407),
.Y(n_468)
);

OR2x6_ASAP7_75t_L g469 ( 
.A(n_451),
.B(n_364),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_427),
.B(n_320),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_385),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_439),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_384),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_427),
.B(n_323),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_390),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_434),
.B(n_325),
.Y(n_476)
);

INVx4_ASAP7_75t_L g477 ( 
.A(n_385),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_417),
.B(n_333),
.Y(n_478)
);

OR2x6_ASAP7_75t_L g479 ( 
.A(n_451),
.B(n_197),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_384),
.Y(n_480)
);

OAI22xp33_ASAP7_75t_L g481 ( 
.A1(n_428),
.A2(n_287),
.B1(n_312),
.B2(n_210),
.Y(n_481)
);

NAND3xp33_ASAP7_75t_L g482 ( 
.A(n_419),
.B(n_217),
.C(n_198),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_434),
.B(n_345),
.Y(n_483)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_385),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_390),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_390),
.Y(n_486)
);

INVx3_ASAP7_75t_L g487 ( 
.A(n_385),
.Y(n_487)
);

INVx2_ASAP7_75t_SL g488 ( 
.A(n_434),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_417),
.B(n_349),
.Y(n_489)
);

INVx4_ASAP7_75t_L g490 ( 
.A(n_385),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_434),
.B(n_353),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_419),
.B(n_354),
.Y(n_492)
);

AND2x6_ASAP7_75t_L g493 ( 
.A(n_413),
.B(n_229),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_388),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_388),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_392),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_434),
.B(n_356),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_392),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_390),
.Y(n_499)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_385),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_448),
.B(n_355),
.Y(n_501)
);

BUFx2_ASAP7_75t_L g502 ( 
.A(n_432),
.Y(n_502)
);

OAI21xp33_ASAP7_75t_SL g503 ( 
.A1(n_419),
.A2(n_266),
.B(n_260),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_394),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_413),
.B(n_362),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_395),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_413),
.B(n_434),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_448),
.B(n_355),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_434),
.B(n_365),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_395),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_451),
.B(n_368),
.Y(n_511)
);

AOI22xp33_ASAP7_75t_L g512 ( 
.A1(n_413),
.A2(n_358),
.B1(n_271),
.B2(n_296),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_413),
.B(n_371),
.Y(n_513)
);

BUFx10_ASAP7_75t_L g514 ( 
.A(n_413),
.Y(n_514)
);

BUFx8_ASAP7_75t_SL g515 ( 
.A(n_404),
.Y(n_515)
);

INVx1_ASAP7_75t_SL g516 ( 
.A(n_432),
.Y(n_516)
);

BUFx3_ASAP7_75t_L g517 ( 
.A(n_407),
.Y(n_517)
);

AOI22xp33_ASAP7_75t_L g518 ( 
.A1(n_397),
.A2(n_277),
.B1(n_292),
.B2(n_278),
.Y(n_518)
);

AND3x2_ASAP7_75t_L g519 ( 
.A(n_432),
.B(n_380),
.C(n_248),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_395),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_395),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_428),
.B(n_375),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_448),
.B(n_312),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_398),
.Y(n_524)
);

AOI22xp33_ASAP7_75t_L g525 ( 
.A1(n_397),
.A2(n_262),
.B1(n_237),
.B2(n_243),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_420),
.A2(n_302),
.B1(n_241),
.B2(n_158),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_451),
.B(n_379),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_398),
.Y(n_528)
);

BUFx3_ASAP7_75t_L g529 ( 
.A(n_407),
.Y(n_529)
);

NAND2xp33_ASAP7_75t_L g530 ( 
.A(n_449),
.B(n_381),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_449),
.B(n_213),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_449),
.B(n_258),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_398),
.Y(n_533)
);

INVx4_ASAP7_75t_L g534 ( 
.A(n_385),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_398),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_386),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_400),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_400),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_400),
.Y(n_539)
);

AOI22x1_ASAP7_75t_L g540 ( 
.A1(n_452),
.A2(n_177),
.B1(n_174),
.B2(n_305),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_394),
.Y(n_541)
);

NAND2xp33_ASAP7_75t_L g542 ( 
.A(n_450),
.B(n_163),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_450),
.B(n_230),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_429),
.Y(n_544)
);

AOI21x1_ASAP7_75t_L g545 ( 
.A1(n_401),
.A2(n_192),
.B(n_274),
.Y(n_545)
);

INVx3_ASAP7_75t_L g546 ( 
.A(n_386),
.Y(n_546)
);

BUFx4f_ASAP7_75t_L g547 ( 
.A(n_407),
.Y(n_547)
);

AOI22xp5_ASAP7_75t_L g548 ( 
.A1(n_420),
.A2(n_286),
.B1(n_174),
.B2(n_177),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_429),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_450),
.B(n_259),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_402),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_402),
.Y(n_552)
);

BUFx2_ASAP7_75t_L g553 ( 
.A(n_440),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_451),
.B(n_377),
.Y(n_554)
);

AND2x6_ASAP7_75t_L g555 ( 
.A(n_420),
.B(n_273),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_399),
.B(n_344),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_429),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_386),
.Y(n_558)
);

INVx5_ASAP7_75t_L g559 ( 
.A(n_386),
.Y(n_559)
);

INVx3_ASAP7_75t_L g560 ( 
.A(n_386),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_429),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_386),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_402),
.Y(n_563)
);

BUFx2_ASAP7_75t_L g564 ( 
.A(n_440),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_402),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g566 ( 
.A(n_452),
.B(n_258),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_397),
.B(n_303),
.Y(n_567)
);

INVx4_ASAP7_75t_L g568 ( 
.A(n_386),
.Y(n_568)
);

AOI22xp33_ASAP7_75t_L g569 ( 
.A1(n_420),
.A2(n_401),
.B1(n_421),
.B2(n_423),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_399),
.B(n_348),
.Y(n_570)
);

OAI21xp33_ASAP7_75t_SL g571 ( 
.A1(n_421),
.A2(n_307),
.B(n_221),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_429),
.Y(n_572)
);

BUFx8_ASAP7_75t_SL g573 ( 
.A(n_440),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_430),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_420),
.B(n_268),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_386),
.Y(n_576)
);

INVx3_ASAP7_75t_L g577 ( 
.A(n_389),
.Y(n_577)
);

AOI22xp33_ASAP7_75t_L g578 ( 
.A1(n_420),
.A2(n_401),
.B1(n_421),
.B2(n_423),
.Y(n_578)
);

BUFx6f_ASAP7_75t_L g579 ( 
.A(n_389),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_405),
.B(n_163),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_389),
.Y(n_581)
);

AOI22xp33_ASAP7_75t_L g582 ( 
.A1(n_401),
.A2(n_192),
.B1(n_258),
.B2(n_304),
.Y(n_582)
);

INVx4_ASAP7_75t_L g583 ( 
.A(n_389),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_389),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_389),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_405),
.B(n_166),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_412),
.B(n_166),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_389),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_412),
.B(n_443),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_430),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_430),
.Y(n_591)
);

INVx3_ASAP7_75t_L g592 ( 
.A(n_389),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_393),
.Y(n_593)
);

INVx4_ASAP7_75t_L g594 ( 
.A(n_393),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_443),
.Y(n_595)
);

INVx6_ASAP7_75t_L g596 ( 
.A(n_407),
.Y(n_596)
);

HB1xp67_ASAP7_75t_L g597 ( 
.A(n_416),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_430),
.Y(n_598)
);

AND2x6_ASAP7_75t_L g599 ( 
.A(n_401),
.B(n_192),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_407),
.B(n_167),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_443),
.B(n_359),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_522),
.B(n_407),
.Y(n_602)
);

INVx2_ASAP7_75t_SL g603 ( 
.A(n_453),
.Y(n_603)
);

AOI22xp5_ASAP7_75t_L g604 ( 
.A1(n_492),
.A2(n_366),
.B1(n_310),
.B2(n_343),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_485),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_455),
.Y(n_606)
);

AOI22xp33_ASAP7_75t_L g607 ( 
.A1(n_482),
.A2(n_423),
.B1(n_430),
.B2(n_435),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_474),
.B(n_410),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_514),
.B(n_410),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_455),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_514),
.B(n_410),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_569),
.B(n_578),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_458),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_514),
.B(n_410),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_470),
.B(n_416),
.Y(n_615)
);

OAI22xp5_ASAP7_75t_L g616 ( 
.A1(n_456),
.A2(n_335),
.B1(n_330),
.B2(n_334),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_514),
.B(n_410),
.Y(n_617)
);

AOI22xp5_ASAP7_75t_L g618 ( 
.A1(n_456),
.A2(n_410),
.B1(n_167),
.B2(n_170),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_478),
.B(n_169),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_489),
.B(n_589),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_527),
.B(n_410),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_505),
.B(n_410),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_580),
.B(n_169),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_485),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_513),
.B(n_435),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_486),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_586),
.B(n_170),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_486),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_458),
.B(n_435),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_461),
.B(n_435),
.Y(n_630)
);

BUFx6f_ASAP7_75t_SL g631 ( 
.A(n_555),
.Y(n_631)
);

INVxp67_ASAP7_75t_L g632 ( 
.A(n_453),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_587),
.B(n_171),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_486),
.Y(n_634)
);

NOR2xp67_ASAP7_75t_SL g635 ( 
.A(n_482),
.B(n_435),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_461),
.B(n_438),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_503),
.B(n_192),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_472),
.B(n_438),
.Y(n_638)
);

INVx4_ASAP7_75t_L g639 ( 
.A(n_467),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_510),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_503),
.B(n_192),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_510),
.Y(n_642)
);

INVx1_ASAP7_75t_SL g643 ( 
.A(n_516),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_472),
.Y(n_644)
);

AOI22xp5_ASAP7_75t_L g645 ( 
.A1(n_555),
.A2(n_171),
.B1(n_173),
.B2(n_175),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_473),
.Y(n_646)
);

AOI22xp5_ASAP7_75t_L g647 ( 
.A1(n_555),
.A2(n_173),
.B1(n_175),
.B2(n_178),
.Y(n_647)
);

BUFx4_ASAP7_75t_L g648 ( 
.A(n_460),
.Y(n_648)
);

AOI22xp33_ASAP7_75t_L g649 ( 
.A1(n_555),
.A2(n_438),
.B1(n_446),
.B2(n_445),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_507),
.B(n_192),
.Y(n_650)
);

BUFx8_ASAP7_75t_L g651 ( 
.A(n_502),
.Y(n_651)
);

INVx2_ASAP7_75t_SL g652 ( 
.A(n_501),
.Y(n_652)
);

AND2x4_ASAP7_75t_L g653 ( 
.A(n_466),
.B(n_422),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_567),
.B(n_178),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_473),
.Y(n_655)
);

OAI22xp5_ASAP7_75t_L g656 ( 
.A1(n_469),
.A2(n_438),
.B1(n_185),
.B2(n_188),
.Y(n_656)
);

OR2x6_ASAP7_75t_L g657 ( 
.A(n_502),
.B(n_553),
.Y(n_657)
);

BUFx6f_ASAP7_75t_L g658 ( 
.A(n_464),
.Y(n_658)
);

HB1xp67_ASAP7_75t_L g659 ( 
.A(n_597),
.Y(n_659)
);

BUFx3_ASAP7_75t_L g660 ( 
.A(n_466),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_555),
.B(n_438),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_555),
.B(n_441),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_555),
.B(n_441),
.Y(n_663)
);

NOR2xp67_ASAP7_75t_L g664 ( 
.A(n_554),
.B(n_422),
.Y(n_664)
);

BUFx3_ASAP7_75t_L g665 ( 
.A(n_466),
.Y(n_665)
);

AND2x4_ASAP7_75t_L g666 ( 
.A(n_466),
.B(n_532),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_510),
.Y(n_667)
);

INVxp67_ASAP7_75t_L g668 ( 
.A(n_553),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_515),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_475),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_480),
.B(n_441),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_544),
.B(n_192),
.Y(n_672)
);

AOI22xp33_ASAP7_75t_L g673 ( 
.A1(n_493),
.A2(n_447),
.B1(n_446),
.B2(n_445),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_544),
.B(n_441),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_454),
.B(n_183),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_480),
.B(n_494),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_494),
.B(n_441),
.Y(n_677)
);

NOR3xp33_ASAP7_75t_L g678 ( 
.A(n_601),
.B(n_433),
.C(n_426),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_549),
.B(n_441),
.Y(n_679)
);

NOR3xp33_ASAP7_75t_L g680 ( 
.A(n_481),
.B(n_433),
.C(n_426),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_495),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_457),
.B(n_183),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_495),
.Y(n_683)
);

INVx2_ASAP7_75t_SL g684 ( 
.A(n_501),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_475),
.Y(n_685)
);

BUFx6f_ASAP7_75t_L g686 ( 
.A(n_464),
.Y(n_686)
);

OR2x2_ASAP7_75t_L g687 ( 
.A(n_564),
.B(n_431),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_549),
.B(n_441),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_496),
.B(n_441),
.Y(n_689)
);

AOI22xp33_ASAP7_75t_L g690 ( 
.A1(n_493),
.A2(n_447),
.B1(n_446),
.B2(n_445),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_496),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_498),
.B(n_424),
.Y(n_692)
);

INVxp67_ASAP7_75t_L g693 ( 
.A(n_564),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_557),
.B(n_185),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_557),
.B(n_188),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_499),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_498),
.B(n_424),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_561),
.B(n_282),
.Y(n_698)
);

NAND2xp33_ASAP7_75t_L g699 ( 
.A(n_493),
.B(n_282),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_523),
.B(n_285),
.Y(n_700)
);

AO22x2_ASAP7_75t_L g701 ( 
.A1(n_459),
.A2(n_447),
.B1(n_418),
.B2(n_442),
.Y(n_701)
);

OR2x2_ASAP7_75t_L g702 ( 
.A(n_523),
.B(n_431),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_504),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_504),
.Y(n_704)
);

INVx3_ASAP7_75t_L g705 ( 
.A(n_537),
.Y(n_705)
);

INVx2_ASAP7_75t_SL g706 ( 
.A(n_508),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_499),
.Y(n_707)
);

AOI22xp33_ASAP7_75t_L g708 ( 
.A1(n_493),
.A2(n_418),
.B1(n_442),
.B2(n_406),
.Y(n_708)
);

A2O1A1Ixp33_ASAP7_75t_L g709 ( 
.A1(n_532),
.A2(n_418),
.B(n_437),
.C(n_436),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_459),
.B(n_285),
.Y(n_710)
);

AOI22xp5_ASAP7_75t_L g711 ( 
.A1(n_530),
.A2(n_290),
.B1(n_295),
.B2(n_300),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_541),
.B(n_424),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_541),
.B(n_424),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_506),
.Y(n_714)
);

CKINVDCx20_ASAP7_75t_R g715 ( 
.A(n_573),
.Y(n_715)
);

INVx2_ASAP7_75t_SL g716 ( 
.A(n_508),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_531),
.B(n_290),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_566),
.B(n_403),
.Y(n_718)
);

INVx2_ASAP7_75t_SL g719 ( 
.A(n_566),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_561),
.Y(n_720)
);

INVxp67_ASAP7_75t_SL g721 ( 
.A(n_467),
.Y(n_721)
);

AOI21xp5_ASAP7_75t_L g722 ( 
.A1(n_600),
.A2(n_444),
.B(n_437),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_556),
.B(n_295),
.Y(n_723)
);

NOR3xp33_ASAP7_75t_L g724 ( 
.A(n_570),
.B(n_191),
.C(n_195),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_572),
.B(n_425),
.Y(n_725)
);

INVx3_ASAP7_75t_L g726 ( 
.A(n_537),
.Y(n_726)
);

INVx3_ASAP7_75t_L g727 ( 
.A(n_538),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_572),
.B(n_425),
.Y(n_728)
);

OR2x2_ASAP7_75t_L g729 ( 
.A(n_543),
.B(n_179),
.Y(n_729)
);

OR2x6_ASAP7_75t_L g730 ( 
.A(n_511),
.B(n_425),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_574),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_506),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_574),
.Y(n_733)
);

AOI22xp5_ASAP7_75t_L g734 ( 
.A1(n_469),
.A2(n_300),
.B1(n_437),
.B2(n_436),
.Y(n_734)
);

AOI22xp5_ASAP7_75t_L g735 ( 
.A1(n_469),
.A2(n_444),
.B1(n_437),
.B2(n_436),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_590),
.Y(n_736)
);

BUFx6f_ASAP7_75t_SL g737 ( 
.A(n_479),
.Y(n_737)
);

OR2x2_ASAP7_75t_L g738 ( 
.A(n_550),
.B(n_179),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_590),
.B(n_425),
.Y(n_739)
);

INVxp67_ASAP7_75t_SL g740 ( 
.A(n_467),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_591),
.B(n_436),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_591),
.B(n_444),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_598),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_598),
.B(n_444),
.Y(n_744)
);

AOI22xp33_ASAP7_75t_L g745 ( 
.A1(n_493),
.A2(n_415),
.B1(n_414),
.B2(n_411),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_538),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_575),
.B(n_393),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_483),
.B(n_393),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_539),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_571),
.B(n_218),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_539),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_551),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_595),
.B(n_403),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_558),
.B(n_393),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_571),
.B(n_224),
.Y(n_755)
);

AOI22xp5_ASAP7_75t_L g756 ( 
.A1(n_469),
.A2(n_415),
.B1(n_414),
.B2(n_411),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_542),
.B(n_227),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_558),
.B(n_393),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_558),
.B(n_393),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_548),
.B(n_231),
.Y(n_760)
);

INVx1_ASAP7_75t_SL g761 ( 
.A(n_465),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_520),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_576),
.B(n_393),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_576),
.B(n_585),
.Y(n_764)
);

INVxp67_ASAP7_75t_L g765 ( 
.A(n_540),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_520),
.Y(n_766)
);

AND2x4_ASAP7_75t_L g767 ( 
.A(n_479),
.B(n_403),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_585),
.B(n_396),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_551),
.Y(n_769)
);

AOI22xp5_ASAP7_75t_L g770 ( 
.A1(n_469),
.A2(n_415),
.B1(n_414),
.B2(n_411),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_562),
.B(n_396),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_521),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_562),
.B(n_396),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_620),
.B(n_512),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_620),
.B(n_525),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_612),
.B(n_562),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_718),
.B(n_493),
.Y(n_777)
);

AOI21xp5_ASAP7_75t_L g778 ( 
.A1(n_621),
.A2(n_547),
.B(n_477),
.Y(n_778)
);

HB1xp67_ASAP7_75t_L g779 ( 
.A(n_657),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_649),
.B(n_673),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_705),
.Y(n_781)
);

O2A1O1Ixp33_ASAP7_75t_L g782 ( 
.A1(n_765),
.A2(n_479),
.B(n_462),
.C(n_491),
.Y(n_782)
);

OAI21xp33_ASAP7_75t_L g783 ( 
.A1(n_760),
.A2(n_548),
.B(n_526),
.Y(n_783)
);

A2O1A1Ixp33_ASAP7_75t_L g784 ( 
.A1(n_654),
.A2(n_526),
.B(n_518),
.C(n_582),
.Y(n_784)
);

HB1xp67_ASAP7_75t_L g785 ( 
.A(n_657),
.Y(n_785)
);

OR2x2_ASAP7_75t_L g786 ( 
.A(n_643),
.B(n_479),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_753),
.B(n_652),
.Y(n_787)
);

AOI21xp5_ASAP7_75t_L g788 ( 
.A1(n_602),
.A2(n_547),
.B(n_583),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_649),
.B(n_581),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_705),
.Y(n_790)
);

BUFx6f_ASAP7_75t_L g791 ( 
.A(n_658),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_654),
.B(n_493),
.Y(n_792)
);

OAI321xp33_ASAP7_75t_L g793 ( 
.A1(n_760),
.A2(n_479),
.A3(n_545),
.B1(n_540),
.B2(n_406),
.C(n_409),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_632),
.B(n_519),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_720),
.Y(n_795)
);

AOI21xp5_ASAP7_75t_L g796 ( 
.A1(n_622),
.A2(n_547),
.B(n_534),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_615),
.B(n_476),
.Y(n_797)
);

OAI21xp33_ASAP7_75t_L g798 ( 
.A1(n_710),
.A2(n_297),
.B(n_294),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_603),
.B(n_497),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_619),
.B(n_509),
.Y(n_800)
);

AOI21xp5_ASAP7_75t_L g801 ( 
.A1(n_608),
.A2(n_534),
.B(n_477),
.Y(n_801)
);

OAI21xp5_ASAP7_75t_L g802 ( 
.A1(n_625),
.A2(n_463),
.B(n_488),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_619),
.B(n_484),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_609),
.A2(n_534),
.B(n_477),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_669),
.Y(n_805)
);

OAI21xp5_ASAP7_75t_L g806 ( 
.A1(n_709),
.A2(n_463),
.B(n_488),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_609),
.A2(n_490),
.B(n_583),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_673),
.B(n_581),
.Y(n_808)
);

AOI21xp5_ASAP7_75t_L g809 ( 
.A1(n_611),
.A2(n_490),
.B(n_583),
.Y(n_809)
);

OAI22xp5_ASAP7_75t_L g810 ( 
.A1(n_666),
.A2(n_529),
.B1(n_517),
.B2(n_464),
.Y(n_810)
);

INVx3_ASAP7_75t_L g811 ( 
.A(n_660),
.Y(n_811)
);

AOI21xp5_ASAP7_75t_L g812 ( 
.A1(n_611),
.A2(n_477),
.B(n_534),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_614),
.A2(n_490),
.B(n_568),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_614),
.A2(n_490),
.B(n_568),
.Y(n_814)
);

INVx2_ASAP7_75t_SL g815 ( 
.A(n_657),
.Y(n_815)
);

A2O1A1Ixp33_ASAP7_75t_L g816 ( 
.A1(n_757),
.A2(n_623),
.B(n_633),
.C(n_627),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_623),
.B(n_484),
.Y(n_817)
);

AOI21xp5_ASAP7_75t_L g818 ( 
.A1(n_617),
.A2(n_568),
.B(n_583),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_690),
.B(n_581),
.Y(n_819)
);

AND2x2_ASAP7_75t_L g820 ( 
.A(n_684),
.B(n_181),
.Y(n_820)
);

OAI21xp5_ASAP7_75t_L g821 ( 
.A1(n_629),
.A2(n_636),
.B(n_630),
.Y(n_821)
);

OAI321xp33_ASAP7_75t_L g822 ( 
.A1(n_750),
.A2(n_755),
.A3(n_723),
.B1(n_675),
.B2(n_757),
.C(n_710),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_731),
.Y(n_823)
);

AO21x1_ASAP7_75t_L g824 ( 
.A1(n_637),
.A2(n_545),
.B(n_588),
.Y(n_824)
);

BUFx12f_ASAP7_75t_L g825 ( 
.A(n_651),
.Y(n_825)
);

AOI21xp5_ASAP7_75t_L g826 ( 
.A1(n_617),
.A2(n_568),
.B(n_517),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_706),
.B(n_181),
.Y(n_827)
);

AOI21xp33_ASAP7_75t_L g828 ( 
.A1(n_723),
.A2(n_269),
.B(n_242),
.Y(n_828)
);

OAI21xp5_ASAP7_75t_L g829 ( 
.A1(n_638),
.A2(n_584),
.B(n_588),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_627),
.B(n_484),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_733),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_633),
.B(n_484),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_747),
.A2(n_529),
.B(n_468),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_646),
.B(n_487),
.Y(n_834)
);

OAI21xp5_ASAP7_75t_L g835 ( 
.A1(n_722),
.A2(n_584),
.B(n_588),
.Y(n_835)
);

OAI21xp33_ASAP7_75t_L g836 ( 
.A1(n_675),
.A2(n_187),
.B(n_283),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_655),
.B(n_487),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_748),
.A2(n_529),
.B(n_468),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_736),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_681),
.B(n_487),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_683),
.B(n_487),
.Y(n_841)
);

AOI22xp5_ASAP7_75t_L g842 ( 
.A1(n_666),
.A2(n_599),
.B1(n_592),
.B2(n_500),
.Y(n_842)
);

A2O1A1Ixp33_ASAP7_75t_L g843 ( 
.A1(n_700),
.A2(n_682),
.B(n_664),
.C(n_719),
.Y(n_843)
);

AND2x4_ASAP7_75t_L g844 ( 
.A(n_660),
.B(n_665),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_716),
.B(n_500),
.Y(n_845)
);

NAND2x1p5_ASAP7_75t_L g846 ( 
.A(n_665),
.B(n_468),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_721),
.A2(n_517),
.B(n_467),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_691),
.B(n_703),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_743),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_704),
.B(n_500),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_606),
.Y(n_851)
);

BUFx6f_ASAP7_75t_L g852 ( 
.A(n_658),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_676),
.B(n_500),
.Y(n_853)
);

NOR2xp67_ASAP7_75t_L g854 ( 
.A(n_604),
.B(n_584),
.Y(n_854)
);

NAND2x1p5_ASAP7_75t_L g855 ( 
.A(n_658),
.B(n_536),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_653),
.B(n_536),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_668),
.B(n_536),
.Y(n_857)
);

AND2x2_ASAP7_75t_L g858 ( 
.A(n_687),
.B(n_187),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_726),
.Y(n_859)
);

BUFx12f_ASAP7_75t_L g860 ( 
.A(n_651),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_653),
.B(n_536),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_693),
.B(n_546),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_740),
.A2(n_471),
.B(n_467),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_610),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_700),
.B(n_546),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_639),
.A2(n_579),
.B(n_471),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_639),
.A2(n_579),
.B(n_471),
.Y(n_867)
);

HB1xp67_ASAP7_75t_L g868 ( 
.A(n_659),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_764),
.A2(n_663),
.B(n_662),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_682),
.B(n_546),
.Y(n_870)
);

INVx2_ASAP7_75t_SL g871 ( 
.A(n_659),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_701),
.B(n_546),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_690),
.B(n_471),
.Y(n_873)
);

BUFx4f_ASAP7_75t_L g874 ( 
.A(n_730),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_613),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_701),
.B(n_560),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_701),
.B(n_560),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_644),
.B(n_560),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_680),
.B(n_560),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_702),
.B(n_283),
.Y(n_880)
);

OAI22xp5_ASAP7_75t_L g881 ( 
.A1(n_756),
.A2(n_596),
.B1(n_577),
.B2(n_592),
.Y(n_881)
);

INVx1_ASAP7_75t_SL g882 ( 
.A(n_648),
.Y(n_882)
);

OAI21xp5_ASAP7_75t_L g883 ( 
.A1(n_661),
.A2(n_577),
.B(n_592),
.Y(n_883)
);

A2O1A1Ixp33_ASAP7_75t_L g884 ( 
.A1(n_750),
.A2(n_592),
.B(n_577),
.C(n_593),
.Y(n_884)
);

BUFx6f_ASAP7_75t_L g885 ( 
.A(n_658),
.Y(n_885)
);

BUFx2_ASAP7_75t_L g886 ( 
.A(n_730),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_726),
.B(n_577),
.Y(n_887)
);

HB1xp67_ASAP7_75t_L g888 ( 
.A(n_767),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_745),
.A2(n_708),
.B(n_771),
.Y(n_889)
);

AND2x4_ASAP7_75t_L g890 ( 
.A(n_767),
.B(n_406),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_745),
.A2(n_579),
.B(n_471),
.Y(n_891)
);

OAI22xp5_ASAP7_75t_L g892 ( 
.A1(n_770),
.A2(n_596),
.B1(n_579),
.B2(n_593),
.Y(n_892)
);

BUFx8_ASAP7_75t_SL g893 ( 
.A(n_715),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_727),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_727),
.B(n_579),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_607),
.B(n_599),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_708),
.A2(n_594),
.B(n_559),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_763),
.A2(n_594),
.B(n_559),
.Y(n_898)
);

OR2x2_ASAP7_75t_L g899 ( 
.A(n_729),
.B(n_289),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_607),
.B(n_599),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_738),
.B(n_599),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_746),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_L g903 ( 
.A(n_761),
.B(n_235),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_768),
.A2(n_594),
.B(n_559),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_749),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_686),
.A2(n_594),
.B(n_559),
.Y(n_906)
);

AND2x2_ASAP7_75t_L g907 ( 
.A(n_755),
.B(n_289),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_751),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_686),
.A2(n_559),
.B(n_593),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_686),
.A2(n_559),
.B(n_552),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_686),
.A2(n_552),
.B(n_563),
.Y(n_911)
);

O2A1O1Ixp33_ASAP7_75t_L g912 ( 
.A1(n_694),
.A2(n_563),
.B(n_565),
.C(n_528),
.Y(n_912)
);

INVx3_ASAP7_75t_L g913 ( 
.A(n_670),
.Y(n_913)
);

INVx3_ASAP7_75t_L g914 ( 
.A(n_685),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_650),
.A2(n_697),
.B(n_692),
.Y(n_915)
);

NOR2xp33_ASAP7_75t_L g916 ( 
.A(n_616),
.B(n_247),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_650),
.A2(n_565),
.B(n_521),
.Y(n_917)
);

AND2x2_ASAP7_75t_SL g918 ( 
.A(n_645),
.B(n_408),
.Y(n_918)
);

INVx1_ASAP7_75t_SL g919 ( 
.A(n_717),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_694),
.B(n_695),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_739),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_712),
.A2(n_528),
.B(n_524),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_713),
.A2(n_689),
.B(n_671),
.Y(n_923)
);

OAI21xp5_ASAP7_75t_L g924 ( 
.A1(n_735),
.A2(n_535),
.B(n_533),
.Y(n_924)
);

A2O1A1Ixp33_ASAP7_75t_L g925 ( 
.A1(n_734),
.A2(n_535),
.B(n_533),
.C(n_524),
.Y(n_925)
);

OAI22xp5_ASAP7_75t_L g926 ( 
.A1(n_730),
.A2(n_631),
.B1(n_618),
.B2(n_647),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_677),
.A2(n_396),
.B(n_596),
.Y(n_927)
);

INVxp67_ASAP7_75t_L g928 ( 
.A(n_695),
.Y(n_928)
);

INVx2_ASAP7_75t_SL g929 ( 
.A(n_698),
.Y(n_929)
);

AND2x2_ASAP7_75t_SL g930 ( 
.A(n_724),
.B(n_699),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_739),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_725),
.A2(n_396),
.B(n_596),
.Y(n_932)
);

O2A1O1Ixp33_ASAP7_75t_L g933 ( 
.A1(n_698),
.A2(n_409),
.B(n_408),
.C(n_599),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_678),
.B(n_599),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_752),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_728),
.A2(n_396),
.B(n_409),
.Y(n_936)
);

INVx3_ASAP7_75t_L g937 ( 
.A(n_696),
.Y(n_937)
);

OAI21xp33_ASAP7_75t_L g938 ( 
.A1(n_711),
.A2(n_291),
.B(n_293),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_L g939 ( 
.A(n_656),
.B(n_251),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_769),
.B(n_599),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_605),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_707),
.B(n_408),
.Y(n_942)
);

HB1xp67_ASAP7_75t_L g943 ( 
.A(n_737),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_737),
.B(n_250),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_741),
.A2(n_396),
.B(n_281),
.Y(n_945)
);

INVx4_ASAP7_75t_L g946 ( 
.A(n_631),
.Y(n_946)
);

INVx3_ASAP7_75t_L g947 ( 
.A(n_714),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_SL g948 ( 
.A(n_742),
.B(n_744),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_754),
.A2(n_396),
.B(n_252),
.Y(n_949)
);

INVx3_ASAP7_75t_L g950 ( 
.A(n_732),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_754),
.A2(n_773),
.B(n_758),
.Y(n_951)
);

NAND3xp33_ASAP7_75t_L g952 ( 
.A(n_635),
.B(n_264),
.C(n_267),
.Y(n_952)
);

OR2x6_ASAP7_75t_L g953 ( 
.A(n_637),
.B(n_304),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_672),
.B(n_305),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_762),
.B(n_270),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_758),
.A2(n_275),
.B(n_280),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_766),
.B(n_276),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_759),
.A2(n_291),
.B(n_299),
.Y(n_958)
);

NOR2xp67_ASAP7_75t_SL g959 ( 
.A(n_641),
.B(n_299),
.Y(n_959)
);

BUFx12f_ASAP7_75t_L g960 ( 
.A(n_641),
.Y(n_960)
);

INVx1_ASAP7_75t_SL g961 ( 
.A(n_672),
.Y(n_961)
);

AOI21x1_ASAP7_75t_L g962 ( 
.A1(n_674),
.A2(n_304),
.B(n_114),
.Y(n_962)
);

AND2x4_ASAP7_75t_L g963 ( 
.A(n_674),
.B(n_154),
.Y(n_963)
);

BUFx6f_ASAP7_75t_L g964 ( 
.A(n_791),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_816),
.A2(n_773),
.B(n_759),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_869),
.A2(n_688),
.B(n_679),
.Y(n_966)
);

AO21x1_ASAP7_75t_L g967 ( 
.A1(n_800),
.A2(n_688),
.B(n_679),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_802),
.A2(n_772),
.B(n_667),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_775),
.B(n_642),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_787),
.B(n_293),
.Y(n_970)
);

AOI22xp5_ASAP7_75t_L g971 ( 
.A1(n_783),
.A2(n_797),
.B1(n_774),
.B2(n_916),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_L g972 ( 
.A(n_822),
.B(n_640),
.Y(n_972)
);

BUFx3_ASAP7_75t_L g973 ( 
.A(n_871),
.Y(n_973)
);

AND2x2_ASAP7_75t_L g974 ( 
.A(n_858),
.B(n_298),
.Y(n_974)
);

INVx3_ASAP7_75t_L g975 ( 
.A(n_791),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_780),
.A2(n_634),
.B(n_628),
.Y(n_976)
);

OA21x2_ASAP7_75t_L g977 ( 
.A1(n_883),
.A2(n_626),
.B(n_624),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_928),
.B(n_298),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_780),
.A2(n_297),
.B(n_294),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_851),
.Y(n_980)
);

OR2x6_ASAP7_75t_L g981 ( 
.A(n_815),
.B(n_138),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_916),
.B(n_14),
.Y(n_982)
);

NOR2x1_ASAP7_75t_R g983 ( 
.A(n_825),
.B(n_21),
.Y(n_983)
);

BUFx12f_ASAP7_75t_L g984 ( 
.A(n_860),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_928),
.B(n_22),
.Y(n_985)
);

AND2x2_ASAP7_75t_L g986 ( 
.A(n_880),
.B(n_26),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_907),
.B(n_26),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_929),
.B(n_27),
.Y(n_988)
);

OAI21xp5_ASAP7_75t_L g989 ( 
.A1(n_896),
.A2(n_136),
.B(n_135),
.Y(n_989)
);

OAI22xp5_ASAP7_75t_SL g990 ( 
.A1(n_882),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_990)
);

NAND3xp33_ASAP7_75t_SL g991 ( 
.A(n_836),
.B(n_29),
.C(n_31),
.Y(n_991)
);

OAI22xp5_ASAP7_75t_L g992 ( 
.A1(n_900),
.A2(n_133),
.B1(n_126),
.B2(n_111),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_941),
.Y(n_993)
);

AOI22x1_ASAP7_75t_L g994 ( 
.A1(n_915),
.A2(n_110),
.B1(n_109),
.B2(n_93),
.Y(n_994)
);

BUFx2_ASAP7_75t_L g995 ( 
.A(n_868),
.Y(n_995)
);

CKINVDCx20_ASAP7_75t_R g996 ( 
.A(n_893),
.Y(n_996)
);

BUFx6f_ASAP7_75t_L g997 ( 
.A(n_791),
.Y(n_997)
);

AOI22x1_ASAP7_75t_L g998 ( 
.A1(n_923),
.A2(n_92),
.B1(n_90),
.B2(n_81),
.Y(n_998)
);

INVx3_ASAP7_75t_L g999 ( 
.A(n_791),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_844),
.B(n_80),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_848),
.B(n_31),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_778),
.A2(n_61),
.B(n_62),
.Y(n_1002)
);

OAI22xp5_ASAP7_75t_SL g1003 ( 
.A1(n_805),
.A2(n_33),
.B1(n_35),
.B2(n_36),
.Y(n_1003)
);

NAND3xp33_ASAP7_75t_SL g1004 ( 
.A(n_784),
.B(n_35),
.C(n_36),
.Y(n_1004)
);

OAI22xp5_ASAP7_75t_L g1005 ( 
.A1(n_874),
.A2(n_37),
.B1(n_38),
.B2(n_41),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_SL g1006 ( 
.A(n_844),
.B(n_42),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_803),
.A2(n_43),
.B(n_44),
.Y(n_1007)
);

AND2x4_ASAP7_75t_L g1008 ( 
.A(n_888),
.B(n_46),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_L g1009 ( 
.A(n_868),
.B(n_47),
.Y(n_1009)
);

A2O1A1Ixp33_ASAP7_75t_L g1010 ( 
.A1(n_797),
.A2(n_939),
.B(n_920),
.C(n_843),
.Y(n_1010)
);

AO32x1_ASAP7_75t_L g1011 ( 
.A1(n_926),
.A2(n_47),
.A3(n_48),
.B1(n_49),
.B2(n_52),
.Y(n_1011)
);

AOI22xp33_ASAP7_75t_L g1012 ( 
.A1(n_939),
.A2(n_953),
.B1(n_828),
.B2(n_930),
.Y(n_1012)
);

BUFx3_ASAP7_75t_L g1013 ( 
.A(n_779),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_905),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_788),
.A2(n_52),
.B(n_54),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_792),
.A2(n_865),
.B(n_830),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_L g1017 ( 
.A(n_903),
.B(n_919),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_864),
.Y(n_1018)
);

NAND2x1p5_ASAP7_75t_L g1019 ( 
.A(n_852),
.B(n_885),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_875),
.B(n_795),
.Y(n_1020)
);

AO22x1_ASAP7_75t_L g1021 ( 
.A1(n_944),
.A2(n_794),
.B1(n_785),
.B2(n_779),
.Y(n_1021)
);

AOI21xp33_ASAP7_75t_L g1022 ( 
.A1(n_899),
.A2(n_901),
.B(n_903),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_823),
.B(n_831),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_839),
.B(n_849),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_817),
.A2(n_832),
.B(n_796),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_799),
.B(n_857),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_874),
.B(n_888),
.Y(n_1027)
);

NOR2xp33_ASAP7_75t_L g1028 ( 
.A(n_786),
.B(n_798),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_SL g1029 ( 
.A(n_799),
.B(n_811),
.Y(n_1029)
);

AOI21x1_ASAP7_75t_L g1030 ( 
.A1(n_776),
.A2(n_879),
.B(n_870),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_L g1031 ( 
.A(n_886),
.B(n_938),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_801),
.A2(n_833),
.B(n_838),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_777),
.A2(n_889),
.B(n_776),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_857),
.B(n_862),
.Y(n_1034)
);

NOR2xp33_ASAP7_75t_L g1035 ( 
.A(n_862),
.B(n_785),
.Y(n_1035)
);

INVx3_ASAP7_75t_L g1036 ( 
.A(n_852),
.Y(n_1036)
);

AOI22xp5_ASAP7_75t_L g1037 ( 
.A1(n_854),
.A2(n_930),
.B1(n_960),
.B2(n_961),
.Y(n_1037)
);

HB1xp67_ASAP7_75t_L g1038 ( 
.A(n_890),
.Y(n_1038)
);

NOR2xp67_ASAP7_75t_L g1039 ( 
.A(n_946),
.B(n_952),
.Y(n_1039)
);

INVxp67_ASAP7_75t_L g1040 ( 
.A(n_820),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_782),
.A2(n_891),
.B(n_853),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_902),
.Y(n_1042)
);

INVx3_ASAP7_75t_L g1043 ( 
.A(n_852),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_908),
.Y(n_1044)
);

INVxp67_ASAP7_75t_L g1045 ( 
.A(n_827),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_R g1046 ( 
.A(n_811),
.B(n_852),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_954),
.B(n_890),
.Y(n_1047)
);

INVx1_ASAP7_75t_SL g1048 ( 
.A(n_943),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_948),
.A2(n_789),
.B(n_873),
.Y(n_1049)
);

OAI22xp5_ASAP7_75t_L g1050 ( 
.A1(n_934),
.A2(n_842),
.B1(n_873),
.B2(n_856),
.Y(n_1050)
);

NAND2x1p5_ASAP7_75t_L g1051 ( 
.A(n_885),
.B(n_963),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_845),
.B(n_957),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_948),
.A2(n_789),
.B(n_821),
.Y(n_1053)
);

O2A1O1Ixp5_ASAP7_75t_L g1054 ( 
.A1(n_959),
.A2(n_824),
.B(n_884),
.C(n_835),
.Y(n_1054)
);

O2A1O1Ixp33_ASAP7_75t_L g1055 ( 
.A1(n_872),
.A2(n_877),
.B(n_876),
.C(n_808),
.Y(n_1055)
);

A2O1A1Ixp33_ASAP7_75t_L g1056 ( 
.A1(n_933),
.A2(n_957),
.B(n_793),
.C(n_845),
.Y(n_1056)
);

BUFx2_ASAP7_75t_L g1057 ( 
.A(n_943),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_SL g1058 ( 
.A(n_885),
.B(n_963),
.Y(n_1058)
);

NOR2xp33_ASAP7_75t_SL g1059 ( 
.A(n_794),
.B(n_944),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_SL g1060 ( 
.A(n_885),
.B(n_955),
.Y(n_1060)
);

A2O1A1Ixp33_ASAP7_75t_L g1061 ( 
.A1(n_921),
.A2(n_931),
.B(n_956),
.C(n_951),
.Y(n_1061)
);

CKINVDCx10_ASAP7_75t_R g1062 ( 
.A(n_953),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_935),
.B(n_918),
.Y(n_1063)
);

INVx2_ASAP7_75t_SL g1064 ( 
.A(n_953),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_829),
.A2(n_940),
.B(n_814),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_L g1066 ( 
.A(n_861),
.B(n_781),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_918),
.B(n_790),
.Y(n_1067)
);

A2O1A1Ixp33_ASAP7_75t_L g1068 ( 
.A1(n_912),
.A2(n_806),
.B(n_958),
.C(n_826),
.Y(n_1068)
);

BUFx3_ASAP7_75t_L g1069 ( 
.A(n_859),
.Y(n_1069)
);

AOI22xp33_ASAP7_75t_L g1070 ( 
.A1(n_894),
.A2(n_937),
.B1(n_950),
.B2(n_914),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_942),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_913),
.Y(n_1072)
);

O2A1O1Ixp33_ASAP7_75t_L g1073 ( 
.A1(n_925),
.A2(n_819),
.B(n_808),
.C(n_850),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_913),
.B(n_937),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_914),
.B(n_947),
.Y(n_1075)
);

OAI21x1_ASAP7_75t_L g1076 ( 
.A1(n_804),
.A2(n_807),
.B(n_809),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_812),
.A2(n_813),
.B(n_818),
.Y(n_1077)
);

BUFx6f_ASAP7_75t_L g1078 ( 
.A(n_846),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_L g1079 ( 
.A(n_947),
.B(n_950),
.Y(n_1079)
);

AND2x2_ASAP7_75t_L g1080 ( 
.A(n_846),
.B(n_924),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_834),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_SL g1082 ( 
.A(n_855),
.B(n_837),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_840),
.B(n_841),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_878),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_855),
.Y(n_1085)
);

O2A1O1Ixp33_ASAP7_75t_L g1086 ( 
.A1(n_819),
.A2(n_810),
.B(n_881),
.C(n_892),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_887),
.B(n_895),
.Y(n_1087)
);

NOR2xp33_ASAP7_75t_SL g1088 ( 
.A(n_949),
.B(n_945),
.Y(n_1088)
);

NOR2xp33_ASAP7_75t_R g1089 ( 
.A(n_962),
.B(n_909),
.Y(n_1089)
);

AND2x2_ASAP7_75t_L g1090 ( 
.A(n_936),
.B(n_917),
.Y(n_1090)
);

OAI22xp5_ASAP7_75t_L g1091 ( 
.A1(n_897),
.A2(n_847),
.B1(n_863),
.B2(n_866),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_922),
.Y(n_1092)
);

OAI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_911),
.A2(n_932),
.B(n_927),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_867),
.A2(n_898),
.B(n_904),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_910),
.Y(n_1095)
);

BUFx2_ASAP7_75t_L g1096 ( 
.A(n_906),
.Y(n_1096)
);

BUFx6f_ASAP7_75t_L g1097 ( 
.A(n_791),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_851),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_851),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_822),
.B(n_620),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_816),
.A2(n_621),
.B(n_869),
.Y(n_1101)
);

INVx3_ASAP7_75t_L g1102 ( 
.A(n_791),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_816),
.A2(n_621),
.B(n_869),
.Y(n_1103)
);

BUFx6f_ASAP7_75t_L g1104 ( 
.A(n_791),
.Y(n_1104)
);

AOI221xp5_ASAP7_75t_L g1105 ( 
.A1(n_783),
.A2(n_822),
.B1(n_620),
.B2(n_774),
.C(n_916),
.Y(n_1105)
);

INVx4_ASAP7_75t_L g1106 ( 
.A(n_791),
.Y(n_1106)
);

NOR2xp33_ASAP7_75t_L g1107 ( 
.A(n_822),
.B(n_620),
.Y(n_1107)
);

O2A1O1Ixp33_ASAP7_75t_L g1108 ( 
.A1(n_816),
.A2(n_822),
.B(n_774),
.C(n_620),
.Y(n_1108)
);

O2A1O1Ixp33_ASAP7_75t_L g1109 ( 
.A1(n_816),
.A2(n_822),
.B(n_774),
.C(n_620),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_787),
.B(n_387),
.Y(n_1110)
);

AO31x2_ASAP7_75t_L g1111 ( 
.A1(n_967),
.A2(n_1100),
.A3(n_1107),
.B(n_1041),
.Y(n_1111)
);

AOI31xp67_ASAP7_75t_L g1112 ( 
.A1(n_971),
.A2(n_1095),
.A3(n_1060),
.B(n_1034),
.Y(n_1112)
);

NAND3xp33_ASAP7_75t_L g1113 ( 
.A(n_982),
.B(n_1105),
.C(n_1012),
.Y(n_1113)
);

O2A1O1Ixp33_ASAP7_75t_SL g1114 ( 
.A1(n_1010),
.A2(n_1105),
.B(n_1108),
.C(n_1109),
.Y(n_1114)
);

OAI21x1_ASAP7_75t_SL g1115 ( 
.A1(n_1055),
.A2(n_1067),
.B(n_1015),
.Y(n_1115)
);

O2A1O1Ixp5_ASAP7_75t_L g1116 ( 
.A1(n_1101),
.A2(n_1103),
.B(n_1032),
.C(n_1052),
.Y(n_1116)
);

AOI221x1_ASAP7_75t_L g1117 ( 
.A1(n_1004),
.A2(n_1015),
.B1(n_1103),
.B2(n_1101),
.C(n_1032),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_1110),
.B(n_1017),
.Y(n_1118)
);

OAI21x1_ASAP7_75t_L g1119 ( 
.A1(n_976),
.A2(n_1094),
.B(n_1076),
.Y(n_1119)
);

BUFx2_ASAP7_75t_L g1120 ( 
.A(n_995),
.Y(n_1120)
);

AO31x2_ASAP7_75t_L g1121 ( 
.A1(n_1041),
.A2(n_1068),
.A3(n_1056),
.B(n_1025),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_1016),
.A2(n_1077),
.B(n_1025),
.Y(n_1122)
);

BUFx6f_ASAP7_75t_L g1123 ( 
.A(n_964),
.Y(n_1123)
);

NOR2xp67_ASAP7_75t_L g1124 ( 
.A(n_1040),
.B(n_1045),
.Y(n_1124)
);

OAI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_1049),
.A2(n_1053),
.B(n_1050),
.Y(n_1125)
);

AOI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_1059),
.A2(n_1037),
.B1(n_1028),
.B2(n_1031),
.Y(n_1126)
);

OA21x2_ASAP7_75t_L g1127 ( 
.A1(n_1054),
.A2(n_1016),
.B(n_1033),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_1077),
.A2(n_1065),
.B(n_1053),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_1065),
.A2(n_1091),
.B(n_1086),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_980),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_1033),
.A2(n_1088),
.B(n_1094),
.Y(n_1131)
);

OR2x2_ASAP7_75t_L g1132 ( 
.A(n_1047),
.B(n_978),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_1018),
.Y(n_1133)
);

AO31x2_ASAP7_75t_L g1134 ( 
.A1(n_972),
.A2(n_1061),
.A3(n_1049),
.B(n_965),
.Y(n_1134)
);

AOI21xp33_ASAP7_75t_L g1135 ( 
.A1(n_1022),
.A2(n_1055),
.B(n_1063),
.Y(n_1135)
);

AO31x2_ASAP7_75t_L g1136 ( 
.A1(n_965),
.A2(n_1092),
.A3(n_968),
.B(n_966),
.Y(n_1136)
);

A2O1A1Ixp33_ASAP7_75t_L g1137 ( 
.A1(n_989),
.A2(n_1026),
.B(n_987),
.C(n_1073),
.Y(n_1137)
);

HB1xp67_ASAP7_75t_L g1138 ( 
.A(n_973),
.Y(n_1138)
);

OAI21x1_ASAP7_75t_L g1139 ( 
.A1(n_976),
.A2(n_1093),
.B(n_966),
.Y(n_1139)
);

AOI221x1_ASAP7_75t_L g1140 ( 
.A1(n_1007),
.A2(n_991),
.B1(n_1002),
.B2(n_1005),
.C(n_1035),
.Y(n_1140)
);

BUFx8_ASAP7_75t_L g1141 ( 
.A(n_984),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1098),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_1099),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_1083),
.A2(n_1087),
.B(n_1058),
.Y(n_1144)
);

AO31x2_ASAP7_75t_L g1145 ( 
.A1(n_968),
.A2(n_1002),
.A3(n_1007),
.B(n_1096),
.Y(n_1145)
);

OAI21x1_ASAP7_75t_L g1146 ( 
.A1(n_1030),
.A2(n_1090),
.B(n_977),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1071),
.B(n_1020),
.Y(n_1147)
);

OA21x2_ASAP7_75t_L g1148 ( 
.A1(n_969),
.A2(n_994),
.B(n_1029),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_1082),
.A2(n_1080),
.B(n_1084),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_974),
.B(n_970),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_1081),
.A2(n_1051),
.B(n_1066),
.Y(n_1151)
);

AO21x2_ASAP7_75t_L g1152 ( 
.A1(n_1089),
.A2(n_1001),
.B(n_1046),
.Y(n_1152)
);

AO32x2_ASAP7_75t_L g1153 ( 
.A1(n_1064),
.A2(n_1003),
.A3(n_992),
.B1(n_1011),
.B2(n_990),
.Y(n_1153)
);

O2A1O1Ixp33_ASAP7_75t_L g1154 ( 
.A1(n_985),
.A2(n_1006),
.B(n_988),
.C(n_1027),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_1042),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1023),
.Y(n_1156)
);

CKINVDCx11_ASAP7_75t_R g1157 ( 
.A(n_996),
.Y(n_1157)
);

AND2x6_ASAP7_75t_L g1158 ( 
.A(n_1078),
.B(n_964),
.Y(n_1158)
);

NOR2xp33_ASAP7_75t_L g1159 ( 
.A(n_1038),
.B(n_1048),
.Y(n_1159)
);

AOI22xp5_ASAP7_75t_L g1160 ( 
.A1(n_1000),
.A2(n_1039),
.B1(n_986),
.B2(n_1021),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1024),
.B(n_979),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_979),
.B(n_1044),
.Y(n_1162)
);

INVx4_ASAP7_75t_L g1163 ( 
.A(n_964),
.Y(n_1163)
);

INVx3_ASAP7_75t_SL g1164 ( 
.A(n_1013),
.Y(n_1164)
);

AOI221xp5_ASAP7_75t_SL g1165 ( 
.A1(n_1009),
.A2(n_1014),
.B1(n_1072),
.B2(n_1070),
.C(n_1057),
.Y(n_1165)
);

AOI21x1_ASAP7_75t_SL g1166 ( 
.A1(n_1008),
.A2(n_1074),
.B(n_1075),
.Y(n_1166)
);

OAI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_1051),
.A2(n_1079),
.B1(n_1078),
.B2(n_993),
.Y(n_1167)
);

BUFx3_ASAP7_75t_L g1168 ( 
.A(n_1008),
.Y(n_1168)
);

HB1xp67_ASAP7_75t_L g1169 ( 
.A(n_1069),
.Y(n_1169)
);

NOR2xp33_ASAP7_75t_L g1170 ( 
.A(n_1062),
.B(n_1085),
.Y(n_1170)
);

INVx4_ASAP7_75t_L g1171 ( 
.A(n_997),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_977),
.A2(n_1019),
.B(n_998),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_1019),
.Y(n_1173)
);

A2O1A1Ixp33_ASAP7_75t_L g1174 ( 
.A1(n_975),
.A2(n_1036),
.B(n_1043),
.C(n_1102),
.Y(n_1174)
);

OR2x6_ASAP7_75t_L g1175 ( 
.A(n_981),
.B(n_1104),
.Y(n_1175)
);

AND2x2_ASAP7_75t_L g1176 ( 
.A(n_981),
.B(n_975),
.Y(n_1176)
);

OAI21x1_ASAP7_75t_L g1177 ( 
.A1(n_999),
.A2(n_1043),
.B(n_1102),
.Y(n_1177)
);

BUFx6f_ASAP7_75t_SL g1178 ( 
.A(n_981),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1106),
.A2(n_1036),
.B(n_997),
.Y(n_1179)
);

BUFx3_ASAP7_75t_L g1180 ( 
.A(n_997),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_1106),
.A2(n_1097),
.B(n_1104),
.Y(n_1181)
);

INVx4_ASAP7_75t_L g1182 ( 
.A(n_1097),
.Y(n_1182)
);

NOR2xp67_ASAP7_75t_L g1183 ( 
.A(n_1097),
.B(n_1104),
.Y(n_1183)
);

OAI21x1_ASAP7_75t_L g1184 ( 
.A1(n_1011),
.A2(n_976),
.B(n_1094),
.Y(n_1184)
);

INVx5_ASAP7_75t_L g1185 ( 
.A(n_1011),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_983),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1101),
.A2(n_1103),
.B(n_816),
.Y(n_1187)
);

O2A1O1Ixp5_ASAP7_75t_SL g1188 ( 
.A1(n_1060),
.A2(n_637),
.B(n_641),
.C(n_828),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_1101),
.A2(n_1103),
.B(n_816),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_SL g1190 ( 
.A(n_1017),
.B(n_1110),
.Y(n_1190)
);

NOR2x1_ASAP7_75t_R g1191 ( 
.A(n_984),
.B(n_669),
.Y(n_1191)
);

NAND2xp33_ASAP7_75t_L g1192 ( 
.A(n_1012),
.B(n_816),
.Y(n_1192)
);

INVx2_ASAP7_75t_L g1193 ( 
.A(n_980),
.Y(n_1193)
);

INVx5_ASAP7_75t_L g1194 ( 
.A(n_964),
.Y(n_1194)
);

AOI31xp67_ASAP7_75t_L g1195 ( 
.A1(n_971),
.A2(n_1095),
.A3(n_637),
.B(n_641),
.Y(n_1195)
);

AO31x2_ASAP7_75t_L g1196 ( 
.A1(n_967),
.A2(n_1107),
.A3(n_1100),
.B(n_1041),
.Y(n_1196)
);

A2O1A1Ixp33_ASAP7_75t_L g1197 ( 
.A1(n_1100),
.A2(n_816),
.B(n_1107),
.C(n_822),
.Y(n_1197)
);

OAI22x1_ASAP7_75t_L g1198 ( 
.A1(n_982),
.A2(n_1100),
.B1(n_1107),
.B2(n_971),
.Y(n_1198)
);

NAND2x1p5_ASAP7_75t_L g1199 ( 
.A(n_973),
.B(n_811),
.Y(n_1199)
);

CKINVDCx11_ASAP7_75t_R g1200 ( 
.A(n_996),
.Y(n_1200)
);

AO31x2_ASAP7_75t_L g1201 ( 
.A1(n_967),
.A2(n_1107),
.A3(n_1100),
.B(n_1041),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1101),
.A2(n_1103),
.B(n_816),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1101),
.A2(n_1103),
.B(n_816),
.Y(n_1203)
);

OAI21x1_ASAP7_75t_L g1204 ( 
.A1(n_976),
.A2(n_1094),
.B(n_1076),
.Y(n_1204)
);

AO31x2_ASAP7_75t_L g1205 ( 
.A1(n_967),
.A2(n_1107),
.A3(n_1100),
.B(n_1041),
.Y(n_1205)
);

OR2x2_ASAP7_75t_L g1206 ( 
.A(n_1110),
.B(n_453),
.Y(n_1206)
);

NAND3xp33_ASAP7_75t_L g1207 ( 
.A(n_982),
.B(n_816),
.C(n_1105),
.Y(n_1207)
);

AO21x1_ASAP7_75t_L g1208 ( 
.A1(n_1100),
.A2(n_1107),
.B(n_1108),
.Y(n_1208)
);

OAI21xp5_ASAP7_75t_SL g1209 ( 
.A1(n_1012),
.A2(n_783),
.B(n_387),
.Y(n_1209)
);

NOR2x1_ASAP7_75t_SL g1210 ( 
.A(n_1058),
.B(n_960),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_980),
.Y(n_1211)
);

OAI22xp5_ASAP7_75t_L g1212 ( 
.A1(n_1012),
.A2(n_816),
.B1(n_1107),
.B2(n_1100),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1101),
.A2(n_1103),
.B(n_816),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_980),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_980),
.Y(n_1215)
);

AOI22xp33_ASAP7_75t_SL g1216 ( 
.A1(n_982),
.A2(n_760),
.B1(n_310),
.B2(n_330),
.Y(n_1216)
);

A2O1A1Ixp33_ASAP7_75t_L g1217 ( 
.A1(n_1100),
.A2(n_816),
.B(n_1107),
.C(n_822),
.Y(n_1217)
);

AO21x1_ASAP7_75t_L g1218 ( 
.A1(n_1100),
.A2(n_1107),
.B(n_1108),
.Y(n_1218)
);

AO21x2_ASAP7_75t_L g1219 ( 
.A1(n_1041),
.A2(n_1016),
.B(n_1025),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_980),
.Y(n_1220)
);

OAI21x1_ASAP7_75t_L g1221 ( 
.A1(n_976),
.A2(n_1094),
.B(n_1076),
.Y(n_1221)
);

OR2x2_ASAP7_75t_L g1222 ( 
.A(n_1110),
.B(n_453),
.Y(n_1222)
);

AO32x2_ASAP7_75t_L g1223 ( 
.A1(n_1050),
.A2(n_1005),
.A3(n_926),
.B1(n_1091),
.B2(n_1064),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_971),
.B(n_620),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_980),
.Y(n_1225)
);

BUFx10_ASAP7_75t_L g1226 ( 
.A(n_1017),
.Y(n_1226)
);

AOI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1101),
.A2(n_1103),
.B(n_816),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1101),
.A2(n_1103),
.B(n_816),
.Y(n_1228)
);

AO31x2_ASAP7_75t_L g1229 ( 
.A1(n_967),
.A2(n_1107),
.A3(n_1100),
.B(n_1041),
.Y(n_1229)
);

OAI22xp5_ASAP7_75t_L g1230 ( 
.A1(n_1012),
.A2(n_816),
.B1(n_1107),
.B2(n_1100),
.Y(n_1230)
);

INVx4_ASAP7_75t_L g1231 ( 
.A(n_964),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1101),
.A2(n_1103),
.B(n_816),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1101),
.A2(n_1103),
.B(n_816),
.Y(n_1233)
);

O2A1O1Ixp33_ASAP7_75t_SL g1234 ( 
.A1(n_1010),
.A2(n_816),
.B(n_1107),
.C(n_1100),
.Y(n_1234)
);

BUFx6f_ASAP7_75t_L g1235 ( 
.A(n_964),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_971),
.B(n_620),
.Y(n_1236)
);

A2O1A1Ixp33_ASAP7_75t_L g1237 ( 
.A1(n_1100),
.A2(n_816),
.B(n_1107),
.C(n_822),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1101),
.A2(n_1103),
.B(n_816),
.Y(n_1238)
);

OR2x2_ASAP7_75t_L g1239 ( 
.A(n_1110),
.B(n_453),
.Y(n_1239)
);

OAI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1100),
.A2(n_816),
.B(n_1107),
.Y(n_1240)
);

CKINVDCx16_ASAP7_75t_R g1241 ( 
.A(n_996),
.Y(n_1241)
);

CKINVDCx20_ASAP7_75t_R g1242 ( 
.A(n_996),
.Y(n_1242)
);

OAI21x1_ASAP7_75t_L g1243 ( 
.A1(n_976),
.A2(n_1094),
.B(n_1076),
.Y(n_1243)
);

OAI21x1_ASAP7_75t_L g1244 ( 
.A1(n_976),
.A2(n_1094),
.B(n_1076),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1101),
.A2(n_1103),
.B(n_816),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_980),
.Y(n_1246)
);

INVxp67_ASAP7_75t_L g1247 ( 
.A(n_995),
.Y(n_1247)
);

OAI21x1_ASAP7_75t_L g1248 ( 
.A1(n_976),
.A2(n_1094),
.B(n_1076),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_980),
.Y(n_1249)
);

INVx4_ASAP7_75t_L g1250 ( 
.A(n_964),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_976),
.A2(n_1094),
.B(n_1076),
.Y(n_1251)
);

BUFx2_ASAP7_75t_L g1252 ( 
.A(n_995),
.Y(n_1252)
);

NAND3xp33_ASAP7_75t_L g1253 ( 
.A(n_982),
.B(n_816),
.C(n_1105),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_980),
.Y(n_1254)
);

AOI22xp33_ASAP7_75t_L g1255 ( 
.A1(n_1113),
.A2(n_1192),
.B1(n_1207),
.B2(n_1253),
.Y(n_1255)
);

BUFx6f_ASAP7_75t_L g1256 ( 
.A(n_1194),
.Y(n_1256)
);

OAI22xp5_ASAP7_75t_L g1257 ( 
.A1(n_1216),
.A2(n_1126),
.B1(n_1118),
.B2(n_1236),
.Y(n_1257)
);

AOI22xp33_ASAP7_75t_L g1258 ( 
.A1(n_1212),
.A2(n_1230),
.B1(n_1198),
.B2(n_1240),
.Y(n_1258)
);

BUFx8_ASAP7_75t_L g1259 ( 
.A(n_1178),
.Y(n_1259)
);

AOI22xp33_ASAP7_75t_L g1260 ( 
.A1(n_1224),
.A2(n_1208),
.B1(n_1218),
.B2(n_1135),
.Y(n_1260)
);

AOI22xp33_ASAP7_75t_L g1261 ( 
.A1(n_1190),
.A2(n_1132),
.B1(n_1125),
.B2(n_1156),
.Y(n_1261)
);

AOI22xp33_ASAP7_75t_SL g1262 ( 
.A1(n_1178),
.A2(n_1226),
.B1(n_1209),
.B2(n_1210),
.Y(n_1262)
);

OAI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1197),
.A2(n_1217),
.B(n_1237),
.Y(n_1263)
);

OAI22xp5_ASAP7_75t_L g1264 ( 
.A1(n_1147),
.A2(n_1206),
.B1(n_1222),
.B2(n_1239),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_SL g1265 ( 
.A1(n_1226),
.A2(n_1150),
.B1(n_1168),
.B2(n_1156),
.Y(n_1265)
);

OAI22xp5_ASAP7_75t_L g1266 ( 
.A1(n_1160),
.A2(n_1137),
.B1(n_1124),
.B2(n_1175),
.Y(n_1266)
);

BUFx2_ASAP7_75t_L g1267 ( 
.A(n_1120),
.Y(n_1267)
);

CKINVDCx6p67_ASAP7_75t_R g1268 ( 
.A(n_1164),
.Y(n_1268)
);

INVx1_ASAP7_75t_SL g1269 ( 
.A(n_1252),
.Y(n_1269)
);

AOI22xp33_ASAP7_75t_SL g1270 ( 
.A1(n_1185),
.A2(n_1187),
.B1(n_1213),
.B2(n_1238),
.Y(n_1270)
);

CKINVDCx11_ASAP7_75t_R g1271 ( 
.A(n_1157),
.Y(n_1271)
);

CKINVDCx11_ASAP7_75t_R g1272 ( 
.A(n_1200),
.Y(n_1272)
);

AOI22xp33_ASAP7_75t_L g1273 ( 
.A1(n_1161),
.A2(n_1162),
.B1(n_1233),
.B2(n_1245),
.Y(n_1273)
);

AOI22xp33_ASAP7_75t_SL g1274 ( 
.A1(n_1185),
.A2(n_1189),
.B1(n_1228),
.B2(n_1232),
.Y(n_1274)
);

BUFx4f_ASAP7_75t_SL g1275 ( 
.A(n_1141),
.Y(n_1275)
);

OAI22xp33_ASAP7_75t_L g1276 ( 
.A1(n_1140),
.A2(n_1175),
.B1(n_1249),
.B2(n_1143),
.Y(n_1276)
);

INVx2_ASAP7_75t_SL g1277 ( 
.A(n_1138),
.Y(n_1277)
);

OAI22xp5_ASAP7_75t_L g1278 ( 
.A1(n_1247),
.A2(n_1159),
.B1(n_1154),
.B2(n_1151),
.Y(n_1278)
);

OAI22xp5_ASAP7_75t_L g1279 ( 
.A1(n_1169),
.A2(n_1149),
.B1(n_1246),
.B2(n_1155),
.Y(n_1279)
);

INVx1_ASAP7_75t_SL g1280 ( 
.A(n_1242),
.Y(n_1280)
);

BUFx6f_ASAP7_75t_L g1281 ( 
.A(n_1194),
.Y(n_1281)
);

BUFx12f_ASAP7_75t_L g1282 ( 
.A(n_1141),
.Y(n_1282)
);

INVx4_ASAP7_75t_L g1283 ( 
.A(n_1194),
.Y(n_1283)
);

CKINVDCx5p33_ASAP7_75t_R g1284 ( 
.A(n_1241),
.Y(n_1284)
);

BUFx2_ASAP7_75t_SL g1285 ( 
.A(n_1183),
.Y(n_1285)
);

BUFx2_ASAP7_75t_L g1286 ( 
.A(n_1180),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1225),
.Y(n_1287)
);

AOI22xp5_ASAP7_75t_L g1288 ( 
.A1(n_1170),
.A2(n_1186),
.B1(n_1234),
.B2(n_1176),
.Y(n_1288)
);

INVx1_ASAP7_75t_SL g1289 ( 
.A(n_1199),
.Y(n_1289)
);

OAI22xp5_ASAP7_75t_L g1290 ( 
.A1(n_1193),
.A2(n_1211),
.B1(n_1254),
.B2(n_1220),
.Y(n_1290)
);

OAI22xp33_ASAP7_75t_L g1291 ( 
.A1(n_1130),
.A2(n_1214),
.B1(n_1215),
.B2(n_1185),
.Y(n_1291)
);

INVx4_ASAP7_75t_L g1292 ( 
.A(n_1158),
.Y(n_1292)
);

INVx6_ASAP7_75t_L g1293 ( 
.A(n_1163),
.Y(n_1293)
);

AOI22xp5_ASAP7_75t_L g1294 ( 
.A1(n_1186),
.A2(n_1152),
.B1(n_1165),
.B2(n_1167),
.Y(n_1294)
);

AOI22xp33_ASAP7_75t_L g1295 ( 
.A1(n_1202),
.A2(n_1227),
.B1(n_1203),
.B2(n_1115),
.Y(n_1295)
);

HB1xp67_ASAP7_75t_L g1296 ( 
.A(n_1134),
.Y(n_1296)
);

AOI22xp5_ASAP7_75t_L g1297 ( 
.A1(n_1114),
.A2(n_1144),
.B1(n_1173),
.B2(n_1158),
.Y(n_1297)
);

BUFx2_ASAP7_75t_L g1298 ( 
.A(n_1123),
.Y(n_1298)
);

CKINVDCx20_ASAP7_75t_R g1299 ( 
.A(n_1235),
.Y(n_1299)
);

AOI22xp33_ASAP7_75t_SL g1300 ( 
.A1(n_1129),
.A2(n_1153),
.B1(n_1131),
.B2(n_1223),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1112),
.Y(n_1301)
);

BUFx2_ASAP7_75t_L g1302 ( 
.A(n_1235),
.Y(n_1302)
);

AOI22xp33_ASAP7_75t_L g1303 ( 
.A1(n_1219),
.A2(n_1127),
.B1(n_1148),
.B2(n_1128),
.Y(n_1303)
);

CKINVDCx6p67_ASAP7_75t_R g1304 ( 
.A(n_1163),
.Y(n_1304)
);

OAI22xp33_ASAP7_75t_L g1305 ( 
.A1(n_1117),
.A2(n_1153),
.B1(n_1148),
.B2(n_1223),
.Y(n_1305)
);

CKINVDCx6p67_ASAP7_75t_R g1306 ( 
.A(n_1171),
.Y(n_1306)
);

CKINVDCx20_ASAP7_75t_R g1307 ( 
.A(n_1171),
.Y(n_1307)
);

CKINVDCx5p33_ASAP7_75t_R g1308 ( 
.A(n_1182),
.Y(n_1308)
);

OAI21xp5_ASAP7_75t_SL g1309 ( 
.A1(n_1122),
.A2(n_1153),
.B(n_1223),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_1177),
.Y(n_1310)
);

BUFx10_ASAP7_75t_L g1311 ( 
.A(n_1191),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_SL g1312 ( 
.A(n_1116),
.B(n_1172),
.Y(n_1312)
);

BUFx6f_ASAP7_75t_L g1313 ( 
.A(n_1182),
.Y(n_1313)
);

OAI22xp33_ASAP7_75t_L g1314 ( 
.A1(n_1127),
.A2(n_1250),
.B1(n_1231),
.B2(n_1179),
.Y(n_1314)
);

AOI22xp5_ASAP7_75t_L g1315 ( 
.A1(n_1231),
.A2(n_1250),
.B1(n_1174),
.B2(n_1181),
.Y(n_1315)
);

BUFx2_ASAP7_75t_L g1316 ( 
.A(n_1134),
.Y(n_1316)
);

BUFx2_ASAP7_75t_L g1317 ( 
.A(n_1111),
.Y(n_1317)
);

BUFx3_ASAP7_75t_L g1318 ( 
.A(n_1196),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_1166),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1196),
.B(n_1201),
.Y(n_1320)
);

INVx6_ASAP7_75t_L g1321 ( 
.A(n_1188),
.Y(n_1321)
);

AOI22xp33_ASAP7_75t_L g1322 ( 
.A1(n_1139),
.A2(n_1184),
.B1(n_1146),
.B2(n_1204),
.Y(n_1322)
);

BUFx6f_ASAP7_75t_L g1323 ( 
.A(n_1119),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1221),
.A2(n_1251),
.B1(n_1248),
.B2(n_1244),
.Y(n_1324)
);

OAI22xp5_ASAP7_75t_L g1325 ( 
.A1(n_1196),
.A2(n_1201),
.B1(n_1229),
.B2(n_1205),
.Y(n_1325)
);

AOI22xp33_ASAP7_75t_L g1326 ( 
.A1(n_1243),
.A2(n_1201),
.B1(n_1205),
.B2(n_1229),
.Y(n_1326)
);

AOI22xp33_ASAP7_75t_L g1327 ( 
.A1(n_1229),
.A2(n_1121),
.B1(n_1145),
.B2(n_1195),
.Y(n_1327)
);

CKINVDCx11_ASAP7_75t_R g1328 ( 
.A(n_1145),
.Y(n_1328)
);

OAI22xp5_ASAP7_75t_L g1329 ( 
.A1(n_1121),
.A2(n_1136),
.B1(n_1216),
.B2(n_1012),
.Y(n_1329)
);

AOI22xp5_ASAP7_75t_L g1330 ( 
.A1(n_1121),
.A2(n_1216),
.B1(n_982),
.B2(n_1059),
.Y(n_1330)
);

AOI22xp33_ASAP7_75t_L g1331 ( 
.A1(n_1113),
.A2(n_783),
.B1(n_982),
.B2(n_1100),
.Y(n_1331)
);

INVx6_ASAP7_75t_L g1332 ( 
.A(n_1194),
.Y(n_1332)
);

AOI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1113),
.A2(n_783),
.B1(n_982),
.B2(n_1100),
.Y(n_1333)
);

AOI22xp33_ASAP7_75t_SL g1334 ( 
.A1(n_1113),
.A2(n_982),
.B1(n_1192),
.B2(n_391),
.Y(n_1334)
);

CKINVDCx20_ASAP7_75t_R g1335 ( 
.A(n_1157),
.Y(n_1335)
);

OAI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1113),
.A2(n_971),
.B1(n_1209),
.B2(n_1253),
.Y(n_1336)
);

OAI22xp5_ASAP7_75t_L g1337 ( 
.A1(n_1216),
.A2(n_1012),
.B1(n_1126),
.B2(n_1113),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1133),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1142),
.Y(n_1339)
);

AOI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1113),
.A2(n_783),
.B1(n_982),
.B2(n_1100),
.Y(n_1340)
);

OAI22xp33_ASAP7_75t_L g1341 ( 
.A1(n_1113),
.A2(n_971),
.B1(n_1209),
.B2(n_1253),
.Y(n_1341)
);

OAI22xp33_ASAP7_75t_L g1342 ( 
.A1(n_1113),
.A2(n_971),
.B1(n_1209),
.B2(n_1253),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1142),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_L g1344 ( 
.A1(n_1113),
.A2(n_783),
.B1(n_982),
.B2(n_1100),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1133),
.Y(n_1345)
);

INVx4_ASAP7_75t_L g1346 ( 
.A(n_1194),
.Y(n_1346)
);

AOI22xp33_ASAP7_75t_L g1347 ( 
.A1(n_1113),
.A2(n_783),
.B1(n_982),
.B2(n_1100),
.Y(n_1347)
);

INVx6_ASAP7_75t_L g1348 ( 
.A(n_1194),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1118),
.B(n_620),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_L g1350 ( 
.A1(n_1113),
.A2(n_783),
.B1(n_982),
.B2(n_1100),
.Y(n_1350)
);

AOI22xp33_ASAP7_75t_L g1351 ( 
.A1(n_1113),
.A2(n_783),
.B1(n_982),
.B2(n_1100),
.Y(n_1351)
);

CKINVDCx20_ASAP7_75t_R g1352 ( 
.A(n_1157),
.Y(n_1352)
);

BUFx3_ASAP7_75t_L g1353 ( 
.A(n_1164),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1118),
.B(n_620),
.Y(n_1354)
);

AOI22xp33_ASAP7_75t_SL g1355 ( 
.A1(n_1113),
.A2(n_982),
.B1(n_1192),
.B2(n_391),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1113),
.A2(n_783),
.B1(n_982),
.B2(n_1100),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_L g1357 ( 
.A1(n_1113),
.A2(n_783),
.B1(n_982),
.B2(n_1100),
.Y(n_1357)
);

AOI22xp33_ASAP7_75t_L g1358 ( 
.A1(n_1113),
.A2(n_783),
.B1(n_982),
.B2(n_1100),
.Y(n_1358)
);

OAI22xp5_ASAP7_75t_L g1359 ( 
.A1(n_1216),
.A2(n_1012),
.B1(n_1126),
.B2(n_1113),
.Y(n_1359)
);

HB1xp67_ASAP7_75t_L g1360 ( 
.A(n_1279),
.Y(n_1360)
);

AND2x4_ASAP7_75t_L g1361 ( 
.A(n_1310),
.B(n_1316),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1296),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1320),
.Y(n_1363)
);

OA21x2_ASAP7_75t_L g1364 ( 
.A1(n_1312),
.A2(n_1309),
.B(n_1303),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1317),
.Y(n_1365)
);

AOI21x1_ASAP7_75t_L g1366 ( 
.A1(n_1312),
.A2(n_1301),
.B(n_1329),
.Y(n_1366)
);

AND2x4_ASAP7_75t_L g1367 ( 
.A(n_1263),
.B(n_1318),
.Y(n_1367)
);

NOR2x1_ASAP7_75t_R g1368 ( 
.A(n_1271),
.B(n_1272),
.Y(n_1368)
);

HB1xp67_ASAP7_75t_L g1369 ( 
.A(n_1267),
.Y(n_1369)
);

HB1xp67_ASAP7_75t_L g1370 ( 
.A(n_1290),
.Y(n_1370)
);

INVxp33_ASAP7_75t_L g1371 ( 
.A(n_1264),
.Y(n_1371)
);

OR2x6_ASAP7_75t_L g1372 ( 
.A(n_1323),
.B(n_1318),
.Y(n_1372)
);

HB1xp67_ASAP7_75t_L g1373 ( 
.A(n_1278),
.Y(n_1373)
);

INVx1_ASAP7_75t_SL g1374 ( 
.A(n_1269),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_L g1375 ( 
.A1(n_1337),
.A2(n_1359),
.B1(n_1334),
.B2(n_1355),
.Y(n_1375)
);

OA21x2_ASAP7_75t_L g1376 ( 
.A1(n_1303),
.A2(n_1327),
.B(n_1326),
.Y(n_1376)
);

INVx3_ASAP7_75t_L g1377 ( 
.A(n_1323),
.Y(n_1377)
);

AOI21x1_ASAP7_75t_L g1378 ( 
.A1(n_1266),
.A2(n_1325),
.B(n_1257),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1287),
.Y(n_1379)
);

INVxp67_ASAP7_75t_R g1380 ( 
.A(n_1275),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1258),
.B(n_1300),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1339),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1343),
.Y(n_1383)
);

OR2x6_ASAP7_75t_L g1384 ( 
.A(n_1292),
.B(n_1321),
.Y(n_1384)
);

OAI21x1_ASAP7_75t_L g1385 ( 
.A1(n_1324),
.A2(n_1322),
.B(n_1295),
.Y(n_1385)
);

BUFx6f_ASAP7_75t_L g1386 ( 
.A(n_1328),
.Y(n_1386)
);

BUFx2_ASAP7_75t_L g1387 ( 
.A(n_1294),
.Y(n_1387)
);

BUFx2_ASAP7_75t_L g1388 ( 
.A(n_1291),
.Y(n_1388)
);

INVx2_ASAP7_75t_SL g1389 ( 
.A(n_1332),
.Y(n_1389)
);

CKINVDCx20_ASAP7_75t_R g1390 ( 
.A(n_1335),
.Y(n_1390)
);

AOI22xp5_ASAP7_75t_L g1391 ( 
.A1(n_1331),
.A2(n_1358),
.B1(n_1356),
.B2(n_1357),
.Y(n_1391)
);

INVx2_ASAP7_75t_L g1392 ( 
.A(n_1321),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1258),
.B(n_1255),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_1321),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1255),
.B(n_1260),
.Y(n_1395)
);

BUFx3_ASAP7_75t_L g1396 ( 
.A(n_1259),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1349),
.B(n_1354),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1305),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1305),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1291),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1273),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1273),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1326),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1295),
.Y(n_1404)
);

BUFx2_ASAP7_75t_L g1405 ( 
.A(n_1276),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1276),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1338),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1345),
.Y(n_1408)
);

OAI21xp5_ASAP7_75t_L g1409 ( 
.A1(n_1333),
.A2(n_1358),
.B(n_1357),
.Y(n_1409)
);

BUFx2_ASAP7_75t_L g1410 ( 
.A(n_1297),
.Y(n_1410)
);

BUFx2_ASAP7_75t_L g1411 ( 
.A(n_1319),
.Y(n_1411)
);

AO21x2_ASAP7_75t_L g1412 ( 
.A1(n_1336),
.A2(n_1342),
.B(n_1341),
.Y(n_1412)
);

HB1xp67_ASAP7_75t_L g1413 ( 
.A(n_1277),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1270),
.Y(n_1414)
);

NAND2x1p5_ASAP7_75t_L g1415 ( 
.A(n_1292),
.B(n_1315),
.Y(n_1415)
);

OR2x2_ASAP7_75t_L g1416 ( 
.A(n_1261),
.B(n_1260),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1274),
.Y(n_1417)
);

AOI21x1_ASAP7_75t_L g1418 ( 
.A1(n_1298),
.A2(n_1302),
.B(n_1286),
.Y(n_1418)
);

INVx4_ASAP7_75t_L g1419 ( 
.A(n_1256),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1314),
.Y(n_1420)
);

BUFx3_ASAP7_75t_L g1421 ( 
.A(n_1259),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1314),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1336),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1341),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1342),
.Y(n_1425)
);

OAI22xp5_ASAP7_75t_L g1426 ( 
.A1(n_1333),
.A2(n_1344),
.B1(n_1340),
.B2(n_1347),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1324),
.Y(n_1427)
);

NAND2x1p5_ASAP7_75t_L g1428 ( 
.A(n_1330),
.B(n_1346),
.Y(n_1428)
);

BUFx2_ASAP7_75t_L g1429 ( 
.A(n_1299),
.Y(n_1429)
);

HB1xp67_ASAP7_75t_L g1430 ( 
.A(n_1289),
.Y(n_1430)
);

AOI21xp5_ASAP7_75t_SL g1431 ( 
.A1(n_1426),
.A2(n_1281),
.B(n_1283),
.Y(n_1431)
);

OR2x6_ASAP7_75t_L g1432 ( 
.A(n_1415),
.B(n_1348),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1367),
.B(n_1265),
.Y(n_1433)
);

NAND3xp33_ASAP7_75t_L g1434 ( 
.A(n_1409),
.B(n_1356),
.C(n_1351),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1373),
.B(n_1351),
.Y(n_1435)
);

AOI221xp5_ASAP7_75t_L g1436 ( 
.A1(n_1375),
.A2(n_1350),
.B1(n_1347),
.B2(n_1344),
.C(n_1340),
.Y(n_1436)
);

OA21x2_ASAP7_75t_L g1437 ( 
.A1(n_1385),
.A2(n_1350),
.B(n_1288),
.Y(n_1437)
);

OAI21xp5_ASAP7_75t_L g1438 ( 
.A1(n_1391),
.A2(n_1424),
.B(n_1423),
.Y(n_1438)
);

A2O1A1Ixp33_ASAP7_75t_L g1439 ( 
.A1(n_1393),
.A2(n_1262),
.B(n_1281),
.C(n_1285),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_1382),
.Y(n_1440)
);

AOI221xp5_ASAP7_75t_L g1441 ( 
.A1(n_1423),
.A2(n_1353),
.B1(n_1280),
.B2(n_1284),
.C(n_1308),
.Y(n_1441)
);

CKINVDCx5p33_ASAP7_75t_R g1442 ( 
.A(n_1390),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1367),
.B(n_1386),
.Y(n_1443)
);

OR2x2_ASAP7_75t_L g1444 ( 
.A(n_1363),
.B(n_1268),
.Y(n_1444)
);

AO32x2_ASAP7_75t_L g1445 ( 
.A1(n_1398),
.A2(n_1399),
.A3(n_1389),
.B1(n_1363),
.B2(n_1419),
.Y(n_1445)
);

NOR2xp33_ASAP7_75t_L g1446 ( 
.A(n_1371),
.B(n_1307),
.Y(n_1446)
);

OAI22xp5_ASAP7_75t_L g1447 ( 
.A1(n_1411),
.A2(n_1306),
.B1(n_1304),
.B2(n_1348),
.Y(n_1447)
);

A2O1A1Ixp33_ASAP7_75t_L g1448 ( 
.A1(n_1393),
.A2(n_1281),
.B(n_1313),
.C(n_1332),
.Y(n_1448)
);

AO32x2_ASAP7_75t_L g1449 ( 
.A1(n_1398),
.A2(n_1346),
.A3(n_1283),
.B1(n_1332),
.B2(n_1348),
.Y(n_1449)
);

OA21x2_ASAP7_75t_L g1450 ( 
.A1(n_1385),
.A2(n_1281),
.B(n_1293),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1386),
.B(n_1293),
.Y(n_1451)
);

BUFx8_ASAP7_75t_SL g1452 ( 
.A(n_1396),
.Y(n_1452)
);

AND2x4_ASAP7_75t_L g1453 ( 
.A(n_1361),
.B(n_1352),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1386),
.B(n_1369),
.Y(n_1454)
);

HB1xp67_ASAP7_75t_L g1455 ( 
.A(n_1362),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1382),
.Y(n_1456)
);

OAI21xp5_ASAP7_75t_L g1457 ( 
.A1(n_1424),
.A2(n_1311),
.B(n_1275),
.Y(n_1457)
);

OAI21xp5_ASAP7_75t_L g1458 ( 
.A1(n_1425),
.A2(n_1311),
.B(n_1282),
.Y(n_1458)
);

OR2x6_ASAP7_75t_L g1459 ( 
.A(n_1415),
.B(n_1428),
.Y(n_1459)
);

AO21x2_ASAP7_75t_L g1460 ( 
.A1(n_1366),
.A2(n_1412),
.B(n_1378),
.Y(n_1460)
);

AND2x4_ASAP7_75t_L g1461 ( 
.A(n_1361),
.B(n_1372),
.Y(n_1461)
);

OA21x2_ASAP7_75t_L g1462 ( 
.A1(n_1366),
.A2(n_1406),
.B(n_1422),
.Y(n_1462)
);

NOR2x1_ASAP7_75t_SL g1463 ( 
.A(n_1412),
.B(n_1418),
.Y(n_1463)
);

NOR2xp33_ASAP7_75t_L g1464 ( 
.A(n_1412),
.B(n_1425),
.Y(n_1464)
);

CKINVDCx5p33_ASAP7_75t_R g1465 ( 
.A(n_1396),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1387),
.B(n_1429),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1387),
.B(n_1429),
.Y(n_1467)
);

CKINVDCx20_ASAP7_75t_R g1468 ( 
.A(n_1396),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1383),
.Y(n_1469)
);

NOR2x1_ASAP7_75t_SL g1470 ( 
.A(n_1372),
.B(n_1384),
.Y(n_1470)
);

A2O1A1Ixp33_ASAP7_75t_L g1471 ( 
.A1(n_1405),
.A2(n_1395),
.B(n_1410),
.C(n_1381),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1381),
.B(n_1413),
.Y(n_1472)
);

A2O1A1Ixp33_ASAP7_75t_L g1473 ( 
.A1(n_1405),
.A2(n_1395),
.B(n_1410),
.C(n_1416),
.Y(n_1473)
);

CKINVDCx20_ASAP7_75t_R g1474 ( 
.A(n_1421),
.Y(n_1474)
);

O2A1O1Ixp33_ASAP7_75t_L g1475 ( 
.A1(n_1416),
.A2(n_1397),
.B(n_1406),
.C(n_1360),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1370),
.B(n_1379),
.Y(n_1476)
);

OAI22xp5_ASAP7_75t_L g1477 ( 
.A1(n_1411),
.A2(n_1415),
.B1(n_1374),
.B2(n_1428),
.Y(n_1477)
);

OAI21xp5_ASAP7_75t_L g1478 ( 
.A1(n_1428),
.A2(n_1402),
.B(n_1401),
.Y(n_1478)
);

AO21x2_ASAP7_75t_L g1479 ( 
.A1(n_1427),
.A2(n_1392),
.B(n_1394),
.Y(n_1479)
);

OR2x6_ASAP7_75t_L g1480 ( 
.A(n_1372),
.B(n_1388),
.Y(n_1480)
);

AOI21xp5_ASAP7_75t_L g1481 ( 
.A1(n_1404),
.A2(n_1401),
.B(n_1402),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1407),
.B(n_1408),
.Y(n_1482)
);

A2O1A1Ixp33_ASAP7_75t_L g1483 ( 
.A1(n_1414),
.A2(n_1417),
.B(n_1388),
.C(n_1400),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1445),
.B(n_1364),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1440),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1440),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1456),
.Y(n_1487)
);

HB1xp67_ASAP7_75t_L g1488 ( 
.A(n_1455),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1445),
.B(n_1364),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1445),
.B(n_1364),
.Y(n_1490)
);

INVx5_ASAP7_75t_L g1491 ( 
.A(n_1459),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1464),
.B(n_1404),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1469),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1464),
.B(n_1420),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1445),
.B(n_1364),
.Y(n_1495)
);

OAI22xp5_ASAP7_75t_L g1496 ( 
.A1(n_1434),
.A2(n_1414),
.B1(n_1417),
.B2(n_1400),
.Y(n_1496)
);

INVx1_ASAP7_75t_SL g1497 ( 
.A(n_1466),
.Y(n_1497)
);

AOI22xp33_ASAP7_75t_L g1498 ( 
.A1(n_1436),
.A2(n_1421),
.B1(n_1420),
.B2(n_1422),
.Y(n_1498)
);

INVxp67_ASAP7_75t_SL g1499 ( 
.A(n_1462),
.Y(n_1499)
);

OR2x6_ASAP7_75t_L g1500 ( 
.A(n_1459),
.B(n_1372),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1479),
.Y(n_1501)
);

INVx1_ASAP7_75t_SL g1502 ( 
.A(n_1467),
.Y(n_1502)
);

CKINVDCx20_ASAP7_75t_R g1503 ( 
.A(n_1452),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1482),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1479),
.Y(n_1505)
);

NOR2xp33_ASAP7_75t_L g1506 ( 
.A(n_1475),
.B(n_1430),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1461),
.B(n_1376),
.Y(n_1507)
);

INVxp67_ASAP7_75t_L g1508 ( 
.A(n_1463),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1462),
.Y(n_1509)
);

HB1xp67_ASAP7_75t_L g1510 ( 
.A(n_1476),
.Y(n_1510)
);

AND2x4_ASAP7_75t_L g1511 ( 
.A(n_1470),
.B(n_1377),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1481),
.B(n_1403),
.Y(n_1512)
);

INVxp67_ASAP7_75t_SL g1513 ( 
.A(n_1450),
.Y(n_1513)
);

BUFx2_ASAP7_75t_L g1514 ( 
.A(n_1511),
.Y(n_1514)
);

OAI21xp33_ASAP7_75t_L g1515 ( 
.A1(n_1506),
.A2(n_1471),
.B(n_1473),
.Y(n_1515)
);

NOR2x1_ASAP7_75t_SL g1516 ( 
.A(n_1500),
.B(n_1459),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1509),
.Y(n_1517)
);

OR2x2_ASAP7_75t_L g1518 ( 
.A(n_1490),
.B(n_1460),
.Y(n_1518)
);

AND2x4_ASAP7_75t_SL g1519 ( 
.A(n_1500),
.B(n_1432),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1509),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1490),
.B(n_1480),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1492),
.B(n_1403),
.Y(n_1522)
);

NOR2xp33_ASAP7_75t_L g1523 ( 
.A(n_1506),
.B(n_1496),
.Y(n_1523)
);

BUFx2_ASAP7_75t_L g1524 ( 
.A(n_1511),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1495),
.B(n_1449),
.Y(n_1525)
);

AND2x4_ASAP7_75t_L g1526 ( 
.A(n_1511),
.B(n_1443),
.Y(n_1526)
);

BUFx2_ASAP7_75t_L g1527 ( 
.A(n_1511),
.Y(n_1527)
);

OR2x2_ASAP7_75t_L g1528 ( 
.A(n_1495),
.B(n_1460),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1495),
.B(n_1449),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1488),
.Y(n_1530)
);

AOI22xp33_ASAP7_75t_L g1531 ( 
.A1(n_1498),
.A2(n_1435),
.B1(n_1438),
.B2(n_1437),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1484),
.B(n_1449),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1484),
.B(n_1437),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1486),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1486),
.Y(n_1535)
);

AO31x2_ASAP7_75t_L g1536 ( 
.A1(n_1505),
.A2(n_1501),
.A3(n_1493),
.B(n_1485),
.Y(n_1536)
);

OAI221xp5_ASAP7_75t_L g1537 ( 
.A1(n_1498),
.A2(n_1471),
.B1(n_1473),
.B2(n_1439),
.C(n_1483),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1486),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1492),
.B(n_1365),
.Y(n_1539)
);

NOR2xp33_ASAP7_75t_L g1540 ( 
.A(n_1496),
.B(n_1444),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1487),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1489),
.B(n_1478),
.Y(n_1542)
);

NAND2x1p5_ASAP7_75t_L g1543 ( 
.A(n_1514),
.B(n_1491),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1534),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1522),
.B(n_1494),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1522),
.B(n_1494),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1539),
.B(n_1504),
.Y(n_1547)
);

NOR4xp25_ASAP7_75t_SL g1548 ( 
.A(n_1515),
.B(n_1465),
.C(n_1513),
.D(n_1442),
.Y(n_1548)
);

OR2x2_ASAP7_75t_L g1549 ( 
.A(n_1518),
.B(n_1489),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1525),
.B(n_1489),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1534),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1539),
.B(n_1504),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1535),
.Y(n_1553)
);

NAND2x1_ASAP7_75t_L g1554 ( 
.A(n_1514),
.B(n_1500),
.Y(n_1554)
);

INVx3_ASAP7_75t_L g1555 ( 
.A(n_1536),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1523),
.B(n_1504),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1525),
.B(n_1507),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1523),
.B(n_1512),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1535),
.Y(n_1559)
);

NOR2x1p5_ASAP7_75t_L g1560 ( 
.A(n_1526),
.B(n_1421),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1517),
.Y(n_1561)
);

OAI222xp33_ASAP7_75t_L g1562 ( 
.A1(n_1537),
.A2(n_1477),
.B1(n_1497),
.B2(n_1502),
.C1(n_1512),
.C2(n_1433),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1517),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1517),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1517),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1525),
.B(n_1507),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1530),
.B(n_1510),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1529),
.B(n_1507),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1529),
.B(n_1507),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1538),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1538),
.Y(n_1571)
);

OR2x2_ASAP7_75t_L g1572 ( 
.A(n_1518),
.B(n_1499),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1520),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1541),
.Y(n_1574)
);

BUFx6f_ASAP7_75t_L g1575 ( 
.A(n_1520),
.Y(n_1575)
);

AND2x4_ASAP7_75t_L g1576 ( 
.A(n_1560),
.B(n_1516),
.Y(n_1576)
);

AOI211xp5_ASAP7_75t_L g1577 ( 
.A1(n_1562),
.A2(n_1515),
.B(n_1537),
.C(n_1540),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1544),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1560),
.B(n_1514),
.Y(n_1579)
);

OAI211xp5_ASAP7_75t_SL g1580 ( 
.A1(n_1558),
.A2(n_1531),
.B(n_1441),
.C(n_1540),
.Y(n_1580)
);

AOI32xp33_ASAP7_75t_L g1581 ( 
.A1(n_1558),
.A2(n_1542),
.A3(n_1531),
.B1(n_1532),
.B2(n_1533),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1556),
.B(n_1542),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1544),
.Y(n_1583)
);

AND2x4_ASAP7_75t_L g1584 ( 
.A(n_1557),
.B(n_1516),
.Y(n_1584)
);

OAI22xp5_ASAP7_75t_L g1585 ( 
.A1(n_1548),
.A2(n_1483),
.B1(n_1556),
.B2(n_1439),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1575),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1575),
.Y(n_1587)
);

OR2x6_ASAP7_75t_L g1588 ( 
.A(n_1554),
.B(n_1431),
.Y(n_1588)
);

INVxp67_ASAP7_75t_SL g1589 ( 
.A(n_1543),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1551),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1575),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1551),
.Y(n_1592)
);

INVx2_ASAP7_75t_SL g1593 ( 
.A(n_1554),
.Y(n_1593)
);

NAND2x1_ASAP7_75t_L g1594 ( 
.A(n_1555),
.B(n_1524),
.Y(n_1594)
);

NOR2xp33_ASAP7_75t_SL g1595 ( 
.A(n_1562),
.B(n_1503),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1553),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1553),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1575),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1559),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1559),
.Y(n_1600)
);

NAND2x1p5_ASAP7_75t_L g1601 ( 
.A(n_1575),
.B(n_1491),
.Y(n_1601)
);

OR2x2_ASAP7_75t_L g1602 ( 
.A(n_1567),
.B(n_1545),
.Y(n_1602)
);

AND2x4_ASAP7_75t_L g1603 ( 
.A(n_1557),
.B(n_1524),
.Y(n_1603)
);

NOR2xp33_ASAP7_75t_L g1604 ( 
.A(n_1545),
.B(n_1368),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1543),
.B(n_1524),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1543),
.B(n_1527),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1570),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1575),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1575),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1543),
.B(n_1527),
.Y(n_1610)
);

INVxp67_ASAP7_75t_L g1611 ( 
.A(n_1567),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1557),
.B(n_1527),
.Y(n_1612)
);

OAI21xp5_ASAP7_75t_L g1613 ( 
.A1(n_1546),
.A2(n_1508),
.B(n_1542),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1574),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1546),
.B(n_1497),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1570),
.Y(n_1616)
);

INVx2_ASAP7_75t_SL g1617 ( 
.A(n_1571),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1577),
.B(n_1547),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1583),
.Y(n_1619)
);

OR2x2_ASAP7_75t_L g1620 ( 
.A(n_1602),
.B(n_1547),
.Y(n_1620)
);

INVx4_ASAP7_75t_L g1621 ( 
.A(n_1576),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1611),
.B(n_1552),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1576),
.B(n_1566),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1576),
.B(n_1566),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1579),
.B(n_1584),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1579),
.B(n_1566),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1604),
.B(n_1552),
.Y(n_1627)
);

AOI211xp5_ASAP7_75t_L g1628 ( 
.A1(n_1580),
.A2(n_1447),
.B(n_1457),
.C(n_1458),
.Y(n_1628)
);

NOR2xp67_ASAP7_75t_SL g1629 ( 
.A(n_1595),
.B(n_1368),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1603),
.Y(n_1630)
);

OR2x2_ASAP7_75t_L g1631 ( 
.A(n_1602),
.B(n_1572),
.Y(n_1631)
);

OR2x2_ASAP7_75t_L g1632 ( 
.A(n_1582),
.B(n_1572),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1583),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1590),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1584),
.B(n_1568),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1581),
.B(n_1472),
.Y(n_1636)
);

INVxp67_ASAP7_75t_L g1637 ( 
.A(n_1585),
.Y(n_1637)
);

INVx1_ASAP7_75t_SL g1638 ( 
.A(n_1605),
.Y(n_1638)
);

OR2x2_ASAP7_75t_L g1639 ( 
.A(n_1615),
.B(n_1572),
.Y(n_1639)
);

NAND2x1_ASAP7_75t_L g1640 ( 
.A(n_1584),
.B(n_1532),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1603),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1588),
.B(n_1568),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1590),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1613),
.B(n_1502),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1588),
.B(n_1568),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1603),
.Y(n_1646)
);

OR2x6_ASAP7_75t_L g1647 ( 
.A(n_1588),
.B(n_1432),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1592),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1588),
.B(n_1569),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1578),
.B(n_1532),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1599),
.B(n_1521),
.Y(n_1651)
);

OR2x2_ASAP7_75t_L g1652 ( 
.A(n_1600),
.B(n_1518),
.Y(n_1652)
);

OR2x2_ASAP7_75t_L g1653 ( 
.A(n_1618),
.B(n_1612),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1619),
.Y(n_1654)
);

OAI21xp33_ASAP7_75t_L g1655 ( 
.A1(n_1637),
.A2(n_1589),
.B(n_1605),
.Y(n_1655)
);

NOR2xp67_ASAP7_75t_L g1656 ( 
.A(n_1621),
.B(n_1593),
.Y(n_1656)
);

AND2x4_ASAP7_75t_L g1657 ( 
.A(n_1625),
.B(n_1593),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1619),
.Y(n_1658)
);

OAI333xp33_ASAP7_75t_L g1659 ( 
.A1(n_1636),
.A2(n_1548),
.A3(n_1508),
.B1(n_1614),
.B2(n_1592),
.B3(n_1596),
.C1(n_1616),
.C2(n_1607),
.C3(n_1597),
.Y(n_1659)
);

OAI22xp33_ASAP7_75t_SL g1660 ( 
.A1(n_1640),
.A2(n_1601),
.B1(n_1594),
.B2(n_1617),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1633),
.Y(n_1661)
);

OAI32xp33_ASAP7_75t_L g1662 ( 
.A1(n_1638),
.A2(n_1601),
.A3(n_1549),
.B1(n_1528),
.B2(n_1610),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1633),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1634),
.Y(n_1664)
);

AOI211xp5_ASAP7_75t_L g1665 ( 
.A1(n_1629),
.A2(n_1610),
.B(n_1606),
.C(n_1446),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1635),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1634),
.Y(n_1667)
);

AOI22xp5_ASAP7_75t_L g1668 ( 
.A1(n_1629),
.A2(n_1606),
.B1(n_1519),
.B2(n_1500),
.Y(n_1668)
);

AOI21xp33_ASAP7_75t_L g1669 ( 
.A1(n_1647),
.A2(n_1617),
.B(n_1601),
.Y(n_1669)
);

OAI22xp33_ASAP7_75t_SL g1670 ( 
.A1(n_1640),
.A2(n_1594),
.B1(n_1528),
.B2(n_1549),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1643),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1643),
.Y(n_1672)
);

NAND2xp33_ASAP7_75t_SL g1673 ( 
.A(n_1621),
.B(n_1503),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1648),
.Y(n_1674)
);

NOR2x1_ASAP7_75t_L g1675 ( 
.A(n_1621),
.B(n_1468),
.Y(n_1675)
);

AOI22xp5_ASAP7_75t_L g1676 ( 
.A1(n_1625),
.A2(n_1519),
.B1(n_1500),
.B2(n_1491),
.Y(n_1676)
);

AOI22xp5_ASAP7_75t_L g1677 ( 
.A1(n_1627),
.A2(n_1519),
.B1(n_1500),
.B2(n_1491),
.Y(n_1677)
);

AOI22xp33_ASAP7_75t_SL g1678 ( 
.A1(n_1659),
.A2(n_1642),
.B1(n_1649),
.B2(n_1645),
.Y(n_1678)
);

OAI22xp33_ASAP7_75t_L g1679 ( 
.A1(n_1668),
.A2(n_1644),
.B1(n_1647),
.B2(n_1641),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1655),
.B(n_1653),
.Y(n_1680)
);

AOI22xp5_ASAP7_75t_L g1681 ( 
.A1(n_1673),
.A2(n_1642),
.B1(n_1645),
.B2(n_1649),
.Y(n_1681)
);

AND2x4_ASAP7_75t_L g1682 ( 
.A(n_1656),
.B(n_1630),
.Y(n_1682)
);

NOR2xp33_ASAP7_75t_L g1683 ( 
.A(n_1675),
.B(n_1452),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1666),
.B(n_1626),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1657),
.Y(n_1685)
);

OAI22xp33_ASAP7_75t_L g1686 ( 
.A1(n_1676),
.A2(n_1647),
.B1(n_1630),
.B2(n_1646),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1654),
.B(n_1648),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1658),
.Y(n_1688)
);

AOI22xp33_ASAP7_75t_L g1689 ( 
.A1(n_1657),
.A2(n_1647),
.B1(n_1646),
.B2(n_1641),
.Y(n_1689)
);

OR2x2_ASAP7_75t_L g1690 ( 
.A(n_1661),
.B(n_1639),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1665),
.B(n_1626),
.Y(n_1691)
);

AOI33xp33_ASAP7_75t_L g1692 ( 
.A1(n_1663),
.A2(n_1628),
.A3(n_1623),
.B1(n_1624),
.B2(n_1635),
.B3(n_1612),
.Y(n_1692)
);

INVx2_ASAP7_75t_L g1693 ( 
.A(n_1664),
.Y(n_1693)
);

NOR2xp33_ASAP7_75t_L g1694 ( 
.A(n_1669),
.B(n_1468),
.Y(n_1694)
);

AOI322xp5_ASAP7_75t_L g1695 ( 
.A1(n_1667),
.A2(n_1550),
.A3(n_1623),
.B1(n_1624),
.B2(n_1622),
.C1(n_1650),
.C2(n_1533),
.Y(n_1695)
);

INVxp67_ASAP7_75t_L g1696 ( 
.A(n_1656),
.Y(n_1696)
);

OAI22xp5_ASAP7_75t_L g1697 ( 
.A1(n_1678),
.A2(n_1677),
.B1(n_1647),
.B2(n_1651),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1687),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1687),
.Y(n_1699)
);

AOI22xp33_ASAP7_75t_SL g1700 ( 
.A1(n_1691),
.A2(n_1660),
.B1(n_1670),
.B2(n_1662),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1685),
.B(n_1671),
.Y(n_1701)
);

AOI221xp5_ASAP7_75t_L g1702 ( 
.A1(n_1680),
.A2(n_1674),
.B1(n_1672),
.B2(n_1631),
.C(n_1632),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1692),
.B(n_1620),
.Y(n_1703)
);

CKINVDCx5p33_ASAP7_75t_R g1704 ( 
.A(n_1683),
.Y(n_1704)
);

INVxp67_ASAP7_75t_L g1705 ( 
.A(n_1694),
.Y(n_1705)
);

AOI221xp5_ASAP7_75t_L g1706 ( 
.A1(n_1679),
.A2(n_1631),
.B1(n_1632),
.B2(n_1620),
.C(n_1639),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1696),
.B(n_1596),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1697),
.B(n_1682),
.Y(n_1708)
);

OR2x2_ASAP7_75t_L g1709 ( 
.A(n_1701),
.B(n_1684),
.Y(n_1709)
);

NAND4xp25_ASAP7_75t_L g1710 ( 
.A(n_1703),
.B(n_1689),
.C(n_1681),
.D(n_1688),
.Y(n_1710)
);

NOR2xp33_ASAP7_75t_L g1711 ( 
.A(n_1704),
.B(n_1686),
.Y(n_1711)
);

AOI221xp5_ASAP7_75t_L g1712 ( 
.A1(n_1700),
.A2(n_1693),
.B1(n_1682),
.B2(n_1690),
.C(n_1695),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1702),
.B(n_1597),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1707),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1698),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1705),
.B(n_1607),
.Y(n_1716)
);

O2A1O1Ixp33_ASAP7_75t_L g1717 ( 
.A1(n_1708),
.A2(n_1699),
.B(n_1706),
.C(n_1652),
.Y(n_1717)
);

NOR2xp67_ASAP7_75t_L g1718 ( 
.A(n_1711),
.B(n_1442),
.Y(n_1718)
);

AOI211xp5_ASAP7_75t_SL g1719 ( 
.A1(n_1712),
.A2(n_1380),
.B(n_1652),
.C(n_1474),
.Y(n_1719)
);

AOI221xp5_ASAP7_75t_L g1720 ( 
.A1(n_1710),
.A2(n_1598),
.B1(n_1586),
.B2(n_1609),
.C(n_1608),
.Y(n_1720)
);

NAND3xp33_ASAP7_75t_SL g1721 ( 
.A(n_1709),
.B(n_1474),
.C(n_1465),
.Y(n_1721)
);

OAI221xp5_ASAP7_75t_SL g1722 ( 
.A1(n_1717),
.A2(n_1713),
.B1(n_1716),
.B2(n_1714),
.C(n_1715),
.Y(n_1722)
);

AOI22xp33_ASAP7_75t_L g1723 ( 
.A1(n_1721),
.A2(n_1587),
.B1(n_1609),
.B2(n_1608),
.Y(n_1723)
);

AOI22xp5_ASAP7_75t_L g1724 ( 
.A1(n_1718),
.A2(n_1586),
.B1(n_1587),
.B2(n_1598),
.Y(n_1724)
);

OAI221xp5_ASAP7_75t_L g1725 ( 
.A1(n_1719),
.A2(n_1591),
.B1(n_1446),
.B2(n_1616),
.C(n_1614),
.Y(n_1725)
);

NOR3xp33_ASAP7_75t_L g1726 ( 
.A(n_1720),
.B(n_1380),
.C(n_1591),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_SL g1727 ( 
.A(n_1718),
.B(n_1453),
.Y(n_1727)
);

HB1xp67_ASAP7_75t_L g1728 ( 
.A(n_1727),
.Y(n_1728)
);

AND2x4_ASAP7_75t_L g1729 ( 
.A(n_1726),
.B(n_1453),
.Y(n_1729)
);

INVx2_ASAP7_75t_SL g1730 ( 
.A(n_1724),
.Y(n_1730)
);

AOI22xp5_ASAP7_75t_L g1731 ( 
.A1(n_1725),
.A2(n_1453),
.B1(n_1454),
.B2(n_1451),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1722),
.Y(n_1732)
);

AOI221xp5_ASAP7_75t_L g1733 ( 
.A1(n_1732),
.A2(n_1730),
.B1(n_1728),
.B2(n_1729),
.C(n_1723),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1729),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1731),
.B(n_1571),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1733),
.B(n_1561),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1736),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1737),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1737),
.Y(n_1739)
);

AOI22x1_ASAP7_75t_L g1740 ( 
.A1(n_1739),
.A2(n_1734),
.B1(n_1735),
.B2(n_1561),
.Y(n_1740)
);

INVxp67_ASAP7_75t_L g1741 ( 
.A(n_1738),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1740),
.Y(n_1742)
);

AO21x2_ASAP7_75t_L g1743 ( 
.A1(n_1741),
.A2(n_1563),
.B(n_1561),
.Y(n_1743)
);

OA21x2_ASAP7_75t_L g1744 ( 
.A1(n_1742),
.A2(n_1743),
.B(n_1564),
.Y(n_1744)
);

NOR2xp67_ASAP7_75t_L g1745 ( 
.A(n_1744),
.B(n_1743),
.Y(n_1745)
);

O2A1O1Ixp33_ASAP7_75t_SL g1746 ( 
.A1(n_1745),
.A2(n_1448),
.B(n_1573),
.C(n_1565),
.Y(n_1746)
);

OAI221xp5_ASAP7_75t_R g1747 ( 
.A1(n_1746),
.A2(n_1555),
.B1(n_1549),
.B2(n_1573),
.C(n_1565),
.Y(n_1747)
);

AOI22xp5_ASAP7_75t_L g1748 ( 
.A1(n_1747),
.A2(n_1565),
.B1(n_1573),
.B2(n_1564),
.Y(n_1748)
);


endmodule