module fake_jpeg_9638_n_329 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_329);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_329;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_10),
.B(n_14),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx24_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

OR2x2_ASAP7_75t_L g29 ( 
.A(n_6),
.B(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_40),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_1),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_34),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_41),
.B(n_42),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g42 ( 
.A(n_22),
.B(n_1),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_43),
.B(n_29),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_38),
.A2(n_32),
.B1(n_19),
.B2(n_17),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_48),
.A2(n_54),
.B1(n_56),
.B2(n_58),
.Y(n_104)
);

CKINVDCx6p67_ASAP7_75t_R g52 ( 
.A(n_35),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_52),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_53),
.B(n_60),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_38),
.A2(n_32),
.B1(n_39),
.B2(n_46),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_43),
.A2(n_32),
.B1(n_33),
.B2(n_21),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_35),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_57),
.B(n_44),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_41),
.A2(n_33),
.B1(n_21),
.B2(n_30),
.Y(n_58)
);

CKINVDCx6p67_ASAP7_75t_R g59 ( 
.A(n_35),
.Y(n_59)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_40),
.A2(n_16),
.B1(n_31),
.B2(n_18),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_62),
.A2(n_65),
.B1(n_72),
.B2(n_24),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_42),
.A2(n_30),
.B1(n_31),
.B2(n_16),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_63),
.A2(n_70),
.B1(n_24),
.B2(n_44),
.Y(n_85)
);

AND2x2_ASAP7_75t_SL g64 ( 
.A(n_44),
.B(n_16),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_64),
.B(n_73),
.C(n_57),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_42),
.A2(n_17),
.B1(n_31),
.B2(n_19),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_36),
.A2(n_17),
.B1(n_18),
.B2(n_28),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_69),
.B(n_27),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_36),
.A2(n_19),
.B1(n_28),
.B2(n_18),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_74),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_37),
.A2(n_28),
.B1(n_26),
.B2(n_25),
.Y(n_72)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_L g75 ( 
.A1(n_45),
.A2(n_27),
.B1(n_23),
.B2(n_20),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_75),
.A2(n_25),
.B1(n_27),
.B2(n_23),
.Y(n_79)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_76),
.B(n_78),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_47),
.B(n_29),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_77),
.B(n_80),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_68),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_79),
.A2(n_85),
.B1(n_93),
.B2(n_96),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_47),
.B(n_29),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

INVx13_ASAP7_75t_L g127 ( 
.A(n_83),
.Y(n_127)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_86),
.Y(n_117)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_87),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_68),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_89),
.B(n_90),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_12),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_64),
.B(n_45),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_91),
.B(n_94),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_102),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_66),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_68),
.Y(n_94)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_95),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_66),
.A2(n_15),
.B1(n_13),
.B2(n_12),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_53),
.B(n_24),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_97),
.B(n_101),
.Y(n_136)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_66),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_64),
.B(n_13),
.Y(n_99)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_99),
.Y(n_133)
);

AO22x1_ASAP7_75t_L g123 ( 
.A1(n_100),
.A2(n_102),
.B1(n_104),
.B2(n_112),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_65),
.B(n_34),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_61),
.A2(n_20),
.B1(n_27),
.B2(n_23),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_103),
.A2(n_108),
.B1(n_112),
.B2(n_59),
.Y(n_124)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_105),
.Y(n_122)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_61),
.Y(n_106)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_106),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_69),
.B(n_1),
.Y(n_107)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_107),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_52),
.A2(n_20),
.B1(n_23),
.B2(n_4),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_72),
.Y(n_109)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_109),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_49),
.B(n_2),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_110),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_48),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_92),
.B(n_59),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_114),
.B(n_119),
.C(n_137),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_91),
.B(n_59),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_123),
.A2(n_104),
.B1(n_76),
.B2(n_109),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_124),
.A2(n_125),
.B1(n_131),
.B2(n_126),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_88),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_125),
.B(n_131),
.Y(n_149)
);

AND2x6_ASAP7_75t_L g129 ( 
.A(n_86),
.B(n_52),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_129),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_88),
.Y(n_131)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_106),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_132),
.B(n_134),
.Y(n_165)
);

INVx13_ASAP7_75t_L g134 ( 
.A(n_111),
.Y(n_134)
);

INVx13_ASAP7_75t_L g135 ( 
.A(n_111),
.Y(n_135)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_135),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_77),
.B(n_59),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_115),
.B(n_80),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_144),
.B(n_151),
.Y(n_190)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_130),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_145),
.B(n_148),
.Y(n_189)
);

MAJx2_ASAP7_75t_L g146 ( 
.A(n_115),
.B(n_101),
.C(n_99),
.Y(n_146)
);

XNOR2x1_ASAP7_75t_L g196 ( 
.A(n_146),
.B(n_34),
.Y(n_196)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_138),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_147),
.B(n_161),
.Y(n_177)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_130),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_136),
.A2(n_107),
.B(n_97),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_150),
.A2(n_154),
.B(n_159),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_115),
.B(n_100),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_113),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_152),
.B(n_155),
.Y(n_201)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_139),
.Y(n_155)
);

OAI21xp33_ASAP7_75t_L g156 ( 
.A1(n_140),
.A2(n_90),
.B(n_84),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_156),
.A2(n_169),
.B(n_67),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_123),
.A2(n_79),
.B1(n_84),
.B2(n_94),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_157),
.A2(n_117),
.B1(n_141),
.B2(n_133),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_128),
.B(n_110),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_158),
.B(n_162),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_138),
.A2(n_82),
.B1(n_98),
.B2(n_106),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_160),
.A2(n_133),
.B1(n_127),
.B2(n_134),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_120),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_139),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_121),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_163),
.B(n_164),
.Y(n_179)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_121),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_124),
.A2(n_78),
.B1(n_89),
.B2(n_87),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_166),
.A2(n_168),
.B1(n_127),
.B2(n_135),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_136),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_167),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_123),
.A2(n_87),
.B1(n_60),
.B2(n_71),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_140),
.A2(n_95),
.B(n_34),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_120),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_170),
.B(n_132),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_128),
.B(n_82),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_171),
.B(n_172),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_116),
.B(n_82),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_114),
.B(n_44),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_173),
.B(n_175),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_119),
.B(n_74),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_174),
.B(n_118),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_137),
.B(n_111),
.C(n_51),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_149),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_176),
.B(n_182),
.Y(n_227)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_180),
.Y(n_210)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_149),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_143),
.B(n_129),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_183),
.B(n_208),
.C(n_175),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_165),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_184),
.B(n_186),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_185),
.A2(n_191),
.B1(n_154),
.B2(n_152),
.Y(n_209)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_172),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_171),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_187),
.B(n_194),
.Y(n_234)
);

AO22x1_ASAP7_75t_SL g188 ( 
.A1(n_157),
.A2(n_141),
.B1(n_117),
.B2(n_116),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_188),
.A2(n_192),
.B1(n_164),
.B2(n_163),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_147),
.B(n_118),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_193),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_158),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_153),
.A2(n_122),
.B1(n_50),
.B2(n_105),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_195),
.A2(n_205),
.B1(n_50),
.B2(n_49),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_196),
.B(n_173),
.Y(n_225)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_168),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_197),
.A2(n_204),
.B1(n_207),
.B2(n_142),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_161),
.B(n_170),
.Y(n_198)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_198),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_166),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_199),
.A2(n_200),
.B(n_174),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_160),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_153),
.A2(n_122),
.B1(n_50),
.B2(n_49),
.Y(n_205)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_145),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_209),
.A2(n_218),
.B1(n_229),
.B2(n_230),
.Y(n_236)
);

INVx13_ASAP7_75t_L g211 ( 
.A(n_177),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_211),
.B(n_222),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_202),
.B(n_143),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_212),
.B(n_217),
.C(n_231),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_178),
.A2(n_151),
.B(n_169),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_214),
.A2(n_219),
.B(n_223),
.Y(n_238)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_189),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_215),
.B(n_216),
.Y(n_258)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_189),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_199),
.A2(n_162),
.B1(n_155),
.B2(n_148),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_178),
.A2(n_144),
.B(n_146),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_221),
.A2(n_191),
.B1(n_188),
.B2(n_185),
.Y(n_252)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_206),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_206),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_225),
.B(n_196),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_226),
.B(n_188),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_194),
.B(n_150),
.Y(n_228)
);

CKINVDCx14_ASAP7_75t_R g247 ( 
.A(n_228),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_204),
.A2(n_142),
.B1(n_67),
.B2(n_51),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_202),
.B(n_146),
.C(n_51),
.Y(n_231)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_232),
.Y(n_248)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_179),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_233),
.B(n_182),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_197),
.A2(n_81),
.B1(n_67),
.B2(n_120),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_235),
.A2(n_186),
.B1(n_187),
.B2(n_176),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_237),
.B(n_240),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_212),
.B(n_183),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_239),
.B(n_243),
.C(n_245),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_219),
.B(n_190),
.Y(n_240)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_242),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_231),
.B(n_190),
.Y(n_243)
);

NOR3xp33_ASAP7_75t_SL g244 ( 
.A(n_218),
.B(n_203),
.C(n_201),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_244),
.B(n_249),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_225),
.B(n_200),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_217),
.B(n_208),
.C(n_181),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_246),
.B(n_250),
.C(n_222),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_211),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_226),
.B(n_181),
.C(n_207),
.Y(n_250)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_251),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_252),
.B(n_256),
.Y(n_272)
);

FAx1_ASAP7_75t_SL g270 ( 
.A(n_253),
.B(n_235),
.CI(n_223),
.CON(n_270),
.SN(n_270)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_215),
.A2(n_188),
.B1(n_192),
.B2(n_205),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_254),
.A2(n_257),
.B1(n_216),
.B2(n_227),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_211),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_209),
.A2(n_203),
.B1(n_201),
.B2(n_195),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_243),
.B(n_214),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_260),
.B(n_262),
.Y(n_282)
);

OR2x2_ASAP7_75t_L g261 ( 
.A(n_255),
.B(n_234),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_261),
.B(n_269),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_241),
.B(n_221),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_241),
.B(n_228),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_263),
.B(n_267),
.C(n_273),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_247),
.B(n_227),
.Y(n_264)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_264),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_266),
.A2(n_274),
.B1(n_250),
.B2(n_258),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_251),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_270),
.A2(n_245),
.B1(n_238),
.B2(n_237),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_239),
.B(n_213),
.C(n_210),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_236),
.A2(n_213),
.B1(n_210),
.B2(n_224),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_246),
.B(n_233),
.Y(n_275)
);

BUFx24_ASAP7_75t_SL g278 ( 
.A(n_275),
.Y(n_278)
);

AOI31xp67_ASAP7_75t_L g277 ( 
.A1(n_261),
.A2(n_244),
.A3(n_254),
.B(n_253),
.Y(n_277)
);

OR2x2_ASAP7_75t_L g294 ( 
.A(n_277),
.B(n_268),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_279),
.B(n_262),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_272),
.A2(n_248),
.B1(n_224),
.B2(n_220),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_280),
.A2(n_287),
.B1(n_264),
.B2(n_271),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_281),
.B(n_285),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_270),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_283),
.B(n_288),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_263),
.B(n_240),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_276),
.A2(n_232),
.B1(n_184),
.B2(n_81),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_267),
.B(n_81),
.C(n_55),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_273),
.B(n_55),
.C(n_3),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_290),
.B(n_291),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_265),
.B(n_2),
.C(n_3),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_292),
.B(n_295),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_294),
.B(n_302),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_289),
.A2(n_274),
.B(n_270),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_296),
.A2(n_304),
.B1(n_3),
.B2(n_5),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_286),
.A2(n_265),
.B1(n_260),
.B2(n_259),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_298),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_278),
.B(n_259),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_299),
.B(n_300),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_288),
.B(n_290),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_291),
.B(n_2),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_284),
.B(n_2),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_303),
.B(n_5),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_284),
.A2(n_3),
.B(n_4),
.Y(n_304)
);

OAI21x1_ASAP7_75t_L g306 ( 
.A1(n_303),
.A2(n_282),
.B(n_4),
.Y(n_306)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_306),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_L g307 ( 
.A1(n_295),
.A2(n_282),
.B1(n_5),
.B2(n_6),
.Y(n_307)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_307),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_308),
.B(n_309),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_294),
.B(n_5),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_310),
.B(n_312),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_305),
.B(n_293),
.C(n_298),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_317),
.B(n_320),
.C(n_11),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_313),
.B(n_301),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_318),
.B(n_10),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_305),
.A2(n_297),
.B1(n_304),
.B2(n_9),
.Y(n_320)
);

NAND3xp33_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_312),
.C(n_313),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_321),
.A2(n_322),
.B1(n_323),
.B2(n_315),
.Y(n_325)
);

AOI322xp5_ASAP7_75t_L g322 ( 
.A1(n_319),
.A2(n_311),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.C1(n_11),
.C2(n_6),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_324),
.B(n_317),
.C(n_314),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_325),
.B(n_326),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_316),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_328),
.B(n_11),
.Y(n_329)
);


endmodule