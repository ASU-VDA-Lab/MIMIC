module fake_jpeg_1917_n_170 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_170);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_170;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

AND2x2_ASAP7_75t_L g12 ( 
.A(n_3),
.B(n_5),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_10),
.B(n_7),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_10),
.B(n_9),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_34),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_35),
.B(n_38),
.Y(n_69)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_36),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_22),
.B(n_8),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_47),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_18),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_40),
.Y(n_83)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_21),
.Y(n_45)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_26),
.B(n_8),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_50),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_12),
.B(n_0),
.C(n_1),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_49),
.B(n_56),
.Y(n_71)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_30),
.B(n_11),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_52),
.B(n_54),
.Y(n_66)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_20),
.B(n_11),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_55),
.B(n_40),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_20),
.B(n_1),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_45),
.A2(n_15),
.B1(n_24),
.B2(n_27),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_57),
.A2(n_68),
.B1(n_70),
.B2(n_73),
.Y(n_108)
);

CKINVDCx6p67_ASAP7_75t_R g60 ( 
.A(n_33),
.Y(n_60)
);

INVx3_ASAP7_75t_SL g102 ( 
.A(n_60),
.Y(n_102)
);

INVx6_ASAP7_75t_SL g64 ( 
.A(n_31),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_64),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_53),
.A2(n_43),
.B1(n_40),
.B2(n_15),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_51),
.A2(n_24),
.B1(n_27),
.B2(n_12),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_L g73 ( 
.A1(n_39),
.A2(n_16),
.B1(n_12),
.B2(n_2),
.Y(n_73)
);

BUFx12_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_74),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_16),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_81),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_41),
.B(n_2),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_46),
.B(n_38),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_84),
.B(n_87),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_35),
.B(n_38),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_88),
.B(n_72),
.Y(n_96)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_66),
.B(n_69),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_92),
.B(n_100),
.Y(n_120)
);

AOI32xp33_ASAP7_75t_L g93 ( 
.A1(n_71),
.A2(n_62),
.A3(n_73),
.B1(n_61),
.B2(n_70),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_93),
.B(n_106),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_57),
.A2(n_68),
.B(n_60),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_94),
.A2(n_79),
.B(n_77),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_95),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_96),
.B(n_109),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_76),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_104),
.Y(n_112)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_59),
.B(n_63),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_80),
.B(n_65),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_101),
.B(n_58),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_83),
.B(n_78),
.Y(n_103)
);

AND2x2_ASAP7_75t_SL g118 ( 
.A(n_103),
.B(n_74),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_85),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_60),
.B(n_85),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_SL g117 ( 
.A(n_105),
.B(n_74),
.C(n_103),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_78),
.B(n_82),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_107),
.Y(n_116)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_105),
.B(n_78),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_113),
.B(n_118),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_115),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_117),
.B(n_102),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_90),
.B(n_89),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_121),
.B(n_124),
.Y(n_133)
);

NOR2x1_ASAP7_75t_L g123 ( 
.A(n_96),
.B(n_108),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_123),
.A2(n_102),
.B(n_91),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_110),
.B(n_96),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_94),
.A2(n_98),
.B1(n_104),
.B2(n_107),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_125),
.A2(n_99),
.B1(n_109),
.B2(n_122),
.Y(n_137)
);

AND2x6_ASAP7_75t_L g126 ( 
.A(n_119),
.B(n_110),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_126),
.B(n_132),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g127 ( 
.A(n_113),
.B(n_103),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_127),
.B(n_128),
.C(n_131),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_119),
.B(n_97),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_116),
.Y(n_129)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_129),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_117),
.B(n_97),
.C(n_102),
.Y(n_131)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_116),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_134),
.B(n_137),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_135),
.B(n_118),
.C(n_112),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_133),
.A2(n_125),
.B1(n_112),
.B2(n_123),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_139),
.A2(n_143),
.B1(n_127),
.B2(n_111),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_142),
.B(n_146),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_136),
.A2(n_115),
.B1(n_120),
.B2(n_122),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_136),
.Y(n_144)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_144),
.Y(n_152)
);

A2O1A1Ixp33_ASAP7_75t_L g146 ( 
.A1(n_126),
.A2(n_122),
.B(n_120),
.C(n_118),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_145),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_147),
.B(n_148),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_146),
.A2(n_128),
.B1(n_135),
.B2(n_131),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_SL g149 ( 
.A(n_140),
.B(n_130),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_149),
.B(n_140),
.C(n_138),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_151),
.B(n_142),
.Y(n_154)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_141),
.Y(n_153)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_153),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_154),
.B(n_149),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_156),
.B(n_150),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_152),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_157),
.B(n_145),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_159),
.B(n_154),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_155),
.A2(n_138),
.B(n_150),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_160),
.B(n_162),
.C(n_156),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_161),
.B(n_158),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_163),
.A2(n_111),
.B(n_148),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_164),
.B(n_165),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_167),
.A2(n_159),
.B(n_164),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_168),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_169),
.B(n_166),
.Y(n_170)
);


endmodule