module fake_jpeg_30997_n_194 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_194);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_194;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_5),
.B(n_10),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_17),
.B(n_13),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_35),
.B(n_50),
.Y(n_64)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_40),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_43),
.Y(n_65)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_17),
.B(n_0),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_45),
.B(n_49),
.Y(n_55)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_14),
.B(n_0),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_31),
.B(n_1),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_52),
.B(n_28),
.Y(n_58)
);

INVx4_ASAP7_75t_SL g53 ( 
.A(n_20),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_53),
.B(n_1),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_14),
.B(n_1),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_54),
.B(n_21),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_36),
.A2(n_28),
.B1(n_18),
.B2(n_24),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_57),
.A2(n_61),
.B1(n_41),
.B2(n_40),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_58),
.B(n_2),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_52),
.A2(n_27),
.B(n_18),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_60),
.B(n_39),
.C(n_43),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_47),
.A2(n_28),
.B1(n_24),
.B2(n_15),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_53),
.A2(n_24),
.B1(n_33),
.B2(n_16),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_66),
.A2(n_81),
.B1(n_83),
.B2(n_42),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_45),
.A2(n_25),
.B1(n_32),
.B2(n_30),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_68),
.A2(n_71),
.B1(n_75),
.B2(n_41),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_49),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_69),
.B(n_78),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_51),
.A2(n_25),
.B1(n_32),
.B2(n_30),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_37),
.A2(n_21),
.B1(n_33),
.B2(n_22),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_29),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_82),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_53),
.A2(n_29),
.B1(n_22),
.B2(n_19),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_48),
.B(n_19),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_44),
.A2(n_16),
.B1(n_2),
.B2(n_4),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_84),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

INVx13_ASAP7_75t_L g114 ( 
.A(n_86),
.Y(n_114)
);

OA22x2_ASAP7_75t_L g87 ( 
.A1(n_57),
.A2(n_61),
.B1(n_60),
.B2(n_74),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_87),
.A2(n_79),
.B1(n_59),
.B2(n_67),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_88),
.A2(n_107),
.B1(n_109),
.B2(n_65),
.Y(n_123)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_89),
.Y(n_121)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_90),
.Y(n_124)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_91),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_92),
.B(n_108),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_64),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_94),
.B(n_99),
.Y(n_122)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g120 ( 
.A(n_96),
.Y(n_120)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_62),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_97),
.Y(n_111)
);

MAJx2_ASAP7_75t_L g98 ( 
.A(n_58),
.B(n_50),
.C(n_46),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_108),
.C(n_87),
.Y(n_116)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_56),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_72),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_101),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_102),
.A2(n_106),
.B1(n_85),
.B2(n_77),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_72),
.Y(n_103)
);

INVxp33_ASAP7_75t_L g115 ( 
.A(n_103),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_79),
.A2(n_34),
.B1(n_38),
.B2(n_6),
.Y(n_106)
);

INVx13_ASAP7_75t_L g107 ( 
.A(n_73),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_69),
.A2(n_65),
.B1(n_59),
.B2(n_70),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_93),
.B(n_55),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_104),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_SL g113 ( 
.A(n_92),
.B(n_55),
.C(n_7),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_113),
.B(n_116),
.C(n_98),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_117),
.A2(n_127),
.B1(n_102),
.B2(n_118),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_89),
.B(n_59),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_119),
.B(n_125),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_123),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_87),
.B(n_59),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_87),
.B(n_70),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_126),
.B(n_77),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_122),
.Y(n_130)
);

NAND3xp33_ASAP7_75t_L g156 ( 
.A(n_130),
.B(n_138),
.C(n_112),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_132),
.B(n_136),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_126),
.A2(n_94),
.B(n_90),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_133),
.A2(n_141),
.B(n_121),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_134),
.B(n_115),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_135),
.A2(n_111),
.B1(n_124),
.B2(n_128),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_129),
.B(n_97),
.C(n_99),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_129),
.B(n_105),
.C(n_96),
.Y(n_137)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_137),
.Y(n_160)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_121),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_125),
.Y(n_139)
);

NOR4xp25_ASAP7_75t_L g157 ( 
.A(n_139),
.B(n_140),
.C(n_142),
.D(n_10),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_110),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_117),
.A2(n_86),
.B(n_103),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_113),
.B(n_100),
.C(n_63),
.Y(n_142)
);

OAI21x1_ASAP7_75t_L g158 ( 
.A1(n_143),
.A2(n_144),
.B(n_12),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_122),
.B(n_95),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_127),
.A2(n_67),
.B1(n_91),
.B2(n_85),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_145),
.A2(n_112),
.B1(n_120),
.B2(n_114),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_119),
.A2(n_63),
.B1(n_107),
.B2(n_8),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_146),
.A2(n_111),
.B1(n_124),
.B2(n_128),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_148),
.B(n_156),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_149),
.A2(n_151),
.B1(n_145),
.B2(n_143),
.Y(n_169)
);

AOI322xp5_ASAP7_75t_SL g150 ( 
.A1(n_137),
.A2(n_114),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.C1(n_4),
.C2(n_12),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_150),
.B(n_152),
.Y(n_168)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_153),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_144),
.B(n_8),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_155),
.B(n_13),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_157),
.B(n_142),
.C(n_147),
.Y(n_165)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_158),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_141),
.A2(n_139),
.B1(n_135),
.B2(n_147),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_159),
.A2(n_132),
.B1(n_131),
.B2(n_133),
.Y(n_164)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_152),
.Y(n_163)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_163),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_164),
.A2(n_169),
.B1(n_160),
.B2(n_154),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_165),
.B(n_167),
.Y(n_174)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_153),
.Y(n_166)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_166),
.Y(n_173)
);

HB1xp67_ASAP7_75t_L g171 ( 
.A(n_161),
.Y(n_171)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_171),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g175 ( 
.A(n_164),
.B(n_154),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_175),
.B(n_160),
.Y(n_179)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_163),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_176),
.B(n_155),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_177),
.A2(n_136),
.B1(n_148),
.B2(n_131),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_171),
.A2(n_166),
.B1(n_161),
.B2(n_159),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_178),
.B(n_182),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_179),
.B(n_181),
.Y(n_186)
);

NOR3xp33_ASAP7_75t_L g184 ( 
.A(n_180),
.B(n_170),
.C(n_162),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_184),
.B(n_170),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_180),
.A2(n_162),
.B1(n_172),
.B2(n_173),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_185),
.B(n_178),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_187),
.B(n_188),
.Y(n_190)
);

NAND4xp25_ASAP7_75t_L g189 ( 
.A(n_186),
.B(n_149),
.C(n_168),
.D(n_174),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_189),
.A2(n_165),
.B(n_183),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_191),
.A2(n_175),
.B(n_179),
.Y(n_192)
);

AOI31xp33_ASAP7_75t_L g193 ( 
.A1(n_192),
.A2(n_190),
.A3(n_187),
.B(n_167),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_193),
.B(n_138),
.Y(n_194)
);


endmodule