module fake_netlist_5_296_n_2001 (n_137, n_168, n_164, n_191, n_91, n_82, n_122, n_194, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_188, n_190, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_196, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_2001);

input n_137;
input n_168;
input n_164;
input n_191;
input n_91;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_188;
input n_190;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_196;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_2001;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_1960;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_1949;
wire n_343;
wire n_1449;
wire n_308;
wire n_1946;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_1948;
wire n_1984;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_798;
wire n_350;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_1931;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1986;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1971;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1978;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_759;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1963;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_1916;
wire n_293;
wire n_677;
wire n_372;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_433;
wire n_604;
wire n_368;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_1874;
wire n_563;
wire n_1987;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_1989;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1980;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_239;
wire n_630;
wire n_1902;
wire n_1941;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1958;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_968;
wire n_315;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_1974;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1966;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1992;
wire n_1643;
wire n_883;
wire n_1983;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1400;
wire n_1342;
wire n_900;
wire n_856;
wire n_1793;
wire n_1976;
wire n_918;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_681;
wire n_584;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_1998;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_1968;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_707;
wire n_1168;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1988;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_1999;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1985;
wire n_1898;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1981;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1995;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_685;
wire n_598;
wire n_928;
wire n_608;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_1975;
wire n_273;
wire n_1937;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_1936;
wire n_1956;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1969;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1990;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx1_ASAP7_75t_L g198 ( 
.A(n_56),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_175),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_162),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_14),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_95),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_88),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_97),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_23),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_189),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_127),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_13),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_89),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_22),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_39),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_41),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_110),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_30),
.Y(n_214)
);

BUFx10_ASAP7_75t_L g215 ( 
.A(n_158),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_112),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_58),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_166),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_174),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_91),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_63),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_136),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g223 ( 
.A(n_44),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_18),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_80),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_13),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_187),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_116),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_98),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_167),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_23),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_42),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_77),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_26),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_1),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_120),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_143),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_177),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_152),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_172),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_27),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_111),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_90),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_118),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_124),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_93),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_74),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_100),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_178),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_161),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_72),
.Y(n_251)
);

BUFx10_ASAP7_75t_L g252 ( 
.A(n_180),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_145),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_20),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_101),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_30),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_115),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_195),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_134),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_140),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_62),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_163),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_103),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_32),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_45),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_135),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_67),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_109),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_156),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_77),
.Y(n_270)
);

BUFx10_ASAP7_75t_L g271 ( 
.A(n_104),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_82),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_99),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_12),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_108),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_58),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_37),
.Y(n_277)
);

INVx2_ASAP7_75t_SL g278 ( 
.A(n_179),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_170),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_69),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_11),
.Y(n_281)
);

BUFx5_ASAP7_75t_L g282 ( 
.A(n_62),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_168),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_86),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_130),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_7),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_68),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_92),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_117),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_173),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_64),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_194),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_121),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_52),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_28),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_150),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_169),
.Y(n_297)
);

BUFx2_ASAP7_75t_L g298 ( 
.A(n_36),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_41),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_27),
.Y(n_300)
);

BUFx10_ASAP7_75t_L g301 ( 
.A(n_26),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_3),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_36),
.Y(n_303)
);

INVx1_ASAP7_75t_SL g304 ( 
.A(n_141),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_122),
.Y(n_305)
);

BUFx2_ASAP7_75t_L g306 ( 
.A(n_128),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_9),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_154),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_126),
.Y(n_309)
);

BUFx2_ASAP7_75t_L g310 ( 
.A(n_159),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_31),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_38),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_59),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_153),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_46),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_125),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_10),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_6),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_72),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_83),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_196),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_42),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_6),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_87),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_142),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_107),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_191),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_47),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_69),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_4),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_61),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_2),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_7),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_35),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g335 ( 
.A(n_11),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_144),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_40),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_131),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_43),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_183),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_149),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_50),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_73),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_20),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_19),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_84),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_68),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_8),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_186),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_57),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_176),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_137),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_9),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_19),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_114),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_57),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_47),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_164),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_73),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_59),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_78),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_76),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_1),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_70),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_74),
.Y(n_365)
);

BUFx5_ASAP7_75t_L g366 ( 
.A(n_96),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_17),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_75),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_22),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_67),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_10),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_61),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_44),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_35),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_182),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_146),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_193),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_190),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_32),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_79),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_33),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_14),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_151),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_113),
.Y(n_384)
);

INVx1_ASAP7_75t_SL g385 ( 
.A(n_147),
.Y(n_385)
);

BUFx2_ASAP7_75t_L g386 ( 
.A(n_132),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_53),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_105),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_60),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_3),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_71),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_21),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_94),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_33),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_282),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_248),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_306),
.B(n_0),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_250),
.Y(n_398)
);

HB1xp67_ASAP7_75t_L g399 ( 
.A(n_335),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_255),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_282),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_207),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_282),
.B(n_0),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_243),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_253),
.Y(n_405)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_223),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_282),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_258),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_282),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_298),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_282),
.Y(n_411)
);

BUFx3_ASAP7_75t_L g412 ( 
.A(n_308),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_259),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_257),
.Y(n_414)
);

INVxp67_ASAP7_75t_SL g415 ( 
.A(n_242),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_260),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_282),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_282),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_262),
.Y(n_419)
);

INVx2_ASAP7_75t_SL g420 ( 
.A(n_301),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_305),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_198),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_201),
.Y(n_423)
);

BUFx2_ASAP7_75t_L g424 ( 
.A(n_205),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_201),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_263),
.Y(n_426)
);

INVxp33_ASAP7_75t_SL g427 ( 
.A(n_205),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_208),
.Y(n_428)
);

NOR2xp67_ASAP7_75t_L g429 ( 
.A(n_210),
.B(n_2),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_266),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_201),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_201),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_268),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_269),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_272),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_366),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_201),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_214),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_324),
.Y(n_439)
);

NOR2xp67_ASAP7_75t_L g440 ( 
.A(n_210),
.B(n_4),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_214),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_338),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_214),
.Y(n_443)
);

NOR2xp67_ASAP7_75t_L g444 ( 
.A(n_270),
.B(n_5),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_273),
.Y(n_445)
);

CKINVDCx14_ASAP7_75t_R g446 ( 
.A(n_310),
.Y(n_446)
);

INVxp67_ASAP7_75t_SL g447 ( 
.A(n_386),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_279),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_366),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_366),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_214),
.Y(n_451)
);

INVxp67_ASAP7_75t_SL g452 ( 
.A(n_308),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_214),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_283),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_312),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_284),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_312),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_341),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_278),
.B(n_5),
.Y(n_459)
);

INVxp67_ASAP7_75t_SL g460 ( 
.A(n_312),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_376),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_288),
.Y(n_462)
);

BUFx2_ASAP7_75t_L g463 ( 
.A(n_211),
.Y(n_463)
);

INVxp67_ASAP7_75t_SL g464 ( 
.A(n_312),
.Y(n_464)
);

INVxp67_ASAP7_75t_SL g465 ( 
.A(n_312),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_270),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_388),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_292),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_277),
.Y(n_469)
);

INVxp67_ASAP7_75t_SL g470 ( 
.A(n_202),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_277),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_278),
.B(n_8),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_297),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_345),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_309),
.Y(n_475)
);

HB1xp67_ASAP7_75t_L g476 ( 
.A(n_211),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_314),
.Y(n_477)
);

INVxp67_ASAP7_75t_L g478 ( 
.A(n_235),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_225),
.B(n_12),
.Y(n_479)
);

NOR2xp67_ASAP7_75t_L g480 ( 
.A(n_345),
.B(n_15),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_316),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_321),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_366),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_325),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_373),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_373),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_326),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_346),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_R g489 ( 
.A(n_349),
.B(n_200),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_247),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_261),
.Y(n_491)
);

HB1xp67_ASAP7_75t_L g492 ( 
.A(n_212),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_379),
.Y(n_493)
);

BUFx2_ASAP7_75t_L g494 ( 
.A(n_212),
.Y(n_494)
);

INVxp33_ASAP7_75t_SL g495 ( 
.A(n_217),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_379),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_470),
.B(n_225),
.Y(n_497)
);

BUFx8_ASAP7_75t_L g498 ( 
.A(n_424),
.Y(n_498)
);

AND2x2_ASAP7_75t_L g499 ( 
.A(n_460),
.B(n_228),
.Y(n_499)
);

NAND2xp33_ASAP7_75t_SL g500 ( 
.A(n_420),
.B(n_217),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_464),
.B(n_228),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_401),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_423),
.Y(n_503)
);

INVxp67_ASAP7_75t_L g504 ( 
.A(n_476),
.Y(n_504)
);

AND2x2_ASAP7_75t_L g505 ( 
.A(n_465),
.B(n_293),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_401),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_452),
.B(n_412),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_401),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_423),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_425),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_395),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_395),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_407),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_407),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_459),
.B(n_200),
.Y(n_515)
);

AND2x4_ASAP7_75t_L g516 ( 
.A(n_425),
.B(n_293),
.Y(n_516)
);

AND2x4_ASAP7_75t_L g517 ( 
.A(n_431),
.B(n_204),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_409),
.Y(n_518)
);

INVx6_ASAP7_75t_L g519 ( 
.A(n_412),
.Y(n_519)
);

AND2x4_ASAP7_75t_L g520 ( 
.A(n_431),
.B(n_213),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_432),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_472),
.B(n_203),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_SL g523 ( 
.A(n_397),
.B(n_301),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_432),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_409),
.Y(n_525)
);

HB1xp67_ASAP7_75t_L g526 ( 
.A(n_399),
.Y(n_526)
);

INVx5_ASAP7_75t_L g527 ( 
.A(n_436),
.Y(n_527)
);

INVx3_ASAP7_75t_L g528 ( 
.A(n_411),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_437),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_411),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_437),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_417),
.Y(n_532)
);

HB1xp67_ASAP7_75t_L g533 ( 
.A(n_492),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_438),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_417),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_438),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_441),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_441),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_443),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_412),
.B(n_392),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_443),
.B(n_203),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_490),
.B(n_215),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_491),
.B(n_215),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_451),
.B(n_453),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_418),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_451),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_453),
.B(n_209),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_447),
.B(n_199),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_455),
.B(n_209),
.Y(n_549)
);

AND2x4_ASAP7_75t_L g550 ( 
.A(n_455),
.B(n_220),
.Y(n_550)
);

BUFx2_ASAP7_75t_L g551 ( 
.A(n_489),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_L g552 ( 
.A1(n_406),
.A2(n_394),
.B1(n_287),
.B2(n_344),
.Y(n_552)
);

INVxp67_ASAP7_75t_L g553 ( 
.A(n_424),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_457),
.B(n_216),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_418),
.Y(n_555)
);

AND2x4_ASAP7_75t_L g556 ( 
.A(n_457),
.B(n_237),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_479),
.B(n_216),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_436),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_466),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_436),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_466),
.Y(n_561)
);

AND2x4_ASAP7_75t_L g562 ( 
.A(n_403),
.B(n_238),
.Y(n_562)
);

INVx3_ASAP7_75t_L g563 ( 
.A(n_449),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_469),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_469),
.Y(n_565)
);

CKINVDCx20_ASAP7_75t_R g566 ( 
.A(n_402),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_471),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_420),
.B(n_215),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_403),
.B(n_218),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_449),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_471),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_474),
.B(n_218),
.Y(n_572)
);

NAND2x1p5_ASAP7_75t_L g573 ( 
.A(n_429),
.B(n_206),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_449),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_450),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_474),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_511),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_507),
.B(n_396),
.Y(n_578)
);

INVx3_ASAP7_75t_L g579 ( 
.A(n_502),
.Y(n_579)
);

AND2x4_ASAP7_75t_L g580 ( 
.A(n_562),
.B(n_244),
.Y(n_580)
);

BUFx2_ASAP7_75t_L g581 ( 
.A(n_526),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_511),
.Y(n_582)
);

INVx3_ASAP7_75t_L g583 ( 
.A(n_502),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_558),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_502),
.Y(n_585)
);

OAI22xp33_ASAP7_75t_L g586 ( 
.A1(n_523),
.A2(n_415),
.B1(n_406),
.B2(n_410),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_507),
.B(n_398),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_507),
.B(n_496),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_558),
.Y(n_589)
);

INVxp33_ASAP7_75t_L g590 ( 
.A(n_526),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_569),
.B(n_400),
.Y(n_591)
);

INVx2_ASAP7_75t_SL g592 ( 
.A(n_519),
.Y(n_592)
);

AOI22xp5_ASAP7_75t_L g593 ( 
.A1(n_523),
.A2(n_356),
.B1(n_347),
.B2(n_224),
.Y(n_593)
);

INVx5_ASAP7_75t_L g594 ( 
.A(n_512),
.Y(n_594)
);

BUFx3_ASAP7_75t_L g595 ( 
.A(n_519),
.Y(n_595)
);

INVx2_ASAP7_75t_SL g596 ( 
.A(n_519),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_558),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_560),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_569),
.B(n_499),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_548),
.B(n_408),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_499),
.B(n_413),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_511),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_560),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_514),
.Y(n_604)
);

INVx3_ASAP7_75t_L g605 ( 
.A(n_502),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_515),
.B(n_416),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_548),
.B(n_419),
.Y(n_607)
);

AND2x6_ASAP7_75t_L g608 ( 
.A(n_562),
.B(n_206),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_514),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_514),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_502),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_560),
.Y(n_612)
);

INVx2_ASAP7_75t_SL g613 ( 
.A(n_519),
.Y(n_613)
);

OR2x6_ASAP7_75t_L g614 ( 
.A(n_562),
.B(n_245),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_530),
.Y(n_615)
);

INVx3_ASAP7_75t_L g616 ( 
.A(n_502),
.Y(n_616)
);

BUFx3_ASAP7_75t_L g617 ( 
.A(n_519),
.Y(n_617)
);

AND2x6_ASAP7_75t_L g618 ( 
.A(n_562),
.B(n_206),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_570),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_551),
.B(n_426),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_499),
.B(n_430),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_568),
.B(n_433),
.Y(n_622)
);

BUFx6f_ASAP7_75t_L g623 ( 
.A(n_502),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_515),
.B(n_434),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_570),
.Y(n_625)
);

AND2x2_ASAP7_75t_L g626 ( 
.A(n_540),
.B(n_485),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_501),
.B(n_435),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_570),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_501),
.B(n_445),
.Y(n_629)
);

BUFx10_ASAP7_75t_L g630 ( 
.A(n_562),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_501),
.B(n_448),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_574),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_574),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_557),
.B(n_454),
.Y(n_634)
);

INVx3_ASAP7_75t_L g635 ( 
.A(n_506),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_574),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_540),
.B(n_485),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_575),
.Y(n_638)
);

BUFx2_ASAP7_75t_L g639 ( 
.A(n_553),
.Y(n_639)
);

AOI22xp33_ASAP7_75t_L g640 ( 
.A1(n_497),
.A2(n_429),
.B1(n_444),
.B2(n_440),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_557),
.B(n_456),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_522),
.B(n_462),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_575),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_522),
.B(n_468),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_575),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_540),
.B(n_496),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_505),
.B(n_473),
.Y(n_647)
);

AND2x6_ASAP7_75t_L g648 ( 
.A(n_497),
.B(n_206),
.Y(n_648)
);

NAND2xp33_ASAP7_75t_L g649 ( 
.A(n_497),
.B(n_477),
.Y(n_649)
);

INVxp33_ASAP7_75t_L g650 ( 
.A(n_552),
.Y(n_650)
);

INVxp33_ASAP7_75t_L g651 ( 
.A(n_552),
.Y(n_651)
);

OAI22x1_ASAP7_75t_L g652 ( 
.A1(n_553),
.A2(n_494),
.B1(n_463),
.B2(n_224),
.Y(n_652)
);

BUFx6f_ASAP7_75t_L g653 ( 
.A(n_506),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_530),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_504),
.B(n_495),
.Y(n_655)
);

NAND3xp33_ASAP7_75t_L g656 ( 
.A(n_504),
.B(n_446),
.C(n_463),
.Y(n_656)
);

BUFx2_ASAP7_75t_L g657 ( 
.A(n_498),
.Y(n_657)
);

INVx3_ASAP7_75t_L g658 ( 
.A(n_506),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_530),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_506),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_542),
.B(n_427),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_543),
.B(n_475),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_505),
.B(n_528),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_505),
.B(n_304),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_532),
.Y(n_665)
);

INVx1_ASAP7_75t_SL g666 ( 
.A(n_566),
.Y(n_666)
);

BUFx6f_ASAP7_75t_L g667 ( 
.A(n_506),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_563),
.Y(n_668)
);

NAND2xp33_ASAP7_75t_L g669 ( 
.A(n_541),
.B(n_206),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_498),
.B(n_481),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_498),
.B(n_482),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_563),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_498),
.B(n_484),
.Y(n_673)
);

NAND2xp33_ASAP7_75t_L g674 ( 
.A(n_541),
.B(n_219),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_532),
.Y(n_675)
);

OR2x6_ASAP7_75t_L g676 ( 
.A(n_572),
.B(n_246),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_532),
.Y(n_677)
);

AOI22xp33_ASAP7_75t_L g678 ( 
.A1(n_517),
.A2(n_440),
.B1(n_444),
.B2(n_480),
.Y(n_678)
);

INVx4_ASAP7_75t_L g679 ( 
.A(n_527),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_528),
.B(n_385),
.Y(n_680)
);

BUFx2_ASAP7_75t_L g681 ( 
.A(n_498),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_528),
.B(n_249),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_500),
.B(n_487),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_572),
.B(n_486),
.Y(n_684)
);

INVx3_ASAP7_75t_L g685 ( 
.A(n_506),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_563),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_563),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_547),
.B(n_488),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_547),
.B(n_494),
.Y(n_689)
);

BUFx6f_ASAP7_75t_SL g690 ( 
.A(n_517),
.Y(n_690)
);

INVx3_ASAP7_75t_L g691 ( 
.A(n_506),
.Y(n_691)
);

INVx4_ASAP7_75t_L g692 ( 
.A(n_527),
.Y(n_692)
);

OR2x6_ASAP7_75t_L g693 ( 
.A(n_549),
.B(n_275),
.Y(n_693)
);

INVx2_ASAP7_75t_SL g694 ( 
.A(n_533),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_528),
.B(n_285),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_508),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_535),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_549),
.B(n_289),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_508),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_508),
.Y(n_700)
);

BUFx6f_ASAP7_75t_L g701 ( 
.A(n_508),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_508),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_554),
.B(n_252),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_554),
.B(n_404),
.Y(n_704)
);

OR2x6_ASAP7_75t_L g705 ( 
.A(n_573),
.B(n_290),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_535),
.Y(n_706)
);

BUFx10_ASAP7_75t_L g707 ( 
.A(n_533),
.Y(n_707)
);

INVx2_ASAP7_75t_SL g708 ( 
.A(n_573),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_535),
.Y(n_709)
);

INVx2_ASAP7_75t_SL g710 ( 
.A(n_573),
.Y(n_710)
);

INVx3_ASAP7_75t_L g711 ( 
.A(n_508),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_508),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_545),
.Y(n_713)
);

INVx2_ASAP7_75t_SL g714 ( 
.A(n_573),
.Y(n_714)
);

BUFx2_ASAP7_75t_L g715 ( 
.A(n_517),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_545),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_545),
.B(n_320),
.Y(n_717)
);

INVx3_ASAP7_75t_L g718 ( 
.A(n_512),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_555),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_517),
.B(n_252),
.Y(n_720)
);

INVx4_ASAP7_75t_L g721 ( 
.A(n_527),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_555),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_555),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_503),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_503),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_512),
.Y(n_726)
);

AOI22xp33_ASAP7_75t_L g727 ( 
.A1(n_517),
.A2(n_520),
.B1(n_556),
.B2(n_550),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_520),
.B(n_252),
.Y(n_728)
);

AND2x6_ASAP7_75t_L g729 ( 
.A(n_580),
.B(n_219),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_606),
.B(n_624),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_626),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_724),
.Y(n_732)
);

BUFx6f_ASAP7_75t_L g733 ( 
.A(n_595),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_694),
.B(n_689),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_644),
.B(n_512),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_599),
.B(n_512),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_708),
.B(n_512),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_708),
.B(n_512),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_724),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_710),
.B(n_513),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_630),
.B(n_513),
.Y(n_741)
);

INVx2_ASAP7_75t_SL g742 ( 
.A(n_707),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_666),
.Y(n_743)
);

AOI22xp5_ASAP7_75t_L g744 ( 
.A1(n_704),
.A2(n_414),
.B1(n_421),
.B2(n_405),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_630),
.B(n_513),
.Y(n_745)
);

BUFx3_ASAP7_75t_L g746 ( 
.A(n_715),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_591),
.B(n_439),
.Y(n_747)
);

HB1xp67_ASAP7_75t_L g748 ( 
.A(n_581),
.Y(n_748)
);

OAI22xp5_ASAP7_75t_L g749 ( 
.A1(n_601),
.A2(n_458),
.B1(n_461),
.B2(n_442),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_710),
.B(n_513),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_725),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_725),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_714),
.B(n_513),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_714),
.B(n_684),
.Y(n_754)
);

OR2x2_ASAP7_75t_L g755 ( 
.A(n_694),
.B(n_422),
.Y(n_755)
);

NAND2xp33_ASAP7_75t_L g756 ( 
.A(n_608),
.B(n_366),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_684),
.B(n_513),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_578),
.B(n_467),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_587),
.B(n_222),
.Y(n_759)
);

INVxp67_ASAP7_75t_L g760 ( 
.A(n_639),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_621),
.B(n_513),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_627),
.B(n_518),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_629),
.B(n_518),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_631),
.B(n_518),
.Y(n_764)
);

INVxp67_ASAP7_75t_L g765 ( 
.A(n_639),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_626),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_SL g767 ( 
.A(n_657),
.B(n_271),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_647),
.B(n_518),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_713),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_630),
.B(n_518),
.Y(n_770)
);

NOR2xp67_ASAP7_75t_L g771 ( 
.A(n_656),
.B(n_422),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_637),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_600),
.B(n_222),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_637),
.Y(n_774)
);

AOI22xp5_ASAP7_75t_L g775 ( 
.A1(n_649),
.A2(n_520),
.B1(n_550),
.B2(n_556),
.Y(n_775)
);

INVx2_ASAP7_75t_SL g776 ( 
.A(n_646),
.Y(n_776)
);

INVx5_ASAP7_75t_L g777 ( 
.A(n_679),
.Y(n_777)
);

HB1xp67_ASAP7_75t_L g778 ( 
.A(n_581),
.Y(n_778)
);

AOI22xp5_ASAP7_75t_L g779 ( 
.A1(n_715),
.A2(n_520),
.B1(n_550),
.B2(n_556),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_630),
.B(n_518),
.Y(n_780)
);

NAND2xp33_ASAP7_75t_L g781 ( 
.A(n_608),
.B(n_366),
.Y(n_781)
);

NOR2xp67_ASAP7_75t_L g782 ( 
.A(n_620),
.B(n_428),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_680),
.B(n_518),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_646),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_663),
.B(n_525),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_580),
.B(n_525),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_580),
.B(n_727),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_607),
.B(n_227),
.Y(n_788)
);

AOI22xp5_ASAP7_75t_L g789 ( 
.A1(n_642),
.A2(n_520),
.B1(n_550),
.B2(n_556),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_580),
.B(n_525),
.Y(n_790)
);

AOI22xp33_ASAP7_75t_L g791 ( 
.A1(n_614),
.A2(n_556),
.B1(n_550),
.B2(n_516),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_664),
.B(n_525),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_698),
.B(n_525),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_588),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_588),
.B(n_525),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_586),
.B(n_525),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_577),
.Y(n_797)
);

OAI22xp33_ASAP7_75t_L g798 ( 
.A1(n_676),
.A2(n_480),
.B1(n_327),
.B2(n_351),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_693),
.B(n_516),
.Y(n_799)
);

BUFx6f_ASAP7_75t_L g800 ( 
.A(n_595),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_693),
.B(n_516),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_693),
.B(n_516),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_634),
.B(n_227),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_693),
.B(n_516),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_641),
.B(n_229),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_693),
.B(n_509),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_676),
.B(n_509),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_726),
.B(n_219),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_577),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_582),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_726),
.B(n_219),
.Y(n_811)
);

INVx2_ASAP7_75t_SL g812 ( 
.A(n_707),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_582),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_602),
.Y(n_814)
);

AND2x4_ASAP7_75t_SL g815 ( 
.A(n_707),
.B(n_271),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_676),
.B(n_510),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_713),
.Y(n_817)
);

OR2x6_ASAP7_75t_L g818 ( 
.A(n_657),
.B(n_392),
.Y(n_818)
);

AND2x6_ASAP7_75t_SL g819 ( 
.A(n_676),
.B(n_241),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_590),
.B(n_229),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_688),
.B(n_230),
.Y(n_821)
);

OR2x2_ASAP7_75t_L g822 ( 
.A(n_655),
.B(n_428),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_602),
.Y(n_823)
);

INVx1_ASAP7_75t_SL g824 ( 
.A(n_707),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_713),
.Y(n_825)
);

BUFx3_ASAP7_75t_L g826 ( 
.A(n_595),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_676),
.B(n_510),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_703),
.B(n_230),
.Y(n_828)
);

INVx3_ASAP7_75t_L g829 ( 
.A(n_617),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_716),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_604),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_640),
.B(n_521),
.Y(n_832)
);

BUFx3_ASAP7_75t_L g833 ( 
.A(n_617),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_678),
.B(n_521),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_716),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_726),
.B(n_219),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_604),
.Y(n_837)
);

INVx3_ASAP7_75t_L g838 ( 
.A(n_617),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_592),
.B(n_524),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_696),
.B(n_699),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_661),
.B(n_236),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_592),
.B(n_596),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_622),
.B(n_236),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_596),
.B(n_524),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_613),
.B(n_529),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_716),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_650),
.B(n_478),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_723),
.Y(n_848)
);

INVx2_ASAP7_75t_SL g849 ( 
.A(n_614),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_723),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_613),
.B(n_529),
.Y(n_851)
);

OAI22xp5_ASAP7_75t_L g852 ( 
.A1(n_614),
.A2(n_380),
.B1(n_336),
.B2(n_393),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_SL g853 ( 
.A(n_696),
.B(n_340),
.Y(n_853)
);

OAI221xp5_ASAP7_75t_L g854 ( 
.A1(n_593),
.A2(n_478),
.B1(n_286),
.B2(n_276),
.C(n_256),
.Y(n_854)
);

AND2x4_ASAP7_75t_L g855 ( 
.A(n_614),
.B(n_559),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_651),
.B(n_683),
.Y(n_856)
);

AOI22xp5_ASAP7_75t_L g857 ( 
.A1(n_614),
.A2(n_239),
.B1(n_240),
.B2(n_296),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_648),
.B(n_696),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_609),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_728),
.B(n_720),
.Y(n_860)
);

AOI22xp33_ASAP7_75t_L g861 ( 
.A1(n_648),
.A2(n_366),
.B1(n_340),
.B2(n_254),
.Y(n_861)
);

BUFx2_ASAP7_75t_L g862 ( 
.A(n_681),
.Y(n_862)
);

A2O1A1Ixp33_ASAP7_75t_L g863 ( 
.A1(n_593),
.A2(n_368),
.B(n_251),
.C(n_295),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_648),
.B(n_531),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_648),
.B(n_531),
.Y(n_865)
);

INVx4_ASAP7_75t_L g866 ( 
.A(n_690),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_699),
.B(n_340),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_648),
.B(n_534),
.Y(n_868)
);

OAI22xp5_ASAP7_75t_L g869 ( 
.A1(n_705),
.A2(n_296),
.B1(n_375),
.B2(n_377),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_609),
.Y(n_870)
);

INVx3_ASAP7_75t_L g871 ( 
.A(n_585),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_699),
.B(n_340),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_648),
.B(n_534),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_723),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_584),
.Y(n_875)
);

OAI22xp33_ASAP7_75t_L g876 ( 
.A1(n_705),
.A2(n_337),
.B1(n_322),
.B2(n_319),
.Y(n_876)
);

INVxp67_ASAP7_75t_L g877 ( 
.A(n_652),
.Y(n_877)
);

INVxp67_ASAP7_75t_L g878 ( 
.A(n_652),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_584),
.Y(n_879)
);

INVxp67_ASAP7_75t_L g880 ( 
.A(n_662),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_610),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_648),
.B(n_536),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_L g883 ( 
.A(n_705),
.B(n_239),
.Y(n_883)
);

O2A1O1Ixp33_ASAP7_75t_L g884 ( 
.A1(n_669),
.A2(n_334),
.B(n_359),
.C(n_362),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_700),
.B(n_536),
.Y(n_885)
);

BUFx6f_ASAP7_75t_L g886 ( 
.A(n_585),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_700),
.B(n_537),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_700),
.B(n_537),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_705),
.B(n_240),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_702),
.B(n_538),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_L g891 ( 
.A(n_705),
.B(n_352),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_670),
.B(n_301),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_610),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_702),
.B(n_538),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_584),
.Y(n_895)
);

AOI22xp33_ASAP7_75t_L g896 ( 
.A1(n_608),
.A2(n_366),
.B1(n_340),
.B2(n_369),
.Y(n_896)
);

OR2x2_ASAP7_75t_L g897 ( 
.A(n_671),
.B(n_221),
.Y(n_897)
);

AOI22xp33_ASAP7_75t_L g898 ( 
.A1(n_608),
.A2(n_370),
.B1(n_374),
.B2(n_300),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_702),
.B(n_352),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_712),
.B(n_355),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_734),
.B(n_847),
.Y(n_901)
);

A2O1A1Ixp33_ASAP7_75t_L g902 ( 
.A1(n_730),
.A2(n_695),
.B(n_682),
.C(n_673),
.Y(n_902)
);

OAI21xp5_ASAP7_75t_L g903 ( 
.A1(n_757),
.A2(n_660),
.B(n_712),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_754),
.B(n_712),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_737),
.A2(n_740),
.B(n_738),
.Y(n_905)
);

OAI21xp33_ASAP7_75t_L g906 ( 
.A1(n_821),
.A2(n_841),
.B(n_755),
.Y(n_906)
);

HB1xp67_ASAP7_75t_L g907 ( 
.A(n_748),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_776),
.B(n_615),
.Y(n_908)
);

BUFx6f_ASAP7_75t_L g909 ( 
.A(n_886),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_750),
.A2(n_753),
.B(n_736),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_776),
.B(n_615),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_759),
.B(n_654),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_746),
.B(n_856),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_735),
.A2(n_623),
.B(n_585),
.Y(n_914)
);

A2O1A1Ixp33_ASAP7_75t_L g915 ( 
.A1(n_860),
.A2(n_660),
.B(n_674),
.C(n_616),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_732),
.B(n_654),
.Y(n_916)
);

OAI21xp5_ASAP7_75t_L g917 ( 
.A1(n_785),
.A2(n_665),
.B(n_659),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_761),
.A2(n_623),
.B(n_585),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_732),
.Y(n_919)
);

O2A1O1Ixp5_ASAP7_75t_L g920 ( 
.A1(n_796),
.A2(n_717),
.B(n_665),
.C(n_719),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_739),
.B(n_659),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_739),
.B(n_675),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_751),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_762),
.A2(n_623),
.B(n_585),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_751),
.B(n_675),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_752),
.B(n_677),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_746),
.B(n_355),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_752),
.B(n_677),
.Y(n_928)
);

OAI21xp5_ASAP7_75t_L g929 ( 
.A1(n_785),
.A2(n_706),
.B(n_697),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_760),
.B(n_718),
.Y(n_930)
);

INVx1_ASAP7_75t_SL g931 ( 
.A(n_778),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_763),
.B(n_697),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_764),
.A2(n_623),
.B(n_585),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_768),
.A2(n_653),
.B(n_623),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_794),
.B(n_706),
.Y(n_935)
);

BUFx6f_ASAP7_75t_L g936 ( 
.A(n_886),
.Y(n_936)
);

NOR2xp67_ASAP7_75t_L g937 ( 
.A(n_880),
.B(n_709),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_743),
.Y(n_938)
);

OAI21xp5_ASAP7_75t_L g939 ( 
.A1(n_795),
.A2(n_719),
.B(n_709),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_731),
.B(n_722),
.Y(n_940)
);

BUFx4f_ASAP7_75t_L g941 ( 
.A(n_862),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_766),
.B(n_722),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_787),
.A2(n_653),
.B(n_623),
.Y(n_943)
);

OAI21x1_ASAP7_75t_L g944 ( 
.A1(n_840),
.A2(n_583),
.B(n_579),
.Y(n_944)
);

O2A1O1Ixp33_ASAP7_75t_L g945 ( 
.A1(n_796),
.A2(n_597),
.B(n_625),
.C(n_628),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_772),
.B(n_579),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_L g947 ( 
.A(n_765),
.B(n_718),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_797),
.Y(n_948)
);

O2A1O1Ixp33_ASAP7_75t_L g949 ( 
.A1(n_787),
.A2(n_597),
.B(n_625),
.C(n_628),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_774),
.B(n_579),
.Y(n_950)
);

INVx2_ASAP7_75t_SL g951 ( 
.A(n_822),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_784),
.B(n_579),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_773),
.B(n_583),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_788),
.B(n_583),
.Y(n_954)
);

OAI22xp5_ASAP7_75t_L g955 ( 
.A1(n_779),
.A2(n_849),
.B1(n_834),
.B2(n_832),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_758),
.B(n_820),
.Y(n_956)
);

OAI21xp5_ASAP7_75t_L g957 ( 
.A1(n_792),
.A2(n_605),
.B(n_583),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_803),
.B(n_805),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_783),
.A2(n_667),
.B(n_653),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_SL g960 ( 
.A(n_743),
.B(n_824),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_747),
.B(n_559),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_741),
.A2(n_770),
.B(n_745),
.Y(n_962)
);

AOI21x1_ASAP7_75t_L g963 ( 
.A1(n_741),
.A2(n_597),
.B(n_589),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_745),
.A2(n_667),
.B(n_653),
.Y(n_964)
);

AND2x4_ASAP7_75t_L g965 ( 
.A(n_855),
.B(n_561),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_770),
.A2(n_667),
.B(n_653),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_806),
.B(n_605),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_807),
.B(n_605),
.Y(n_968)
);

BUFx3_ASAP7_75t_L g969 ( 
.A(n_742),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_816),
.B(n_605),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_827),
.B(n_829),
.Y(n_971)
);

OAI321xp33_ASAP7_75t_L g972 ( 
.A1(n_854),
.A2(n_381),
.A3(n_363),
.B1(n_360),
.B2(n_353),
.C(n_348),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_L g973 ( 
.A(n_877),
.B(n_878),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_780),
.A2(n_667),
.B(n_653),
.Y(n_974)
);

INVx3_ASAP7_75t_L g975 ( 
.A(n_826),
.Y(n_975)
);

AND2x4_ASAP7_75t_L g976 ( 
.A(n_855),
.B(n_561),
.Y(n_976)
);

NOR2xp67_ASAP7_75t_L g977 ( 
.A(n_812),
.B(n_668),
.Y(n_977)
);

BUFx6f_ASAP7_75t_L g978 ( 
.A(n_886),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_829),
.B(n_611),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_L g980 ( 
.A(n_749),
.B(n_897),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_780),
.A2(n_701),
.B(n_667),
.Y(n_981)
);

O2A1O1Ixp33_ASAP7_75t_L g982 ( 
.A1(n_863),
.A2(n_900),
.B(n_899),
.C(n_801),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_809),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_792),
.A2(n_701),
.B(n_667),
.Y(n_984)
);

BUFx6f_ASAP7_75t_L g985 ( 
.A(n_886),
.Y(n_985)
);

AND2x4_ASAP7_75t_L g986 ( 
.A(n_855),
.B(n_849),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_829),
.B(n_611),
.Y(n_987)
);

OAI21xp5_ASAP7_75t_L g988 ( 
.A1(n_793),
.A2(n_616),
.B(n_611),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_838),
.A2(n_701),
.B(n_616),
.Y(n_989)
);

OAI21xp5_ASAP7_75t_L g990 ( 
.A1(n_793),
.A2(n_616),
.B(n_611),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_838),
.B(n_635),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_838),
.B(n_635),
.Y(n_992)
);

HB1xp67_ASAP7_75t_L g993 ( 
.A(n_799),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_786),
.A2(n_701),
.B(n_658),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_810),
.B(n_635),
.Y(n_995)
);

AO21x1_ASAP7_75t_L g996 ( 
.A1(n_883),
.A2(n_364),
.B(n_668),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_786),
.A2(n_701),
.B(n_658),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_790),
.A2(n_842),
.B(n_777),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_813),
.Y(n_999)
);

NOR2xp33_ASAP7_75t_SL g1000 ( 
.A(n_767),
.B(n_271),
.Y(n_1000)
);

O2A1O1Ixp33_ASAP7_75t_SL g1001 ( 
.A1(n_790),
.A2(n_685),
.B(n_711),
.C(n_691),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_814),
.B(n_635),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_823),
.B(n_831),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_777),
.A2(n_701),
.B(n_685),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_892),
.B(n_718),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_837),
.B(n_658),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_859),
.B(n_658),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_870),
.Y(n_1008)
);

INVx3_ASAP7_75t_L g1009 ( 
.A(n_826),
.Y(n_1009)
);

INVx3_ASAP7_75t_L g1010 ( 
.A(n_833),
.Y(n_1010)
);

OAI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_840),
.A2(n_691),
.B(n_685),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_881),
.B(n_685),
.Y(n_1012)
);

AOI22xp5_ASAP7_75t_L g1013 ( 
.A1(n_889),
.A2(n_690),
.B1(n_618),
.B2(n_608),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_769),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_893),
.B(n_691),
.Y(n_1015)
);

BUFx2_ASAP7_75t_SL g1016 ( 
.A(n_866),
.Y(n_1016)
);

INVxp67_ASAP7_75t_L g1017 ( 
.A(n_771),
.Y(n_1017)
);

OAI22xp5_ASAP7_75t_L g1018 ( 
.A1(n_775),
.A2(n_690),
.B1(n_711),
.B2(n_691),
.Y(n_1018)
);

INVxp67_ASAP7_75t_L g1019 ( 
.A(n_782),
.Y(n_1019)
);

OAI22xp5_ASAP7_75t_L g1020 ( 
.A1(n_789),
.A2(n_690),
.B1(n_711),
.B2(n_718),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_833),
.B(n_711),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_769),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_777),
.A2(n_721),
.B(n_692),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_828),
.B(n_608),
.Y(n_1024)
);

OAI22xp5_ASAP7_75t_L g1025 ( 
.A1(n_891),
.A2(n_378),
.B1(n_358),
.B2(n_383),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_777),
.A2(n_692),
.B(n_679),
.Y(n_1026)
);

OAI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_858),
.A2(n_598),
.B(n_589),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_777),
.A2(n_692),
.B(n_679),
.Y(n_1028)
);

AND2x2_ASAP7_75t_L g1029 ( 
.A(n_815),
.B(n_564),
.Y(n_1029)
);

CKINVDCx8_ASAP7_75t_R g1030 ( 
.A(n_819),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_815),
.B(n_564),
.Y(n_1031)
);

OR2x2_ASAP7_75t_L g1032 ( 
.A(n_744),
.B(n_565),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_802),
.A2(n_721),
.B(n_692),
.Y(n_1033)
);

INVxp67_ASAP7_75t_L g1034 ( 
.A(n_804),
.Y(n_1034)
);

A2O1A1Ixp33_ASAP7_75t_L g1035 ( 
.A1(n_843),
.A2(n_668),
.B(n_687),
.C(n_686),
.Y(n_1035)
);

NOR2x2_ASAP7_75t_L g1036 ( 
.A(n_818),
.B(n_221),
.Y(n_1036)
);

A2O1A1Ixp33_ASAP7_75t_L g1037 ( 
.A1(n_857),
.A2(n_672),
.B(n_687),
.C(n_686),
.Y(n_1037)
);

BUFx4f_ASAP7_75t_L g1038 ( 
.A(n_818),
.Y(n_1038)
);

O2A1O1Ixp33_ASAP7_75t_SL g1039 ( 
.A1(n_798),
.A2(n_687),
.B(n_686),
.C(n_672),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_817),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_L g1041 ( 
.A(n_869),
.B(n_672),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_825),
.B(n_830),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_825),
.B(n_608),
.Y(n_1043)
);

AOI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_899),
.A2(n_900),
.B1(n_791),
.B2(n_852),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_839),
.A2(n_721),
.B(n_679),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_844),
.A2(n_721),
.B(n_594),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_830),
.Y(n_1047)
);

OAI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_866),
.A2(n_375),
.B1(n_377),
.B2(n_378),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_835),
.B(n_618),
.Y(n_1049)
);

NAND2x1p5_ASAP7_75t_L g1050 ( 
.A(n_866),
.B(n_594),
.Y(n_1050)
);

A2O1A1Ixp33_ASAP7_75t_L g1051 ( 
.A1(n_863),
.A2(n_598),
.B(n_643),
.C(n_638),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_SL g1052 ( 
.A(n_733),
.B(n_589),
.Y(n_1052)
);

O2A1O1Ixp33_ASAP7_75t_L g1053 ( 
.A1(n_876),
.A2(n_645),
.B(n_643),
.C(n_638),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_835),
.B(n_618),
.Y(n_1054)
);

BUFx8_ASAP7_75t_L g1055 ( 
.A(n_729),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_846),
.B(n_618),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_846),
.B(n_618),
.Y(n_1057)
);

OAI21x1_ASAP7_75t_SL g1058 ( 
.A1(n_884),
.A2(n_603),
.B(n_598),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_848),
.B(n_618),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_845),
.A2(n_851),
.B(n_871),
.Y(n_1060)
);

O2A1O1Ixp33_ASAP7_75t_L g1061 ( 
.A1(n_808),
.A2(n_645),
.B(n_643),
.C(n_638),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_871),
.A2(n_594),
.B(n_527),
.Y(n_1062)
);

OAI21xp33_ASAP7_75t_L g1063 ( 
.A1(n_818),
.A2(n_231),
.B(n_226),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_848),
.B(n_618),
.Y(n_1064)
);

AO21x1_ASAP7_75t_L g1065 ( 
.A1(n_885),
.A2(n_612),
.B(n_603),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_SL g1066 ( 
.A(n_733),
.B(n_383),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_871),
.A2(n_594),
.B(n_527),
.Y(n_1067)
);

O2A1O1Ixp33_ASAP7_75t_L g1068 ( 
.A1(n_808),
.A2(n_645),
.B(n_636),
.C(n_633),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_733),
.A2(n_594),
.B(n_527),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_L g1070 ( 
.A(n_818),
.B(n_264),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_850),
.B(n_874),
.Y(n_1071)
);

NOR2xp33_ASAP7_75t_L g1072 ( 
.A(n_850),
.B(n_265),
.Y(n_1072)
);

NAND2xp33_ASAP7_75t_L g1073 ( 
.A(n_733),
.B(n_384),
.Y(n_1073)
);

AND2x4_ASAP7_75t_L g1074 ( 
.A(n_800),
.B(n_874),
.Y(n_1074)
);

AOI22xp5_ASAP7_75t_L g1075 ( 
.A1(n_864),
.A2(n_384),
.B1(n_633),
.B2(n_632),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_800),
.A2(n_594),
.B(n_527),
.Y(n_1076)
);

BUFx6f_ASAP7_75t_L g1077 ( 
.A(n_800),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_SL g1078 ( 
.A(n_800),
.B(n_565),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_L g1079 ( 
.A(n_875),
.B(n_267),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_887),
.A2(n_527),
.B(n_633),
.Y(n_1080)
);

A2O1A1Ixp33_ASAP7_75t_L g1081 ( 
.A1(n_888),
.A2(n_636),
.B(n_632),
.C(n_628),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_SL g1082 ( 
.A(n_865),
.B(n_567),
.Y(n_1082)
);

NOR2xp33_ASAP7_75t_L g1083 ( 
.A(n_875),
.B(n_274),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_890),
.A2(n_636),
.B(n_632),
.Y(n_1084)
);

INVx1_ASAP7_75t_SL g1085 ( 
.A(n_811),
.Y(n_1085)
);

NOR2xp33_ASAP7_75t_L g1086 ( 
.A(n_879),
.B(n_895),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_L g1087 ( 
.A(n_879),
.B(n_280),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_895),
.B(n_603),
.Y(n_1088)
);

AOI22xp33_ASAP7_75t_L g1089 ( 
.A1(n_756),
.A2(n_226),
.B1(n_231),
.B2(n_232),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_894),
.B(n_612),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_868),
.Y(n_1091)
);

OAI22xp5_ASAP7_75t_L g1092 ( 
.A1(n_861),
.A2(n_625),
.B1(n_619),
.B2(n_612),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_L g1093 ( 
.A(n_956),
.B(n_873),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_958),
.B(n_898),
.Y(n_1094)
);

HB1xp67_ASAP7_75t_L g1095 ( 
.A(n_907),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_901),
.B(n_729),
.Y(n_1096)
);

BUFx3_ASAP7_75t_L g1097 ( 
.A(n_938),
.Y(n_1097)
);

AOI22xp33_ASAP7_75t_L g1098 ( 
.A1(n_980),
.A2(n_729),
.B1(n_781),
.B2(n_756),
.Y(n_1098)
);

BUFx2_ASAP7_75t_L g1099 ( 
.A(n_907),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_961),
.B(n_729),
.Y(n_1100)
);

O2A1O1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_955),
.A2(n_811),
.B(n_836),
.C(n_872),
.Y(n_1101)
);

A2O1A1Ixp33_ASAP7_75t_L g1102 ( 
.A1(n_906),
.A2(n_980),
.B(n_982),
.C(n_1044),
.Y(n_1102)
);

A2O1A1Ixp33_ASAP7_75t_L g1103 ( 
.A1(n_962),
.A2(n_882),
.B(n_781),
.C(n_896),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_1014),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_919),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_910),
.A2(n_872),
.B(n_867),
.Y(n_1106)
);

O2A1O1Ixp33_ASAP7_75t_L g1107 ( 
.A1(n_902),
.A2(n_836),
.B(n_867),
.C(n_853),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_993),
.B(n_729),
.Y(n_1108)
);

AOI21xp33_ASAP7_75t_L g1109 ( 
.A1(n_951),
.A2(n_232),
.B(n_233),
.Y(n_1109)
);

BUFx3_ASAP7_75t_L g1110 ( 
.A(n_941),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_SL g1111 ( 
.A(n_986),
.B(n_571),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_1040),
.Y(n_1112)
);

OAI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_920),
.A2(n_853),
.B(n_619),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_993),
.B(n_729),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_1022),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_905),
.A2(n_619),
.B(n_544),
.Y(n_1116)
);

HB1xp67_ASAP7_75t_L g1117 ( 
.A(n_931),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_1034),
.B(n_576),
.Y(n_1118)
);

BUFx3_ASAP7_75t_L g1119 ( 
.A(n_941),
.Y(n_1119)
);

O2A1O1Ixp33_ASAP7_75t_L g1120 ( 
.A1(n_1034),
.A2(n_546),
.B(n_539),
.C(n_544),
.Y(n_1120)
);

BUFx6f_ASAP7_75t_L g1121 ( 
.A(n_909),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_937),
.B(n_576),
.Y(n_1122)
);

OAI22xp5_ASAP7_75t_L g1123 ( 
.A1(n_1005),
.A2(n_339),
.B1(n_281),
.B2(n_291),
.Y(n_1123)
);

NOR2xp33_ASAP7_75t_R g1124 ( 
.A(n_960),
.B(n_233),
.Y(n_1124)
);

AOI22xp5_ASAP7_75t_L g1125 ( 
.A1(n_913),
.A2(n_1017),
.B1(n_1005),
.B2(n_1019),
.Y(n_1125)
);

OR2x6_ASAP7_75t_L g1126 ( 
.A(n_1016),
.B(n_486),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_948),
.B(n_539),
.Y(n_1127)
);

NAND3xp33_ASAP7_75t_SL g1128 ( 
.A(n_1000),
.B(n_234),
.C(n_302),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_923),
.Y(n_1129)
);

INVx4_ASAP7_75t_L g1130 ( 
.A(n_1077),
.Y(n_1130)
);

INVx3_ASAP7_75t_L g1131 ( 
.A(n_1077),
.Y(n_1131)
);

BUFx12f_ASAP7_75t_L g1132 ( 
.A(n_1055),
.Y(n_1132)
);

NOR2xp33_ASAP7_75t_L g1133 ( 
.A(n_1019),
.B(n_294),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_1047),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_983),
.B(n_546),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_999),
.Y(n_1136)
);

INVx3_ASAP7_75t_L g1137 ( 
.A(n_1077),
.Y(n_1137)
);

O2A1O1Ixp33_ASAP7_75t_L g1138 ( 
.A1(n_912),
.A2(n_483),
.B(n_450),
.C(n_493),
.Y(n_1138)
);

AO32x2_ASAP7_75t_L g1139 ( 
.A1(n_1020),
.A2(n_15),
.A3(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_1139)
);

CKINVDCx16_ASAP7_75t_R g1140 ( 
.A(n_969),
.Y(n_1140)
);

OAI22xp5_ASAP7_75t_L g1141 ( 
.A1(n_1024),
.A2(n_342),
.B1(n_307),
.B2(n_311),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1008),
.B(n_299),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_1030),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_930),
.B(n_313),
.Y(n_1144)
);

AO21x1_ASAP7_75t_L g1145 ( 
.A1(n_953),
.A2(n_483),
.B(n_450),
.Y(n_1145)
);

BUFx6f_ASAP7_75t_L g1146 ( 
.A(n_909),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_SL g1147 ( 
.A(n_1038),
.B(n_315),
.Y(n_1147)
);

O2A1O1Ixp33_ASAP7_75t_L g1148 ( 
.A1(n_935),
.A2(n_483),
.B(n_493),
.C(n_317),
.Y(n_1148)
);

O2A1O1Ixp33_ASAP7_75t_L g1149 ( 
.A1(n_940),
.A2(n_350),
.B(n_318),
.C(n_323),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_954),
.A2(n_328),
.B(n_329),
.Y(n_1150)
);

AO22x1_ASAP7_75t_L g1151 ( 
.A1(n_973),
.A2(n_391),
.B1(n_390),
.B2(n_389),
.Y(n_1151)
);

OAI22x1_ASAP7_75t_L g1152 ( 
.A1(n_973),
.A2(n_391),
.B1(n_390),
.B2(n_389),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_930),
.B(n_330),
.Y(n_1153)
);

A2O1A1Ixp33_ASAP7_75t_L g1154 ( 
.A1(n_1041),
.A2(n_331),
.B(n_332),
.C(n_333),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_1074),
.Y(n_1155)
);

OAI22xp5_ASAP7_75t_L g1156 ( 
.A1(n_1091),
.A2(n_343),
.B1(n_382),
.B2(n_372),
.Y(n_1156)
);

OR2x2_ASAP7_75t_L g1157 ( 
.A(n_1032),
.B(n_302),
.Y(n_1157)
);

AOI21x1_ASAP7_75t_L g1158 ( 
.A1(n_971),
.A2(n_197),
.B(n_192),
.Y(n_1158)
);

INVxp67_ASAP7_75t_L g1159 ( 
.A(n_1029),
.Y(n_1159)
);

AND2x2_ASAP7_75t_L g1160 ( 
.A(n_1031),
.B(n_303),
.Y(n_1160)
);

NAND3xp33_ASAP7_75t_SL g1161 ( 
.A(n_1070),
.B(n_387),
.C(n_382),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_932),
.A2(n_387),
.B(n_372),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_908),
.Y(n_1163)
);

NOR2xp33_ASAP7_75t_L g1164 ( 
.A(n_1017),
.B(n_371),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_939),
.A2(n_371),
.B(n_367),
.Y(n_1165)
);

NOR2xp33_ASAP7_75t_L g1166 ( 
.A(n_1063),
.B(n_367),
.Y(n_1166)
);

OAI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_1003),
.A2(n_361),
.B1(n_357),
.B2(n_354),
.Y(n_1167)
);

OAI22xp5_ASAP7_75t_L g1168 ( 
.A1(n_975),
.A2(n_361),
.B1(n_357),
.B2(n_354),
.Y(n_1168)
);

INVx5_ASAP7_75t_L g1169 ( 
.A(n_909),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_911),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_947),
.B(n_365),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_946),
.Y(n_1172)
);

INVxp67_ASAP7_75t_L g1173 ( 
.A(n_927),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_950),
.Y(n_1174)
);

BUFx2_ASAP7_75t_L g1175 ( 
.A(n_965),
.Y(n_1175)
);

OAI22xp5_ASAP7_75t_L g1176 ( 
.A1(n_975),
.A2(n_365),
.B1(n_303),
.B2(n_188),
.Y(n_1176)
);

NOR2xp33_ASAP7_75t_L g1177 ( 
.A(n_1070),
.B(n_16),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_947),
.B(n_21),
.Y(n_1178)
);

O2A1O1Ixp33_ASAP7_75t_L g1179 ( 
.A1(n_942),
.A2(n_24),
.B(n_25),
.C(n_28),
.Y(n_1179)
);

OR2x6_ASAP7_75t_L g1180 ( 
.A(n_976),
.B(n_185),
.Y(n_1180)
);

OAI21x1_ASAP7_75t_L g1181 ( 
.A1(n_944),
.A2(n_184),
.B(n_181),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_952),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_916),
.Y(n_1183)
);

AOI21x1_ASAP7_75t_L g1184 ( 
.A1(n_914),
.A2(n_171),
.B(n_165),
.Y(n_1184)
);

INVx3_ASAP7_75t_L g1185 ( 
.A(n_1077),
.Y(n_1185)
);

AOI221xp5_ASAP7_75t_L g1186 ( 
.A1(n_1089),
.A2(n_24),
.B1(n_25),
.B2(n_29),
.C(n_31),
.Y(n_1186)
);

O2A1O1Ixp33_ASAP7_75t_SL g1187 ( 
.A1(n_1037),
.A2(n_160),
.B(n_157),
.C(n_155),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_1042),
.Y(n_1188)
);

NAND3xp33_ASAP7_75t_SL g1189 ( 
.A(n_1025),
.B(n_29),
.C(n_34),
.Y(n_1189)
);

BUFx2_ASAP7_75t_SL g1190 ( 
.A(n_976),
.Y(n_1190)
);

AO221x2_ASAP7_75t_L g1191 ( 
.A1(n_1048),
.A2(n_972),
.B1(n_1036),
.B2(n_38),
.C(n_39),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_918),
.A2(n_148),
.B(n_139),
.Y(n_1192)
);

AND2x2_ASAP7_75t_SL g1193 ( 
.A(n_1038),
.B(n_34),
.Y(n_1193)
);

AOI22xp33_ASAP7_75t_L g1194 ( 
.A1(n_996),
.A2(n_37),
.B1(n_40),
.B2(n_43),
.Y(n_1194)
);

BUFx2_ASAP7_75t_L g1195 ( 
.A(n_1009),
.Y(n_1195)
);

NOR2xp33_ASAP7_75t_L g1196 ( 
.A(n_1009),
.B(n_45),
.Y(n_1196)
);

A2O1A1Ixp33_ASAP7_75t_L g1197 ( 
.A1(n_1041),
.A2(n_46),
.B(n_48),
.C(n_49),
.Y(n_1197)
);

AOI22xp5_ASAP7_75t_L g1198 ( 
.A1(n_1066),
.A2(n_138),
.B1(n_133),
.B2(n_129),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_924),
.A2(n_119),
.B(n_106),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_SL g1200 ( 
.A(n_1010),
.B(n_123),
.Y(n_1200)
);

O2A1O1Ixp33_ASAP7_75t_L g1201 ( 
.A1(n_1051),
.A2(n_915),
.B(n_904),
.C(n_1035),
.Y(n_1201)
);

A2O1A1Ixp33_ASAP7_75t_L g1202 ( 
.A1(n_1072),
.A2(n_48),
.B(n_49),
.C(n_50),
.Y(n_1202)
);

BUFx2_ASAP7_75t_L g1203 ( 
.A(n_1010),
.Y(n_1203)
);

HB1xp67_ASAP7_75t_L g1204 ( 
.A(n_977),
.Y(n_1204)
);

AO32x1_ASAP7_75t_L g1205 ( 
.A1(n_1018),
.A2(n_51),
.A3(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_1205)
);

INVxp67_ASAP7_75t_SL g1206 ( 
.A(n_909),
.Y(n_1206)
);

BUFx2_ASAP7_75t_L g1207 ( 
.A(n_936),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_933),
.A2(n_85),
.B(n_81),
.Y(n_1208)
);

A2O1A1Ixp33_ASAP7_75t_L g1209 ( 
.A1(n_1072),
.A2(n_51),
.B(n_54),
.C(n_55),
.Y(n_1209)
);

BUFx6f_ASAP7_75t_L g1210 ( 
.A(n_936),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_934),
.A2(n_102),
.B(n_56),
.Y(n_1211)
);

A2O1A1Ixp33_ASAP7_75t_SL g1212 ( 
.A1(n_1079),
.A2(n_55),
.B(n_60),
.C(n_63),
.Y(n_1212)
);

A2O1A1Ixp33_ASAP7_75t_L g1213 ( 
.A1(n_1079),
.A2(n_64),
.B(n_65),
.C(n_66),
.Y(n_1213)
);

AOI22xp33_ASAP7_75t_L g1214 ( 
.A1(n_1083),
.A2(n_65),
.B1(n_66),
.B2(n_70),
.Y(n_1214)
);

AOI22xp33_ASAP7_75t_L g1215 ( 
.A1(n_1083),
.A2(n_71),
.B1(n_75),
.B2(n_76),
.Y(n_1215)
);

AOI22xp33_ASAP7_75t_L g1216 ( 
.A1(n_1087),
.A2(n_78),
.B1(n_1082),
.B2(n_970),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_921),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1087),
.B(n_967),
.Y(n_1218)
);

CKINVDCx11_ASAP7_75t_R g1219 ( 
.A(n_936),
.Y(n_1219)
);

NOR2xp33_ASAP7_75t_L g1220 ( 
.A(n_1085),
.B(n_968),
.Y(n_1220)
);

BUFx6f_ASAP7_75t_L g1221 ( 
.A(n_936),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1086),
.B(n_922),
.Y(n_1222)
);

INVx3_ASAP7_75t_L g1223 ( 
.A(n_978),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_959),
.A2(n_903),
.B(n_943),
.Y(n_1224)
);

O2A1O1Ixp5_ASAP7_75t_SL g1225 ( 
.A1(n_1052),
.A2(n_1078),
.B(n_917),
.C(n_929),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_1071),
.Y(n_1226)
);

AOI21x1_ASAP7_75t_L g1227 ( 
.A1(n_963),
.A2(n_1052),
.B(n_984),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_1058),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_SL g1229 ( 
.A(n_978),
.B(n_985),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_979),
.A2(n_987),
.B(n_991),
.Y(n_1230)
);

CKINVDCx14_ASAP7_75t_R g1231 ( 
.A(n_978),
.Y(n_1231)
);

O2A1O1Ixp5_ASAP7_75t_L g1232 ( 
.A1(n_1065),
.A2(n_920),
.B(n_1060),
.C(n_998),
.Y(n_1232)
);

NOR2x1_ASAP7_75t_L g1233 ( 
.A(n_1073),
.B(n_1021),
.Y(n_1233)
);

NOR2xp33_ASAP7_75t_R g1234 ( 
.A(n_1055),
.B(n_978),
.Y(n_1234)
);

CKINVDCx20_ASAP7_75t_R g1235 ( 
.A(n_985),
.Y(n_1235)
);

BUFx4f_ASAP7_75t_L g1236 ( 
.A(n_985),
.Y(n_1236)
);

NOR3xp33_ASAP7_75t_SL g1237 ( 
.A(n_994),
.B(n_997),
.C(n_1011),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1088),
.Y(n_1238)
);

NOR2xp33_ASAP7_75t_L g1239 ( 
.A(n_1089),
.B(n_1002),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_992),
.A2(n_1090),
.B(n_1027),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_925),
.A2(n_926),
.B(n_928),
.Y(n_1241)
);

O2A1O1Ixp33_ASAP7_75t_L g1242 ( 
.A1(n_1039),
.A2(n_1081),
.B(n_1053),
.C(n_945),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_989),
.A2(n_949),
.B(n_957),
.Y(n_1243)
);

HB1xp67_ASAP7_75t_L g1244 ( 
.A(n_985),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_995),
.Y(n_1245)
);

A2O1A1Ixp33_ASAP7_75t_L g1246 ( 
.A1(n_1013),
.A2(n_1075),
.B(n_1086),
.C(n_990),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1006),
.B(n_1012),
.Y(n_1247)
);

A2O1A1Ixp33_ASAP7_75t_L g1248 ( 
.A1(n_988),
.A2(n_964),
.B(n_966),
.C(n_974),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1007),
.Y(n_1249)
);

A2O1A1Ixp33_ASAP7_75t_L g1250 ( 
.A1(n_981),
.A2(n_1015),
.B(n_1068),
.C(n_1061),
.Y(n_1250)
);

O2A1O1Ixp33_ASAP7_75t_L g1251 ( 
.A1(n_1001),
.A2(n_1092),
.B(n_1056),
.C(n_1057),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1084),
.B(n_1064),
.Y(n_1252)
);

OAI22xp5_ASAP7_75t_L g1253 ( 
.A1(n_1043),
.A2(n_1059),
.B1(n_1054),
.B2(n_1049),
.Y(n_1253)
);

BUFx2_ASAP7_75t_L g1254 ( 
.A(n_1050),
.Y(n_1254)
);

OAI21x1_ASAP7_75t_L g1255 ( 
.A1(n_1227),
.A2(n_1004),
.B(n_1080),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1218),
.A2(n_1224),
.B(n_1241),
.Y(n_1256)
);

INVx2_ASAP7_75t_SL g1257 ( 
.A(n_1110),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1136),
.Y(n_1258)
);

AOI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1224),
.A2(n_1033),
.B(n_1045),
.Y(n_1259)
);

AOI22xp5_ASAP7_75t_L g1260 ( 
.A1(n_1177),
.A2(n_1046),
.B1(n_1050),
.B2(n_1076),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1105),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1129),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1241),
.A2(n_1023),
.B(n_1026),
.Y(n_1263)
);

OA21x2_ASAP7_75t_L g1264 ( 
.A1(n_1232),
.A2(n_1062),
.B(n_1067),
.Y(n_1264)
);

OAI22xp5_ASAP7_75t_L g1265 ( 
.A1(n_1102),
.A2(n_1028),
.B1(n_1069),
.B2(n_1098),
.Y(n_1265)
);

INVx2_ASAP7_75t_SL g1266 ( 
.A(n_1119),
.Y(n_1266)
);

A2O1A1Ixp33_ASAP7_75t_L g1267 ( 
.A1(n_1093),
.A2(n_1166),
.B(n_1125),
.C(n_1239),
.Y(n_1267)
);

INVx3_ASAP7_75t_L g1268 ( 
.A(n_1169),
.Y(n_1268)
);

INVx1_ASAP7_75t_SL g1269 ( 
.A(n_1099),
.Y(n_1269)
);

INVx3_ASAP7_75t_L g1270 ( 
.A(n_1169),
.Y(n_1270)
);

BUFx10_ASAP7_75t_L g1271 ( 
.A(n_1143),
.Y(n_1271)
);

AND2x2_ASAP7_75t_L g1272 ( 
.A(n_1160),
.B(n_1175),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1134),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1222),
.A2(n_1240),
.B(n_1246),
.Y(n_1274)
);

NOR2xp33_ASAP7_75t_L g1275 ( 
.A(n_1159),
.B(n_1117),
.Y(n_1275)
);

NOR2xp33_ASAP7_75t_L g1276 ( 
.A(n_1173),
.B(n_1161),
.Y(n_1276)
);

A2O1A1Ixp33_ASAP7_75t_L g1277 ( 
.A1(n_1149),
.A2(n_1216),
.B(n_1094),
.C(n_1154),
.Y(n_1277)
);

AOI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1240),
.A2(n_1243),
.B(n_1248),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1163),
.B(n_1170),
.Y(n_1279)
);

AOI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1243),
.A2(n_1201),
.B(n_1106),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1104),
.Y(n_1281)
);

OAI21x1_ASAP7_75t_L g1282 ( 
.A1(n_1230),
.A2(n_1116),
.B(n_1181),
.Y(n_1282)
);

BUFx10_ASAP7_75t_L g1283 ( 
.A(n_1164),
.Y(n_1283)
);

BUFx10_ASAP7_75t_L g1284 ( 
.A(n_1133),
.Y(n_1284)
);

AO21x1_ASAP7_75t_L g1285 ( 
.A1(n_1211),
.A2(n_1178),
.B(n_1242),
.Y(n_1285)
);

AOI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1201),
.A2(n_1106),
.B(n_1247),
.Y(n_1286)
);

O2A1O1Ixp33_ASAP7_75t_L g1287 ( 
.A1(n_1189),
.A2(n_1197),
.B(n_1209),
.C(n_1213),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1157),
.B(n_1193),
.Y(n_1288)
);

AOI22xp5_ASAP7_75t_L g1289 ( 
.A1(n_1191),
.A2(n_1189),
.B1(n_1128),
.B2(n_1186),
.Y(n_1289)
);

OAI22xp5_ASAP7_75t_L g1290 ( 
.A1(n_1183),
.A2(n_1217),
.B1(n_1214),
.B2(n_1215),
.Y(n_1290)
);

AOI22xp5_ASAP7_75t_L g1291 ( 
.A1(n_1191),
.A2(n_1128),
.B1(n_1220),
.B2(n_1152),
.Y(n_1291)
);

BUFx12f_ASAP7_75t_L g1292 ( 
.A(n_1132),
.Y(n_1292)
);

OAI21x1_ASAP7_75t_L g1293 ( 
.A1(n_1230),
.A2(n_1116),
.B(n_1242),
.Y(n_1293)
);

AOI22x1_ASAP7_75t_L g1294 ( 
.A1(n_1150),
.A2(n_1211),
.B1(n_1228),
.B2(n_1208),
.Y(n_1294)
);

AO22x2_ASAP7_75t_L g1295 ( 
.A1(n_1139),
.A2(n_1165),
.B1(n_1205),
.B2(n_1176),
.Y(n_1295)
);

NAND3xp33_ASAP7_75t_L g1296 ( 
.A(n_1202),
.B(n_1165),
.C(n_1149),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1112),
.Y(n_1297)
);

AOI31xp67_ASAP7_75t_L g1298 ( 
.A1(n_1252),
.A2(n_1200),
.A3(n_1238),
.B(n_1188),
.Y(n_1298)
);

BUFx12f_ASAP7_75t_L g1299 ( 
.A(n_1219),
.Y(n_1299)
);

OAI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1225),
.A2(n_1251),
.B(n_1107),
.Y(n_1300)
);

OAI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1251),
.A2(n_1107),
.B(n_1103),
.Y(n_1301)
);

O2A1O1Ixp33_ASAP7_75t_L g1302 ( 
.A1(n_1212),
.A2(n_1109),
.B(n_1179),
.C(n_1123),
.Y(n_1302)
);

O2A1O1Ixp33_ASAP7_75t_SL g1303 ( 
.A1(n_1096),
.A2(n_1100),
.B(n_1229),
.C(n_1182),
.Y(n_1303)
);

BUFx2_ASAP7_75t_L g1304 ( 
.A(n_1235),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1127),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1135),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1118),
.Y(n_1307)
);

AOI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1250),
.A2(n_1101),
.B(n_1169),
.Y(n_1308)
);

OR2x2_ASAP7_75t_L g1309 ( 
.A(n_1095),
.B(n_1171),
.Y(n_1309)
);

OAI22xp5_ASAP7_75t_L g1310 ( 
.A1(n_1226),
.A2(n_1194),
.B1(n_1231),
.B2(n_1172),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1174),
.B(n_1144),
.Y(n_1311)
);

AOI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1101),
.A2(n_1169),
.B(n_1245),
.Y(n_1312)
);

NAND2x1p5_ASAP7_75t_L g1313 ( 
.A(n_1236),
.B(n_1130),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_1140),
.Y(n_1314)
);

A2O1A1Ixp33_ASAP7_75t_L g1315 ( 
.A1(n_1148),
.A2(n_1150),
.B(n_1162),
.C(n_1153),
.Y(n_1315)
);

OAI22xp5_ASAP7_75t_SL g1316 ( 
.A1(n_1180),
.A2(n_1196),
.B1(n_1167),
.B2(n_1198),
.Y(n_1316)
);

O2A1O1Ixp33_ASAP7_75t_L g1317 ( 
.A1(n_1179),
.A2(n_1147),
.B(n_1162),
.C(n_1141),
.Y(n_1317)
);

INVx3_ASAP7_75t_L g1318 ( 
.A(n_1130),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1122),
.Y(n_1319)
);

NOR2xp33_ASAP7_75t_L g1320 ( 
.A(n_1142),
.B(n_1190),
.Y(n_1320)
);

AOI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1249),
.A2(n_1233),
.B(n_1113),
.Y(n_1321)
);

AOI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1253),
.A2(n_1236),
.B(n_1126),
.Y(n_1322)
);

AO31x2_ASAP7_75t_L g1323 ( 
.A1(n_1145),
.A2(n_1208),
.A3(n_1192),
.B(n_1199),
.Y(n_1323)
);

OAI22xp5_ASAP7_75t_L g1324 ( 
.A1(n_1180),
.A2(n_1126),
.B1(n_1203),
.B2(n_1195),
.Y(n_1324)
);

OA21x2_ASAP7_75t_L g1325 ( 
.A1(n_1237),
.A2(n_1192),
.B(n_1199),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1120),
.Y(n_1326)
);

AOI21xp33_ASAP7_75t_L g1327 ( 
.A1(n_1148),
.A2(n_1111),
.B(n_1108),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1120),
.Y(n_1328)
);

AO31x2_ASAP7_75t_L g1329 ( 
.A1(n_1114),
.A2(n_1155),
.A3(n_1156),
.B(n_1205),
.Y(n_1329)
);

A2O1A1Ixp33_ASAP7_75t_L g1330 ( 
.A1(n_1138),
.A2(n_1204),
.B(n_1185),
.C(n_1137),
.Y(n_1330)
);

OA21x2_ASAP7_75t_L g1331 ( 
.A1(n_1184),
.A2(n_1158),
.B(n_1206),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1244),
.Y(n_1332)
);

A2O1A1Ixp33_ASAP7_75t_L g1333 ( 
.A1(n_1138),
.A2(n_1131),
.B(n_1137),
.C(n_1185),
.Y(n_1333)
);

OR2x2_ASAP7_75t_L g1334 ( 
.A(n_1168),
.B(n_1151),
.Y(n_1334)
);

OAI21xp5_ASAP7_75t_L g1335 ( 
.A1(n_1187),
.A2(n_1126),
.B(n_1131),
.Y(n_1335)
);

BUFx2_ASAP7_75t_L g1336 ( 
.A(n_1234),
.Y(n_1336)
);

AOI21x1_ASAP7_75t_L g1337 ( 
.A1(n_1254),
.A2(n_1207),
.B(n_1180),
.Y(n_1337)
);

AOI31xp67_ASAP7_75t_L g1338 ( 
.A1(n_1205),
.A2(n_1139),
.A3(n_1223),
.B(n_1121),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1223),
.B(n_1124),
.Y(n_1339)
);

BUFx2_ASAP7_75t_R g1340 ( 
.A(n_1121),
.Y(n_1340)
);

O2A1O1Ixp33_ASAP7_75t_SL g1341 ( 
.A1(n_1139),
.A2(n_1146),
.B(n_1210),
.C(n_1221),
.Y(n_1341)
);

INVx6_ASAP7_75t_L g1342 ( 
.A(n_1146),
.Y(n_1342)
);

BUFx3_ASAP7_75t_L g1343 ( 
.A(n_1221),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1163),
.B(n_730),
.Y(n_1344)
);

OAI21xp5_ASAP7_75t_L g1345 ( 
.A1(n_1102),
.A2(n_730),
.B(n_1246),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1163),
.B(n_730),
.Y(n_1346)
);

AO32x2_ASAP7_75t_L g1347 ( 
.A1(n_1141),
.A2(n_955),
.A3(n_1139),
.B1(n_1123),
.B2(n_852),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1163),
.B(n_730),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1177),
.A2(n_730),
.B1(n_958),
.B2(n_980),
.Y(n_1349)
);

AO32x2_ASAP7_75t_L g1350 ( 
.A1(n_1141),
.A2(n_955),
.A3(n_1139),
.B1(n_1123),
.B2(n_852),
.Y(n_1350)
);

A2O1A1Ixp33_ASAP7_75t_L g1351 ( 
.A1(n_1102),
.A2(n_730),
.B(n_958),
.C(n_906),
.Y(n_1351)
);

OAI21x1_ASAP7_75t_L g1352 ( 
.A1(n_1227),
.A2(n_1230),
.B(n_963),
.Y(n_1352)
);

AOI21x1_ASAP7_75t_L g1353 ( 
.A1(n_1227),
.A2(n_1243),
.B(n_1240),
.Y(n_1353)
);

O2A1O1Ixp33_ASAP7_75t_L g1354 ( 
.A1(n_1177),
.A2(n_730),
.B(n_958),
.C(n_906),
.Y(n_1354)
);

NOR2xp33_ASAP7_75t_L g1355 ( 
.A(n_1159),
.B(n_730),
.Y(n_1355)
);

OAI22x1_ASAP7_75t_L g1356 ( 
.A1(n_1177),
.A2(n_730),
.B1(n_593),
.B2(n_1125),
.Y(n_1356)
);

OA21x2_ASAP7_75t_L g1357 ( 
.A1(n_1232),
.A2(n_1224),
.B(n_1243),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1136),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1163),
.B(n_730),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1163),
.B(n_730),
.Y(n_1360)
);

AO31x2_ASAP7_75t_L g1361 ( 
.A1(n_1145),
.A2(n_1102),
.A3(n_1065),
.B(n_1224),
.Y(n_1361)
);

O2A1O1Ixp33_ASAP7_75t_SL g1362 ( 
.A1(n_1102),
.A2(n_958),
.B(n_730),
.C(n_1197),
.Y(n_1362)
);

OR2x2_ASAP7_75t_L g1363 ( 
.A(n_1157),
.B(n_666),
.Y(n_1363)
);

OAI21x1_ASAP7_75t_L g1364 ( 
.A1(n_1227),
.A2(n_1230),
.B(n_963),
.Y(n_1364)
);

INVxp67_ASAP7_75t_SL g1365 ( 
.A(n_1095),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_SL g1366 ( 
.A(n_1140),
.B(n_730),
.Y(n_1366)
);

OAI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1227),
.A2(n_1230),
.B(n_963),
.Y(n_1367)
);

AOI22xp5_ASAP7_75t_L g1368 ( 
.A1(n_1177),
.A2(n_730),
.B1(n_958),
.B2(n_980),
.Y(n_1368)
);

AOI21xp5_ASAP7_75t_L g1369 ( 
.A1(n_1218),
.A2(n_730),
.B(n_958),
.Y(n_1369)
);

A2O1A1Ixp33_ASAP7_75t_L g1370 ( 
.A1(n_1102),
.A2(n_730),
.B(n_958),
.C(n_906),
.Y(n_1370)
);

AOI21xp5_ASAP7_75t_L g1371 ( 
.A1(n_1218),
.A2(n_730),
.B(n_958),
.Y(n_1371)
);

AOI21xp5_ASAP7_75t_L g1372 ( 
.A1(n_1218),
.A2(n_730),
.B(n_958),
.Y(n_1372)
);

AO31x2_ASAP7_75t_L g1373 ( 
.A1(n_1145),
.A2(n_1102),
.A3(n_1065),
.B(n_1224),
.Y(n_1373)
);

A2O1A1Ixp33_ASAP7_75t_L g1374 ( 
.A1(n_1102),
.A2(n_730),
.B(n_958),
.C(n_906),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1163),
.B(n_730),
.Y(n_1375)
);

NOR2xp33_ASAP7_75t_SL g1376 ( 
.A(n_1193),
.B(n_730),
.Y(n_1376)
);

AO31x2_ASAP7_75t_L g1377 ( 
.A1(n_1145),
.A2(n_1102),
.A3(n_1065),
.B(n_1224),
.Y(n_1377)
);

AOI21xp5_ASAP7_75t_L g1378 ( 
.A1(n_1218),
.A2(n_730),
.B(n_958),
.Y(n_1378)
);

BUFx6f_ASAP7_75t_L g1379 ( 
.A(n_1219),
.Y(n_1379)
);

A2O1A1Ixp33_ASAP7_75t_L g1380 ( 
.A1(n_1102),
.A2(n_730),
.B(n_958),
.C(n_906),
.Y(n_1380)
);

A2O1A1Ixp33_ASAP7_75t_L g1381 ( 
.A1(n_1102),
.A2(n_730),
.B(n_958),
.C(n_906),
.Y(n_1381)
);

OAI21x1_ASAP7_75t_L g1382 ( 
.A1(n_1227),
.A2(n_1230),
.B(n_963),
.Y(n_1382)
);

BUFx6f_ASAP7_75t_L g1383 ( 
.A(n_1219),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1160),
.B(n_901),
.Y(n_1384)
);

OAI21x1_ASAP7_75t_L g1385 ( 
.A1(n_1227),
.A2(n_1230),
.B(n_963),
.Y(n_1385)
);

NAND2x1p5_ASAP7_75t_L g1386 ( 
.A(n_1169),
.B(n_1236),
.Y(n_1386)
);

NOR2xp33_ASAP7_75t_L g1387 ( 
.A(n_1159),
.B(n_730),
.Y(n_1387)
);

OAI22xp33_ASAP7_75t_L g1388 ( 
.A1(n_1177),
.A2(n_730),
.B1(n_1000),
.B2(n_958),
.Y(n_1388)
);

BUFx3_ASAP7_75t_L g1389 ( 
.A(n_1110),
.Y(n_1389)
);

INVx3_ASAP7_75t_L g1390 ( 
.A(n_1169),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1136),
.Y(n_1391)
);

NOR4xp25_ASAP7_75t_L g1392 ( 
.A(n_1189),
.B(n_1179),
.C(n_1197),
.D(n_1102),
.Y(n_1392)
);

AOI31xp67_ASAP7_75t_L g1393 ( 
.A1(n_1228),
.A2(n_1218),
.A3(n_1252),
.B(n_732),
.Y(n_1393)
);

BUFx2_ASAP7_75t_L g1394 ( 
.A(n_1117),
.Y(n_1394)
);

BUFx6f_ASAP7_75t_L g1395 ( 
.A(n_1219),
.Y(n_1395)
);

OAI22x1_ASAP7_75t_L g1396 ( 
.A1(n_1177),
.A2(n_730),
.B1(n_593),
.B2(n_1125),
.Y(n_1396)
);

CKINVDCx20_ASAP7_75t_R g1397 ( 
.A(n_1140),
.Y(n_1397)
);

NAND3xp33_ASAP7_75t_L g1398 ( 
.A(n_1177),
.B(n_730),
.C(n_958),
.Y(n_1398)
);

AOI221x1_ASAP7_75t_L g1399 ( 
.A1(n_1102),
.A2(n_730),
.B1(n_1177),
.B2(n_958),
.C(n_1189),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1163),
.B(n_730),
.Y(n_1400)
);

AOI21xp5_ASAP7_75t_L g1401 ( 
.A1(n_1218),
.A2(n_730),
.B(n_958),
.Y(n_1401)
);

INVx2_ASAP7_75t_L g1402 ( 
.A(n_1115),
.Y(n_1402)
);

CKINVDCx5p33_ASAP7_75t_R g1403 ( 
.A(n_1097),
.Y(n_1403)
);

OAI21x1_ASAP7_75t_SL g1404 ( 
.A1(n_1211),
.A2(n_982),
.B(n_996),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_L g1405 ( 
.A1(n_1227),
.A2(n_1230),
.B(n_963),
.Y(n_1405)
);

CKINVDCx5p33_ASAP7_75t_R g1406 ( 
.A(n_1097),
.Y(n_1406)
);

OA21x2_ASAP7_75t_L g1407 ( 
.A1(n_1232),
.A2(n_1224),
.B(n_1243),
.Y(n_1407)
);

BUFx10_ASAP7_75t_L g1408 ( 
.A(n_1177),
.Y(n_1408)
);

AO31x2_ASAP7_75t_L g1409 ( 
.A1(n_1145),
.A2(n_1102),
.A3(n_1065),
.B(n_1224),
.Y(n_1409)
);

OAI22xp33_ASAP7_75t_L g1410 ( 
.A1(n_1177),
.A2(n_730),
.B1(n_1000),
.B2(n_958),
.Y(n_1410)
);

O2A1O1Ixp5_ASAP7_75t_SL g1411 ( 
.A1(n_1178),
.A2(n_958),
.B(n_703),
.C(n_900),
.Y(n_1411)
);

OR2x2_ASAP7_75t_L g1412 ( 
.A(n_1157),
.B(n_666),
.Y(n_1412)
);

AOI22xp33_ASAP7_75t_L g1413 ( 
.A1(n_1349),
.A2(n_1398),
.B1(n_1396),
.B2(n_1356),
.Y(n_1413)
);

BUFx4f_ASAP7_75t_SL g1414 ( 
.A(n_1397),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1258),
.Y(n_1415)
);

BUFx12f_ASAP7_75t_L g1416 ( 
.A(n_1314),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1358),
.Y(n_1417)
);

AOI22xp5_ASAP7_75t_L g1418 ( 
.A1(n_1376),
.A2(n_1368),
.B1(n_1388),
.B2(n_1410),
.Y(n_1418)
);

BUFx4f_ASAP7_75t_L g1419 ( 
.A(n_1379),
.Y(n_1419)
);

CKINVDCx20_ASAP7_75t_R g1420 ( 
.A(n_1403),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_SL g1421 ( 
.A1(n_1376),
.A2(n_1345),
.B1(n_1398),
.B2(n_1288),
.Y(n_1421)
);

AOI22xp33_ASAP7_75t_L g1422 ( 
.A1(n_1316),
.A2(n_1368),
.B1(n_1289),
.B2(n_1345),
.Y(n_1422)
);

INVx6_ASAP7_75t_L g1423 ( 
.A(n_1379),
.Y(n_1423)
);

BUFx2_ASAP7_75t_L g1424 ( 
.A(n_1272),
.Y(n_1424)
);

OAI22x1_ASAP7_75t_L g1425 ( 
.A1(n_1289),
.A2(n_1291),
.B1(n_1296),
.B2(n_1276),
.Y(n_1425)
);

OAI22xp33_ASAP7_75t_L g1426 ( 
.A1(n_1291),
.A2(n_1399),
.B1(n_1375),
.B2(n_1360),
.Y(n_1426)
);

AOI22xp33_ASAP7_75t_L g1427 ( 
.A1(n_1316),
.A2(n_1296),
.B1(n_1371),
.B2(n_1401),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_SL g1428 ( 
.A1(n_1310),
.A2(n_1408),
.B1(n_1290),
.B2(n_1295),
.Y(n_1428)
);

AOI22xp33_ASAP7_75t_L g1429 ( 
.A1(n_1369),
.A2(n_1378),
.B1(n_1372),
.B2(n_1290),
.Y(n_1429)
);

CKINVDCx6p67_ASAP7_75t_R g1430 ( 
.A(n_1292),
.Y(n_1430)
);

CKINVDCx6p67_ASAP7_75t_R g1431 ( 
.A(n_1299),
.Y(n_1431)
);

BUFx2_ASAP7_75t_L g1432 ( 
.A(n_1304),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1344),
.B(n_1346),
.Y(n_1433)
);

BUFx3_ASAP7_75t_L g1434 ( 
.A(n_1389),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1391),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1348),
.B(n_1359),
.Y(n_1436)
);

OAI22xp5_ASAP7_75t_L g1437 ( 
.A1(n_1400),
.A2(n_1267),
.B1(n_1354),
.B2(n_1355),
.Y(n_1437)
);

AOI22xp33_ASAP7_75t_L g1438 ( 
.A1(n_1408),
.A2(n_1310),
.B1(n_1328),
.B2(n_1326),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1261),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1262),
.Y(n_1440)
);

OAI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1334),
.A2(n_1307),
.B1(n_1311),
.B2(n_1279),
.Y(n_1441)
);

AOI22xp33_ASAP7_75t_L g1442 ( 
.A1(n_1295),
.A2(n_1319),
.B1(n_1305),
.B2(n_1306),
.Y(n_1442)
);

BUFx12f_ASAP7_75t_L g1443 ( 
.A(n_1379),
.Y(n_1443)
);

AOI22xp5_ASAP7_75t_L g1444 ( 
.A1(n_1320),
.A2(n_1366),
.B1(n_1387),
.B2(n_1384),
.Y(n_1444)
);

INVx6_ASAP7_75t_L g1445 ( 
.A(n_1383),
.Y(n_1445)
);

INVxp67_ASAP7_75t_L g1446 ( 
.A(n_1365),
.Y(n_1446)
);

INVx4_ASAP7_75t_L g1447 ( 
.A(n_1386),
.Y(n_1447)
);

CKINVDCx11_ASAP7_75t_R g1448 ( 
.A(n_1271),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1273),
.Y(n_1449)
);

BUFx12f_ASAP7_75t_L g1450 ( 
.A(n_1383),
.Y(n_1450)
);

OAI21xp5_ASAP7_75t_SL g1451 ( 
.A1(n_1287),
.A2(n_1317),
.B(n_1381),
.Y(n_1451)
);

OR2x6_ASAP7_75t_L g1452 ( 
.A(n_1322),
.B(n_1337),
.Y(n_1452)
);

BUFx3_ASAP7_75t_L g1453 ( 
.A(n_1383),
.Y(n_1453)
);

OAI22xp5_ASAP7_75t_L g1454 ( 
.A1(n_1351),
.A2(n_1374),
.B1(n_1380),
.B2(n_1370),
.Y(n_1454)
);

INVx6_ASAP7_75t_L g1455 ( 
.A(n_1395),
.Y(n_1455)
);

HB1xp67_ASAP7_75t_L g1456 ( 
.A(n_1329),
.Y(n_1456)
);

AOI22xp33_ASAP7_75t_L g1457 ( 
.A1(n_1285),
.A2(n_1301),
.B1(n_1284),
.B2(n_1283),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1281),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1309),
.B(n_1275),
.Y(n_1459)
);

BUFx8_ASAP7_75t_L g1460 ( 
.A(n_1395),
.Y(n_1460)
);

BUFx12f_ASAP7_75t_L g1461 ( 
.A(n_1395),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1297),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1298),
.Y(n_1463)
);

OAI22xp33_ASAP7_75t_L g1464 ( 
.A1(n_1363),
.A2(n_1412),
.B1(n_1324),
.B2(n_1301),
.Y(n_1464)
);

OAI22xp5_ASAP7_75t_L g1465 ( 
.A1(n_1269),
.A2(n_1324),
.B1(n_1339),
.B2(n_1277),
.Y(n_1465)
);

INVx1_ASAP7_75t_SL g1466 ( 
.A(n_1269),
.Y(n_1466)
);

CKINVDCx20_ASAP7_75t_R g1467 ( 
.A(n_1406),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1332),
.Y(n_1468)
);

CKINVDCx11_ASAP7_75t_R g1469 ( 
.A(n_1271),
.Y(n_1469)
);

BUFx4f_ASAP7_75t_SL g1470 ( 
.A(n_1336),
.Y(n_1470)
);

INVx1_ASAP7_75t_SL g1471 ( 
.A(n_1340),
.Y(n_1471)
);

BUFx2_ASAP7_75t_L g1472 ( 
.A(n_1343),
.Y(n_1472)
);

OAI21xp5_ASAP7_75t_SL g1473 ( 
.A1(n_1302),
.A2(n_1315),
.B(n_1308),
.Y(n_1473)
);

BUFx3_ASAP7_75t_L g1474 ( 
.A(n_1257),
.Y(n_1474)
);

NAND2x1p5_ASAP7_75t_L g1475 ( 
.A(n_1270),
.B(n_1390),
.Y(n_1475)
);

AOI22xp5_ASAP7_75t_L g1476 ( 
.A1(n_1284),
.A2(n_1283),
.B1(n_1362),
.B2(n_1266),
.Y(n_1476)
);

AOI22xp33_ASAP7_75t_SL g1477 ( 
.A1(n_1300),
.A2(n_1294),
.B1(n_1392),
.B2(n_1404),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_SL g1478 ( 
.A1(n_1300),
.A2(n_1392),
.B1(n_1280),
.B2(n_1341),
.Y(n_1478)
);

OAI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1274),
.A2(n_1286),
.B1(n_1321),
.B2(n_1256),
.Y(n_1479)
);

OAI22xp33_ASAP7_75t_R g1480 ( 
.A1(n_1347),
.A2(n_1350),
.B1(n_1338),
.B2(n_1411),
.Y(n_1480)
);

OAI21xp5_ASAP7_75t_L g1481 ( 
.A1(n_1327),
.A2(n_1312),
.B(n_1265),
.Y(n_1481)
);

BUFx6f_ASAP7_75t_L g1482 ( 
.A(n_1342),
.Y(n_1482)
);

OAI22xp5_ASAP7_75t_L g1483 ( 
.A1(n_1330),
.A2(n_1313),
.B1(n_1335),
.B2(n_1333),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1329),
.Y(n_1484)
);

AOI22xp33_ASAP7_75t_L g1485 ( 
.A1(n_1278),
.A2(n_1325),
.B1(n_1357),
.B2(n_1407),
.Y(n_1485)
);

AOI22xp33_ASAP7_75t_L g1486 ( 
.A1(n_1325),
.A2(n_1407),
.B1(n_1357),
.B2(n_1265),
.Y(n_1486)
);

CKINVDCx20_ASAP7_75t_R g1487 ( 
.A(n_1342),
.Y(n_1487)
);

AOI22xp33_ASAP7_75t_L g1488 ( 
.A1(n_1293),
.A2(n_1335),
.B1(n_1350),
.B2(n_1347),
.Y(n_1488)
);

OAI22xp5_ASAP7_75t_SL g1489 ( 
.A1(n_1318),
.A2(n_1260),
.B1(n_1331),
.B2(n_1350),
.Y(n_1489)
);

AOI22xp33_ASAP7_75t_L g1490 ( 
.A1(n_1347),
.A2(n_1259),
.B1(n_1264),
.B2(n_1260),
.Y(n_1490)
);

AOI22xp5_ASAP7_75t_L g1491 ( 
.A1(n_1303),
.A2(n_1331),
.B1(n_1264),
.B2(n_1263),
.Y(n_1491)
);

INVx4_ASAP7_75t_L g1492 ( 
.A(n_1329),
.Y(n_1492)
);

AOI22xp33_ASAP7_75t_SL g1493 ( 
.A1(n_1282),
.A2(n_1405),
.B1(n_1385),
.B2(n_1352),
.Y(n_1493)
);

AOI22xp5_ASAP7_75t_L g1494 ( 
.A1(n_1255),
.A2(n_1382),
.B1(n_1367),
.B2(n_1364),
.Y(n_1494)
);

BUFx6f_ASAP7_75t_SL g1495 ( 
.A(n_1393),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1361),
.B(n_1409),
.Y(n_1496)
);

OAI22x1_ASAP7_75t_L g1497 ( 
.A1(n_1353),
.A2(n_1361),
.B1(n_1373),
.B2(n_1377),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1361),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1373),
.Y(n_1499)
);

INVx1_ASAP7_75t_SL g1500 ( 
.A(n_1377),
.Y(n_1500)
);

INVx4_ASAP7_75t_L g1501 ( 
.A(n_1377),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1409),
.Y(n_1502)
);

BUFx6f_ASAP7_75t_L g1503 ( 
.A(n_1323),
.Y(n_1503)
);

AOI22xp33_ASAP7_75t_L g1504 ( 
.A1(n_1323),
.A2(n_730),
.B1(n_1177),
.B2(n_1356),
.Y(n_1504)
);

AOI22xp33_ASAP7_75t_L g1505 ( 
.A1(n_1349),
.A2(n_730),
.B1(n_1191),
.B2(n_1398),
.Y(n_1505)
);

CKINVDCx20_ASAP7_75t_R g1506 ( 
.A(n_1397),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1402),
.Y(n_1507)
);

OAI22xp5_ASAP7_75t_L g1508 ( 
.A1(n_1368),
.A2(n_730),
.B1(n_1349),
.B2(n_1398),
.Y(n_1508)
);

AOI22xp33_ASAP7_75t_L g1509 ( 
.A1(n_1349),
.A2(n_730),
.B1(n_1191),
.B2(n_1398),
.Y(n_1509)
);

BUFx2_ASAP7_75t_SL g1510 ( 
.A(n_1397),
.Y(n_1510)
);

BUFx2_ASAP7_75t_SL g1511 ( 
.A(n_1397),
.Y(n_1511)
);

INVx5_ASAP7_75t_L g1512 ( 
.A(n_1268),
.Y(n_1512)
);

AOI22xp33_ASAP7_75t_SL g1513 ( 
.A1(n_1376),
.A2(n_730),
.B1(n_1000),
.B2(n_1191),
.Y(n_1513)
);

AOI22xp33_ASAP7_75t_L g1514 ( 
.A1(n_1349),
.A2(n_730),
.B1(n_1191),
.B2(n_1398),
.Y(n_1514)
);

CKINVDCx5p33_ASAP7_75t_R g1515 ( 
.A(n_1403),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1258),
.Y(n_1516)
);

AOI22xp33_ASAP7_75t_L g1517 ( 
.A1(n_1349),
.A2(n_730),
.B1(n_1191),
.B2(n_1398),
.Y(n_1517)
);

OAI22xp5_ASAP7_75t_L g1518 ( 
.A1(n_1368),
.A2(n_730),
.B1(n_1349),
.B2(n_1398),
.Y(n_1518)
);

BUFx6f_ASAP7_75t_L g1519 ( 
.A(n_1386),
.Y(n_1519)
);

BUFx2_ASAP7_75t_SL g1520 ( 
.A(n_1397),
.Y(n_1520)
);

AOI22xp33_ASAP7_75t_L g1521 ( 
.A1(n_1349),
.A2(n_730),
.B1(n_1191),
.B2(n_1398),
.Y(n_1521)
);

OAI21xp5_ASAP7_75t_SL g1522 ( 
.A1(n_1368),
.A2(n_730),
.B(n_593),
.Y(n_1522)
);

BUFx3_ASAP7_75t_L g1523 ( 
.A(n_1389),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1344),
.B(n_730),
.Y(n_1524)
);

BUFx6f_ASAP7_75t_L g1525 ( 
.A(n_1386),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1258),
.Y(n_1526)
);

CKINVDCx20_ASAP7_75t_R g1527 ( 
.A(n_1397),
.Y(n_1527)
);

AOI22xp33_ASAP7_75t_L g1528 ( 
.A1(n_1349),
.A2(n_730),
.B1(n_1191),
.B2(n_1398),
.Y(n_1528)
);

OAI22xp5_ASAP7_75t_L g1529 ( 
.A1(n_1368),
.A2(n_730),
.B1(n_1349),
.B2(n_1398),
.Y(n_1529)
);

BUFx3_ASAP7_75t_L g1530 ( 
.A(n_1389),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1344),
.B(n_730),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1258),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1258),
.Y(n_1533)
);

INVxp67_ASAP7_75t_L g1534 ( 
.A(n_1394),
.Y(n_1534)
);

OAI22xp33_ASAP7_75t_L g1535 ( 
.A1(n_1368),
.A2(n_1376),
.B1(n_1289),
.B2(n_730),
.Y(n_1535)
);

OAI22xp5_ASAP7_75t_L g1536 ( 
.A1(n_1368),
.A2(n_730),
.B1(n_1349),
.B2(n_1398),
.Y(n_1536)
);

BUFx10_ASAP7_75t_L g1537 ( 
.A(n_1379),
.Y(n_1537)
);

BUFx2_ASAP7_75t_SL g1538 ( 
.A(n_1397),
.Y(n_1538)
);

CKINVDCx5p33_ASAP7_75t_R g1539 ( 
.A(n_1403),
.Y(n_1539)
);

AOI22xp33_ASAP7_75t_SL g1540 ( 
.A1(n_1376),
.A2(n_730),
.B1(n_1000),
.B2(n_1191),
.Y(n_1540)
);

AOI22xp33_ASAP7_75t_SL g1541 ( 
.A1(n_1376),
.A2(n_730),
.B1(n_1000),
.B2(n_1191),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1258),
.Y(n_1542)
);

AOI22xp33_ASAP7_75t_L g1543 ( 
.A1(n_1349),
.A2(n_730),
.B1(n_1191),
.B2(n_1398),
.Y(n_1543)
);

AOI22xp33_ASAP7_75t_SL g1544 ( 
.A1(n_1376),
.A2(n_730),
.B1(n_1000),
.B2(n_1191),
.Y(n_1544)
);

INVx1_ASAP7_75t_SL g1545 ( 
.A(n_1269),
.Y(n_1545)
);

AOI22xp33_ASAP7_75t_L g1546 ( 
.A1(n_1349),
.A2(n_730),
.B1(n_1191),
.B2(n_1398),
.Y(n_1546)
);

AOI22xp33_ASAP7_75t_SL g1547 ( 
.A1(n_1376),
.A2(n_730),
.B1(n_1000),
.B2(n_1191),
.Y(n_1547)
);

OAI22xp33_ASAP7_75t_L g1548 ( 
.A1(n_1368),
.A2(n_1376),
.B1(n_1289),
.B2(n_730),
.Y(n_1548)
);

OAI22xp33_ASAP7_75t_L g1549 ( 
.A1(n_1368),
.A2(n_1376),
.B1(n_1289),
.B2(n_730),
.Y(n_1549)
);

INVx6_ASAP7_75t_L g1550 ( 
.A(n_1379),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1384),
.B(n_1288),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1258),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1437),
.B(n_1524),
.Y(n_1553)
);

AO21x2_ASAP7_75t_L g1554 ( 
.A1(n_1481),
.A2(n_1479),
.B(n_1491),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1531),
.B(n_1433),
.Y(n_1555)
);

AO21x2_ASAP7_75t_L g1556 ( 
.A1(n_1479),
.A2(n_1473),
.B(n_1494),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1415),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1442),
.B(n_1428),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1484),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1436),
.B(n_1459),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1498),
.Y(n_1561)
);

OAI21xp5_ASAP7_75t_L g1562 ( 
.A1(n_1508),
.A2(n_1529),
.B(n_1518),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1499),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1502),
.Y(n_1564)
);

BUFx2_ASAP7_75t_L g1565 ( 
.A(n_1452),
.Y(n_1565)
);

OA21x2_ASAP7_75t_L g1566 ( 
.A1(n_1488),
.A2(n_1490),
.B(n_1486),
.Y(n_1566)
);

AOI221xp5_ASAP7_75t_L g1567 ( 
.A1(n_1522),
.A2(n_1536),
.B1(n_1549),
.B2(n_1548),
.C(n_1535),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1456),
.Y(n_1568)
);

NOR2x1_ASAP7_75t_R g1569 ( 
.A(n_1448),
.B(n_1469),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1442),
.B(n_1428),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1425),
.B(n_1496),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1456),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1478),
.B(n_1422),
.Y(n_1573)
);

BUFx2_ASAP7_75t_L g1574 ( 
.A(n_1452),
.Y(n_1574)
);

AO21x2_ASAP7_75t_L g1575 ( 
.A1(n_1463),
.A2(n_1451),
.B(n_1454),
.Y(n_1575)
);

OA21x2_ASAP7_75t_L g1576 ( 
.A1(n_1488),
.A2(n_1490),
.B(n_1486),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1503),
.Y(n_1577)
);

BUFx3_ASAP7_75t_L g1578 ( 
.A(n_1452),
.Y(n_1578)
);

OR2x6_ASAP7_75t_L g1579 ( 
.A(n_1489),
.B(n_1483),
.Y(n_1579)
);

OR2x2_ASAP7_75t_L g1580 ( 
.A(n_1500),
.B(n_1492),
.Y(n_1580)
);

AOI21xp5_ASAP7_75t_L g1581 ( 
.A1(n_1427),
.A2(n_1429),
.B(n_1535),
.Y(n_1581)
);

OR2x2_ASAP7_75t_L g1582 ( 
.A(n_1492),
.B(n_1501),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1478),
.B(n_1413),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1480),
.Y(n_1584)
);

BUFx2_ASAP7_75t_L g1585 ( 
.A(n_1446),
.Y(n_1585)
);

OAI21x1_ASAP7_75t_L g1586 ( 
.A1(n_1485),
.A2(n_1429),
.B(n_1427),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1426),
.B(n_1505),
.Y(n_1587)
);

AOI21x1_ASAP7_75t_L g1588 ( 
.A1(n_1497),
.A2(n_1465),
.B(n_1435),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_1417),
.Y(n_1589)
);

HB1xp67_ASAP7_75t_SL g1590 ( 
.A(n_1460),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1413),
.B(n_1421),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1495),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1495),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1426),
.B(n_1505),
.Y(n_1594)
);

AO21x1_ASAP7_75t_L g1595 ( 
.A1(n_1548),
.A2(n_1549),
.B(n_1441),
.Y(n_1595)
);

INVx1_ASAP7_75t_SL g1596 ( 
.A(n_1466),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_1439),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1421),
.B(n_1477),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1477),
.B(n_1504),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1440),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1516),
.Y(n_1601)
);

OR2x2_ASAP7_75t_L g1602 ( 
.A(n_1464),
.B(n_1441),
.Y(n_1602)
);

HB1xp67_ASAP7_75t_L g1603 ( 
.A(n_1534),
.Y(n_1603)
);

HB1xp67_ASAP7_75t_L g1604 ( 
.A(n_1534),
.Y(n_1604)
);

AOI22xp5_ASAP7_75t_L g1605 ( 
.A1(n_1513),
.A2(n_1540),
.B1(n_1544),
.B2(n_1541),
.Y(n_1605)
);

BUFx3_ASAP7_75t_L g1606 ( 
.A(n_1432),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1526),
.Y(n_1607)
);

NOR2xp33_ASAP7_75t_L g1608 ( 
.A(n_1551),
.B(n_1444),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1532),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1533),
.Y(n_1610)
);

AOI22xp33_ASAP7_75t_L g1611 ( 
.A1(n_1513),
.A2(n_1540),
.B1(n_1544),
.B2(n_1541),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1542),
.Y(n_1612)
);

OR2x2_ASAP7_75t_L g1613 ( 
.A(n_1464),
.B(n_1438),
.Y(n_1613)
);

INVx3_ASAP7_75t_L g1614 ( 
.A(n_1512),
.Y(n_1614)
);

NAND2x1p5_ASAP7_75t_L g1615 ( 
.A(n_1512),
.B(n_1418),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1509),
.B(n_1514),
.Y(n_1616)
);

INVx3_ASAP7_75t_L g1617 ( 
.A(n_1512),
.Y(n_1617)
);

AOI21xp5_ASAP7_75t_L g1618 ( 
.A1(n_1485),
.A2(n_1493),
.B(n_1509),
.Y(n_1618)
);

BUFx6f_ASAP7_75t_L g1619 ( 
.A(n_1512),
.Y(n_1619)
);

HB1xp67_ASAP7_75t_L g1620 ( 
.A(n_1545),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1514),
.B(n_1517),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1457),
.B(n_1552),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1457),
.B(n_1458),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1547),
.B(n_1438),
.Y(n_1624)
);

BUFx3_ASAP7_75t_L g1625 ( 
.A(n_1475),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1449),
.Y(n_1626)
);

HB1xp67_ASAP7_75t_L g1627 ( 
.A(n_1424),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1462),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1493),
.Y(n_1629)
);

OAI22xp33_ASAP7_75t_L g1630 ( 
.A1(n_1476),
.A2(n_1470),
.B1(n_1414),
.B2(n_1471),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1547),
.B(n_1507),
.Y(n_1631)
);

BUFx2_ASAP7_75t_L g1632 ( 
.A(n_1468),
.Y(n_1632)
);

BUFx2_ASAP7_75t_L g1633 ( 
.A(n_1472),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1521),
.Y(n_1634)
);

OAI21x1_ASAP7_75t_L g1635 ( 
.A1(n_1521),
.A2(n_1528),
.B(n_1546),
.Y(n_1635)
);

OAI21xp5_ASAP7_75t_L g1636 ( 
.A1(n_1528),
.A2(n_1543),
.B(n_1546),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1543),
.B(n_1511),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1510),
.B(n_1538),
.Y(n_1638)
);

AO21x2_ASAP7_75t_L g1639 ( 
.A1(n_1519),
.A2(n_1525),
.B(n_1447),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1520),
.B(n_1525),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1482),
.Y(n_1641)
);

AOI322xp5_ASAP7_75t_L g1642 ( 
.A1(n_1506),
.A2(n_1527),
.A3(n_1443),
.B1(n_1461),
.B2(n_1450),
.C1(n_1453),
.C2(n_1487),
.Y(n_1642)
);

OAI21x1_ASAP7_75t_L g1643 ( 
.A1(n_1423),
.A2(n_1550),
.B(n_1455),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1474),
.Y(n_1644)
);

AOI21x1_ASAP7_75t_L g1645 ( 
.A1(n_1470),
.A2(n_1455),
.B(n_1550),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1423),
.Y(n_1646)
);

AO31x2_ASAP7_75t_L g1647 ( 
.A1(n_1423),
.A2(n_1455),
.A3(n_1550),
.B(n_1445),
.Y(n_1647)
);

AOI211xp5_ASAP7_75t_L g1648 ( 
.A1(n_1434),
.A2(n_1530),
.B(n_1523),
.C(n_1539),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1445),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1537),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1537),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1419),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1419),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1460),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1414),
.B(n_1515),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1416),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1431),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1430),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1420),
.Y(n_1659)
);

INVx2_ASAP7_75t_SL g1660 ( 
.A(n_1467),
.Y(n_1660)
);

BUFx3_ASAP7_75t_L g1661 ( 
.A(n_1452),
.Y(n_1661)
);

OAI21xp5_ASAP7_75t_L g1662 ( 
.A1(n_1562),
.A2(n_1581),
.B(n_1567),
.Y(n_1662)
);

AO21x1_ASAP7_75t_L g1663 ( 
.A1(n_1605),
.A2(n_1553),
.B(n_1636),
.Y(n_1663)
);

AND2x4_ASAP7_75t_L g1664 ( 
.A(n_1578),
.B(n_1661),
.Y(n_1664)
);

OAI21xp5_ASAP7_75t_L g1665 ( 
.A1(n_1605),
.A2(n_1635),
.B(n_1594),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1637),
.B(n_1571),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1597),
.B(n_1601),
.Y(n_1667)
);

NOR2xp33_ASAP7_75t_L g1668 ( 
.A(n_1555),
.B(n_1560),
.Y(n_1668)
);

OAI21xp5_ASAP7_75t_L g1669 ( 
.A1(n_1635),
.A2(n_1587),
.B(n_1611),
.Y(n_1669)
);

A2O1A1Ixp33_ASAP7_75t_L g1670 ( 
.A1(n_1573),
.A2(n_1602),
.B(n_1598),
.C(n_1624),
.Y(n_1670)
);

A2O1A1Ixp33_ASAP7_75t_L g1671 ( 
.A1(n_1573),
.A2(n_1602),
.B(n_1598),
.C(n_1624),
.Y(n_1671)
);

OAI211xp5_ASAP7_75t_L g1672 ( 
.A1(n_1583),
.A2(n_1616),
.B(n_1621),
.C(n_1591),
.Y(n_1672)
);

AND2x4_ASAP7_75t_L g1673 ( 
.A(n_1578),
.B(n_1661),
.Y(n_1673)
);

AOI21xp5_ASAP7_75t_L g1674 ( 
.A1(n_1595),
.A2(n_1554),
.B(n_1556),
.Y(n_1674)
);

A2O1A1Ixp33_ASAP7_75t_L g1675 ( 
.A1(n_1613),
.A2(n_1591),
.B(n_1583),
.C(n_1599),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1607),
.B(n_1612),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1566),
.B(n_1576),
.Y(n_1677)
);

BUFx3_ASAP7_75t_L g1678 ( 
.A(n_1647),
.Y(n_1678)
);

OR2x2_ASAP7_75t_L g1679 ( 
.A(n_1632),
.B(n_1627),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1566),
.B(n_1576),
.Y(n_1680)
);

AO32x2_ASAP7_75t_L g1681 ( 
.A1(n_1584),
.A2(n_1595),
.A3(n_1572),
.B1(n_1568),
.B2(n_1566),
.Y(n_1681)
);

OR2x2_ASAP7_75t_L g1682 ( 
.A(n_1585),
.B(n_1557),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1576),
.B(n_1631),
.Y(n_1683)
);

CKINVDCx5p33_ASAP7_75t_R g1684 ( 
.A(n_1590),
.Y(n_1684)
);

BUFx2_ASAP7_75t_L g1685 ( 
.A(n_1633),
.Y(n_1685)
);

NOR2x1_ASAP7_75t_L g1686 ( 
.A(n_1639),
.B(n_1630),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1589),
.Y(n_1687)
);

AO21x1_ASAP7_75t_L g1688 ( 
.A1(n_1584),
.A2(n_1634),
.B(n_1599),
.Y(n_1688)
);

OR2x6_ASAP7_75t_L g1689 ( 
.A(n_1578),
.B(n_1661),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1620),
.B(n_1603),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1604),
.B(n_1631),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_SL g1692 ( 
.A(n_1613),
.B(n_1615),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1609),
.B(n_1610),
.Y(n_1693)
);

OAI22xp5_ASAP7_75t_L g1694 ( 
.A1(n_1579),
.A2(n_1608),
.B1(n_1634),
.B2(n_1615),
.Y(n_1694)
);

A2O1A1Ixp33_ASAP7_75t_L g1695 ( 
.A1(n_1618),
.A2(n_1586),
.B(n_1570),
.C(n_1558),
.Y(n_1695)
);

A2O1A1Ixp33_ASAP7_75t_L g1696 ( 
.A1(n_1586),
.A2(n_1570),
.B(n_1558),
.C(n_1622),
.Y(n_1696)
);

O2A1O1Ixp33_ASAP7_75t_SL g1697 ( 
.A1(n_1642),
.A2(n_1592),
.B(n_1593),
.C(n_1653),
.Y(n_1697)
);

OAI22xp5_ASAP7_75t_L g1698 ( 
.A1(n_1579),
.A2(n_1615),
.B1(n_1653),
.B2(n_1652),
.Y(n_1698)
);

AO32x2_ASAP7_75t_L g1699 ( 
.A1(n_1568),
.A2(n_1572),
.A3(n_1588),
.B1(n_1622),
.B2(n_1559),
.Y(n_1699)
);

AO21x2_ASAP7_75t_L g1700 ( 
.A1(n_1592),
.A2(n_1593),
.B(n_1554),
.Y(n_1700)
);

OA21x2_ASAP7_75t_L g1701 ( 
.A1(n_1629),
.A2(n_1559),
.B(n_1564),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1606),
.B(n_1640),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1600),
.Y(n_1703)
);

OAI22xp5_ASAP7_75t_L g1704 ( 
.A1(n_1579),
.A2(n_1652),
.B1(n_1606),
.B2(n_1633),
.Y(n_1704)
);

AOI221xp5_ASAP7_75t_L g1705 ( 
.A1(n_1623),
.A2(n_1596),
.B1(n_1644),
.B2(n_1629),
.C(n_1575),
.Y(n_1705)
);

CKINVDCx5p33_ASAP7_75t_R g1706 ( 
.A(n_1660),
.Y(n_1706)
);

A2O1A1Ixp33_ASAP7_75t_L g1707 ( 
.A1(n_1579),
.A2(n_1565),
.B(n_1574),
.C(n_1642),
.Y(n_1707)
);

OAI22xp5_ASAP7_75t_L g1708 ( 
.A1(n_1644),
.A2(n_1648),
.B1(n_1650),
.B2(n_1651),
.Y(n_1708)
);

HB1xp67_ASAP7_75t_L g1709 ( 
.A(n_1575),
.Y(n_1709)
);

OAI22xp5_ASAP7_75t_L g1710 ( 
.A1(n_1650),
.A2(n_1651),
.B1(n_1654),
.B2(n_1658),
.Y(n_1710)
);

AOI21xp5_ASAP7_75t_L g1711 ( 
.A1(n_1554),
.A2(n_1619),
.B(n_1617),
.Y(n_1711)
);

A2O1A1Ixp33_ASAP7_75t_L g1712 ( 
.A1(n_1643),
.A2(n_1619),
.B(n_1628),
.C(n_1614),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1628),
.B(n_1626),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1683),
.B(n_1564),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1667),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1683),
.B(n_1561),
.Y(n_1716)
);

AOI22xp33_ASAP7_75t_L g1717 ( 
.A1(n_1662),
.A2(n_1656),
.B1(n_1659),
.B2(n_1657),
.Y(n_1717)
);

NOR3xp33_ASAP7_75t_L g1718 ( 
.A(n_1672),
.B(n_1638),
.C(n_1569),
.Y(n_1718)
);

OR2x2_ASAP7_75t_L g1719 ( 
.A(n_1701),
.B(n_1580),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1677),
.B(n_1563),
.Y(n_1720)
);

HB1xp67_ASAP7_75t_L g1721 ( 
.A(n_1701),
.Y(n_1721)
);

AOI22xp33_ASAP7_75t_L g1722 ( 
.A1(n_1663),
.A2(n_1656),
.B1(n_1659),
.B2(n_1657),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1676),
.Y(n_1723)
);

INVx2_ASAP7_75t_SL g1724 ( 
.A(n_1689),
.Y(n_1724)
);

NOR2x1_ASAP7_75t_L g1725 ( 
.A(n_1686),
.B(n_1625),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1687),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1687),
.Y(n_1727)
);

AOI22xp33_ASAP7_75t_SL g1728 ( 
.A1(n_1665),
.A2(n_1619),
.B1(n_1660),
.B2(n_1654),
.Y(n_1728)
);

HB1xp67_ASAP7_75t_L g1729 ( 
.A(n_1701),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1703),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1680),
.B(n_1577),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1680),
.B(n_1577),
.Y(n_1732)
);

AOI22xp33_ASAP7_75t_L g1733 ( 
.A1(n_1669),
.A2(n_1656),
.B1(n_1658),
.B2(n_1649),
.Y(n_1733)
);

NOR2xp33_ASAP7_75t_L g1734 ( 
.A(n_1675),
.B(n_1641),
.Y(n_1734)
);

CKINVDCx20_ASAP7_75t_R g1735 ( 
.A(n_1684),
.Y(n_1735)
);

INVx2_ASAP7_75t_L g1736 ( 
.A(n_1693),
.Y(n_1736)
);

OR2x2_ASAP7_75t_L g1737 ( 
.A(n_1709),
.B(n_1582),
.Y(n_1737)
);

INVx1_ASAP7_75t_SL g1738 ( 
.A(n_1679),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1713),
.B(n_1588),
.Y(n_1739)
);

AOI211xp5_ASAP7_75t_L g1740 ( 
.A1(n_1697),
.A2(n_1569),
.B(n_1646),
.C(n_1649),
.Y(n_1740)
);

AND2x4_ASAP7_75t_L g1741 ( 
.A(n_1724),
.B(n_1678),
.Y(n_1741)
);

AOI221xp5_ASAP7_75t_L g1742 ( 
.A1(n_1722),
.A2(n_1675),
.B1(n_1671),
.B2(n_1670),
.C(n_1695),
.Y(n_1742)
);

BUFx3_ASAP7_75t_L g1743 ( 
.A(n_1724),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1714),
.B(n_1666),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1726),
.Y(n_1745)
);

NAND3xp33_ASAP7_75t_SL g1746 ( 
.A(n_1722),
.B(n_1671),
.C(n_1670),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1721),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1714),
.B(n_1716),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1716),
.B(n_1699),
.Y(n_1749)
);

OAI322xp33_ASAP7_75t_L g1750 ( 
.A1(n_1734),
.A2(n_1668),
.A3(n_1674),
.B1(n_1694),
.B2(n_1691),
.C1(n_1690),
.C2(n_1692),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1721),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1715),
.B(n_1699),
.Y(n_1752)
);

NAND3xp33_ASAP7_75t_L g1753 ( 
.A(n_1717),
.B(n_1695),
.C(n_1705),
.Y(n_1753)
);

OR2x2_ASAP7_75t_L g1754 ( 
.A(n_1719),
.B(n_1700),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1715),
.B(n_1699),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1726),
.Y(n_1756)
);

NOR2x1p5_ASAP7_75t_L g1757 ( 
.A(n_1739),
.B(n_1684),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1726),
.Y(n_1758)
);

NAND3xp33_ASAP7_75t_L g1759 ( 
.A(n_1717),
.B(n_1740),
.C(n_1733),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1727),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1729),
.Y(n_1761)
);

OR2x2_ASAP7_75t_L g1762 ( 
.A(n_1719),
.B(n_1700),
.Y(n_1762)
);

INVx3_ASAP7_75t_L g1763 ( 
.A(n_1730),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1715),
.B(n_1681),
.Y(n_1764)
);

OAI221xp5_ASAP7_75t_L g1765 ( 
.A1(n_1733),
.A2(n_1707),
.B1(n_1696),
.B2(n_1697),
.C(n_1692),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_SL g1766 ( 
.A(n_1728),
.B(n_1688),
.Y(n_1766)
);

OAI211xp5_ASAP7_75t_L g1767 ( 
.A1(n_1740),
.A2(n_1696),
.B(n_1707),
.C(n_1712),
.Y(n_1767)
);

OAI221xp5_ASAP7_75t_L g1768 ( 
.A1(n_1718),
.A2(n_1708),
.B1(n_1698),
.B2(n_1704),
.C(n_1712),
.Y(n_1768)
);

INVx2_ASAP7_75t_L g1769 ( 
.A(n_1729),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1727),
.Y(n_1770)
);

AOI31xp33_ASAP7_75t_L g1771 ( 
.A1(n_1728),
.A2(n_1710),
.A3(n_1706),
.B(n_1711),
.Y(n_1771)
);

BUFx3_ASAP7_75t_L g1772 ( 
.A(n_1724),
.Y(n_1772)
);

INVx4_ASAP7_75t_L g1773 ( 
.A(n_1737),
.Y(n_1773)
);

INVx4_ASAP7_75t_L g1774 ( 
.A(n_1737),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1723),
.B(n_1681),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1723),
.B(n_1681),
.Y(n_1776)
);

INVx3_ASAP7_75t_L g1777 ( 
.A(n_1736),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1723),
.B(n_1681),
.Y(n_1778)
);

OR2x2_ASAP7_75t_L g1779 ( 
.A(n_1719),
.B(n_1682),
.Y(n_1779)
);

INVx2_ASAP7_75t_L g1780 ( 
.A(n_1777),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1749),
.B(n_1720),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1745),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1749),
.B(n_1720),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1749),
.B(n_1731),
.Y(n_1784)
);

OR2x2_ASAP7_75t_L g1785 ( 
.A(n_1754),
.B(n_1739),
.Y(n_1785)
);

INVx1_ASAP7_75t_SL g1786 ( 
.A(n_1743),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1756),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1756),
.Y(n_1788)
);

BUFx2_ASAP7_75t_L g1789 ( 
.A(n_1743),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1752),
.B(n_1755),
.Y(n_1790)
);

OAI211xp5_ASAP7_75t_SL g1791 ( 
.A1(n_1742),
.A2(n_1718),
.B(n_1725),
.C(n_1734),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_SL g1792 ( 
.A(n_1753),
.B(n_1725),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1758),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1764),
.B(n_1720),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1777),
.Y(n_1795)
);

INVx1_ASAP7_75t_SL g1796 ( 
.A(n_1743),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1777),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1777),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1777),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_1763),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1760),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1760),
.Y(n_1802)
);

INVx2_ASAP7_75t_L g1803 ( 
.A(n_1763),
.Y(n_1803)
);

INVxp67_ASAP7_75t_L g1804 ( 
.A(n_1766),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1770),
.Y(n_1805)
);

OR2x2_ASAP7_75t_L g1806 ( 
.A(n_1754),
.B(n_1736),
.Y(n_1806)
);

NOR2x1p5_ASAP7_75t_L g1807 ( 
.A(n_1746),
.B(n_1706),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1764),
.B(n_1775),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1770),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1764),
.B(n_1732),
.Y(n_1810)
);

AND2x4_ASAP7_75t_L g1811 ( 
.A(n_1763),
.B(n_1725),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1782),
.Y(n_1812)
);

INVx2_ASAP7_75t_L g1813 ( 
.A(n_1800),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1782),
.Y(n_1814)
);

OR2x2_ASAP7_75t_L g1815 ( 
.A(n_1785),
.B(n_1779),
.Y(n_1815)
);

INVx1_ASAP7_75t_SL g1816 ( 
.A(n_1789),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1804),
.B(n_1738),
.Y(n_1817)
);

INVxp67_ASAP7_75t_SL g1818 ( 
.A(n_1792),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1790),
.B(n_1744),
.Y(n_1819)
);

AND2x4_ASAP7_75t_L g1820 ( 
.A(n_1789),
.B(n_1773),
.Y(n_1820)
);

BUFx3_ASAP7_75t_L g1821 ( 
.A(n_1789),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1782),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1787),
.Y(n_1823)
);

INVx2_ASAP7_75t_L g1824 ( 
.A(n_1800),
.Y(n_1824)
);

INVx1_ASAP7_75t_SL g1825 ( 
.A(n_1792),
.Y(n_1825)
);

AND2x2_ASAP7_75t_L g1826 ( 
.A(n_1790),
.B(n_1744),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1800),
.Y(n_1827)
);

INVx2_ASAP7_75t_L g1828 ( 
.A(n_1800),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1803),
.Y(n_1829)
);

OR2x2_ASAP7_75t_L g1830 ( 
.A(n_1785),
.B(n_1794),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1787),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1790),
.B(n_1744),
.Y(n_1832)
);

NOR3xp33_ASAP7_75t_L g1833 ( 
.A(n_1804),
.B(n_1753),
.C(n_1746),
.Y(n_1833)
);

AND2x2_ASAP7_75t_L g1834 ( 
.A(n_1784),
.B(n_1757),
.Y(n_1834)
);

INVx2_ASAP7_75t_SL g1835 ( 
.A(n_1786),
.Y(n_1835)
);

BUFx3_ASAP7_75t_L g1836 ( 
.A(n_1786),
.Y(n_1836)
);

INVx2_ASAP7_75t_L g1837 ( 
.A(n_1803),
.Y(n_1837)
);

INVx2_ASAP7_75t_L g1838 ( 
.A(n_1803),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1787),
.Y(n_1839)
);

AOI22xp5_ASAP7_75t_L g1840 ( 
.A1(n_1791),
.A2(n_1759),
.B1(n_1742),
.B2(n_1767),
.Y(n_1840)
);

INVx2_ASAP7_75t_L g1841 ( 
.A(n_1803),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1788),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1788),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1784),
.B(n_1757),
.Y(n_1844)
);

AOI21x1_ASAP7_75t_L g1845 ( 
.A1(n_1788),
.A2(n_1766),
.B(n_1751),
.Y(n_1845)
);

OR2x2_ASAP7_75t_L g1846 ( 
.A(n_1785),
.B(n_1779),
.Y(n_1846)
);

OAI21xp33_ASAP7_75t_L g1847 ( 
.A1(n_1791),
.A2(n_1759),
.B(n_1771),
.Y(n_1847)
);

NAND2xp33_ASAP7_75t_SL g1848 ( 
.A(n_1807),
.B(n_1735),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1801),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1807),
.B(n_1738),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1801),
.Y(n_1851)
);

AOI22xp5_ASAP7_75t_L g1852 ( 
.A1(n_1796),
.A2(n_1767),
.B1(n_1765),
.B2(n_1768),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1784),
.B(n_1743),
.Y(n_1853)
);

NOR2xp33_ASAP7_75t_L g1854 ( 
.A(n_1796),
.B(n_1735),
.Y(n_1854)
);

OR2x2_ASAP7_75t_L g1855 ( 
.A(n_1794),
.B(n_1779),
.Y(n_1855)
);

OR2x2_ASAP7_75t_L g1856 ( 
.A(n_1781),
.B(n_1748),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1801),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1834),
.B(n_1808),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1812),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_SL g1860 ( 
.A(n_1847),
.B(n_1771),
.Y(n_1860)
);

OR2x2_ASAP7_75t_L g1861 ( 
.A(n_1825),
.B(n_1781),
.Y(n_1861)
);

INVx2_ASAP7_75t_L g1862 ( 
.A(n_1845),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1834),
.B(n_1808),
.Y(n_1863)
);

HB1xp67_ASAP7_75t_L g1864 ( 
.A(n_1821),
.Y(n_1864)
);

NOR2xp33_ASAP7_75t_L g1865 ( 
.A(n_1854),
.B(n_1655),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1812),
.Y(n_1866)
);

INVx2_ASAP7_75t_SL g1867 ( 
.A(n_1821),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1814),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1814),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1822),
.Y(n_1870)
);

OAI22xp5_ASAP7_75t_SL g1871 ( 
.A1(n_1840),
.A2(n_1765),
.B1(n_1768),
.B2(n_1750),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1833),
.B(n_1847),
.Y(n_1872)
);

INVx1_ASAP7_75t_SL g1873 ( 
.A(n_1825),
.Y(n_1873)
);

AND2x2_ASAP7_75t_L g1874 ( 
.A(n_1844),
.B(n_1819),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1840),
.B(n_1773),
.Y(n_1875)
);

BUFx2_ASAP7_75t_L g1876 ( 
.A(n_1821),
.Y(n_1876)
);

INVx2_ASAP7_75t_L g1877 ( 
.A(n_1845),
.Y(n_1877)
);

XOR2xp5_ASAP7_75t_L g1878 ( 
.A(n_1852),
.B(n_1645),
.Y(n_1878)
);

AND2x4_ASAP7_75t_L g1879 ( 
.A(n_1819),
.B(n_1811),
.Y(n_1879)
);

BUFx2_ASAP7_75t_L g1880 ( 
.A(n_1836),
.Y(n_1880)
);

CKINVDCx16_ASAP7_75t_R g1881 ( 
.A(n_1852),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1822),
.Y(n_1882)
);

INVx1_ASAP7_75t_SL g1883 ( 
.A(n_1848),
.Y(n_1883)
);

NOR3xp33_ASAP7_75t_L g1884 ( 
.A(n_1818),
.B(n_1750),
.C(n_1646),
.Y(n_1884)
);

HB1xp67_ASAP7_75t_L g1885 ( 
.A(n_1836),
.Y(n_1885)
);

AND2x2_ASAP7_75t_L g1886 ( 
.A(n_1844),
.B(n_1808),
.Y(n_1886)
);

NOR2xp33_ASAP7_75t_SL g1887 ( 
.A(n_1817),
.B(n_1773),
.Y(n_1887)
);

OR2x6_ASAP7_75t_L g1888 ( 
.A(n_1836),
.B(n_1689),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1826),
.B(n_1810),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1823),
.Y(n_1890)
);

OR2x2_ASAP7_75t_L g1891 ( 
.A(n_1830),
.B(n_1783),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_L g1892 ( 
.A(n_1835),
.B(n_1773),
.Y(n_1892)
);

OAI22xp5_ASAP7_75t_L g1893 ( 
.A1(n_1850),
.A2(n_1783),
.B1(n_1748),
.B2(n_1689),
.Y(n_1893)
);

AND2x2_ASAP7_75t_L g1894 ( 
.A(n_1826),
.B(n_1810),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1835),
.B(n_1773),
.Y(n_1895)
);

AOI22xp5_ASAP7_75t_L g1896 ( 
.A1(n_1860),
.A2(n_1820),
.B1(n_1853),
.B2(n_1832),
.Y(n_1896)
);

OAI32xp33_ASAP7_75t_L g1897 ( 
.A1(n_1881),
.A2(n_1816),
.A3(n_1830),
.B1(n_1815),
.B2(n_1846),
.Y(n_1897)
);

INVxp67_ASAP7_75t_L g1898 ( 
.A(n_1880),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_1881),
.B(n_1832),
.Y(n_1899)
);

AOI221xp5_ASAP7_75t_L g1900 ( 
.A1(n_1872),
.A2(n_1816),
.B1(n_1820),
.B2(n_1823),
.C(n_1857),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1880),
.Y(n_1901)
);

OAI21xp5_ASAP7_75t_L g1902 ( 
.A1(n_1884),
.A2(n_1820),
.B(n_1853),
.Y(n_1902)
);

AND2x2_ASAP7_75t_L g1903 ( 
.A(n_1858),
.B(n_1820),
.Y(n_1903)
);

XNOR2xp5_ASAP7_75t_L g1904 ( 
.A(n_1871),
.B(n_1702),
.Y(n_1904)
);

NAND2x1_ASAP7_75t_L g1905 ( 
.A(n_1876),
.B(n_1811),
.Y(n_1905)
);

INVx2_ASAP7_75t_L g1906 ( 
.A(n_1876),
.Y(n_1906)
);

OAI21xp33_ASAP7_75t_L g1907 ( 
.A1(n_1875),
.A2(n_1846),
.B(n_1815),
.Y(n_1907)
);

HB1xp67_ASAP7_75t_L g1908 ( 
.A(n_1885),
.Y(n_1908)
);

NOR2xp33_ASAP7_75t_L g1909 ( 
.A(n_1871),
.B(n_1856),
.Y(n_1909)
);

AOI22xp33_ASAP7_75t_L g1910 ( 
.A1(n_1883),
.A2(n_1762),
.B1(n_1842),
.B2(n_1831),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1859),
.Y(n_1911)
);

AOI22xp5_ASAP7_75t_L g1912 ( 
.A1(n_1878),
.A2(n_1664),
.B1(n_1673),
.B2(n_1741),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1859),
.Y(n_1913)
);

OAI21xp5_ASAP7_75t_L g1914 ( 
.A1(n_1878),
.A2(n_1839),
.B(n_1831),
.Y(n_1914)
);

AOI221xp5_ASAP7_75t_L g1915 ( 
.A1(n_1873),
.A2(n_1857),
.B1(n_1839),
.B2(n_1842),
.C(n_1851),
.Y(n_1915)
);

AOI322xp5_ASAP7_75t_L g1916 ( 
.A1(n_1858),
.A2(n_1863),
.A3(n_1886),
.B1(n_1877),
.B2(n_1862),
.C1(n_1889),
.C2(n_1894),
.Y(n_1916)
);

NAND4xp25_ASAP7_75t_L g1917 ( 
.A(n_1865),
.B(n_1887),
.C(n_1874),
.D(n_1861),
.Y(n_1917)
);

AOI22xp33_ASAP7_75t_L g1918 ( 
.A1(n_1863),
.A2(n_1762),
.B1(n_1849),
.B2(n_1851),
.Y(n_1918)
);

INVx2_ASAP7_75t_L g1919 ( 
.A(n_1886),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1866),
.Y(n_1920)
);

OAI32xp33_ASAP7_75t_L g1921 ( 
.A1(n_1862),
.A2(n_1856),
.A3(n_1855),
.B1(n_1774),
.B2(n_1843),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1864),
.B(n_1855),
.Y(n_1922)
);

AOI21xp5_ASAP7_75t_L g1923 ( 
.A1(n_1867),
.A2(n_1849),
.B(n_1843),
.Y(n_1923)
);

AOI222xp33_ASAP7_75t_L g1924 ( 
.A1(n_1909),
.A2(n_1862),
.B1(n_1877),
.B2(n_1867),
.C1(n_1868),
.C2(n_1890),
.Y(n_1924)
);

OR2x2_ASAP7_75t_L g1925 ( 
.A(n_1899),
.B(n_1861),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1909),
.B(n_1874),
.Y(n_1926)
);

AOI21xp33_ASAP7_75t_SL g1927 ( 
.A1(n_1914),
.A2(n_1888),
.B(n_1892),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1901),
.B(n_1889),
.Y(n_1928)
);

NOR2xp67_ASAP7_75t_SL g1929 ( 
.A(n_1908),
.B(n_1877),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1906),
.B(n_1894),
.Y(n_1930)
);

OAI22xp5_ASAP7_75t_L g1931 ( 
.A1(n_1896),
.A2(n_1888),
.B1(n_1895),
.B2(n_1891),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1908),
.Y(n_1932)
);

NAND3xp33_ASAP7_75t_L g1933 ( 
.A(n_1900),
.B(n_1868),
.C(n_1866),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1898),
.Y(n_1934)
);

AOI21xp33_ASAP7_75t_L g1935 ( 
.A1(n_1897),
.A2(n_1888),
.B(n_1893),
.Y(n_1935)
);

OAI222xp33_ASAP7_75t_L g1936 ( 
.A1(n_1912),
.A2(n_1888),
.B1(n_1891),
.B2(n_1879),
.C1(n_1774),
.C2(n_1890),
.Y(n_1936)
);

NOR2xp33_ASAP7_75t_L g1937 ( 
.A(n_1917),
.B(n_1888),
.Y(n_1937)
);

OAI22xp5_ASAP7_75t_L g1938 ( 
.A1(n_1904),
.A2(n_1879),
.B1(n_1882),
.B2(n_1870),
.Y(n_1938)
);

OAI21xp33_ASAP7_75t_SL g1939 ( 
.A1(n_1916),
.A2(n_1910),
.B(n_1915),
.Y(n_1939)
);

NOR2x1_ASAP7_75t_L g1940 ( 
.A(n_1911),
.B(n_1869),
.Y(n_1940)
);

OAI22xp33_ASAP7_75t_L g1941 ( 
.A1(n_1902),
.A2(n_1774),
.B1(n_1772),
.B2(n_1879),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1898),
.Y(n_1942)
);

NOR3xp33_ASAP7_75t_L g1943 ( 
.A(n_1907),
.B(n_1870),
.C(n_1869),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1913),
.Y(n_1944)
);

AND2x2_ASAP7_75t_L g1945 ( 
.A(n_1934),
.B(n_1903),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1940),
.Y(n_1946)
);

INVx2_ASAP7_75t_L g1947 ( 
.A(n_1932),
.Y(n_1947)
);

XNOR2xp5_ASAP7_75t_L g1948 ( 
.A(n_1938),
.B(n_1922),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1942),
.Y(n_1949)
);

INVx2_ASAP7_75t_L g1950 ( 
.A(n_1925),
.Y(n_1950)
);

BUFx2_ASAP7_75t_L g1951 ( 
.A(n_1930),
.Y(n_1951)
);

NOR2x1_ASAP7_75t_L g1952 ( 
.A(n_1933),
.B(n_1920),
.Y(n_1952)
);

AOI21xp5_ASAP7_75t_L g1953 ( 
.A1(n_1939),
.A2(n_1923),
.B(n_1921),
.Y(n_1953)
);

INVx2_ASAP7_75t_L g1954 ( 
.A(n_1928),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1926),
.B(n_1919),
.Y(n_1955)
);

NAND3xp33_ASAP7_75t_SL g1956 ( 
.A(n_1953),
.B(n_1924),
.C(n_1927),
.Y(n_1956)
);

AOI211xp5_ASAP7_75t_L g1957 ( 
.A1(n_1948),
.A2(n_1935),
.B(n_1929),
.C(n_1937),
.Y(n_1957)
);

AOI21xp5_ASAP7_75t_L g1958 ( 
.A1(n_1952),
.A2(n_1924),
.B(n_1931),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_SL g1959 ( 
.A(n_1950),
.B(n_1941),
.Y(n_1959)
);

NOR3xp33_ASAP7_75t_L g1960 ( 
.A(n_1950),
.B(n_1944),
.C(n_1936),
.Y(n_1960)
);

AND2x4_ASAP7_75t_L g1961 ( 
.A(n_1945),
.B(n_1943),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1945),
.B(n_1910),
.Y(n_1962)
);

NAND4xp25_ASAP7_75t_L g1963 ( 
.A(n_1955),
.B(n_1918),
.C(n_1882),
.D(n_1879),
.Y(n_1963)
);

XNOR2x1_ASAP7_75t_L g1964 ( 
.A(n_1954),
.B(n_1905),
.Y(n_1964)
);

NOR2xp33_ASAP7_75t_L g1965 ( 
.A(n_1951),
.B(n_1918),
.Y(n_1965)
);

O2A1O1Ixp33_ASAP7_75t_SL g1966 ( 
.A1(n_1956),
.A2(n_1946),
.B(n_1947),
.C(n_1949),
.Y(n_1966)
);

AO32x1_ASAP7_75t_L g1967 ( 
.A1(n_1960),
.A2(n_1947),
.A3(n_1954),
.B1(n_1841),
.B2(n_1838),
.Y(n_1967)
);

AOI211xp5_ASAP7_75t_L g1968 ( 
.A1(n_1958),
.A2(n_1811),
.B(n_1838),
.C(n_1837),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1961),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1962),
.Y(n_1970)
);

AOI211xp5_ASAP7_75t_L g1971 ( 
.A1(n_1965),
.A2(n_1811),
.B(n_1838),
.C(n_1837),
.Y(n_1971)
);

OAI221xp5_ASAP7_75t_SL g1972 ( 
.A1(n_1968),
.A2(n_1957),
.B1(n_1963),
.B2(n_1964),
.C(n_1959),
.Y(n_1972)
);

OA22x2_ASAP7_75t_L g1973 ( 
.A1(n_1969),
.A2(n_1841),
.B1(n_1837),
.B2(n_1829),
.Y(n_1973)
);

AOI221x1_ASAP7_75t_L g1974 ( 
.A1(n_1970),
.A2(n_1841),
.B1(n_1829),
.B2(n_1828),
.C(n_1827),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1967),
.Y(n_1975)
);

OAI22xp5_ASAP7_75t_L g1976 ( 
.A1(n_1971),
.A2(n_1811),
.B1(n_1769),
.B2(n_1751),
.Y(n_1976)
);

XNOR2xp5_ASAP7_75t_L g1977 ( 
.A(n_1966),
.B(n_1685),
.Y(n_1977)
);

OAI221xp5_ASAP7_75t_L g1978 ( 
.A1(n_1966),
.A2(n_1813),
.B1(n_1828),
.B2(n_1827),
.C(n_1824),
.Y(n_1978)
);

AOI22xp5_ASAP7_75t_SL g1979 ( 
.A1(n_1977),
.A2(n_1811),
.B1(n_1747),
.B2(n_1761),
.Y(n_1979)
);

XOR2xp5_ASAP7_75t_L g1980 ( 
.A(n_1975),
.B(n_1973),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_L g1981 ( 
.A(n_1976),
.B(n_1802),
.Y(n_1981)
);

OA22x2_ASAP7_75t_L g1982 ( 
.A1(n_1974),
.A2(n_1829),
.B1(n_1828),
.B2(n_1827),
.Y(n_1982)
);

INVx1_ASAP7_75t_SL g1983 ( 
.A(n_1972),
.Y(n_1983)
);

NAND4xp75_ASAP7_75t_L g1984 ( 
.A(n_1978),
.B(n_1824),
.C(n_1813),
.D(n_1761),
.Y(n_1984)
);

NAND4xp75_ASAP7_75t_L g1985 ( 
.A(n_1980),
.B(n_1824),
.C(n_1813),
.D(n_1761),
.Y(n_1985)
);

INVx2_ASAP7_75t_L g1986 ( 
.A(n_1982),
.Y(n_1986)
);

AOI322xp5_ASAP7_75t_L g1987 ( 
.A1(n_1983),
.A2(n_1747),
.A3(n_1751),
.B1(n_1769),
.B2(n_1778),
.C1(n_1776),
.C2(n_1775),
.Y(n_1987)
);

OAI22xp5_ASAP7_75t_L g1988 ( 
.A1(n_1979),
.A2(n_1799),
.B1(n_1797),
.B2(n_1798),
.Y(n_1988)
);

INVxp67_ASAP7_75t_SL g1989 ( 
.A(n_1986),
.Y(n_1989)
);

OAI22x1_ASAP7_75t_L g1990 ( 
.A1(n_1989),
.A2(n_1985),
.B1(n_1981),
.B2(n_1984),
.Y(n_1990)
);

XNOR2xp5_ASAP7_75t_L g1991 ( 
.A(n_1990),
.B(n_1988),
.Y(n_1991)
);

AOI22x1_ASAP7_75t_L g1992 ( 
.A1(n_1990),
.A2(n_1987),
.B1(n_1769),
.B2(n_1747),
.Y(n_1992)
);

OAI31xp33_ASAP7_75t_L g1993 ( 
.A1(n_1991),
.A2(n_1769),
.A3(n_1780),
.B(n_1795),
.Y(n_1993)
);

OAI22x1_ASAP7_75t_L g1994 ( 
.A1(n_1992),
.A2(n_1780),
.B1(n_1795),
.B2(n_1797),
.Y(n_1994)
);

AOI221xp5_ASAP7_75t_L g1995 ( 
.A1(n_1994),
.A2(n_1802),
.B1(n_1805),
.B2(n_1809),
.C(n_1793),
.Y(n_1995)
);

OAI22xp5_ASAP7_75t_L g1996 ( 
.A1(n_1993),
.A2(n_1795),
.B1(n_1797),
.B2(n_1798),
.Y(n_1996)
);

AOI21xp5_ASAP7_75t_L g1997 ( 
.A1(n_1996),
.A2(n_1795),
.B(n_1780),
.Y(n_1997)
);

AND2x2_ASAP7_75t_L g1998 ( 
.A(n_1997),
.B(n_1995),
.Y(n_1998)
);

AOI21xp5_ASAP7_75t_L g1999 ( 
.A1(n_1998),
.A2(n_1797),
.B(n_1780),
.Y(n_1999)
);

OAI221xp5_ASAP7_75t_R g2000 ( 
.A1(n_1999),
.A2(n_1647),
.B1(n_1798),
.B2(n_1799),
.C(n_1806),
.Y(n_2000)
);

AOI22xp33_ASAP7_75t_L g2001 ( 
.A1(n_2000),
.A2(n_1799),
.B1(n_1798),
.B2(n_1802),
.Y(n_2001)
);


endmodule