module fake_jpeg_22349_n_186 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_186);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_186;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_122;
wire n_75;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_14),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx5_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx14_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx5p33_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_14),
.B(n_2),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_0),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_32),
.B(n_18),
.Y(n_66)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

BUFx24_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

INVxp67_ASAP7_75t_SL g68 ( 
.A(n_34),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_35),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_37),
.A2(n_44),
.B1(n_17),
.B2(n_28),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_30),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_38),
.B(n_41),
.Y(n_71)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_43),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_40),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_30),
.B(n_22),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_15),
.B(n_0),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_45),
.B(n_23),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_32),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_48),
.B(n_57),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_34),
.A2(n_19),
.B(n_28),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_51),
.A2(n_53),
.B(n_4),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_22),
.Y(n_52)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_34),
.A2(n_33),
.B(n_35),
.Y(n_53)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_58),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_56),
.B(n_64),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_32),
.B(n_15),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_34),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_35),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_59),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_16),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_63),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_21),
.Y(n_62)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_62),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_24),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

NOR2x1_ASAP7_75t_R g88 ( 
.A(n_66),
.B(n_1),
.Y(n_88)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_67),
.B(n_70),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_42),
.A2(n_27),
.B1(n_26),
.B2(n_29),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_69),
.A2(n_74),
.B1(n_25),
.B2(n_16),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_40),
.B(n_21),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_40),
.B(n_29),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_72),
.B(n_4),
.Y(n_92)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_73),
.B(n_8),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_39),
.A2(n_27),
.B1(n_26),
.B2(n_25),
.Y(n_74)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_76),
.B(n_93),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_80),
.A2(n_91),
.B1(n_69),
.B2(n_56),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_73),
.B(n_23),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_83),
.B(n_85),
.Y(n_102)
);

BUFx24_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_59),
.B(n_1),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_88),
.A2(n_47),
.B1(n_55),
.B2(n_6),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

INVx13_ASAP7_75t_L g112 ( 
.A(n_89),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_49),
.B(n_2),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_90),
.B(n_92),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_51),
.A2(n_48),
.B1(n_53),
.B2(n_60),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_94),
.A2(n_65),
.B1(n_71),
.B2(n_55),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_66),
.B(n_72),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_95),
.B(n_63),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_63),
.B(n_4),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_96),
.B(n_100),
.Y(n_118)
);

BUFx4f_ASAP7_75t_L g97 ( 
.A(n_46),
.Y(n_97)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

AND2x4_ASAP7_75t_L g99 ( 
.A(n_66),
.B(n_5),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_58),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_57),
.B(n_5),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_101),
.A2(n_111),
.B1(n_92),
.B2(n_88),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_116),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_99),
.B(n_74),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_105),
.B(n_122),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_94),
.A2(n_67),
.B1(n_61),
.B2(n_64),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_106),
.A2(n_113),
.B1(n_120),
.B2(n_91),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_86),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_107),
.B(n_117),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_108),
.B(n_119),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_82),
.A2(n_47),
.B1(n_46),
.B2(n_58),
.Y(n_113)
);

AND2x6_ASAP7_75t_L g115 ( 
.A(n_99),
.B(n_12),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_115),
.B(n_99),
.C(n_78),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_79),
.B(n_54),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_82),
.A2(n_46),
.B1(n_54),
.B2(n_10),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_79),
.B(n_77),
.Y(n_121)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_121),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_78),
.B(n_8),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_124),
.B(n_134),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_103),
.A2(n_95),
.B(n_116),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_125),
.B(n_135),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_126),
.A2(n_127),
.B1(n_137),
.B2(n_138),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_106),
.A2(n_80),
.B1(n_86),
.B2(n_76),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_113),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_128),
.B(n_133),
.Y(n_142)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_110),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g134 ( 
.A(n_104),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_107),
.B(n_87),
.Y(n_136)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_136),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_112),
.A2(n_84),
.B1(n_97),
.B2(n_81),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_109),
.B(n_98),
.Y(n_139)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_139),
.Y(n_154)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_120),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_140),
.B(n_141),
.Y(n_151)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_101),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_130),
.B(n_119),
.C(n_114),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_143),
.B(n_152),
.C(n_123),
.Y(n_159)
);

OAI22x1_ASAP7_75t_L g144 ( 
.A1(n_134),
.A2(n_84),
.B1(n_105),
.B2(n_115),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_144),
.A2(n_127),
.B1(n_140),
.B2(n_126),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_134),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_145),
.A2(n_112),
.B(n_89),
.Y(n_166)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_129),
.Y(n_146)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_146),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_135),
.A2(n_81),
.B1(n_109),
.B2(n_117),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_150),
.A2(n_128),
.B1(n_104),
.B2(n_84),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_130),
.B(n_75),
.C(n_98),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_123),
.B(n_118),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_155),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_157),
.A2(n_153),
.B1(n_150),
.B2(n_144),
.Y(n_168)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_151),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_158),
.B(n_155),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_159),
.B(n_160),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_148),
.A2(n_125),
.B(n_124),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_143),
.B(n_141),
.C(n_132),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_162),
.B(n_152),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_163),
.B(n_166),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_142),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_164),
.B(n_165),
.Y(n_167)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_151),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_168),
.B(n_170),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_161),
.B(n_147),
.Y(n_171)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_171),
.Y(n_178)
);

A2O1A1Ixp33_ASAP7_75t_SL g173 ( 
.A1(n_158),
.A2(n_148),
.B(n_149),
.C(n_131),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_163),
.B(n_146),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_174),
.B(n_166),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_176),
.B(n_177),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_169),
.A2(n_156),
.B1(n_160),
.B2(n_162),
.Y(n_177)
);

AOI322xp5_ASAP7_75t_L g180 ( 
.A1(n_173),
.A2(n_156),
.A3(n_159),
.B1(n_154),
.B2(n_122),
.C1(n_102),
.C2(n_145),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_180),
.B(n_167),
.C(n_172),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_181),
.B(n_179),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_178),
.A2(n_175),
.B1(n_54),
.B2(n_11),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_184),
.B(n_182),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_185),
.B(n_183),
.Y(n_186)
);


endmodule