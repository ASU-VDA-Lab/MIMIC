module fake_jpeg_2075_n_501 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_501);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_501;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

BUFx8_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

INVx11_ASAP7_75t_SL g45 ( 
.A(n_4),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_10),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_56),
.Y(n_125)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_57),
.Y(n_131)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_58),
.Y(n_151)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_59),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_60),
.Y(n_137)
);

BUFx16f_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g184 ( 
.A(n_61),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_62),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_63),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_64),
.Y(n_123)
);

AOI21xp33_ASAP7_75t_L g65 ( 
.A1(n_21),
.A2(n_17),
.B(n_16),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_65),
.B(n_3),
.Y(n_197)
);

BUFx12_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g135 ( 
.A(n_66),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_38),
.B(n_17),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_67),
.B(n_68),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_24),
.B(n_16),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_69),
.Y(n_150)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_70),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_24),
.B(n_16),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_71),
.B(n_82),
.Y(n_129)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g172 ( 
.A(n_72),
.Y(n_172)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_20),
.Y(n_73)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_73),
.Y(n_145)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_74),
.Y(n_173)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_31),
.Y(n_75)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_75),
.Y(n_183)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_76),
.Y(n_141)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_31),
.Y(n_77)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_77),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_45),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_78),
.B(n_79),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_22),
.Y(n_79)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_80),
.Y(n_138)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_26),
.Y(n_81)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_81),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_36),
.B(n_0),
.Y(n_82)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_35),
.Y(n_83)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_83),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_22),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_84),
.B(n_90),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_26),
.B(n_0),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_85),
.B(n_88),
.Y(n_142)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_39),
.Y(n_86)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_86),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_28),
.Y(n_87)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_87),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_34),
.B(n_1),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_29),
.Y(n_89)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_89),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_22),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_91),
.Y(n_153)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_36),
.Y(n_92)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_92),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_29),
.Y(n_93)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_93),
.Y(n_147)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_28),
.Y(n_94)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_94),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_19),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_95),
.B(n_106),
.Y(n_146)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_18),
.Y(n_96)
);

INVx5_ASAP7_75t_SL g175 ( 
.A(n_96),
.Y(n_175)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_97),
.Y(n_163)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_34),
.Y(n_98)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_98),
.Y(n_192)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_50),
.Y(n_99)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_99),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_32),
.B(n_14),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_100),
.B(n_110),
.Y(n_152)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_50),
.Y(n_101)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_101),
.Y(n_155)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_53),
.Y(n_102)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_102),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_52),
.Y(n_103)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_103),
.Y(n_160)
);

BUFx12_ASAP7_75t_L g104 ( 
.A(n_19),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_104),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_29),
.Y(n_105)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_105),
.Y(n_167)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_37),
.Y(n_106)
);

BUFx16f_ASAP7_75t_L g107 ( 
.A(n_19),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g159 ( 
.A(n_107),
.Y(n_159)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_37),
.Y(n_108)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_108),
.Y(n_165)
);

BUFx16f_ASAP7_75t_L g109 ( 
.A(n_25),
.Y(n_109)
);

INVx8_ASAP7_75t_L g182 ( 
.A(n_109),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_32),
.B(n_33),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_49),
.Y(n_111)
);

INVx6_ASAP7_75t_L g201 ( 
.A(n_111),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_53),
.Y(n_112)
);

NAND2xp33_ASAP7_75t_SL g136 ( 
.A(n_112),
.B(n_55),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_49),
.Y(n_113)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_113),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_49),
.Y(n_114)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_114),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g115 ( 
.A(n_25),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_115),
.B(n_120),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_47),
.Y(n_116)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_116),
.Y(n_170)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_53),
.Y(n_117)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_117),
.Y(n_171)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_41),
.Y(n_118)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_118),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_47),
.Y(n_119)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_119),
.Y(n_177)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_41),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_58),
.A2(n_40),
.B1(n_30),
.B2(n_53),
.Y(n_122)
);

OA22x2_ASAP7_75t_L g209 ( 
.A1(n_122),
.A2(n_140),
.B1(n_174),
.B2(n_186),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_72),
.B(n_26),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_126),
.B(n_132),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_73),
.B(n_55),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_112),
.B(n_26),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_133),
.B(n_143),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_136),
.B(n_144),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_58),
.A2(n_40),
.B1(n_30),
.B2(n_48),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_107),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_91),
.B(n_54),
.C(n_51),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_62),
.A2(n_18),
.B1(n_54),
.B2(n_46),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_149),
.A2(n_164),
.B1(n_179),
.B2(n_185),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_117),
.B(n_51),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_161),
.B(n_162),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_103),
.B(n_46),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_63),
.A2(n_48),
.B1(n_42),
.B2(n_33),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_74),
.A2(n_42),
.B1(n_44),
.B2(n_43),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_61),
.B(n_47),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_178),
.B(n_190),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_64),
.A2(n_43),
.B1(n_25),
.B2(n_44),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_74),
.B(n_1),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_180),
.B(n_195),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_89),
.A2(n_43),
.B1(n_25),
.B2(n_5),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_56),
.A2(n_86),
.B1(n_83),
.B2(n_76),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_119),
.A2(n_43),
.B1(n_25),
.B2(n_5),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_189),
.A2(n_175),
.B1(n_191),
.B2(n_125),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_116),
.B(n_2),
.Y(n_190)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_114),
.Y(n_193)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_193),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_109),
.B(n_3),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_94),
.A2(n_43),
.B1(n_5),
.B2(n_6),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_196),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_197),
.B(n_198),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_93),
.B(n_3),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_60),
.B(n_14),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_200),
.B(n_202),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_111),
.Y(n_202)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_139),
.Y(n_205)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_205),
.Y(n_276)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_165),
.Y(n_207)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_207),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_124),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_208),
.Y(n_314)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_182),
.Y(n_212)
);

INVx4_ASAP7_75t_SL g304 ( 
.A(n_212),
.Y(n_304)
);

AND2x2_ASAP7_75t_SL g213 ( 
.A(n_180),
.B(n_87),
.Y(n_213)
);

CKINVDCx14_ASAP7_75t_R g291 ( 
.A(n_213),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_129),
.B(n_113),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_216),
.B(n_227),
.Y(n_282)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_168),
.Y(n_217)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_217),
.Y(n_272)
);

INVx13_ASAP7_75t_L g218 ( 
.A(n_159),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_218),
.Y(n_317)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_169),
.Y(n_219)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_219),
.Y(n_287)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_176),
.Y(n_220)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_220),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_195),
.A2(n_134),
.B(n_152),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_221),
.A2(n_258),
.B(n_211),
.Y(n_296)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_182),
.Y(n_223)
);

BUFx2_ASAP7_75t_L g288 ( 
.A(n_223),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_124),
.Y(n_224)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_224),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_159),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_225),
.B(n_232),
.Y(n_273)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_138),
.Y(n_226)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_226),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_142),
.B(n_105),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_146),
.B(n_102),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_229),
.B(n_242),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_121),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_230),
.Y(n_280)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_138),
.Y(n_231)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_231),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_133),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_L g233 ( 
.A1(n_163),
.A2(n_101),
.B1(n_99),
.B2(n_80),
.Y(n_233)
);

OAI22xp33_ASAP7_75t_SL g308 ( 
.A1(n_233),
.A2(n_261),
.B1(n_203),
.B2(n_247),
.Y(n_308)
);

INVx8_ASAP7_75t_L g234 ( 
.A(n_184),
.Y(n_234)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_234),
.Y(n_302)
);

OAI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_149),
.A2(n_66),
.B1(n_104),
.B2(n_8),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g279 ( 
.A1(n_236),
.A2(n_151),
.B1(n_173),
.B2(n_191),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_127),
.B(n_6),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_237),
.B(n_239),
.Y(n_285)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_130),
.Y(n_238)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_238),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_181),
.B(n_6),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_183),
.B(n_7),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_240),
.B(n_243),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_241),
.A2(n_246),
.B1(n_255),
.B2(n_257),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_188),
.B(n_11),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_192),
.B(n_11),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_194),
.B(n_13),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_244),
.B(n_251),
.Y(n_275)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_170),
.Y(n_245)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_245),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_196),
.A2(n_66),
.B1(n_14),
.B2(n_13),
.Y(n_246)
);

OR2x2_ASAP7_75t_SL g247 ( 
.A(n_153),
.B(n_104),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_247),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g248 ( 
.A(n_141),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_248),
.Y(n_281)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_172),
.Y(n_249)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_249),
.Y(n_319)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_158),
.Y(n_250)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_250),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_145),
.B(n_148),
.Y(n_251)
);

O2A1O1Ixp33_ASAP7_75t_L g252 ( 
.A1(n_174),
.A2(n_186),
.B(n_175),
.C(n_140),
.Y(n_252)
);

O2A1O1Ixp33_ASAP7_75t_L g283 ( 
.A1(n_252),
.A2(n_135),
.B(n_166),
.C(n_184),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_187),
.B(n_172),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_253),
.B(n_254),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_126),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_122),
.A2(n_177),
.B1(n_123),
.B2(n_201),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_131),
.B(n_154),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_256),
.B(n_260),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_121),
.A2(n_123),
.B1(n_201),
.B2(n_128),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_171),
.A2(n_150),
.B(n_157),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_160),
.B(n_157),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_259),
.B(n_263),
.Y(n_301)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_199),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_261),
.A2(n_258),
.B1(n_235),
.B2(n_265),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_128),
.B(n_147),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_262),
.B(n_208),
.Y(n_300)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_199),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_147),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_264),
.B(n_268),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_141),
.B(n_125),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_265),
.B(n_266),
.Y(n_305)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_155),
.Y(n_266)
);

AND2x2_ASAP7_75t_SL g267 ( 
.A(n_137),
.B(n_156),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_267),
.B(n_265),
.C(n_256),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_184),
.B(n_156),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_155),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_269),
.B(n_270),
.Y(n_310)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_158),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_216),
.A2(n_167),
.B1(n_137),
.B2(n_166),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_274),
.A2(n_290),
.B1(n_294),
.B2(n_267),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_279),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_283),
.A2(n_286),
.B(n_209),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_252),
.A2(n_167),
.B(n_222),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_222),
.A2(n_227),
.B1(n_204),
.B2(n_213),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_296),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_206),
.B(n_222),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_297),
.B(n_312),
.C(n_293),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_300),
.B(n_311),
.Y(n_321)
);

AOI22x1_ASAP7_75t_SL g303 ( 
.A1(n_213),
.A2(n_240),
.B1(n_239),
.B2(n_243),
.Y(n_303)
);

AOI211xp5_ASAP7_75t_L g322 ( 
.A1(n_303),
.A2(n_267),
.B(n_260),
.C(n_218),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_L g339 ( 
.A1(n_308),
.A2(n_226),
.B1(n_245),
.B2(n_215),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_228),
.B(n_237),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_221),
.B(n_210),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_214),
.B(n_205),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_313),
.B(n_223),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_262),
.B(n_256),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_316),
.B(n_271),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_318),
.B(n_305),
.Y(n_356)
);

NAND3xp33_ASAP7_75t_L g374 ( 
.A(n_322),
.B(n_324),
.C(n_330),
.Y(n_374)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_276),
.Y(n_323)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_323),
.Y(n_365)
);

AOI21x1_ASAP7_75t_L g360 ( 
.A1(n_325),
.A2(n_320),
.B(n_298),
.Y(n_360)
);

INVx3_ASAP7_75t_L g326 ( 
.A(n_306),
.Y(n_326)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_326),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_291),
.A2(n_209),
.B1(n_266),
.B2(n_269),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_327),
.A2(n_346),
.B(n_350),
.Y(n_362)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_276),
.Y(n_328)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_328),
.Y(n_378)
);

AOI22xp33_ASAP7_75t_SL g329 ( 
.A1(n_317),
.A2(n_209),
.B1(n_250),
.B2(n_270),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_329),
.A2(n_336),
.B1(n_338),
.B2(n_341),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_292),
.B(n_207),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_275),
.B(n_220),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_331),
.B(n_349),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_332),
.A2(n_343),
.B1(n_345),
.B2(n_348),
.Y(n_364)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_304),
.Y(n_334)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_334),
.Y(n_384)
);

INVx5_ASAP7_75t_L g335 ( 
.A(n_314),
.Y(n_335)
);

HB1xp67_ASAP7_75t_L g387 ( 
.A(n_335),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_294),
.A2(n_209),
.B1(n_264),
.B2(n_230),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_286),
.A2(n_212),
.B(n_231),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_337),
.A2(n_347),
.B(n_281),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_282),
.A2(n_215),
.B1(n_217),
.B2(n_219),
.Y(n_338)
);

OR2x2_ASAP7_75t_L g381 ( 
.A(n_339),
.B(n_304),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_314),
.Y(n_340)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_340),
.Y(n_382)
);

AOI22x1_ASAP7_75t_L g341 ( 
.A1(n_290),
.A2(n_224),
.B1(n_234),
.B2(n_283),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_278),
.Y(n_342)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_342),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_282),
.A2(n_277),
.B1(n_316),
.B2(n_300),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_277),
.A2(n_299),
.B1(n_284),
.B2(n_303),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_296),
.A2(n_273),
.B(n_289),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_317),
.A2(n_318),
.B(n_309),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_274),
.A2(n_299),
.B1(n_297),
.B2(n_285),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_348),
.A2(n_353),
.B1(n_295),
.B2(n_315),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_307),
.B(n_301),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_SL g350 ( 
.A1(n_285),
.A2(n_271),
.B(n_311),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_278),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_351),
.B(n_352),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_307),
.B(n_319),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_271),
.A2(n_305),
.B1(n_310),
.B2(n_312),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_293),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_354),
.B(n_358),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_355),
.B(n_357),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_356),
.B(n_272),
.C(n_287),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_319),
.B(n_305),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_SL g400 ( 
.A1(n_360),
.A2(n_371),
.B(n_373),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_364),
.B(n_367),
.Y(n_393)
);

AO21x2_ASAP7_75t_L g366 ( 
.A1(n_336),
.A2(n_320),
.B(n_298),
.Y(n_366)
);

BUFx4f_ASAP7_75t_SL g404 ( 
.A(n_366),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_SL g406 ( 
.A(n_367),
.B(n_379),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_343),
.A2(n_280),
.B1(n_306),
.B2(n_295),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_368),
.A2(n_385),
.B1(n_342),
.B2(n_354),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_332),
.A2(n_280),
.B1(n_304),
.B2(n_315),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_370),
.A2(n_337),
.B1(n_323),
.B2(n_328),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_L g371 ( 
.A1(n_344),
.A2(n_302),
.B(n_281),
.Y(n_371)
);

BUFx24_ASAP7_75t_SL g375 ( 
.A(n_346),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_375),
.B(n_324),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_350),
.B(n_288),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_SL g403 ( 
.A(n_377),
.B(n_330),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_357),
.B(n_288),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_380),
.B(n_386),
.C(n_388),
.Y(n_408)
);

CKINVDCx14_ASAP7_75t_R g414 ( 
.A(n_381),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_345),
.A2(n_302),
.B1(n_272),
.B2(n_287),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_356),
.B(n_353),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_347),
.B(n_355),
.C(n_321),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_389),
.A2(n_393),
.B1(n_370),
.B2(n_366),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_L g390 ( 
.A1(n_360),
.A2(n_373),
.B(n_374),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_390),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_SL g424 ( 
.A(n_391),
.B(n_407),
.Y(n_424)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_392),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_362),
.A2(n_325),
.B(n_341),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g426 ( 
.A1(n_394),
.A2(n_395),
.B(n_396),
.Y(n_426)
);

AOI22xp33_ASAP7_75t_SL g395 ( 
.A1(n_361),
.A2(n_334),
.B1(n_333),
.B2(n_341),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_SL g396 ( 
.A1(n_362),
.A2(n_322),
.B(n_358),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_376),
.B(n_352),
.Y(n_397)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_397),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_386),
.B(n_372),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_398),
.B(n_405),
.Y(n_417)
);

AOI21xp5_ASAP7_75t_L g399 ( 
.A1(n_364),
.A2(n_327),
.B(n_321),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_399),
.B(n_413),
.Y(n_430)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_365),
.Y(n_401)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_401),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_369),
.B(n_331),
.Y(n_402)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_402),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_403),
.B(n_410),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_372),
.B(n_349),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_376),
.B(n_338),
.Y(n_407)
);

INVx4_ASAP7_75t_L g409 ( 
.A(n_363),
.Y(n_409)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_409),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_SL g410 ( 
.A1(n_371),
.A2(n_351),
.B(n_326),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_379),
.B(n_340),
.C(n_335),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_411),
.B(n_380),
.C(n_384),
.Y(n_416)
);

CKINVDCx14_ASAP7_75t_R g412 ( 
.A(n_359),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_412),
.Y(n_432)
);

CKINVDCx14_ASAP7_75t_R g413 ( 
.A(n_385),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_393),
.A2(n_366),
.B1(n_368),
.B2(n_381),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_415),
.A2(n_429),
.B1(n_404),
.B2(n_414),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_416),
.B(n_421),
.C(n_434),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_398),
.B(n_388),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_419),
.B(n_427),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_408),
.B(n_378),
.C(n_383),
.Y(n_421)
);

HB1xp67_ASAP7_75t_L g437 ( 
.A(n_423),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_SL g427 ( 
.A(n_408),
.B(n_384),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_399),
.A2(n_366),
.B1(n_382),
.B2(n_387),
.Y(n_429)
);

NOR3xp33_ASAP7_75t_SL g431 ( 
.A(n_391),
.B(n_366),
.C(n_363),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_431),
.B(n_410),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_SL g434 ( 
.A(n_406),
.B(n_340),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_397),
.B(n_402),
.Y(n_436)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_436),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g455 ( 
.A1(n_439),
.A2(n_441),
.B1(n_449),
.B2(n_450),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_432),
.B(n_403),
.Y(n_440)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_440),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_418),
.A2(n_394),
.B1(n_390),
.B2(n_414),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_425),
.B(n_407),
.Y(n_442)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_442),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_L g444 ( 
.A1(n_426),
.A2(n_400),
.B(n_396),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_444),
.B(n_447),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_425),
.B(n_392),
.Y(n_446)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_446),
.Y(n_465)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_422),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_420),
.B(n_411),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g464 ( 
.A(n_448),
.Y(n_464)
);

OR2x2_ASAP7_75t_L g450 ( 
.A(n_433),
.B(n_389),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_427),
.B(n_406),
.C(n_405),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_451),
.B(n_453),
.Y(n_461)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_422),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_452),
.B(n_409),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_424),
.B(n_401),
.Y(n_453)
);

XOR2x2_ASAP7_75t_L g454 ( 
.A(n_443),
.B(n_426),
.Y(n_454)
);

INVxp67_ASAP7_75t_L g471 ( 
.A(n_454),
.Y(n_471)
);

A2O1A1O1Ixp25_ASAP7_75t_L g456 ( 
.A1(n_444),
.A2(n_436),
.B(n_430),
.C(n_428),
.D(n_434),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_L g467 ( 
.A1(n_456),
.A2(n_428),
.B(n_450),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_443),
.B(n_419),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_457),
.B(n_463),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_448),
.B(n_421),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_462),
.B(n_466),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_438),
.B(n_417),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_L g480 ( 
.A1(n_467),
.A2(n_468),
.B(n_445),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_L g468 ( 
.A1(n_461),
.A2(n_451),
.B(n_416),
.Y(n_468)
);

BUFx24_ASAP7_75t_SL g469 ( 
.A(n_459),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_SL g483 ( 
.A(n_469),
.B(n_470),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_457),
.B(n_438),
.C(n_417),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_454),
.B(n_441),
.C(n_437),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_472),
.B(n_473),
.C(n_475),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_464),
.B(n_463),
.C(n_455),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_458),
.B(n_445),
.C(n_418),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_471),
.B(n_456),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_477),
.B(n_484),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_SL g478 ( 
.A1(n_471),
.A2(n_458),
.B(n_460),
.Y(n_478)
);

AOI21xp33_ASAP7_75t_L g485 ( 
.A1(n_478),
.A2(n_480),
.B(n_439),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_474),
.A2(n_460),
.B1(n_465),
.B2(n_446),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_481),
.A2(n_447),
.B1(n_415),
.B2(n_435),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_476),
.B(n_430),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_482),
.B(n_479),
.Y(n_490)
);

AOI22xp33_ASAP7_75t_L g484 ( 
.A1(n_475),
.A2(n_404),
.B1(n_465),
.B2(n_442),
.Y(n_484)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_485),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_479),
.B(n_423),
.C(n_429),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_486),
.B(n_487),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_483),
.B(n_435),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_489),
.B(n_490),
.Y(n_494)
);

HB1xp67_ASAP7_75t_L g492 ( 
.A(n_488),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_492),
.B(n_486),
.Y(n_495)
);

OAI321xp33_ASAP7_75t_L g497 ( 
.A1(n_495),
.A2(n_496),
.A3(n_493),
.B1(n_494),
.B2(n_431),
.C(n_482),
.Y(n_497)
);

OAI21xp5_ASAP7_75t_SL g496 ( 
.A1(n_491),
.A2(n_477),
.B(n_484),
.Y(n_496)
);

BUFx24_ASAP7_75t_SL g498 ( 
.A(n_497),
.Y(n_498)
);

BUFx24_ASAP7_75t_SL g499 ( 
.A(n_498),
.Y(n_499)
);

FAx1_ASAP7_75t_SL g500 ( 
.A(n_499),
.B(n_404),
.CI(n_396),
.CON(n_500),
.SN(n_500)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_500),
.B(n_400),
.C(n_404),
.Y(n_501)
);


endmodule