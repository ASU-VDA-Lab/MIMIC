module fake_jpeg_20598_n_167 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_167);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_167;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_17),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_31),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_42),
.Y(n_52)
);

INVx6_ASAP7_75t_SL g53 ( 
.A(n_44),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

BUFx24_ASAP7_75t_L g55 ( 
.A(n_3),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_40),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_5),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_14),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_15),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_4),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_8),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_11),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_39),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_5),
.Y(n_65)
);

BUFx12_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_38),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_9),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_11),
.Y(n_69)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_12),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_18),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_7),
.Y(n_74)
);

BUFx16f_ASAP7_75t_L g75 ( 
.A(n_9),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_28),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_54),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_79),
.Y(n_87)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_81),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_83),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_77),
.B(n_57),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_85),
.A2(n_89),
.B1(n_66),
.B2(n_47),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_82),
.A2(n_70),
.B1(n_55),
.B2(n_74),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_83),
.A2(n_63),
.B1(n_53),
.B2(n_76),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_91),
.B(n_59),
.Y(n_96)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_92),
.Y(n_97)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_94),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_96),
.A2(n_62),
.B1(n_1),
.B2(n_3),
.Y(n_122)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_86),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_98),
.Y(n_124)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_99),
.Y(n_110)
);

BUFx2_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_100),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_101),
.Y(n_119)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_93),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_105),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_69),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_103),
.B(n_104),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_88),
.B(n_46),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_89),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_65),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_107),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_68),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_101),
.A2(n_50),
.B(n_48),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_109),
.A2(n_117),
.B(n_120),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_97),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_111),
.B(n_112),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_95),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_97),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_113),
.B(n_123),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_98),
.A2(n_84),
.B1(n_73),
.B2(n_52),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_114),
.A2(n_118),
.B1(n_0),
.B2(n_1),
.Y(n_135)
);

MAJx3_ASAP7_75t_L g115 ( 
.A(n_100),
.B(n_66),
.C(n_75),
.Y(n_115)
);

HAxp5_ASAP7_75t_SL g127 ( 
.A(n_115),
.B(n_59),
.CON(n_127),
.SN(n_127)
);

NAND2x1_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_47),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_105),
.A2(n_84),
.B1(n_64),
.B2(n_56),
.Y(n_118)
);

OAI21xp33_ASAP7_75t_L g120 ( 
.A1(n_105),
.A2(n_67),
.B(n_71),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_122),
.A2(n_125),
.B1(n_110),
.B2(n_108),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_95),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_127),
.A2(n_134),
.B1(n_135),
.B2(n_137),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_121),
.Y(n_128)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_128),
.Y(n_146)
);

OAI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_119),
.A2(n_73),
.B1(n_72),
.B2(n_49),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_130),
.A2(n_131),
.B1(n_0),
.B2(n_4),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_120),
.B(n_75),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_132),
.B(n_136),
.C(n_139),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_119),
.A2(n_30),
.B(n_43),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_111),
.B(n_60),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_116),
.A2(n_72),
.B1(n_32),
.B2(n_33),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_115),
.A2(n_60),
.B1(n_49),
.B2(n_51),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_138),
.A2(n_10),
.B1(n_13),
.B2(n_20),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_117),
.B(n_24),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_141),
.A2(n_144),
.B1(n_145),
.B2(n_147),
.Y(n_151)
);

A2O1A1Ixp33_ASAP7_75t_L g142 ( 
.A1(n_127),
.A2(n_6),
.B(n_7),
.C(n_8),
.Y(n_142)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_142),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_126),
.A2(n_129),
.B1(n_133),
.B2(n_135),
.Y(n_144)
);

OA21x2_ASAP7_75t_L g145 ( 
.A1(n_138),
.A2(n_124),
.B(n_35),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_137),
.A2(n_124),
.B1(n_10),
.B2(n_6),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g153 ( 
.A(n_148),
.B(n_21),
.Y(n_153)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_146),
.Y(n_149)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_149),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_140),
.B(n_139),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_152),
.B(n_153),
.C(n_145),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_154),
.A2(n_150),
.B(n_142),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_156),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_157),
.A2(n_150),
.B(n_155),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_145),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_143),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_151),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_161),
.B(n_146),
.Y(n_162)
);

NOR3xp33_ASAP7_75t_SL g163 ( 
.A(n_162),
.B(n_147),
.C(n_23),
.Y(n_163)
);

INVxp33_ASAP7_75t_SL g164 ( 
.A(n_163),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_164),
.A2(n_22),
.B(n_25),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_27),
.C(n_36),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_37),
.Y(n_167)
);


endmodule