module fake_ariane_1453_n_108 (n_8, n_3, n_2, n_11, n_7, n_16, n_5, n_14, n_1, n_0, n_12, n_15, n_6, n_13, n_9, n_17, n_4, n_10, n_108);

input n_8;
input n_3;
input n_2;
input n_11;
input n_7;
input n_16;
input n_5;
input n_14;
input n_1;
input n_0;
input n_12;
input n_15;
input n_6;
input n_13;
input n_9;
input n_17;
input n_4;
input n_10;

output n_108;

wire n_83;
wire n_56;
wire n_60;
wire n_64;
wire n_90;
wire n_38;
wire n_47;
wire n_18;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_34;
wire n_69;
wire n_95;
wire n_92;
wire n_98;
wire n_74;
wire n_33;
wire n_19;
wire n_40;
wire n_106;
wire n_53;
wire n_21;
wire n_66;
wire n_71;
wire n_24;
wire n_96;
wire n_49;
wire n_20;
wire n_100;
wire n_50;
wire n_62;
wire n_51;
wire n_76;
wire n_103;
wire n_79;
wire n_26;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_107;
wire n_72;
wire n_105;
wire n_44;
wire n_30;
wire n_82;
wire n_31;
wire n_42;
wire n_57;
wire n_70;
wire n_85;
wire n_48;
wire n_94;
wire n_101;
wire n_32;
wire n_37;
wire n_58;
wire n_65;
wire n_45;
wire n_52;
wire n_73;
wire n_77;
wire n_93;
wire n_23;
wire n_61;
wire n_102;
wire n_22;
wire n_43;
wire n_81;
wire n_87;
wire n_27;
wire n_29;
wire n_41;
wire n_55;
wire n_28;
wire n_80;
wire n_97;
wire n_88;
wire n_68;
wire n_104;
wire n_78;
wire n_39;
wire n_59;
wire n_63;
wire n_99;
wire n_35;
wire n_54;
wire n_25;

INVxp67_ASAP7_75t_SL g18 ( 
.A(n_17),
.Y(n_18)
);

HB1xp67_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

NOR2xp67_ASAP7_75t_L g22 ( 
.A(n_11),
.B(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVxp67_ASAP7_75t_SL g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx2_ASAP7_75t_SL g34 ( 
.A(n_20),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_21),
.B(n_0),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_27),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_21),
.B(n_3),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

NAND2xp33_ASAP7_75t_SL g39 ( 
.A(n_27),
.B(n_4),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_19),
.B(n_5),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_25),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

OAI221xp5_ASAP7_75t_L g46 ( 
.A1(n_42),
.A2(n_43),
.B1(n_41),
.B2(n_37),
.C(n_35),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

NAND2x1p5_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_22),
.Y(n_48)
);

AO22x2_ASAP7_75t_L g49 ( 
.A1(n_35),
.A2(n_30),
.B1(n_29),
.B2(n_26),
.Y(n_49)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_24),
.Y(n_50)
);

AND2x4_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_18),
.Y(n_51)
);

AO22x2_ASAP7_75t_L g52 ( 
.A1(n_34),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_34),
.Y(n_55)
);

CKINVDCx5p33_ASAP7_75t_R g56 ( 
.A(n_51),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_46),
.A2(n_39),
.B1(n_36),
.B2(n_32),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_32),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

O2A1O1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_58),
.A2(n_53),
.B(n_44),
.C(n_46),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_59),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_55),
.Y(n_62)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_44),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_59),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_49),
.Y(n_65)
);

OA21x2_ASAP7_75t_L g66 ( 
.A1(n_54),
.A2(n_52),
.B(n_49),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_65),
.B(n_54),
.Y(n_68)
);

AND2x2_ASAP7_75t_SL g69 ( 
.A(n_66),
.B(n_28),
.Y(n_69)
);

AND2x4_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_9),
.Y(n_70)
);

AND2x4_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_10),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_70),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_70),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_67),
.B(n_63),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_73),
.Y(n_75)
);

AO21x2_ASAP7_75t_L g76 ( 
.A1(n_72),
.A2(n_64),
.B(n_71),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_73),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_74),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_77),
.B(n_78),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_78),
.B(n_71),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_77),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_75),
.B(n_67),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_75),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_79),
.B(n_82),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_76),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_81),
.B(n_76),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_83),
.A2(n_69),
.B1(n_68),
.B2(n_36),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_76),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_79),
.B(n_70),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_84),
.B(n_71),
.Y(n_90)
);

NOR3xp33_ASAP7_75t_L g91 ( 
.A(n_86),
.B(n_71),
.C(n_70),
.Y(n_91)
);

OAI32xp33_ASAP7_75t_L g92 ( 
.A1(n_87),
.A2(n_48),
.A3(n_65),
.B1(n_52),
.B2(n_63),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_89),
.B(n_71),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_90),
.B(n_85),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_93),
.Y(n_95)
);

AOI22x1_ASAP7_75t_L g96 ( 
.A1(n_95),
.A2(n_70),
.B1(n_48),
.B2(n_88),
.Y(n_96)
);

NOR3x1_ASAP7_75t_L g97 ( 
.A(n_94),
.B(n_10),
.C(n_64),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_95),
.B(n_91),
.Y(n_98)
);

NAND4xp25_ASAP7_75t_L g99 ( 
.A(n_97),
.B(n_92),
.C(n_62),
.D(n_60),
.Y(n_99)
);

NAND4xp25_ASAP7_75t_L g100 ( 
.A(n_98),
.B(n_60),
.C(n_68),
.D(n_66),
.Y(n_100)
);

NOR2x1_ASAP7_75t_L g101 ( 
.A(n_98),
.B(n_66),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_96),
.A2(n_66),
.B1(n_69),
.B2(n_68),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_101),
.B(n_66),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_102),
.A2(n_69),
.B1(n_28),
.B2(n_61),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_103),
.B(n_100),
.Y(n_105)
);

OAI322xp33_ASAP7_75t_L g106 ( 
.A1(n_104),
.A2(n_14),
.A3(n_28),
.B1(n_33),
.B2(n_99),
.C1(n_36),
.C2(n_21),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_105),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_107),
.A2(n_106),
.B1(n_28),
.B2(n_33),
.Y(n_108)
);


endmodule