module real_aes_8897_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_504;
wire n_455;
wire n_310;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_417;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_505;
wire n_502;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_713;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_719;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g107 ( .A(n_0), .B(n_86), .C(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g435 ( .A(n_0), .Y(n_435) );
A2O1A1Ixp33_ASAP7_75t_L g182 ( .A1(n_1), .A2(n_141), .B(n_146), .C(n_183), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_2), .A2(n_136), .B(n_206), .Y(n_205) );
INVx1_ASAP7_75t_L g453 ( .A(n_3), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_4), .B(n_160), .Y(n_213) );
AOI22xp5_ASAP7_75t_L g713 ( .A1(n_5), .A2(n_15), .B1(n_714), .B2(n_715), .Y(n_713) );
CKINVDCx20_ASAP7_75t_R g715 ( .A(n_5), .Y(n_715) );
AOI21xp33_ASAP7_75t_L g470 ( .A1(n_6), .A2(n_136), .B(n_471), .Y(n_470) );
AND2x6_ASAP7_75t_L g141 ( .A(n_7), .B(n_142), .Y(n_141) );
INVx1_ASAP7_75t_L g170 ( .A(n_8), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_9), .B(n_106), .Y(n_105) );
NOR2xp33_ASAP7_75t_L g436 ( .A(n_9), .B(n_44), .Y(n_436) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_10), .A2(n_248), .B(n_531), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_11), .B(n_151), .Y(n_187) );
INVx1_ASAP7_75t_L g475 ( .A(n_12), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_13), .B(n_150), .Y(n_523) );
INVx1_ASAP7_75t_L g134 ( .A(n_14), .Y(n_134) );
CKINVDCx20_ASAP7_75t_R g714 ( .A(n_15), .Y(n_714) );
INVx1_ASAP7_75t_L g535 ( .A(n_16), .Y(n_535) );
A2O1A1Ixp33_ASAP7_75t_L g195 ( .A1(n_17), .A2(n_171), .B(n_196), .C(n_198), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_18), .B(n_160), .Y(n_199) );
AOI22xp5_ASAP7_75t_L g101 ( .A1(n_19), .A2(n_102), .B1(n_111), .B2(n_725), .Y(n_101) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_20), .B(n_464), .Y(n_514) );
AOI222xp33_ASAP7_75t_L g440 ( .A1(n_21), .A2(n_441), .B1(n_713), .B2(n_716), .C1(n_719), .C2(n_723), .Y(n_440) );
NAND2xp5_ASAP7_75t_SL g501 ( .A(n_22), .B(n_136), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_23), .B(n_256), .Y(n_255) );
A2O1A1Ixp33_ASAP7_75t_L g149 ( .A1(n_24), .A2(n_150), .B(n_152), .C(n_156), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_25), .B(n_160), .Y(n_467) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_26), .B(n_151), .Y(n_220) );
A2O1A1Ixp33_ASAP7_75t_L g533 ( .A1(n_27), .A2(n_154), .B(n_198), .C(n_534), .Y(n_533) );
NAND2xp5_ASAP7_75t_SL g232 ( .A(n_28), .B(n_151), .Y(n_232) );
CKINVDCx16_ASAP7_75t_R g216 ( .A(n_29), .Y(n_216) );
INVx1_ASAP7_75t_L g230 ( .A(n_30), .Y(n_230) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_31), .Y(n_140) );
CKINVDCx20_ASAP7_75t_R g180 ( .A(n_32), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_33), .B(n_151), .Y(n_454) );
INVx1_ASAP7_75t_L g253 ( .A(n_34), .Y(n_253) );
INVx1_ASAP7_75t_L g488 ( .A(n_35), .Y(n_488) );
INVx2_ASAP7_75t_L g139 ( .A(n_36), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g190 ( .A(n_37), .Y(n_190) );
A2O1A1Ixp33_ASAP7_75t_L g208 ( .A1(n_38), .A2(n_150), .B(n_209), .C(n_211), .Y(n_208) );
INVxp67_ASAP7_75t_L g254 ( .A(n_39), .Y(n_254) );
CKINVDCx14_ASAP7_75t_R g207 ( .A(n_40), .Y(n_207) );
A2O1A1Ixp33_ASAP7_75t_L g228 ( .A1(n_41), .A2(n_146), .B(n_229), .C(n_235), .Y(n_228) );
A2O1A1Ixp33_ASAP7_75t_L g502 ( .A1(n_42), .A2(n_141), .B(n_146), .C(n_503), .Y(n_502) );
OAI22xp5_ASAP7_75t_SL g118 ( .A1(n_43), .A2(n_90), .B1(n_119), .B2(n_120), .Y(n_118) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_43), .Y(n_120) );
INVx1_ASAP7_75t_L g106 ( .A(n_44), .Y(n_106) );
INVx1_ASAP7_75t_L g487 ( .A(n_45), .Y(n_487) );
A2O1A1Ixp33_ASAP7_75t_L g167 ( .A1(n_46), .A2(n_168), .B(n_169), .C(n_172), .Y(n_167) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_47), .B(n_151), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_48), .B(n_438), .Y(n_437) );
CKINVDCx20_ASAP7_75t_R g237 ( .A(n_49), .Y(n_237) );
CKINVDCx20_ASAP7_75t_R g250 ( .A(n_50), .Y(n_250) );
INVx1_ASAP7_75t_L g144 ( .A(n_51), .Y(n_144) );
CKINVDCx16_ASAP7_75t_R g489 ( .A(n_52), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_53), .B(n_136), .Y(n_525) );
AOI22xp5_ASAP7_75t_L g485 ( .A1(n_54), .A2(n_146), .B1(n_156), .B2(n_486), .Y(n_485) );
CKINVDCx20_ASAP7_75t_R g507 ( .A(n_55), .Y(n_507) );
CKINVDCx16_ASAP7_75t_R g450 ( .A(n_56), .Y(n_450) );
CKINVDCx14_ASAP7_75t_R g166 ( .A(n_57), .Y(n_166) );
A2O1A1Ixp33_ASAP7_75t_L g473 ( .A1(n_58), .A2(n_168), .B(n_211), .C(n_474), .Y(n_473) );
CKINVDCx20_ASAP7_75t_R g516 ( .A(n_59), .Y(n_516) );
INVx1_ASAP7_75t_L g472 ( .A(n_60), .Y(n_472) );
INVx1_ASAP7_75t_L g142 ( .A(n_61), .Y(n_142) );
INVx1_ASAP7_75t_L g133 ( .A(n_62), .Y(n_133) );
INVx1_ASAP7_75t_SL g210 ( .A(n_63), .Y(n_210) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_64), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_65), .B(n_160), .Y(n_159) );
INVx1_ASAP7_75t_L g219 ( .A(n_66), .Y(n_219) );
A2O1A1Ixp33_ASAP7_75t_SL g463 ( .A1(n_67), .A2(n_211), .B(n_464), .C(n_465), .Y(n_463) );
INVxp67_ASAP7_75t_L g466 ( .A(n_68), .Y(n_466) );
INVx1_ASAP7_75t_L g110 ( .A(n_69), .Y(n_110) );
AOI21xp5_ASAP7_75t_L g164 ( .A1(n_70), .A2(n_136), .B(n_165), .Y(n_164) );
CKINVDCx20_ASAP7_75t_R g223 ( .A(n_71), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_72), .A2(n_136), .B(n_193), .Y(n_192) );
CKINVDCx20_ASAP7_75t_R g491 ( .A(n_73), .Y(n_491) );
INVx1_ASAP7_75t_L g510 ( .A(n_74), .Y(n_510) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_75), .A2(n_248), .B(n_249), .Y(n_247) );
INVx1_ASAP7_75t_L g194 ( .A(n_76), .Y(n_194) );
CKINVDCx16_ASAP7_75t_R g227 ( .A(n_77), .Y(n_227) );
A2O1A1Ixp33_ASAP7_75t_L g511 ( .A1(n_78), .A2(n_141), .B(n_146), .C(n_512), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g135 ( .A1(n_79), .A2(n_136), .B(n_143), .Y(n_135) );
INVx1_ASAP7_75t_L g197 ( .A(n_80), .Y(n_197) );
NAND2xp5_ASAP7_75t_SL g504 ( .A(n_81), .B(n_231), .Y(n_504) );
INVx2_ASAP7_75t_L g131 ( .A(n_82), .Y(n_131) );
INVx1_ASAP7_75t_L g184 ( .A(n_83), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_84), .B(n_464), .Y(n_505) );
A2O1A1Ixp33_ASAP7_75t_L g451 ( .A1(n_85), .A2(n_141), .B(n_146), .C(n_452), .Y(n_451) );
OR2x2_ASAP7_75t_L g432 ( .A(n_86), .B(n_433), .Y(n_432) );
INVx2_ASAP7_75t_L g711 ( .A(n_86), .Y(n_711) );
OR2x2_ASAP7_75t_L g712 ( .A(n_86), .B(n_434), .Y(n_712) );
A2O1A1Ixp33_ASAP7_75t_L g217 ( .A1(n_87), .A2(n_146), .B(n_218), .C(n_221), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_88), .B(n_163), .Y(n_476) );
CKINVDCx20_ASAP7_75t_R g457 ( .A(n_89), .Y(n_457) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_90), .Y(n_119) );
A2O1A1Ixp33_ASAP7_75t_L g520 ( .A1(n_91), .A2(n_141), .B(n_146), .C(n_521), .Y(n_520) );
CKINVDCx20_ASAP7_75t_R g527 ( .A(n_92), .Y(n_527) );
INVx1_ASAP7_75t_L g462 ( .A(n_93), .Y(n_462) );
CKINVDCx16_ASAP7_75t_R g532 ( .A(n_94), .Y(n_532) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_95), .B(n_231), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_96), .B(n_129), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_97), .B(n_129), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_98), .B(n_110), .Y(n_109) );
INVx2_ASAP7_75t_L g153 ( .A(n_99), .Y(n_153) );
AOI21xp5_ASAP7_75t_L g460 ( .A1(n_100), .A2(n_136), .B(n_461), .Y(n_460) );
INVx1_ASAP7_75t_SL g102 ( .A(n_103), .Y(n_102) );
BUFx4f_ASAP7_75t_SL g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_SL g726 ( .A(n_104), .Y(n_726) );
OR2x2_ASAP7_75t_L g104 ( .A(n_105), .B(n_107), .Y(n_104) );
INVx1_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
AO21x2_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_116), .B(n_439), .Y(n_111) );
INVx1_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
BUFx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
INVx1_ASAP7_75t_L g724 ( .A(n_114), .Y(n_724) );
INVx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
OAI21xp5_ASAP7_75t_SL g116 ( .A1(n_117), .A2(n_429), .B(n_437), .Y(n_116) );
AOI22xp5_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_121), .B1(n_427), .B2(n_428), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g427 ( .A(n_118), .Y(n_427) );
OAI22xp5_ASAP7_75t_L g719 ( .A1(n_121), .A2(n_710), .B1(n_720), .B2(n_721), .Y(n_719) );
BUFx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx1_ASAP7_75t_L g428 ( .A(n_122), .Y(n_428) );
AND2x2_ASAP7_75t_L g122 ( .A(n_123), .B(n_353), .Y(n_122) );
NOR4xp25_ASAP7_75t_L g123 ( .A(n_124), .B(n_295), .C(n_325), .D(n_335), .Y(n_123) );
OAI211xp5_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_200), .B(n_258), .C(n_285), .Y(n_124) );
OAI222xp33_ASAP7_75t_L g380 ( .A1(n_125), .A2(n_300), .B1(n_381), .B2(n_382), .C1(n_383), .C2(n_384), .Y(n_380) );
OR2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_175), .Y(n_125) );
AOI33xp33_ASAP7_75t_L g306 ( .A1(n_126), .A2(n_293), .A3(n_294), .B1(n_307), .B2(n_312), .B3(n_314), .Y(n_306) );
OAI211xp5_ASAP7_75t_SL g363 ( .A1(n_126), .A2(n_364), .B(n_366), .C(n_368), .Y(n_363) );
OR2x2_ASAP7_75t_L g379 ( .A(n_126), .B(n_365), .Y(n_379) );
INVx1_ASAP7_75t_L g412 ( .A(n_126), .Y(n_412) );
OR2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_162), .Y(n_126) );
INVx2_ASAP7_75t_L g289 ( .A(n_127), .Y(n_289) );
AND2x2_ASAP7_75t_L g305 ( .A(n_127), .B(n_191), .Y(n_305) );
HB1xp67_ASAP7_75t_L g340 ( .A(n_127), .Y(n_340) );
AND2x2_ASAP7_75t_L g369 ( .A(n_127), .B(n_162), .Y(n_369) );
OA21x2_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_135), .B(n_159), .Y(n_127) );
OA21x2_ASAP7_75t_L g191 ( .A1(n_128), .A2(n_192), .B(n_199), .Y(n_191) );
OA21x2_ASAP7_75t_L g204 ( .A1(n_128), .A2(n_205), .B(n_213), .Y(n_204) );
HB1xp67_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx4_ASAP7_75t_L g161 ( .A(n_129), .Y(n_161) );
OA21x2_ASAP7_75t_L g459 ( .A1(n_129), .A2(n_460), .B(n_467), .Y(n_459) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx1_ASAP7_75t_L g246 ( .A(n_130), .Y(n_246) );
AND2x2_ASAP7_75t_L g130 ( .A(n_131), .B(n_132), .Y(n_130) );
AND2x2_ASAP7_75t_SL g163 ( .A(n_131), .B(n_132), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_133), .B(n_134), .Y(n_132) );
BUFx2_ASAP7_75t_L g248 ( .A(n_136), .Y(n_248) );
AND2x4_ASAP7_75t_L g136 ( .A(n_137), .B(n_141), .Y(n_136) );
NAND2x1p5_ASAP7_75t_L g181 ( .A(n_137), .B(n_141), .Y(n_181) );
AND2x2_ASAP7_75t_L g137 ( .A(n_138), .B(n_140), .Y(n_137) );
INVx1_ASAP7_75t_L g234 ( .A(n_138), .Y(n_234) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx2_ASAP7_75t_L g147 ( .A(n_139), .Y(n_147) );
INVx1_ASAP7_75t_L g157 ( .A(n_139), .Y(n_157) );
INVx1_ASAP7_75t_L g148 ( .A(n_140), .Y(n_148) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_140), .Y(n_151) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_140), .Y(n_155) );
INVx3_ASAP7_75t_L g171 ( .A(n_140), .Y(n_171) );
INVx1_ASAP7_75t_L g464 ( .A(n_140), .Y(n_464) );
INVx4_ASAP7_75t_SL g158 ( .A(n_141), .Y(n_158) );
BUFx3_ASAP7_75t_L g235 ( .A(n_141), .Y(n_235) );
O2A1O1Ixp33_ASAP7_75t_SL g143 ( .A1(n_144), .A2(n_145), .B(n_149), .C(n_158), .Y(n_143) );
O2A1O1Ixp33_ASAP7_75t_SL g165 ( .A1(n_145), .A2(n_158), .B(n_166), .C(n_167), .Y(n_165) );
O2A1O1Ixp33_ASAP7_75t_SL g193 ( .A1(n_145), .A2(n_158), .B(n_194), .C(n_195), .Y(n_193) );
O2A1O1Ixp33_ASAP7_75t_L g206 ( .A1(n_145), .A2(n_158), .B(n_207), .C(n_208), .Y(n_206) );
O2A1O1Ixp33_ASAP7_75t_SL g249 ( .A1(n_145), .A2(n_158), .B(n_250), .C(n_251), .Y(n_249) );
O2A1O1Ixp33_ASAP7_75t_L g461 ( .A1(n_145), .A2(n_158), .B(n_462), .C(n_463), .Y(n_461) );
O2A1O1Ixp33_ASAP7_75t_L g471 ( .A1(n_145), .A2(n_158), .B(n_472), .C(n_473), .Y(n_471) );
O2A1O1Ixp33_ASAP7_75t_L g531 ( .A1(n_145), .A2(n_158), .B(n_532), .C(n_533), .Y(n_531) );
INVx5_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AND2x6_ASAP7_75t_L g146 ( .A(n_147), .B(n_148), .Y(n_146) );
BUFx3_ASAP7_75t_L g173 ( .A(n_147), .Y(n_173) );
BUFx6f_ASAP7_75t_L g212 ( .A(n_147), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_150), .B(n_210), .Y(n_209) );
INVx4_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g168 ( .A(n_151), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g152 ( .A(n_153), .B(n_154), .Y(n_152) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_154), .B(n_197), .Y(n_196) );
OAI22xp33_ASAP7_75t_L g252 ( .A1(n_154), .A2(n_231), .B1(n_253), .B2(n_254), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g534 ( .A(n_154), .B(n_535), .Y(n_534) );
INVx4_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx2_ASAP7_75t_L g186 ( .A(n_155), .Y(n_186) );
OAI22xp5_ASAP7_75t_SL g486 ( .A1(n_155), .A2(n_186), .B1(n_487), .B2(n_488), .Y(n_486) );
INVx2_ASAP7_75t_L g455 ( .A(n_156), .Y(n_455) );
INVx3_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx1_ASAP7_75t_L g221 ( .A(n_158), .Y(n_221) );
OAI22xp33_ASAP7_75t_L g484 ( .A1(n_158), .A2(n_181), .B1(n_485), .B2(n_489), .Y(n_484) );
OA21x2_ASAP7_75t_L g469 ( .A1(n_160), .A2(n_470), .B(n_476), .Y(n_469) );
INVx3_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_161), .B(n_190), .Y(n_189) );
AO21x2_ASAP7_75t_L g214 ( .A1(n_161), .A2(n_215), .B(n_222), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_161), .B(n_237), .Y(n_236) );
NOR2xp33_ASAP7_75t_SL g506 ( .A(n_161), .B(n_507), .Y(n_506) );
INVx2_ASAP7_75t_L g269 ( .A(n_162), .Y(n_269) );
BUFx3_ASAP7_75t_L g277 ( .A(n_162), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_162), .B(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g288 ( .A(n_162), .B(n_289), .Y(n_288) );
NOR2xp33_ASAP7_75t_L g317 ( .A(n_162), .B(n_176), .Y(n_317) );
AND2x2_ASAP7_75t_L g386 ( .A(n_162), .B(n_320), .Y(n_386) );
OA21x2_ASAP7_75t_L g162 ( .A1(n_163), .A2(n_164), .B(n_174), .Y(n_162) );
INVx1_ASAP7_75t_L g178 ( .A(n_163), .Y(n_178) );
INVx2_ASAP7_75t_L g224 ( .A(n_163), .Y(n_224) );
O2A1O1Ixp33_ASAP7_75t_L g226 ( .A1(n_163), .A2(n_181), .B(n_227), .C(n_228), .Y(n_226) );
OA21x2_ASAP7_75t_L g529 ( .A1(n_163), .A2(n_530), .B(n_536), .Y(n_529) );
NOR2xp33_ASAP7_75t_L g169 ( .A(n_170), .B(n_171), .Y(n_169) );
INVx5_ASAP7_75t_L g231 ( .A(n_171), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_171), .B(n_466), .Y(n_465) );
NOR2xp33_ASAP7_75t_L g474 ( .A(n_171), .B(n_475), .Y(n_474) );
INVx2_ASAP7_75t_L g188 ( .A(n_172), .Y(n_188) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx1_ASAP7_75t_L g198 ( .A(n_173), .Y(n_198) );
INVx2_ASAP7_75t_SL g280 ( .A(n_175), .Y(n_280) );
OR2x2_ASAP7_75t_L g175 ( .A(n_176), .B(n_191), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_176), .B(n_269), .Y(n_268) );
INVx1_ASAP7_75t_L g322 ( .A(n_176), .Y(n_322) );
AND2x2_ASAP7_75t_L g333 ( .A(n_176), .B(n_289), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_176), .B(n_318), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_176), .B(n_320), .Y(n_365) );
AND2x2_ASAP7_75t_L g424 ( .A(n_176), .B(n_369), .Y(n_424) );
INVx4_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
AND2x2_ASAP7_75t_L g294 ( .A(n_177), .B(n_191), .Y(n_294) );
AND2x2_ASAP7_75t_L g304 ( .A(n_177), .B(n_305), .Y(n_304) );
BUFx3_ASAP7_75t_L g326 ( .A(n_177), .Y(n_326) );
AND3x2_ASAP7_75t_L g385 ( .A(n_177), .B(n_386), .C(n_387), .Y(n_385) );
AO21x2_ASAP7_75t_L g177 ( .A1(n_178), .A2(n_179), .B(n_189), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_178), .B(n_457), .Y(n_456) );
NOR2xp33_ASAP7_75t_L g515 ( .A(n_178), .B(n_516), .Y(n_515) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_178), .B(n_527), .Y(n_526) );
OAI21xp5_ASAP7_75t_L g179 ( .A1(n_180), .A2(n_181), .B(n_182), .Y(n_179) );
OAI21xp5_ASAP7_75t_L g215 ( .A1(n_181), .A2(n_216), .B(n_217), .Y(n_215) );
OAI21xp5_ASAP7_75t_L g449 ( .A1(n_181), .A2(n_450), .B(n_451), .Y(n_449) );
OAI21xp5_ASAP7_75t_L g509 ( .A1(n_181), .A2(n_510), .B(n_511), .Y(n_509) );
O2A1O1Ixp5_ASAP7_75t_L g183 ( .A1(n_184), .A2(n_185), .B(n_187), .C(n_188), .Y(n_183) );
O2A1O1Ixp33_ASAP7_75t_L g218 ( .A1(n_185), .A2(n_188), .B(n_219), .C(n_220), .Y(n_218) );
INVx2_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_188), .A2(n_504), .B(n_505), .Y(n_503) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_188), .A2(n_513), .B(n_514), .Y(n_512) );
HB1xp67_ASAP7_75t_L g276 ( .A(n_191), .Y(n_276) );
INVx1_ASAP7_75t_SL g320 ( .A(n_191), .Y(n_320) );
NAND3xp33_ASAP7_75t_L g332 ( .A(n_191), .B(n_269), .C(n_333), .Y(n_332) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_201), .B(n_238), .Y(n_200) );
A2O1A1Ixp33_ASAP7_75t_L g355 ( .A1(n_201), .A2(n_304), .B(n_356), .C(n_358), .Y(n_355) );
INVx1_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_203), .B(n_225), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_203), .B(n_362), .Y(n_361) );
INVx2_ASAP7_75t_SL g372 ( .A(n_203), .Y(n_372) );
AND2x2_ASAP7_75t_L g393 ( .A(n_203), .B(n_240), .Y(n_393) );
NOR2xp33_ASAP7_75t_L g421 ( .A(n_203), .B(n_302), .Y(n_421) );
AND2x2_ASAP7_75t_L g203 ( .A(n_204), .B(n_214), .Y(n_203) );
AND2x2_ASAP7_75t_L g266 ( .A(n_204), .B(n_257), .Y(n_266) );
INVx2_ASAP7_75t_L g273 ( .A(n_204), .Y(n_273) );
AND2x2_ASAP7_75t_L g293 ( .A(n_204), .B(n_240), .Y(n_293) );
AND2x2_ASAP7_75t_L g343 ( .A(n_204), .B(n_225), .Y(n_343) );
INVx1_ASAP7_75t_L g347 ( .A(n_204), .Y(n_347) );
INVx3_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
HB1xp67_ASAP7_75t_L g524 ( .A(n_212), .Y(n_524) );
INVx2_ASAP7_75t_SL g257 ( .A(n_214), .Y(n_257) );
BUFx2_ASAP7_75t_L g283 ( .A(n_214), .Y(n_283) );
AND2x2_ASAP7_75t_L g410 ( .A(n_214), .B(n_225), .Y(n_410) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_223), .B(n_224), .Y(n_222) );
INVx1_ASAP7_75t_L g256 ( .A(n_224), .Y(n_256) );
AO21x2_ASAP7_75t_L g518 ( .A1(n_224), .A2(n_519), .B(n_526), .Y(n_518) );
INVx3_ASAP7_75t_SL g240 ( .A(n_225), .Y(n_240) );
AND2x2_ASAP7_75t_L g265 ( .A(n_225), .B(n_266), .Y(n_265) );
AND2x4_ASAP7_75t_L g272 ( .A(n_225), .B(n_273), .Y(n_272) );
OR2x2_ASAP7_75t_L g302 ( .A(n_225), .B(n_262), .Y(n_302) );
OR2x2_ASAP7_75t_L g311 ( .A(n_225), .B(n_257), .Y(n_311) );
HB1xp67_ASAP7_75t_L g329 ( .A(n_225), .Y(n_329) );
AND2x2_ASAP7_75t_L g334 ( .A(n_225), .B(n_287), .Y(n_334) );
AND2x2_ASAP7_75t_L g362 ( .A(n_225), .B(n_242), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_225), .B(n_398), .Y(n_397) );
OR2x2_ASAP7_75t_L g400 ( .A(n_225), .B(n_241), .Y(n_400) );
OR2x6_ASAP7_75t_L g225 ( .A(n_226), .B(n_236), .Y(n_225) );
O2A1O1Ixp33_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_231), .B(n_232), .C(n_233), .Y(n_229) );
O2A1O1Ixp33_ASAP7_75t_L g452 ( .A1(n_231), .A2(n_453), .B(n_454), .C(n_455), .Y(n_452) );
INVx2_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
NAND2xp5_ASAP7_75t_SL g251 ( .A(n_234), .B(n_252), .Y(n_251) );
INVx1_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
OR2x2_ASAP7_75t_L g239 ( .A(n_240), .B(n_241), .Y(n_239) );
AND2x2_ASAP7_75t_L g324 ( .A(n_240), .B(n_273), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_240), .B(n_266), .Y(n_352) );
AND2x2_ASAP7_75t_L g370 ( .A(n_240), .B(n_287), .Y(n_370) );
OR2x2_ASAP7_75t_L g241 ( .A(n_242), .B(n_257), .Y(n_241) );
AND2x2_ASAP7_75t_L g271 ( .A(n_242), .B(n_257), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_242), .B(n_300), .Y(n_299) );
BUFx3_ASAP7_75t_L g309 ( .A(n_242), .Y(n_309) );
OR2x2_ASAP7_75t_L g357 ( .A(n_242), .B(n_277), .Y(n_357) );
OA21x2_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_247), .B(n_255), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
AO21x2_ASAP7_75t_L g262 ( .A1(n_244), .A2(n_263), .B(n_264), .Y(n_262) );
AO21x2_ASAP7_75t_L g508 ( .A1(n_244), .A2(n_509), .B(n_515), .Y(n_508) );
INVx1_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
AOI21xp5_ASAP7_75t_SL g500 ( .A1(n_245), .A2(n_501), .B(n_502), .Y(n_500) );
INVx2_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
AO21x2_ASAP7_75t_L g448 ( .A1(n_246), .A2(n_449), .B(n_456), .Y(n_448) );
AO21x2_ASAP7_75t_L g483 ( .A1(n_246), .A2(n_484), .B(n_490), .Y(n_483) );
NOR2xp33_ASAP7_75t_L g490 ( .A(n_246), .B(n_491), .Y(n_490) );
INVx1_ASAP7_75t_L g263 ( .A(n_247), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_255), .Y(n_264) );
AND2x2_ASAP7_75t_L g292 ( .A(n_257), .B(n_262), .Y(n_292) );
INVx1_ASAP7_75t_L g300 ( .A(n_257), .Y(n_300) );
AND2x2_ASAP7_75t_L g395 ( .A(n_257), .B(n_273), .Y(n_395) );
AOI222xp33_ASAP7_75t_L g258 ( .A1(n_259), .A2(n_267), .B1(n_270), .B2(n_274), .C1(n_278), .C2(n_281), .Y(n_258) );
INVx1_ASAP7_75t_L g390 ( .A(n_259), .Y(n_390) );
AND2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_265), .Y(n_259) );
AND2x2_ASAP7_75t_L g286 ( .A(n_260), .B(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g297 ( .A(n_260), .B(n_266), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_260), .B(n_288), .Y(n_313) );
OAI222xp33_ASAP7_75t_L g335 ( .A1(n_260), .A2(n_336), .B1(n_341), .B2(n_342), .C1(n_350), .C2(n_352), .Y(n_335) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVx1_ASAP7_75t_SL g261 ( .A(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g323 ( .A(n_262), .B(n_324), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_262), .B(n_343), .Y(n_383) );
AND2x2_ASAP7_75t_L g394 ( .A(n_262), .B(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g402 ( .A(n_265), .Y(n_402) );
NAND2xp5_ASAP7_75t_SL g381 ( .A(n_267), .B(n_318), .Y(n_381) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
NOR2xp33_ASAP7_75t_L g321 ( .A(n_269), .B(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g339 ( .A(n_269), .B(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g270 ( .A(n_271), .B(n_272), .Y(n_270) );
INVx3_ASAP7_75t_L g284 ( .A(n_272), .Y(n_284) );
O2A1O1Ixp33_ASAP7_75t_L g374 ( .A1(n_272), .A2(n_375), .B(n_378), .C(n_380), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_272), .B(n_309), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_272), .B(n_292), .Y(n_414) );
AND2x2_ASAP7_75t_L g287 ( .A(n_273), .B(n_283), .Y(n_287) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_276), .B(n_277), .Y(n_275) );
INVx1_ASAP7_75t_L g314 ( .A(n_276), .Y(n_314) );
NAND2xp5_ASAP7_75t_SL g303 ( .A(n_277), .B(n_304), .Y(n_303) );
OR2x2_ASAP7_75t_L g366 ( .A(n_277), .B(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g405 ( .A(n_277), .B(n_305), .Y(n_405) );
INVx1_ASAP7_75t_L g417 ( .A(n_277), .Y(n_417) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_280), .B(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
OR2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_284), .Y(n_282) );
INVx1_ASAP7_75t_L g398 ( .A(n_283), .Y(n_398) );
A2O1A1Ixp33_ASAP7_75t_SL g285 ( .A1(n_286), .A2(n_288), .B(n_290), .C(n_294), .Y(n_285) );
AOI22xp33_ASAP7_75t_L g330 ( .A1(n_286), .A2(n_316), .B1(n_331), .B2(n_334), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_287), .B(n_301), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_287), .B(n_309), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_288), .B(n_346), .Y(n_345) );
INVx1_ASAP7_75t_SL g351 ( .A(n_288), .Y(n_351) );
AND2x2_ASAP7_75t_L g358 ( .A(n_288), .B(n_338), .Y(n_358) );
INVx2_ASAP7_75t_L g319 ( .A(n_289), .Y(n_319) );
INVxp67_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
NOR4xp25_ASAP7_75t_L g296 ( .A(n_293), .B(n_297), .C(n_298), .D(n_301), .Y(n_296) );
INVx1_ASAP7_75t_SL g367 ( .A(n_294), .Y(n_367) );
AND2x2_ASAP7_75t_L g411 ( .A(n_294), .B(n_412), .Y(n_411) );
OAI211xp5_ASAP7_75t_SL g295 ( .A1(n_296), .A2(n_303), .B(n_306), .C(n_315), .Y(n_295) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx1_ASAP7_75t_SL g301 ( .A(n_302), .Y(n_301) );
NOR2xp33_ASAP7_75t_L g423 ( .A(n_302), .B(n_372), .Y(n_423) );
AOI22xp5_ASAP7_75t_L g422 ( .A1(n_304), .A2(n_423), .B1(n_424), .B2(n_425), .Y(n_422) );
INVx1_ASAP7_75t_SL g377 ( .A(n_305), .Y(n_377) );
AND2x2_ASAP7_75t_L g416 ( .A(n_305), .B(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
NAND2xp5_ASAP7_75t_SL g409 ( .A(n_309), .B(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
NOR2xp33_ASAP7_75t_L g328 ( .A(n_313), .B(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_314), .B(n_339), .Y(n_399) );
OAI21xp5_ASAP7_75t_SL g315 ( .A1(n_316), .A2(n_321), .B(n_323), .Y(n_315) );
AND2x2_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
INVx1_ASAP7_75t_L g391 ( .A(n_318), .Y(n_391) );
AND2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
INVx2_ASAP7_75t_L g419 ( .A(n_319), .Y(n_419) );
HB1xp67_ASAP7_75t_L g346 ( .A(n_320), .Y(n_346) );
OAI21xp33_ASAP7_75t_L g325 ( .A1(n_326), .A2(n_327), .B(n_330), .Y(n_325) );
CKINVDCx16_ASAP7_75t_R g338 ( .A(n_326), .Y(n_338) );
OR2x2_ASAP7_75t_L g376 ( .A(n_326), .B(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
AOI21xp33_ASAP7_75t_SL g371 ( .A1(n_329), .A2(n_372), .B(n_373), .Y(n_371) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
AOI221xp5_ASAP7_75t_L g359 ( .A1(n_333), .A2(n_360), .B1(n_363), .B2(n_370), .C(n_371), .Y(n_359) );
INVx1_ASAP7_75t_SL g403 ( .A(n_334), .Y(n_403) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g337 ( .A(n_338), .B(n_339), .Y(n_337) );
OR2x2_ASAP7_75t_L g350 ( .A(n_338), .B(n_351), .Y(n_350) );
INVxp67_ASAP7_75t_L g387 ( .A(n_340), .Y(n_387) );
AOI22xp5_ASAP7_75t_L g342 ( .A1(n_343), .A2(n_344), .B1(n_347), .B2(n_348), .Y(n_342) );
INVx1_ASAP7_75t_L g382 ( .A(n_343), .Y(n_382) );
INVxp67_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_346), .B(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
NOR4xp25_ASAP7_75t_L g353 ( .A(n_354), .B(n_388), .C(n_401), .D(n_413), .Y(n_353) );
NAND3xp33_ASAP7_75t_SL g354 ( .A(n_355), .B(n_359), .C(n_374), .Y(n_354) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
NOR2xp33_ASAP7_75t_L g375 ( .A(n_357), .B(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_364), .B(n_369), .Y(n_373) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
OAI221xp5_ASAP7_75t_SL g401 ( .A1(n_376), .A2(n_402), .B1(n_403), .B2(n_404), .C(n_406), .Y(n_401) );
O2A1O1Ixp33_ASAP7_75t_L g392 ( .A1(n_378), .A2(n_393), .B(n_394), .C(n_396), .Y(n_392) );
INVx2_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
OAI22xp5_ASAP7_75t_L g396 ( .A1(n_379), .A2(n_397), .B1(n_399), .B2(n_400), .Y(n_396) );
INVx2_ASAP7_75t_SL g384 ( .A(n_385), .Y(n_384) );
A2O1A1Ixp33_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_390), .B(n_391), .C(n_392), .Y(n_388) );
INVx1_ASAP7_75t_L g407 ( .A(n_400), .Y(n_407) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
OAI21xp5_ASAP7_75t_SL g406 ( .A1(n_407), .A2(n_408), .B(n_411), .Y(n_406) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
OAI221xp5_ASAP7_75t_SL g413 ( .A1(n_414), .A2(n_415), .B1(n_418), .B2(n_420), .C(n_422), .Y(n_413) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVxp67_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
OAI22xp5_ASAP7_75t_SL g441 ( .A1(n_428), .A2(n_442), .B1(n_710), .B2(n_712), .Y(n_441) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_SL g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_SL g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_SL g438 ( .A(n_432), .Y(n_438) );
NOR2x2_ASAP7_75t_L g718 ( .A(n_433), .B(n_711), .Y(n_718) );
INVx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
OR2x2_ASAP7_75t_L g710 ( .A(n_434), .B(n_711), .Y(n_710) );
AND2x2_ASAP7_75t_L g434 ( .A(n_435), .B(n_436), .Y(n_434) );
AOI21xp33_ASAP7_75t_L g439 ( .A1(n_437), .A2(n_440), .B(n_724), .Y(n_439) );
INVx1_ASAP7_75t_L g720 ( .A(n_442), .Y(n_720) );
NAND2x1_ASAP7_75t_L g442 ( .A(n_443), .B(n_626), .Y(n_442) );
NOR5xp2_ASAP7_75t_L g443 ( .A(n_444), .B(n_549), .C(n_581), .D(n_596), .E(n_613), .Y(n_443) );
A2O1A1Ixp33_ASAP7_75t_L g444 ( .A1(n_445), .A2(n_477), .B(n_496), .C(n_537), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_446), .B(n_458), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_446), .B(n_649), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_446), .B(n_601), .Y(n_664) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_447), .B(n_546), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_447), .B(n_493), .Y(n_550) );
AND2x2_ASAP7_75t_L g591 ( .A(n_447), .B(n_592), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_447), .B(n_560), .Y(n_595) );
OR2x2_ASAP7_75t_L g632 ( .A(n_447), .B(n_483), .Y(n_632) );
INVx3_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
AND2x2_ASAP7_75t_L g482 ( .A(n_448), .B(n_483), .Y(n_482) );
INVx3_ASAP7_75t_L g540 ( .A(n_448), .Y(n_540) );
OR2x2_ASAP7_75t_L g703 ( .A(n_448), .B(n_543), .Y(n_703) );
AOI22xp5_ASAP7_75t_L g605 ( .A1(n_458), .A2(n_606), .B1(n_607), .B2(n_610), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_458), .B(n_540), .Y(n_689) );
AND2x2_ASAP7_75t_L g458 ( .A(n_459), .B(n_468), .Y(n_458) );
AND2x2_ASAP7_75t_L g495 ( .A(n_459), .B(n_483), .Y(n_495) );
AND2x2_ASAP7_75t_L g542 ( .A(n_459), .B(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g547 ( .A(n_459), .Y(n_547) );
INVx3_ASAP7_75t_L g560 ( .A(n_459), .Y(n_560) );
OR2x2_ASAP7_75t_L g580 ( .A(n_459), .B(n_543), .Y(n_580) );
AND2x2_ASAP7_75t_L g599 ( .A(n_459), .B(n_469), .Y(n_599) );
BUFx2_ASAP7_75t_L g631 ( .A(n_459), .Y(n_631) );
AND2x4_ASAP7_75t_L g546 ( .A(n_468), .B(n_547), .Y(n_546) );
INVx1_ASAP7_75t_SL g468 ( .A(n_469), .Y(n_468) );
BUFx2_ASAP7_75t_L g481 ( .A(n_469), .Y(n_481) );
INVx2_ASAP7_75t_L g494 ( .A(n_469), .Y(n_494) );
OR2x2_ASAP7_75t_L g562 ( .A(n_469), .B(n_543), .Y(n_562) );
AND2x2_ASAP7_75t_L g592 ( .A(n_469), .B(n_483), .Y(n_592) );
AND2x2_ASAP7_75t_L g609 ( .A(n_469), .B(n_540), .Y(n_609) );
AND2x2_ASAP7_75t_L g649 ( .A(n_469), .B(n_560), .Y(n_649) );
AND2x2_ASAP7_75t_SL g685 ( .A(n_469), .B(n_495), .Y(n_685) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
NAND2xp33_ASAP7_75t_SL g478 ( .A(n_479), .B(n_492), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_480), .B(n_482), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g663 ( .A(n_480), .B(n_664), .Y(n_663) );
INVx1_ASAP7_75t_SL g480 ( .A(n_481), .Y(n_480) );
OAI21xp33_ASAP7_75t_L g623 ( .A1(n_481), .A2(n_495), .B(n_624), .Y(n_623) );
NOR2xp33_ASAP7_75t_L g679 ( .A(n_481), .B(n_483), .Y(n_679) );
AND2x2_ASAP7_75t_L g615 ( .A(n_482), .B(n_616), .Y(n_615) );
INVx3_ASAP7_75t_L g543 ( .A(n_483), .Y(n_543) );
HB1xp67_ASAP7_75t_L g641 ( .A(n_483), .Y(n_641) );
NOR2xp33_ASAP7_75t_L g708 ( .A(n_492), .B(n_540), .Y(n_708) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_493), .A2(n_651), .B1(n_652), .B2(n_657), .Y(n_650) );
AND2x2_ASAP7_75t_L g493 ( .A(n_494), .B(n_495), .Y(n_493) );
AND2x2_ASAP7_75t_L g541 ( .A(n_494), .B(n_542), .Y(n_541) );
OR2x2_ASAP7_75t_L g579 ( .A(n_494), .B(n_580), .Y(n_579) );
INVx1_ASAP7_75t_SL g616 ( .A(n_494), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_495), .B(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g670 ( .A(n_495), .Y(n_670) );
CKINVDCx16_ASAP7_75t_R g496 ( .A(n_497), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_498), .B(n_517), .Y(n_497) );
INVx4_ASAP7_75t_L g556 ( .A(n_498), .Y(n_556) );
AND2x2_ASAP7_75t_L g634 ( .A(n_498), .B(n_601), .Y(n_634) );
AND2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_508), .Y(n_498) );
INVx3_ASAP7_75t_L g553 ( .A(n_499), .Y(n_553) );
AND2x2_ASAP7_75t_L g567 ( .A(n_499), .B(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g571 ( .A(n_499), .Y(n_571) );
INVx2_ASAP7_75t_L g585 ( .A(n_499), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_499), .B(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g642 ( .A(n_499), .B(n_637), .Y(n_642) );
AND2x2_ASAP7_75t_L g707 ( .A(n_499), .B(n_677), .Y(n_707) );
OR2x6_ASAP7_75t_L g499 ( .A(n_500), .B(n_506), .Y(n_499) );
AND2x2_ASAP7_75t_L g548 ( .A(n_508), .B(n_529), .Y(n_548) );
INVx2_ASAP7_75t_L g568 ( .A(n_508), .Y(n_568) );
INVx1_ASAP7_75t_L g573 ( .A(n_517), .Y(n_573) );
AND2x2_ASAP7_75t_L g619 ( .A(n_517), .B(n_567), .Y(n_619) );
AND2x2_ASAP7_75t_L g517 ( .A(n_518), .B(n_528), .Y(n_517) );
INVx2_ASAP7_75t_L g558 ( .A(n_518), .Y(n_558) );
INVx1_ASAP7_75t_L g566 ( .A(n_518), .Y(n_566) );
AND2x2_ASAP7_75t_L g584 ( .A(n_518), .B(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_518), .B(n_568), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_520), .B(n_525), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_522), .A2(n_523), .B(n_524), .Y(n_521) );
AND2x2_ASAP7_75t_L g601 ( .A(n_528), .B(n_558), .Y(n_601) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx2_ASAP7_75t_L g554 ( .A(n_529), .Y(n_554) );
AND2x2_ASAP7_75t_L g637 ( .A(n_529), .B(n_568), .Y(n_637) );
OAI21xp5_ASAP7_75t_SL g537 ( .A1(n_538), .A2(n_544), .B(n_548), .Y(n_537) );
INVx1_ASAP7_75t_SL g582 ( .A(n_538), .Y(n_582) );
AND2x2_ASAP7_75t_L g538 ( .A(n_539), .B(n_541), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_539), .B(n_546), .Y(n_639) );
INVx1_ASAP7_75t_SL g539 ( .A(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g588 ( .A(n_540), .B(n_543), .Y(n_588) );
AND2x2_ASAP7_75t_L g617 ( .A(n_540), .B(n_561), .Y(n_617) );
OR2x2_ASAP7_75t_L g620 ( .A(n_540), .B(n_580), .Y(n_620) );
AOI222xp33_ASAP7_75t_L g684 ( .A1(n_541), .A2(n_633), .B1(n_685), .B2(n_686), .C1(n_688), .C2(n_690), .Y(n_684) );
BUFx2_ASAP7_75t_L g598 ( .A(n_543), .Y(n_598) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
AND2x2_ASAP7_75t_L g587 ( .A(n_546), .B(n_588), .Y(n_587) );
INVx3_ASAP7_75t_SL g604 ( .A(n_546), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_546), .B(n_598), .Y(n_658) );
AND2x2_ASAP7_75t_L g593 ( .A(n_548), .B(n_553), .Y(n_593) );
INVx1_ASAP7_75t_L g612 ( .A(n_548), .Y(n_612) );
OAI221xp5_ASAP7_75t_SL g549 ( .A1(n_550), .A2(n_551), .B1(n_555), .B2(n_559), .C(n_563), .Y(n_549) );
OR2x2_ASAP7_75t_L g621 ( .A(n_551), .B(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_553), .B(n_554), .Y(n_552) );
AND2x2_ASAP7_75t_L g606 ( .A(n_553), .B(n_576), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_553), .B(n_566), .Y(n_646) );
AND2x2_ASAP7_75t_L g651 ( .A(n_553), .B(n_601), .Y(n_651) );
HB1xp67_ASAP7_75t_L g661 ( .A(n_553), .Y(n_661) );
NAND2x1_ASAP7_75t_SL g672 ( .A(n_553), .B(n_673), .Y(n_672) );
OR2x2_ASAP7_75t_L g557 ( .A(n_554), .B(n_558), .Y(n_557) );
INVx2_ASAP7_75t_L g577 ( .A(n_554), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_554), .B(n_572), .Y(n_603) );
INVx1_ASAP7_75t_L g669 ( .A(n_554), .Y(n_669) );
INVx1_ASAP7_75t_L g644 ( .A(n_555), .Y(n_644) );
OR2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_557), .Y(n_555) );
INVx1_ASAP7_75t_L g656 ( .A(n_556), .Y(n_656) );
NOR2xp67_ASAP7_75t_L g668 ( .A(n_556), .B(n_669), .Y(n_668) );
INVx2_ASAP7_75t_L g673 ( .A(n_557), .Y(n_673) );
NOR2xp33_ASAP7_75t_L g680 ( .A(n_557), .B(n_681), .Y(n_680) );
AND2x2_ASAP7_75t_L g576 ( .A(n_558), .B(n_577), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_558), .B(n_568), .Y(n_589) );
INVx1_ASAP7_75t_L g655 ( .A(n_558), .Y(n_655) );
INVx1_ASAP7_75t_L g676 ( .A(n_559), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_560), .B(n_561), .Y(n_559) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
OAI21xp5_ASAP7_75t_SL g563 ( .A1(n_564), .A2(n_569), .B(n_578), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_565), .B(n_567), .Y(n_564) );
AND2x2_ASAP7_75t_L g709 ( .A(n_565), .B(n_642), .Y(n_709) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g677 ( .A(n_566), .B(n_637), .Y(n_677) );
AOI32xp33_ASAP7_75t_L g590 ( .A1(n_567), .A2(n_573), .A3(n_591), .B1(n_593), .B2(n_594), .Y(n_590) );
AOI322xp5_ASAP7_75t_L g692 ( .A1(n_567), .A2(n_599), .A3(n_682), .B1(n_693), .B2(n_694), .C1(n_695), .C2(n_697), .Y(n_692) );
INVx2_ASAP7_75t_L g572 ( .A(n_568), .Y(n_572) );
INVx1_ASAP7_75t_L g682 ( .A(n_568), .Y(n_682) );
OAI22xp5_ASAP7_75t_L g569 ( .A1(n_570), .A2(n_573), .B1(n_574), .B2(n_575), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_570), .B(n_576), .Y(n_625) );
AND2x2_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_571), .B(n_637), .Y(n_687) );
INVx1_ASAP7_75t_L g574 ( .A(n_572), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_572), .B(n_601), .Y(n_691) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx1_ASAP7_75t_SL g578 ( .A(n_579), .Y(n_578) );
NOR2xp33_ASAP7_75t_L g674 ( .A(n_580), .B(n_675), .Y(n_674) );
OAI221xp5_ASAP7_75t_SL g581 ( .A1(n_582), .A2(n_583), .B1(n_586), .B2(n_589), .C(n_590), .Y(n_581) );
OR2x2_ASAP7_75t_L g602 ( .A(n_583), .B(n_603), .Y(n_602) );
OR2x2_ASAP7_75t_L g611 ( .A(n_583), .B(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g636 ( .A(n_584), .B(n_637), .Y(n_636) );
INVx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g640 ( .A(n_594), .B(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
OAI221xp5_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_600), .B1(n_602), .B2(n_604), .C(n_605), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_598), .B(n_599), .Y(n_597) );
AOI22xp5_ASAP7_75t_L g628 ( .A1(n_598), .A2(n_629), .B1(n_633), .B2(n_634), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_599), .B(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g704 ( .A(n_599), .Y(n_704) );
INVx1_ASAP7_75t_L g698 ( .A(n_601), .Y(n_698) );
INVx1_ASAP7_75t_SL g633 ( .A(n_602), .Y(n_633) );
NOR2xp33_ASAP7_75t_L g694 ( .A(n_604), .B(n_632), .Y(n_694) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_609), .B(n_668), .Y(n_667) );
INVx1_ASAP7_75t_SL g675 ( .A(n_609), .Y(n_675) );
INVx1_ASAP7_75t_SL g610 ( .A(n_611), .Y(n_610) );
OAI221xp5_ASAP7_75t_SL g613 ( .A1(n_614), .A2(n_618), .B1(n_620), .B2(n_621), .C(n_623), .Y(n_613) );
NOR2xp33_ASAP7_75t_SL g614 ( .A(n_615), .B(n_617), .Y(n_614) );
AOI22xp5_ASAP7_75t_L g678 ( .A1(n_615), .A2(n_633), .B1(n_679), .B2(n_680), .Y(n_678) );
CKINVDCx14_ASAP7_75t_R g618 ( .A(n_619), .Y(n_618) );
OAI21xp33_ASAP7_75t_L g697 ( .A1(n_620), .A2(n_698), .B(n_699), .Y(n_697) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
NOR3xp33_ASAP7_75t_SL g626 ( .A(n_627), .B(n_659), .C(n_683), .Y(n_626) );
NAND4xp25_ASAP7_75t_L g627 ( .A(n_628), .B(n_635), .C(n_643), .D(n_650), .Y(n_627) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
OR2x2_ASAP7_75t_L g630 ( .A(n_631), .B(n_632), .Y(n_630) );
INVx1_ASAP7_75t_L g706 ( .A(n_631), .Y(n_706) );
INVx3_ASAP7_75t_SL g700 ( .A(n_632), .Y(n_700) );
OR2x2_ASAP7_75t_L g705 ( .A(n_632), .B(n_706), .Y(n_705) );
AOI22xp5_ASAP7_75t_L g635 ( .A1(n_636), .A2(n_638), .B1(n_640), .B2(n_642), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_637), .B(n_655), .Y(n_696) );
INVxp67_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
OAI21xp5_ASAP7_75t_SL g643 ( .A1(n_644), .A2(n_645), .B(n_647), .Y(n_643) );
INVxp67_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_654), .B(n_656), .Y(n_653) );
INVxp67_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
OAI211xp5_ASAP7_75t_SL g659 ( .A1(n_660), .A2(n_662), .B(n_665), .C(n_678), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g693 ( .A(n_664), .Y(n_693) );
AOI222xp33_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_670), .B1(n_671), .B2(n_674), .C1(n_676), .C2(n_677), .Y(n_665) );
INVxp67_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
NAND4xp25_ASAP7_75t_SL g702 ( .A(n_675), .B(n_703), .C(n_704), .D(n_705), .Y(n_702) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
NAND3xp33_ASAP7_75t_SL g683 ( .A(n_684), .B(n_692), .C(n_701), .Y(n_683) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_707), .B1(n_708), .B2(n_709), .Y(n_701) );
INVx1_ASAP7_75t_L g722 ( .A(n_712), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_713), .Y(n_723) );
INVx1_ASAP7_75t_SL g716 ( .A(n_717), .Y(n_716) );
INVx3_ASAP7_75t_SL g717 ( .A(n_718), .Y(n_717) );
INVx2_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_SL g725 ( .A(n_726), .Y(n_725) );
endmodule