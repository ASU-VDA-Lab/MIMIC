module real_aes_6030_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_800;
wire n_778;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_943;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_905;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_852;
wire n_766;
wire n_132;
wire n_857;
wire n_919;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_923;
wire n_952;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_937;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_889;
wire n_955;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_958;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_953;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_356;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_938;
wire n_121;
wire n_352;
wire n_935;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_951;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_872;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_909;
wire n_298;
wire n_523;
wire n_860;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_950;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_936;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_142;
wire n_561;
wire n_947;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_913;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_917;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_957;
wire n_296;
wire n_954;
wire n_702;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_945;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_133;
wire n_934;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_927;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_291;
wire n_907;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_939;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_928;
wire n_155;
wire n_637;
wire n_243;
wire n_899;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_922;
wire n_520;
wire n_482;
wire n_633;
wire n_679;
wire n_926;
wire n_149;
wire n_942;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_946;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_888;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_929;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_949;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_921;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
NAND2xp5_ASAP7_75t_L g125 ( .A(n_0), .B(n_126), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g153 ( .A(n_1), .Y(n_153) );
INVx1_ASAP7_75t_L g648 ( .A(n_2), .Y(n_648) );
AOI22xp5_ASAP7_75t_L g101 ( .A1(n_3), .A2(n_102), .B1(n_946), .B2(n_956), .Y(n_101) );
O2A1O1Ixp33_ASAP7_75t_SL g201 ( .A1(n_4), .A2(n_148), .B(n_202), .C(n_204), .Y(n_201) );
OAI22xp33_ASAP7_75t_L g138 ( .A1(n_5), .A2(n_84), .B1(n_133), .B2(n_139), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_6), .B(n_537), .Y(n_603) );
INVx1_ASAP7_75t_L g514 ( .A(n_7), .Y(n_514) );
INVx1_ASAP7_75t_L g524 ( .A(n_7), .Y(n_524) );
INVxp67_ASAP7_75t_L g921 ( .A(n_7), .Y(n_921) );
BUFx2_ASAP7_75t_L g952 ( .A(n_7), .Y(n_952) );
NAND2xp5_ASAP7_75t_SL g604 ( .A(n_8), .B(n_296), .Y(n_604) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_9), .A2(n_35), .B1(n_536), .B2(n_587), .Y(n_586) );
AOI22xp5_ASAP7_75t_L g671 ( .A1(n_10), .A2(n_41), .B1(n_559), .B2(n_672), .Y(n_671) );
AOI22xp5_ASAP7_75t_L g633 ( .A1(n_11), .A2(n_68), .B1(n_625), .B2(n_627), .Y(n_633) );
INVx1_ASAP7_75t_L g643 ( .A(n_12), .Y(n_643) );
CKINVDCx5p33_ASAP7_75t_R g181 ( .A(n_13), .Y(n_181) );
OAI22xp5_ASAP7_75t_L g192 ( .A1(n_14), .A2(n_74), .B1(n_139), .B2(n_193), .Y(n_192) );
CKINVDCx5p33_ASAP7_75t_R g223 ( .A(n_15), .Y(n_223) );
INVx1_ASAP7_75t_L g646 ( .A(n_16), .Y(n_646) );
AOI22xp5_ASAP7_75t_L g191 ( .A1(n_17), .A2(n_64), .B1(n_133), .B2(n_154), .Y(n_191) );
OA21x2_ASAP7_75t_L g128 ( .A1(n_18), .A2(n_73), .B(n_129), .Y(n_128) );
OA21x2_ASAP7_75t_L g168 ( .A1(n_18), .A2(n_73), .B(n_129), .Y(n_168) );
AOI22xp5_ASAP7_75t_L g624 ( .A1(n_19), .A2(n_71), .B1(n_625), .B2(n_627), .Y(n_624) );
INVx1_ASAP7_75t_L g640 ( .A(n_20), .Y(n_640) );
CKINVDCx5p33_ASAP7_75t_R g172 ( .A(n_21), .Y(n_172) );
BUFx3_ASAP7_75t_L g106 ( .A(n_22), .Y(n_106) );
O2A1O1Ixp33_ASAP7_75t_L g208 ( .A1(n_23), .A2(n_140), .B(n_209), .C(n_210), .Y(n_208) );
OAI22xp33_ASAP7_75t_SL g132 ( .A1(n_24), .A2(n_46), .B1(n_133), .B2(n_134), .Y(n_132) );
AOI22xp33_ASAP7_75t_L g254 ( .A1(n_25), .A2(n_33), .B1(n_134), .B2(n_179), .Y(n_254) );
AO22x1_ASAP7_75t_L g599 ( .A1(n_26), .A2(n_81), .B1(n_548), .B2(n_600), .Y(n_599) );
CKINVDCx5p33_ASAP7_75t_R g540 ( .A(n_27), .Y(n_540) );
AND2x2_ASAP7_75t_L g558 ( .A(n_28), .B(n_559), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_29), .B(n_548), .Y(n_547) );
O2A1O1Ixp5_ASAP7_75t_L g291 ( .A1(n_30), .A2(n_148), .B(n_292), .C(n_293), .Y(n_291) );
INVx1_ASAP7_75t_L g519 ( .A(n_31), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g955 ( .A(n_31), .B(n_83), .Y(n_955) );
AOI22x1_ASAP7_75t_L g674 ( .A1(n_32), .A2(n_96), .B1(n_583), .B2(n_625), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_34), .B(n_590), .Y(n_589) );
OAI22xp5_ASAP7_75t_SL g943 ( .A1(n_36), .A2(n_56), .B1(n_944), .B2(n_945), .Y(n_943) );
INVx1_ASAP7_75t_L g945 ( .A(n_36), .Y(n_945) );
AND2x2_ASAP7_75t_L g953 ( .A(n_37), .B(n_954), .Y(n_953) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_38), .B(n_218), .Y(n_258) );
CKINVDCx5p33_ASAP7_75t_R g294 ( .A(n_39), .Y(n_294) );
NAND2xp5_ASAP7_75t_SL g568 ( .A(n_40), .B(n_569), .Y(n_568) );
CKINVDCx5p33_ASAP7_75t_R g206 ( .A(n_42), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_43), .B(n_616), .Y(n_615) );
AOI22xp5_ASAP7_75t_L g110 ( .A1(n_44), .A2(n_58), .B1(n_111), .B2(n_112), .Y(n_110) );
INVx1_ASAP7_75t_L g112 ( .A(n_44), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_45), .B(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g129 ( .A(n_47), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g923 ( .A(n_48), .Y(n_923) );
AND2x4_ASAP7_75t_L g142 ( .A(n_49), .B(n_143), .Y(n_142) );
AND2x4_ASAP7_75t_L g166 ( .A(n_49), .B(n_143), .Y(n_166) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_50), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g151 ( .A(n_51), .Y(n_151) );
INVx2_ASAP7_75t_L g629 ( .A(n_52), .Y(n_629) );
O2A1O1Ixp33_ASAP7_75t_L g175 ( .A1(n_53), .A2(n_148), .B(n_176), .C(n_178), .Y(n_175) );
INVx2_ASAP7_75t_L g228 ( .A(n_54), .Y(n_228) );
CKINVDCx5p33_ASAP7_75t_R g300 ( .A(n_55), .Y(n_300) );
CKINVDCx5p33_ASAP7_75t_R g944 ( .A(n_56), .Y(n_944) );
CKINVDCx5p33_ASAP7_75t_R g150 ( .A(n_57), .Y(n_150) );
INVx1_ASAP7_75t_L g111 ( .A(n_58), .Y(n_111) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_59), .A2(n_76), .B1(n_536), .B2(n_583), .Y(n_582) );
CKINVDCx5p33_ASAP7_75t_R g915 ( .A(n_60), .Y(n_915) );
CKINVDCx14_ASAP7_75t_R g606 ( .A(n_61), .Y(n_606) );
AND2x2_ASAP7_75t_L g566 ( .A(n_62), .B(n_548), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_63), .B(n_157), .Y(n_156) );
AOI22xp5_ASAP7_75t_L g255 ( .A1(n_65), .A2(n_82), .B1(n_203), .B2(n_256), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_66), .B(n_618), .Y(n_617) );
CKINVDCx5p33_ASAP7_75t_R g155 ( .A(n_67), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_69), .B(n_157), .Y(n_609) );
NAND2xp33_ASAP7_75t_R g196 ( .A(n_70), .B(n_168), .Y(n_196) );
AOI22xp33_ASAP7_75t_L g265 ( .A1(n_70), .A2(n_99), .B1(n_218), .B2(n_266), .Y(n_265) );
NAND2x1p5_ASAP7_75t_L g570 ( .A(n_72), .B(n_553), .Y(n_570) );
CKINVDCx14_ASAP7_75t_R g677 ( .A(n_75), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_77), .B(n_537), .Y(n_613) );
OR2x6_ASAP7_75t_L g516 ( .A(n_78), .B(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g950 ( .A(n_78), .Y(n_950) );
CKINVDCx5p33_ASAP7_75t_R g227 ( .A(n_79), .Y(n_227) );
CKINVDCx5p33_ASAP7_75t_R g224 ( .A(n_80), .Y(n_224) );
INVx1_ASAP7_75t_L g518 ( .A(n_83), .Y(n_518) );
INVx1_ASAP7_75t_L g954 ( .A(n_85), .Y(n_954) );
BUFx5_ASAP7_75t_L g133 ( .A(n_86), .Y(n_133) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_86), .Y(n_135) );
INVx1_ASAP7_75t_L g180 ( .A(n_86), .Y(n_180) );
INVx2_ASAP7_75t_L g215 ( .A(n_87), .Y(n_215) );
INVx2_ASAP7_75t_L g650 ( .A(n_88), .Y(n_650) );
INVx2_ASAP7_75t_L g183 ( .A(n_89), .Y(n_183) );
CKINVDCx5p33_ASAP7_75t_R g211 ( .A(n_90), .Y(n_211) );
NAND2xp33_ASAP7_75t_L g562 ( .A(n_91), .B(n_563), .Y(n_562) );
INVx2_ASAP7_75t_SL g143 ( .A(n_92), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_93), .B(n_543), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_94), .B(n_569), .Y(n_612) );
INVx1_ASAP7_75t_L g298 ( .A(n_95), .Y(n_298) );
INVx2_ASAP7_75t_L g302 ( .A(n_97), .Y(n_302) );
OAI21xp33_ASAP7_75t_SL g170 ( .A1(n_98), .A2(n_133), .B(n_171), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_99), .B(n_218), .Y(n_217) );
INVxp67_ASAP7_75t_SL g244 ( .A(n_99), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_100), .B(n_551), .Y(n_550) );
AO21x2_ASAP7_75t_L g102 ( .A1(n_103), .A2(n_107), .B(n_937), .Y(n_102) );
BUFx4_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
BUFx8_ASAP7_75t_L g938 ( .A(n_104), .Y(n_938) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
CKINVDCx6p67_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_108), .B(n_927), .Y(n_107) );
AOI211xp5_ASAP7_75t_L g108 ( .A1(n_109), .A2(n_113), .B(n_914), .C(n_922), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g927 ( .A(n_110), .B(n_928), .Y(n_927) );
OAI21xp5_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_511), .B(n_520), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx2_ASAP7_75t_L g933 ( .A(n_115), .Y(n_933) );
OR2x2_ASAP7_75t_L g115 ( .A(n_116), .B(n_425), .Y(n_115) );
NAND4xp25_ASAP7_75t_L g116 ( .A(n_117), .B(n_322), .C(n_377), .D(n_406), .Y(n_116) );
NOR2xp67_ASAP7_75t_L g117 ( .A(n_118), .B(n_231), .Y(n_117) );
AND2x2_ASAP7_75t_L g118 ( .A(n_119), .B(n_184), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OAI221xp5_ASAP7_75t_SL g323 ( .A1(n_120), .A2(n_324), .B1(n_330), .B2(n_332), .C(n_335), .Y(n_323) );
OR2x2_ASAP7_75t_L g120 ( .A(n_121), .B(n_159), .Y(n_120) );
INVx1_ASAP7_75t_SL g121 ( .A(n_122), .Y(n_121) );
AND2x2_ASAP7_75t_L g407 ( .A(n_122), .B(n_408), .Y(n_407) );
OAI21xp33_ASAP7_75t_L g507 ( .A1(n_122), .A2(n_508), .B(n_510), .Y(n_507) );
AND2x4_ASAP7_75t_L g122 ( .A(n_123), .B(n_144), .Y(n_122) );
AND2x2_ASAP7_75t_L g309 ( .A(n_123), .B(n_163), .Y(n_309) );
INVx1_ASAP7_75t_L g402 ( .A(n_123), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_123), .B(n_287), .Y(n_444) );
INVx3_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
HB1xp67_ASAP7_75t_L g270 ( .A(n_124), .Y(n_270) );
INVx2_ASAP7_75t_L g281 ( .A(n_124), .Y(n_281) );
NAND2xp33_ASAP7_75t_R g340 ( .A(n_124), .B(n_163), .Y(n_340) );
INVx1_ASAP7_75t_L g363 ( .A(n_124), .Y(n_363) );
AND2x2_ASAP7_75t_L g370 ( .A(n_124), .B(n_144), .Y(n_370) );
AND2x2_ASAP7_75t_L g382 ( .A(n_124), .B(n_163), .Y(n_382) );
AND2x4_ASAP7_75t_L g124 ( .A(n_125), .B(n_130), .Y(n_124) );
INVx2_ASAP7_75t_L g146 ( .A(n_126), .Y(n_146) );
NOR2xp33_ASAP7_75t_SL g212 ( .A(n_126), .B(n_213), .Y(n_212) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_127), .B(n_142), .Y(n_141) );
NOR2xp33_ASAP7_75t_SL g214 ( .A(n_127), .B(n_215), .Y(n_214) );
INVx2_ASAP7_75t_L g218 ( .A(n_127), .Y(n_218) );
INVx3_ASAP7_75t_L g553 ( .A(n_127), .Y(n_553) );
INVx4_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx2_ASAP7_75t_L g158 ( .A(n_128), .Y(n_158) );
BUFx3_ASAP7_75t_L g315 ( .A(n_128), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_131), .B(n_137), .Y(n_130) );
NAND2xp5_ASAP7_75t_SL g131 ( .A(n_132), .B(n_136), .Y(n_131) );
AOI22xp33_ASAP7_75t_SL g149 ( .A1(n_133), .A2(n_134), .B1(n_150), .B2(n_151), .Y(n_149) );
AOI22xp33_ASAP7_75t_L g152 ( .A1(n_133), .A2(n_153), .B1(n_154), .B2(n_155), .Y(n_152) );
NAND2xp5_ASAP7_75t_SL g171 ( .A(n_133), .B(n_172), .Y(n_171) );
AOI22xp5_ASAP7_75t_L g222 ( .A1(n_133), .A2(n_134), .B1(n_223), .B2(n_224), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_133), .B(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_133), .B(n_300), .Y(n_299) );
INVx2_ASAP7_75t_L g537 ( .A(n_133), .Y(n_537) );
INVx2_ASAP7_75t_L g548 ( .A(n_133), .Y(n_548) );
INVx2_ASAP7_75t_L g618 ( .A(n_133), .Y(n_618) );
INVx2_ASAP7_75t_L g626 ( .A(n_133), .Y(n_626) );
INVx2_ASAP7_75t_L g205 ( .A(n_134), .Y(n_205) );
INVx2_ASAP7_75t_SL g256 ( .A(n_134), .Y(n_256) );
INVx2_ASAP7_75t_L g560 ( .A(n_134), .Y(n_560) );
INVx1_ASAP7_75t_L g563 ( .A(n_134), .Y(n_563) );
INVx1_ASAP7_75t_L g569 ( .A(n_134), .Y(n_569) );
INVx6_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g139 ( .A(n_135), .Y(n_139) );
INVx2_ASAP7_75t_L g154 ( .A(n_135), .Y(n_154) );
INVx3_ASAP7_75t_L g177 ( .A(n_135), .Y(n_177) );
INVx3_ASAP7_75t_L g140 ( .A(n_136), .Y(n_140) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_136), .Y(n_148) );
INVx4_ASAP7_75t_L g174 ( .A(n_136), .Y(n_174) );
BUFx6f_ASAP7_75t_L g253 ( .A(n_136), .Y(n_253) );
INVx1_ASAP7_75t_L g257 ( .A(n_136), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_136), .B(n_298), .Y(n_297) );
INVxp67_ASAP7_75t_L g564 ( .A(n_136), .Y(n_564) );
NOR2xp33_ASAP7_75t_L g639 ( .A(n_136), .B(n_640), .Y(n_639) );
NOR2xp33_ASAP7_75t_L g642 ( .A(n_136), .B(n_643), .Y(n_642) );
AOI21xp5_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_140), .B(n_141), .Y(n_137) );
INVx1_ASAP7_75t_L g543 ( .A(n_139), .Y(n_543) );
OAI221xp5_ASAP7_75t_L g147 ( .A1(n_140), .A2(n_142), .B1(n_148), .B2(n_149), .C(n_152), .Y(n_147) );
INVx3_ASAP7_75t_L g632 ( .A(n_140), .Y(n_632) );
INVx1_ASAP7_75t_L g195 ( .A(n_142), .Y(n_195) );
BUFx6f_ASAP7_75t_L g239 ( .A(n_142), .Y(n_239) );
INVx3_ASAP7_75t_L g575 ( .A(n_142), .Y(n_575) );
INVx3_ASAP7_75t_L g581 ( .A(n_142), .Y(n_581) );
AND2x2_ASAP7_75t_L g248 ( .A(n_144), .B(n_249), .Y(n_248) );
OR2x2_ASAP7_75t_L g311 ( .A(n_144), .B(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g350 ( .A(n_144), .B(n_351), .Y(n_350) );
OA21x2_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_147), .B(n_156), .Y(n_144) );
OA21x2_ASAP7_75t_L g273 ( .A1(n_145), .A2(n_147), .B(n_156), .Y(n_273) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
OR2x2_ASAP7_75t_L g243 ( .A(n_146), .B(n_244), .Y(n_243) );
AOI21xp33_ASAP7_75t_SL g573 ( .A1(n_146), .A2(n_574), .B(n_576), .Y(n_573) );
AOI22xp5_ASAP7_75t_L g190 ( .A1(n_148), .A2(n_174), .B1(n_191), .B2(n_192), .Y(n_190) );
INVx1_ASAP7_75t_L g229 ( .A(n_148), .Y(n_229) );
OAI22xp33_ASAP7_75t_L g242 ( .A1(n_148), .A2(n_174), .B1(n_222), .B2(n_226), .Y(n_242) );
INVxp67_ASAP7_75t_L g549 ( .A(n_148), .Y(n_549) );
INVx2_ASAP7_75t_SL g572 ( .A(n_148), .Y(n_572) );
INVx1_ASAP7_75t_L g598 ( .A(n_148), .Y(n_598) );
INVx1_ASAP7_75t_L g209 ( .A(n_154), .Y(n_209) );
AOI22xp5_ASAP7_75t_L g226 ( .A1(n_154), .A2(n_179), .B1(n_227), .B2(n_228), .Y(n_226) );
INVx2_ASAP7_75t_L g546 ( .A(n_154), .Y(n_546) );
NOR2xp67_ASAP7_75t_L g194 ( .A(n_157), .B(n_195), .Y(n_194) );
NOR2x1_ASAP7_75t_L g619 ( .A(n_157), .B(n_575), .Y(n_619) );
INVx3_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_158), .B(n_183), .Y(n_182) );
BUFx3_ASAP7_75t_L g230 ( .A(n_158), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g649 ( .A(n_158), .B(n_650), .Y(n_649) );
OR2x2_ASAP7_75t_L g404 ( .A(n_159), .B(n_405), .Y(n_404) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
NAND2x1p5_ASAP7_75t_L g279 ( .A(n_160), .B(n_280), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_160), .B(n_331), .Y(n_414) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx1_ASAP7_75t_L g260 ( .A(n_162), .Y(n_260) );
AND2x2_ASAP7_75t_L g485 ( .A(n_162), .B(n_370), .Y(n_485) );
AND2x2_ASAP7_75t_L g508 ( .A(n_162), .B(n_509), .Y(n_508) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx1_ASAP7_75t_L g274 ( .A(n_163), .Y(n_274) );
INVx2_ASAP7_75t_L g287 ( .A(n_163), .Y(n_287) );
OR2x2_ASAP7_75t_L g375 ( .A(n_163), .B(n_281), .Y(n_375) );
AND2x2_ASAP7_75t_L g422 ( .A(n_163), .B(n_272), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_163), .B(n_273), .Y(n_440) );
BUFx2_ASAP7_75t_L g472 ( .A(n_163), .Y(n_472) );
INVx3_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
AOI21x1_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_169), .B(n_182), .Y(n_164) );
AND2x2_ASAP7_75t_L g165 ( .A(n_166), .B(n_167), .Y(n_165) );
INVx4_ASAP7_75t_L g213 ( .A(n_166), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_166), .B(n_240), .Y(n_251) );
INVx1_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
BUFx3_ASAP7_75t_L g241 ( .A(n_168), .Y(n_241) );
INVx2_ASAP7_75t_L g267 ( .A(n_168), .Y(n_267) );
INVx1_ASAP7_75t_L g303 ( .A(n_168), .Y(n_303) );
NOR2xp33_ASAP7_75t_L g580 ( .A(n_168), .B(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g591 ( .A(n_168), .Y(n_591) );
AOI21xp5_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_173), .B(n_175), .Y(n_169) );
AOI221xp5_ASAP7_75t_L g220 ( .A1(n_173), .A2(n_213), .B1(n_221), .B2(n_225), .C(n_229), .Y(n_220) );
INVx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
OAI22xp5_ASAP7_75t_L g295 ( .A1(n_174), .A2(n_296), .B1(n_297), .B2(n_299), .Y(n_295) );
NAND3xp33_ASAP7_75t_SL g623 ( .A(n_174), .B(n_267), .C(n_574), .Y(n_623) );
NOR2xp33_ASAP7_75t_SL g645 ( .A(n_174), .B(n_646), .Y(n_645) );
NOR2xp33_ASAP7_75t_L g647 ( .A(n_174), .B(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx1_ASAP7_75t_L g292 ( .A(n_177), .Y(n_292) );
INVx1_ASAP7_75t_L g296 ( .A(n_177), .Y(n_296) );
INVx2_ASAP7_75t_L g588 ( .A(n_177), .Y(n_588) );
INVx2_ASAP7_75t_L g616 ( .A(n_177), .Y(n_616) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_179), .B(n_181), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_179), .B(n_211), .Y(n_210) );
INVx2_ASAP7_75t_L g601 ( .A(n_179), .Y(n_601) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx2_ASAP7_75t_L g193 ( .A(n_180), .Y(n_193) );
AOI221xp5_ASAP7_75t_L g406 ( .A1(n_184), .A2(n_407), .B1(n_409), .B2(n_412), .C(n_415), .Y(n_406) );
INVx2_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_186), .B(n_197), .Y(n_185) );
OR2x2_ASAP7_75t_L g234 ( .A(n_186), .B(n_235), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_186), .B(n_236), .Y(n_434) );
OR2x2_ASAP7_75t_L g467 ( .A(n_186), .B(n_342), .Y(n_467) );
INVx2_ASAP7_75t_SL g186 ( .A(n_187), .Y(n_186) );
HB1xp67_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
AND2x2_ASAP7_75t_L g278 ( .A(n_188), .B(n_237), .Y(n_278) );
INVx2_ASAP7_75t_L g329 ( .A(n_188), .Y(n_329) );
AND2x2_ASAP7_75t_L g373 ( .A(n_188), .B(n_334), .Y(n_373) );
INVx1_ASAP7_75t_L g387 ( .A(n_188), .Y(n_387) );
AND2x2_ASAP7_75t_L g188 ( .A(n_189), .B(n_196), .Y(n_188) );
AND2x2_ASAP7_75t_L g264 ( .A(n_189), .B(n_265), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_190), .B(n_194), .Y(n_189) );
INVx2_ASAP7_75t_L g203 ( .A(n_193), .Y(n_203) );
OR2x2_ASAP7_75t_L g596 ( .A(n_195), .B(n_551), .Y(n_596) );
NOR2xp33_ASAP7_75t_L g636 ( .A(n_195), .B(n_266), .Y(n_636) );
INVxp67_ASAP7_75t_SL g430 ( .A(n_197), .Y(n_430) );
BUFx6f_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
AND2x2_ASAP7_75t_L g424 ( .A(n_198), .B(n_328), .Y(n_424) );
AND2x2_ASAP7_75t_L g497 ( .A(n_198), .B(n_386), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_198), .B(n_501), .Y(n_500) );
AND2x2_ASAP7_75t_L g198 ( .A(n_199), .B(n_216), .Y(n_198) );
AND2x4_ASAP7_75t_L g236 ( .A(n_199), .B(n_237), .Y(n_236) );
INVx1_ASAP7_75t_L g277 ( .A(n_199), .Y(n_277) );
INVx1_ASAP7_75t_L g327 ( .A(n_199), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_199), .B(n_289), .Y(n_338) );
INVx2_ASAP7_75t_L g344 ( .A(n_199), .Y(n_344) );
HB1xp67_ASAP7_75t_L g390 ( .A(n_199), .Y(n_390) );
OR2x2_ASAP7_75t_L g411 ( .A(n_199), .B(n_216), .Y(n_411) );
HB1xp67_ASAP7_75t_L g505 ( .A(n_199), .Y(n_505) );
AO31x2_ASAP7_75t_L g199 ( .A1(n_200), .A2(n_207), .A3(n_212), .B(n_214), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
INVx3_ASAP7_75t_L g672 ( .A(n_203), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_205), .B(n_206), .Y(n_204) );
INVx1_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
NOR3xp33_ASAP7_75t_L g290 ( .A(n_213), .B(n_291), .C(n_295), .Y(n_290) );
AND2x2_ASAP7_75t_L g305 ( .A(n_216), .B(n_277), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_216), .B(n_288), .Y(n_345) );
NOR2xp33_ASAP7_75t_L g459 ( .A(n_216), .B(n_460), .Y(n_459) );
AND2x2_ASAP7_75t_L g216 ( .A(n_217), .B(n_219), .Y(n_216) );
AND2x2_ASAP7_75t_L g263 ( .A(n_219), .B(n_264), .Y(n_263) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_220), .B(n_230), .Y(n_219) );
INVx1_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVx1_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g614 ( .A1(n_229), .A2(n_615), .B(n_617), .Y(n_614) );
AO21x2_ASAP7_75t_L g289 ( .A1(n_230), .A2(n_290), .B(n_301), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_232), .B(n_283), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_233), .A2(n_245), .B(n_261), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
INVx2_ASAP7_75t_SL g235 ( .A(n_236), .Y(n_235) );
OAI21xp33_ASAP7_75t_L g391 ( .A1(n_236), .A2(n_392), .B(n_394), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_236), .B(n_386), .Y(n_394) );
AND2x2_ASAP7_75t_L g486 ( .A(n_236), .B(n_328), .Y(n_486) );
AND2x2_ASAP7_75t_L g510 ( .A(n_236), .B(n_373), .Y(n_510) );
INVx1_ASAP7_75t_L g318 ( .A(n_237), .Y(n_318) );
OAI21x1_ASAP7_75t_L g237 ( .A1(n_238), .A2(n_242), .B(n_243), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_239), .B(n_240), .Y(n_238) );
OAI21x1_ASAP7_75t_L g534 ( .A1(n_239), .A2(n_535), .B(n_544), .Y(n_534) );
AO31x2_ASAP7_75t_L g669 ( .A1(n_239), .A2(n_670), .A3(n_675), .B(n_676), .Y(n_669) );
AO31x2_ASAP7_75t_L g690 ( .A1(n_239), .A2(n_670), .A3(n_675), .B(n_676), .Y(n_690) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
OR2x2_ASAP7_75t_L g246 ( .A(n_247), .B(n_259), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_248), .B(n_285), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_248), .B(n_358), .Y(n_357) );
AOI21xp5_ASAP7_75t_L g461 ( .A1(n_248), .A2(n_374), .B(n_420), .Y(n_461) );
INVx1_ASAP7_75t_L g351 ( .A(n_249), .Y(n_351) );
INVx3_ASAP7_75t_L g369 ( .A(n_249), .Y(n_369) );
AND2x2_ASAP7_75t_L g509 ( .A(n_249), .B(n_281), .Y(n_509) );
INVx2_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
INVx1_ASAP7_75t_L g365 ( .A(n_250), .Y(n_365) );
OAI21x1_ASAP7_75t_L g250 ( .A1(n_251), .A2(n_252), .B(n_258), .Y(n_250) );
INVx1_ASAP7_75t_L g313 ( .A(n_252), .Y(n_313) );
OA22x2_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_254), .B1(n_255), .B2(n_257), .Y(n_252) );
OAI22xp5_ASAP7_75t_L g535 ( .A1(n_253), .A2(n_536), .B1(n_538), .B2(n_542), .Y(n_535) );
INVx4_ASAP7_75t_L g541 ( .A(n_253), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_253), .B(n_580), .Y(n_579) );
AOI21xp5_ASAP7_75t_L g611 ( .A1(n_253), .A2(n_612), .B(n_613), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_257), .B(n_580), .Y(n_585) );
INVx1_ASAP7_75t_L g673 ( .A(n_257), .Y(n_673) );
INVx1_ASAP7_75t_L g316 ( .A(n_258), .Y(n_316) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_260), .B(n_407), .Y(n_489) );
OAI22x1_ASAP7_75t_L g261 ( .A1(n_262), .A2(n_268), .B1(n_275), .B2(n_279), .Y(n_261) );
OR2x2_ASAP7_75t_L g332 ( .A(n_262), .B(n_333), .Y(n_332) );
OR2x2_ASAP7_75t_L g399 ( .A(n_262), .B(n_400), .Y(n_399) );
OR2x2_ASAP7_75t_L g454 ( .A(n_262), .B(n_338), .Y(n_454) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g376 ( .A(n_263), .B(n_334), .Y(n_376) );
INVx1_ASAP7_75t_L g504 ( .A(n_263), .Y(n_504) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
NAND3xp33_ASAP7_75t_L g631 ( .A(n_267), .B(n_574), .C(n_632), .Y(n_631) );
OR2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_271), .Y(n_268) );
INVxp67_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_270), .B(n_365), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_272), .B(n_274), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
INVx2_ASAP7_75t_L g282 ( .A(n_273), .Y(n_282) );
INVx1_ASAP7_75t_L g348 ( .A(n_274), .Y(n_348) );
OAI221xp5_ASAP7_75t_L g448 ( .A1(n_275), .A2(n_379), .B1(n_394), .B2(n_449), .C(n_451), .Y(n_448) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
AND2x4_ASAP7_75t_L g336 ( .A(n_278), .B(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g360 ( .A(n_278), .B(n_361), .Y(n_360) );
AND2x4_ASAP7_75t_L g380 ( .A(n_280), .B(n_364), .Y(n_380) );
NAND2x1p5_ASAP7_75t_L g495 ( .A(n_280), .B(n_472), .Y(n_495) );
AND2x4_ASAP7_75t_L g280 ( .A(n_281), .B(n_282), .Y(n_280) );
AND2x4_ASAP7_75t_L g383 ( .A(n_282), .B(n_312), .Y(n_383) );
OA21x2_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_304), .B(n_306), .Y(n_283) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
OR2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
BUFx2_ASAP7_75t_L g358 ( .A(n_287), .Y(n_358) );
AND2x4_ASAP7_75t_L g328 ( .A(n_288), .B(n_329), .Y(n_328) );
INVx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
HB1xp67_ASAP7_75t_L g321 ( .A(n_289), .Y(n_321) );
INVx2_ASAP7_75t_L g334 ( .A(n_289), .Y(n_334) );
AND2x2_ASAP7_75t_L g361 ( .A(n_289), .B(n_344), .Y(n_361) );
AND2x2_ASAP7_75t_L g386 ( .A(n_289), .B(n_387), .Y(n_386) );
BUFx2_ASAP7_75t_R g501 ( .A(n_289), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_305), .B(n_386), .Y(n_416) );
NAND4xp75_ASAP7_75t_L g306 ( .A(n_307), .B(n_310), .C(n_317), .D(n_319), .Y(n_306) );
INVx2_ASAP7_75t_SL g307 ( .A(n_308), .Y(n_307) );
OR2x2_ASAP7_75t_L g330 ( .A(n_308), .B(n_331), .Y(n_330) );
INVx2_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_309), .B(n_369), .Y(n_450) );
OAI32xp33_ASAP7_75t_L g398 ( .A1(n_310), .A2(n_399), .A3(n_401), .B1(n_403), .B2(n_404), .Y(n_398) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx2_ASAP7_75t_L g331 ( .A(n_311), .Y(n_331) );
AOI21xp5_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_314), .B(n_316), .Y(n_312) );
OR2x2_ASAP7_75t_L g605 ( .A(n_314), .B(n_606), .Y(n_605) );
NOR2xp67_ASAP7_75t_SL g676 ( .A(n_314), .B(n_677), .Y(n_676) );
INVx3_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
OA21x2_ASAP7_75t_L g533 ( .A1(n_315), .A2(n_534), .B(n_550), .Y(n_533) );
OA21x2_ASAP7_75t_L g659 ( .A1(n_315), .A2(n_534), .B(n_550), .Y(n_659) );
INVx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AND3x1_ASAP7_75t_L g446 ( .A(n_320), .B(n_429), .C(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_323), .B(n_352), .Y(n_322) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_328), .Y(n_325) );
INVx2_ASAP7_75t_SL g326 ( .A(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g480 ( .A(n_327), .Y(n_480) );
AND2x2_ASAP7_75t_L g428 ( .A(n_328), .B(n_348), .Y(n_428) );
AND2x2_ASAP7_75t_L g355 ( .A(n_329), .B(n_344), .Y(n_355) );
INVx1_ASAP7_75t_L g483 ( .A(n_329), .Y(n_483) );
NOR2xp33_ASAP7_75t_L g339 ( .A(n_331), .B(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g436 ( .A(n_331), .B(n_402), .Y(n_436) );
AND2x2_ASAP7_75t_L g478 ( .A(n_331), .B(n_374), .Y(n_478) );
HB1xp67_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g460 ( .A(n_334), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g335 ( .A1(n_336), .A2(n_339), .B1(n_341), .B2(n_346), .Y(n_335) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx2_ASAP7_75t_L g403 ( .A(n_341), .Y(n_403) );
INVx2_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
OR2x2_ASAP7_75t_L g342 ( .A(n_343), .B(n_345), .Y(n_342) );
INVx1_ASAP7_75t_L g372 ( .A(n_343), .Y(n_372) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g356 ( .A(n_345), .Y(n_356) );
NOR2x1_ASAP7_75t_L g346 ( .A(n_347), .B(n_349), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
OR2x2_ASAP7_75t_L g396 ( .A(n_348), .B(n_397), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_348), .B(n_349), .Y(n_456) );
INVxp67_ASAP7_75t_SL g452 ( .A(n_349), .Y(n_452) );
INVx3_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g447 ( .A(n_350), .B(n_358), .Y(n_447) );
NOR3xp33_ASAP7_75t_L g469 ( .A(n_350), .B(n_465), .C(n_470), .Y(n_469) );
OAI221xp5_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_357), .B1(n_359), .B2(n_362), .C(n_366), .Y(n_352) );
INVxp67_ASAP7_75t_SL g353 ( .A(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_355), .B(n_356), .Y(n_354) );
AND2x2_ASAP7_75t_L g458 ( .A(n_355), .B(n_459), .Y(n_458) );
OAI22xp5_ASAP7_75t_L g455 ( .A1(n_359), .A2(n_456), .B1(n_457), .B2(n_461), .Y(n_455) );
INVx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g400 ( .A(n_361), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_363), .B(n_364), .Y(n_362) );
INVx1_ASAP7_75t_L g421 ( .A(n_363), .Y(n_421) );
NOR2xp67_ASAP7_75t_L g439 ( .A(n_363), .B(n_440), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_364), .B(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
AOI22xp5_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_371), .B1(n_374), .B2(n_376), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_369), .B(n_370), .Y(n_368) );
INVx3_ASAP7_75t_L g408 ( .A(n_369), .Y(n_408) );
AND2x2_ASAP7_75t_L g492 ( .A(n_369), .B(n_485), .Y(n_492) );
AND2x2_ASAP7_75t_L g506 ( .A(n_369), .B(n_382), .Y(n_506) );
AND2x2_ASAP7_75t_L g418 ( .A(n_370), .B(n_408), .Y(n_418) );
AND2x2_ASAP7_75t_L g371 ( .A(n_372), .B(n_373), .Y(n_371) );
OR2x2_ASAP7_75t_L g474 ( .A(n_372), .B(n_385), .Y(n_474) );
BUFx2_ASAP7_75t_L g393 ( .A(n_373), .Y(n_393) );
AND2x2_ASAP7_75t_L g476 ( .A(n_374), .B(n_383), .Y(n_476) );
INVx2_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AOI221xp5_ASAP7_75t_L g377 ( .A1(n_378), .A2(n_384), .B1(n_391), .B2(n_395), .C(n_398), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_379), .B(n_381), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_382), .B(n_383), .Y(n_381) );
INVx2_ASAP7_75t_L g397 ( .A(n_383), .Y(n_397) );
INVx2_ASAP7_75t_SL g466 ( .A(n_383), .Y(n_466) );
NOR2xp33_ASAP7_75t_L g384 ( .A(n_385), .B(n_388), .Y(n_384) );
OR2x2_ASAP7_75t_L g441 ( .A(n_385), .B(n_388), .Y(n_441) );
INVx2_ASAP7_75t_SL g385 ( .A(n_386), .Y(n_385) );
AND2x4_ASAP7_75t_L g409 ( .A(n_386), .B(n_410), .Y(n_409) );
INVxp67_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVxp67_ASAP7_75t_SL g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
BUFx3_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_403), .B(n_432), .Y(n_431) );
AND2x2_ASAP7_75t_L g427 ( .A(n_408), .B(n_428), .Y(n_427) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_408), .B(n_471), .Y(n_470) );
OAI21xp5_ASAP7_75t_L g442 ( .A1(n_409), .A2(n_424), .B(n_443), .Y(n_442) );
INVx2_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
BUFx2_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
OAI22xp5_ASAP7_75t_L g415 ( .A1(n_416), .A2(n_417), .B1(n_419), .B2(n_423), .Y(n_415) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
AND2x4_ASAP7_75t_L g420 ( .A(n_421), .B(n_422), .Y(n_420) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
NAND4xp25_ASAP7_75t_L g425 ( .A(n_426), .B(n_445), .C(n_462), .D(n_487), .Y(n_425) );
AOI221x1_ASAP7_75t_L g426 ( .A1(n_427), .A2(n_429), .B1(n_431), .B2(n_435), .C(n_437), .Y(n_426) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
OAI21xp5_ASAP7_75t_L g437 ( .A1(n_438), .A2(n_441), .B(n_442), .Y(n_437) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
NOR3xp33_ASAP7_75t_L g445 ( .A(n_446), .B(n_448), .C(n_455), .Y(n_445) );
BUFx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_452), .B(n_453), .Y(n_451) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
OAI21xp33_ASAP7_75t_SL g463 ( .A1(n_457), .A2(n_464), .B(n_467), .Y(n_463) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
HB1xp67_ASAP7_75t_L g493 ( .A(n_459), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_460), .B(n_483), .Y(n_482) );
AOI21xp33_ASAP7_75t_L g462 ( .A1(n_463), .A2(n_468), .B(n_473), .Y(n_462) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVxp67_ASAP7_75t_SL g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
OAI221xp5_ASAP7_75t_L g473 ( .A1(n_474), .A2(n_475), .B1(n_477), .B2(n_479), .C(n_484), .Y(n_473) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx2_ASAP7_75t_SL g477 ( .A(n_478), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_480), .B(n_481), .Y(n_479) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_485), .B(n_486), .Y(n_484) );
O2A1O1Ixp5_ASAP7_75t_L g487 ( .A1(n_488), .A2(n_490), .B(n_493), .C(n_494), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
OAI211xp5_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_496), .B(n_498), .C(n_507), .Y(n_494) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
OAI21xp5_ASAP7_75t_L g498 ( .A1(n_499), .A2(n_502), .B(n_506), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
OR2x2_ASAP7_75t_L g503 ( .A(n_504), .B(n_505), .Y(n_503) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
CKINVDCx5p33_ASAP7_75t_R g512 ( .A(n_513), .Y(n_512) );
INVx2_ASAP7_75t_L g931 ( .A(n_513), .Y(n_931) );
OR2x6_ASAP7_75t_L g513 ( .A(n_514), .B(n_515), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g920 ( .A(n_515), .B(n_921), .Y(n_920) );
INVx8_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
AND2x2_ASAP7_75t_L g523 ( .A(n_516), .B(n_524), .Y(n_523) );
OR2x6_ASAP7_75t_L g926 ( .A(n_516), .B(n_524), .Y(n_926) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_518), .B(n_519), .Y(n_517) );
NAND2xp33_ASAP7_75t_L g520 ( .A(n_521), .B(n_525), .Y(n_520) );
BUFx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
HB1xp67_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx2_ASAP7_75t_L g936 ( .A(n_523), .Y(n_936) );
INVx2_ASAP7_75t_L g935 ( .A(n_525), .Y(n_935) );
XNOR2xp5_ASAP7_75t_L g942 ( .A(n_525), .B(n_943), .Y(n_942) );
NAND3x1_ASAP7_75t_L g525 ( .A(n_526), .B(n_777), .C(n_853), .Y(n_525) );
NOR2x1_ASAP7_75t_L g526 ( .A(n_527), .B(n_706), .Y(n_526) );
NAND3xp33_ASAP7_75t_L g527 ( .A(n_528), .B(n_660), .C(n_686), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
OAI22xp5_ASAP7_75t_L g529 ( .A1(n_530), .A2(n_592), .B1(n_651), .B2(n_655), .Y(n_529) );
OR2x2_ASAP7_75t_L g530 ( .A(n_531), .B(n_554), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g875 ( .A(n_531), .B(n_725), .Y(n_875) );
AND3x2_ASAP7_75t_L g881 ( .A(n_531), .B(n_657), .C(n_761), .Y(n_881) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
AND2x2_ASAP7_75t_L g714 ( .A(n_532), .B(n_669), .Y(n_714) );
AND2x2_ASAP7_75t_L g751 ( .A(n_532), .B(n_577), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g829 ( .A(n_532), .B(n_794), .Y(n_829) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx2_ASAP7_75t_L g701 ( .A(n_533), .Y(n_701) );
INVx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_539), .B(n_541), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
OAI22x1_ASAP7_75t_L g670 ( .A1(n_541), .A2(n_671), .B1(n_673), .B2(n_674), .Y(n_670) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_545), .A2(n_547), .B(n_549), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_546), .B(n_642), .Y(n_641) );
AOI22xp5_ASAP7_75t_L g644 ( .A1(n_546), .A2(n_548), .B1(n_645), .B2(n_647), .Y(n_644) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
OR2x2_ASAP7_75t_L g628 ( .A(n_552), .B(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_555), .B(n_577), .Y(n_554) );
INVx1_ASAP7_75t_L g912 ( .A(n_555), .Y(n_912) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVxp67_ASAP7_75t_L g657 ( .A(n_556), .Y(n_657) );
AND2x2_ASAP7_75t_L g667 ( .A(n_556), .B(n_668), .Y(n_667) );
INVx2_ASAP7_75t_L g713 ( .A(n_556), .Y(n_713) );
AO21x2_ASAP7_75t_L g556 ( .A1(n_557), .A2(n_565), .B(n_573), .Y(n_556) );
AO21x2_ASAP7_75t_L g693 ( .A1(n_557), .A2(n_565), .B(n_573), .Y(n_693) );
OAI21x1_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_561), .B(n_564), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_559), .B(n_639), .Y(n_638) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx2_ASAP7_75t_L g583 ( .A(n_563), .Y(n_583) );
OAI21x1_ASAP7_75t_SL g565 ( .A1(n_566), .A2(n_567), .B(n_571), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_568), .B(n_570), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_570), .B(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g576 ( .A(n_570), .Y(n_576) );
AOI21x1_ASAP7_75t_L g602 ( .A1(n_572), .A2(n_603), .B(n_604), .Y(n_602) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g658 ( .A(n_577), .B(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g698 ( .A(n_577), .Y(n_698) );
INVx1_ASAP7_75t_L g738 ( .A(n_577), .Y(n_738) );
INVx2_ASAP7_75t_L g794 ( .A(n_577), .Y(n_794) );
NAND2x1p5_ASAP7_75t_L g577 ( .A(n_578), .B(n_584), .Y(n_577) );
AND2x2_ASAP7_75t_L g665 ( .A(n_578), .B(n_584), .Y(n_665) );
OR2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_582), .Y(n_578) );
OA21x2_ASAP7_75t_L g584 ( .A1(n_585), .A2(n_586), .B(n_589), .Y(n_584) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g627 ( .A(n_588), .Y(n_627) );
INVx1_ASAP7_75t_L g675 ( .A(n_590), .Y(n_675) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
INVx2_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_594), .B(n_620), .Y(n_593) );
INVx2_ASAP7_75t_L g721 ( .A(n_594), .Y(n_721) );
AND2x4_ASAP7_75t_L g757 ( .A(n_594), .B(n_758), .Y(n_757) );
AND2x2_ASAP7_75t_L g843 ( .A(n_594), .B(n_742), .Y(n_843) );
AND2x2_ASAP7_75t_L g594 ( .A(n_595), .B(n_607), .Y(n_594) );
AND2x2_ASAP7_75t_L g653 ( .A(n_595), .B(n_608), .Y(n_653) );
INVx2_ASAP7_75t_SL g685 ( .A(n_595), .Y(n_685) );
OAI21x1_ASAP7_75t_L g595 ( .A1(n_596), .A2(n_597), .B(n_605), .Y(n_595) );
OAI21xp5_ASAP7_75t_L g800 ( .A1(n_596), .A2(n_597), .B(n_605), .Y(n_800) );
AOI21x1_ASAP7_75t_L g597 ( .A1(n_598), .A2(n_599), .B(n_602), .Y(n_597) );
INVx2_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g730 ( .A(n_607), .Y(n_730) );
AND2x2_ASAP7_75t_L g852 ( .A(n_607), .B(n_621), .Y(n_852) );
INVx3_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx2_ASAP7_75t_L g681 ( .A(n_608), .Y(n_681) );
AND2x2_ASAP7_75t_L g773 ( .A(n_608), .B(n_685), .Y(n_773) );
AND2x4_ASAP7_75t_L g608 ( .A(n_609), .B(n_610), .Y(n_608) );
OAI21x1_ASAP7_75t_L g610 ( .A1(n_611), .A2(n_614), .B(n_619), .Y(n_610) );
INVx2_ASAP7_75t_L g654 ( .A(n_620), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_620), .B(n_764), .Y(n_763) );
HB1xp67_ASAP7_75t_L g808 ( .A(n_620), .Y(n_808) );
NAND2xp5_ASAP7_75t_L g906 ( .A(n_620), .B(n_907), .Y(n_906) );
AND2x2_ASAP7_75t_L g620 ( .A(n_621), .B(n_634), .Y(n_620) );
INVx1_ASAP7_75t_L g682 ( .A(n_621), .Y(n_682) );
INVx1_ASAP7_75t_L g720 ( .A(n_621), .Y(n_720) );
INVx1_ASAP7_75t_L g728 ( .A(n_621), .Y(n_728) );
INVx2_ASAP7_75t_L g743 ( .A(n_621), .Y(n_743) );
NOR2x1_ASAP7_75t_L g758 ( .A(n_621), .B(n_759), .Y(n_758) );
AND2x2_ASAP7_75t_L g769 ( .A(n_621), .B(n_635), .Y(n_769) );
OR2x6_ASAP7_75t_L g621 ( .A(n_622), .B(n_630), .Y(n_621) );
OAI21x1_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_624), .B(n_628), .Y(n_622) );
INVx2_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
NOR2xp67_ASAP7_75t_L g630 ( .A(n_631), .B(n_633), .Y(n_630) );
AND2x2_ASAP7_75t_L g742 ( .A(n_634), .B(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g684 ( .A(n_635), .B(n_685), .Y(n_684) );
INVxp67_ASAP7_75t_L g705 ( .A(n_635), .Y(n_705) );
INVx1_ASAP7_75t_L g754 ( .A(n_635), .Y(n_754) );
INVx1_ASAP7_75t_L g759 ( .A(n_635), .Y(n_759) );
OR2x2_ASAP7_75t_L g799 ( .A(n_635), .B(n_800), .Y(n_799) );
AO21x2_ASAP7_75t_L g635 ( .A1(n_636), .A2(n_637), .B(n_649), .Y(n_635) );
NAND3xp33_ASAP7_75t_SL g637 ( .A(n_638), .B(n_641), .C(n_644), .Y(n_637) );
NAND2xp33_ASAP7_75t_SL g824 ( .A(n_651), .B(n_825), .Y(n_824) );
OR2x2_ASAP7_75t_L g651 ( .A(n_652), .B(n_654), .Y(n_651) );
INVx2_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
AND2x2_ASAP7_75t_L g776 ( .A(n_653), .B(n_769), .Y(n_776) );
AND2x2_ASAP7_75t_L g791 ( .A(n_653), .B(n_719), .Y(n_791) );
AND2x2_ASAP7_75t_L g804 ( .A(n_653), .B(n_805), .Y(n_804) );
HB1xp67_ASAP7_75t_L g899 ( .A(n_654), .Y(n_899) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_655), .B(n_662), .Y(n_661) );
INVx2_ASAP7_75t_SL g655 ( .A(n_656), .Y(n_655) );
AND2x2_ASAP7_75t_L g656 ( .A(n_657), .B(n_658), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_658), .B(n_716), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g848 ( .A(n_658), .B(n_849), .Y(n_848) );
AND2x2_ASAP7_75t_L g908 ( .A(n_658), .B(n_909), .Y(n_908) );
AND2x2_ASAP7_75t_L g664 ( .A(n_659), .B(n_665), .Y(n_664) );
AND2x2_ASAP7_75t_L g692 ( .A(n_659), .B(n_693), .Y(n_692) );
NAND2x1_ASAP7_75t_L g735 ( .A(n_659), .B(n_668), .Y(n_735) );
NAND2xp5_ASAP7_75t_SL g660 ( .A(n_661), .B(n_678), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_663), .B(n_666), .Y(n_662) );
HB1xp67_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
AND2x4_ASAP7_75t_L g724 ( .A(n_664), .B(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g817 ( .A(n_664), .Y(n_817) );
AND2x2_ASAP7_75t_L g837 ( .A(n_664), .B(n_716), .Y(n_837) );
INVx2_ASAP7_75t_SL g695 ( .A(n_665), .Y(n_695) );
BUFx3_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_667), .B(n_811), .Y(n_810) );
AND2x2_ASAP7_75t_L g867 ( .A(n_667), .B(n_761), .Y(n_867) );
AOI32xp33_ASAP7_75t_L g877 ( .A1(n_667), .A2(n_798), .A3(n_878), .B1(n_879), .B2(n_881), .Y(n_877) );
INVx2_ASAP7_75t_L g703 ( .A(n_668), .Y(n_703) );
INVx1_ASAP7_75t_L g909 ( .A(n_668), .Y(n_909) );
INVx3_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
OAI321xp33_ASAP7_75t_L g896 ( .A1(n_679), .A2(n_897), .A3(n_899), .B1(n_900), .B2(n_902), .C(n_903), .Y(n_896) );
NAND2x2_ASAP7_75t_L g679 ( .A(n_680), .B(n_683), .Y(n_679) );
AND2x2_ASAP7_75t_L g860 ( .A(n_680), .B(n_798), .Y(n_860) );
AND2x2_ASAP7_75t_L g680 ( .A(n_681), .B(n_682), .Y(n_680) );
NOR2xp33_ASAP7_75t_L g704 ( .A(n_681), .B(n_705), .Y(n_704) );
INVx2_ASAP7_75t_L g741 ( .A(n_681), .Y(n_741) );
HB1xp67_ASAP7_75t_L g797 ( .A(n_681), .Y(n_797) );
OR2x2_ASAP7_75t_L g816 ( .A(n_681), .B(n_799), .Y(n_816) );
OR2x2_ASAP7_75t_L g839 ( .A(n_682), .B(n_721), .Y(n_839) );
AND2x2_ASAP7_75t_L g887 ( .A(n_682), .B(n_773), .Y(n_887) );
BUFx3_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_684), .B(n_728), .Y(n_747) );
AND2x4_ASAP7_75t_L g851 ( .A(n_684), .B(n_852), .Y(n_851) );
INVx1_ASAP7_75t_L g731 ( .A(n_685), .Y(n_731) );
INVx1_ASAP7_75t_L g764 ( .A(n_685), .Y(n_764) );
OAI21xp5_ASAP7_75t_L g686 ( .A1(n_687), .A2(n_696), .B(n_704), .Y(n_686) );
AND2x2_ASAP7_75t_L g687 ( .A(n_688), .B(n_691), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g832 ( .A(n_689), .B(n_701), .Y(n_832) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
OR2x2_ASAP7_75t_L g717 ( .A(n_690), .B(n_693), .Y(n_717) );
AND2x4_ASAP7_75t_L g725 ( .A(n_690), .B(n_713), .Y(n_725) );
AND2x2_ASAP7_75t_L g739 ( .A(n_690), .B(n_693), .Y(n_739) );
INVx2_ASAP7_75t_L g774 ( .A(n_691), .Y(n_774) );
AND2x2_ASAP7_75t_L g691 ( .A(n_692), .B(n_694), .Y(n_691) );
INVx2_ASAP7_75t_L g822 ( .A(n_692), .Y(n_822) );
AND2x2_ASAP7_75t_L g840 ( .A(n_692), .B(n_702), .Y(n_840) );
AND2x4_ASAP7_75t_L g700 ( .A(n_693), .B(n_701), .Y(n_700) );
INVx2_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
OR2x2_ASAP7_75t_L g734 ( .A(n_695), .B(n_735), .Y(n_734) );
INVx2_ASAP7_75t_L g761 ( .A(n_695), .Y(n_761) );
AND2x2_ASAP7_75t_L g823 ( .A(n_695), .B(n_703), .Y(n_823) );
AND2x2_ASAP7_75t_L g696 ( .A(n_697), .B(n_699), .Y(n_696) );
AND2x2_ASAP7_75t_L g878 ( .A(n_697), .B(n_752), .Y(n_878) );
INVx2_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
AOI221xp5_ASAP7_75t_L g756 ( .A1(n_699), .A2(n_757), .B1(n_760), .B2(n_762), .C(n_765), .Y(n_756) );
AND2x2_ASAP7_75t_L g699 ( .A(n_700), .B(n_702), .Y(n_699) );
AND2x2_ASAP7_75t_L g793 ( .A(n_700), .B(n_794), .Y(n_793) );
BUFx3_ASAP7_75t_L g834 ( .A(n_700), .Y(n_834) );
INVxp67_ASAP7_75t_SL g857 ( .A(n_701), .Y(n_857) );
INVx1_ASAP7_75t_L g889 ( .A(n_702), .Y(n_889) );
INVx2_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g782 ( .A(n_703), .Y(n_782) );
AND2x2_ASAP7_75t_L g885 ( .A(n_704), .B(n_864), .Y(n_885) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_707), .B(n_756), .Y(n_706) );
NOR3xp33_ASAP7_75t_L g707 ( .A(n_708), .B(n_722), .C(n_744), .Y(n_707) );
NOR2xp33_ASAP7_75t_L g708 ( .A(n_709), .B(n_718), .Y(n_708) );
AND2x2_ASAP7_75t_L g709 ( .A(n_710), .B(n_715), .Y(n_709) );
OAI21xp33_ASAP7_75t_L g744 ( .A1(n_710), .A2(n_745), .B(n_748), .Y(n_744) );
NAND2x1p5_ASAP7_75t_L g710 ( .A(n_711), .B(n_714), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g902 ( .A(n_714), .Y(n_902) );
INVx2_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx2_ASAP7_75t_L g767 ( .A(n_717), .Y(n_767) );
INVx1_ASAP7_75t_L g819 ( .A(n_718), .Y(n_819) );
OR2x2_ASAP7_75t_SL g718 ( .A(n_719), .B(n_721), .Y(n_718) );
INVx2_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
AND2x2_ASAP7_75t_L g904 ( .A(n_720), .B(n_895), .Y(n_904) );
OR2x2_ASAP7_75t_L g785 ( .A(n_721), .B(n_786), .Y(n_785) );
OAI21xp33_ASAP7_75t_L g722 ( .A1(n_723), .A2(n_726), .B(n_732), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
BUFx3_ASAP7_75t_L g755 ( .A(n_725), .Y(n_755) );
AND2x2_ASAP7_75t_L g760 ( .A(n_725), .B(n_761), .Y(n_760) );
NOR2xp67_ASAP7_75t_L g789 ( .A(n_725), .B(n_750), .Y(n_789) );
INVx3_ASAP7_75t_L g849 ( .A(n_725), .Y(n_849) );
OR2x2_ASAP7_75t_L g726 ( .A(n_727), .B(n_729), .Y(n_726) );
HB1xp67_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
AND2x2_ASAP7_75t_L g864 ( .A(n_728), .B(n_865), .Y(n_864) );
OR2x2_ASAP7_75t_L g729 ( .A(n_730), .B(n_731), .Y(n_729) );
INVx1_ASAP7_75t_L g752 ( .A(n_730), .Y(n_752) );
INVxp67_ASAP7_75t_SL g814 ( .A(n_731), .Y(n_814) );
OAI21xp33_ASAP7_75t_L g732 ( .A1(n_733), .A2(n_736), .B(n_740), .Y(n_732) );
INVx2_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
AND2x2_ASAP7_75t_L g736 ( .A(n_737), .B(n_739), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g805 ( .A(n_738), .Y(n_805) );
INVx1_ASAP7_75t_L g883 ( .A(n_738), .Y(n_883) );
NOR3xp33_ASAP7_75t_L g845 ( .A(n_739), .B(n_767), .C(n_823), .Y(n_845) );
INVx2_ASAP7_75t_L g884 ( .A(n_739), .Y(n_884) );
AOI22xp5_ASAP7_75t_L g886 ( .A1(n_739), .A2(n_887), .B1(n_888), .B2(n_891), .Y(n_886) );
AND2x2_ASAP7_75t_L g901 ( .A(n_739), .B(n_761), .Y(n_901) );
INVx2_ASAP7_75t_L g870 ( .A(n_740), .Y(n_870) );
AND2x2_ASAP7_75t_L g740 ( .A(n_741), .B(n_742), .Y(n_740) );
AND2x2_ASAP7_75t_L g863 ( .A(n_741), .B(n_754), .Y(n_863) );
INVx1_ASAP7_75t_L g907 ( .A(n_741), .Y(n_907) );
AND2x2_ASAP7_75t_L g847 ( .A(n_742), .B(n_773), .Y(n_847) );
INVx1_ASAP7_75t_L g880 ( .A(n_742), .Y(n_880) );
OAI21xp33_ASAP7_75t_L g910 ( .A1(n_745), .A2(n_911), .B(n_913), .Y(n_910) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
NAND4xp25_ASAP7_75t_L g748 ( .A(n_749), .B(n_752), .C(n_753), .D(n_755), .Y(n_748) );
INVx2_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx2_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx1_ASAP7_75t_L g783 ( .A(n_751), .Y(n_783) );
INVx1_ASAP7_75t_L g898 ( .A(n_752), .Y(n_898) );
INVx2_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx2_ASAP7_75t_L g825 ( .A(n_757), .Y(n_825) );
NAND2x1_ASAP7_75t_L g766 ( .A(n_761), .B(n_767), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g913 ( .A(n_762), .B(n_793), .Y(n_913) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
OAI32xp33_ASAP7_75t_L g765 ( .A1(n_766), .A2(n_768), .A3(n_770), .B1(n_774), .B2(n_775), .Y(n_765) );
INVx1_ASAP7_75t_L g779 ( .A(n_766), .Y(n_779) );
A2O1A1Ixp33_ASAP7_75t_L g882 ( .A1(n_767), .A2(n_883), .B(n_884), .C(n_885), .Y(n_882) );
HB1xp67_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
INVx1_ASAP7_75t_L g786 ( .A(n_769), .Y(n_786) );
AND2x2_ASAP7_75t_L g813 ( .A(n_769), .B(n_814), .Y(n_813) );
NAND2x1_ASAP7_75t_SL g835 ( .A(n_769), .B(n_773), .Y(n_835) );
NAND2xp5_ASAP7_75t_L g871 ( .A(n_769), .B(n_872), .Y(n_871) );
INVx1_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVx1_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
INVx2_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
INVx2_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
AND4x1_ASAP7_75t_L g777 ( .A(n_778), .B(n_801), .C(n_818), .D(n_836), .Y(n_777) );
O2A1O1Ixp5_ASAP7_75t_L g778 ( .A1(n_779), .A2(n_780), .B(n_784), .C(n_787), .Y(n_778) );
INVx1_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
OR2x2_ASAP7_75t_L g781 ( .A(n_782), .B(n_783), .Y(n_781) );
NAND2xp5_ASAP7_75t_SL g803 ( .A(n_782), .B(n_804), .Y(n_803) );
INVx2_ASAP7_75t_SL g784 ( .A(n_785), .Y(n_784) );
OAI22xp5_ASAP7_75t_L g787 ( .A1(n_788), .A2(n_790), .B1(n_792), .B2(n_795), .Y(n_787) );
INVx1_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
INVx1_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
INVx2_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
INVx1_ASAP7_75t_L g811 ( .A(n_794), .Y(n_811) );
INVx1_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
AND2x2_ASAP7_75t_L g796 ( .A(n_797), .B(n_798), .Y(n_796) );
INVx1_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
INVx2_ASAP7_75t_L g895 ( .A(n_799), .Y(n_895) );
BUFx2_ASAP7_75t_L g865 ( .A(n_800), .Y(n_865) );
AOI21xp5_ASAP7_75t_L g801 ( .A1(n_802), .A2(n_806), .B(n_809), .Y(n_801) );
INVx1_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
OR2x2_ASAP7_75t_L g831 ( .A(n_805), .B(n_832), .Y(n_831) );
INVx1_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
INVx1_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
OAI22xp5_ASAP7_75t_SL g809 ( .A1(n_810), .A2(n_812), .B1(n_815), .B2(n_817), .Y(n_809) );
INVx1_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
HB1xp67_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
AOI221xp5_ASAP7_75t_L g818 ( .A1(n_819), .A2(n_820), .B1(n_824), .B2(n_826), .C(n_830), .Y(n_818) );
AND2x4_ASAP7_75t_L g820 ( .A(n_821), .B(n_823), .Y(n_820) );
INVx1_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
INVx1_ASAP7_75t_L g890 ( .A(n_822), .Y(n_890) );
INVx1_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
INVx1_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
INVx1_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
OR2x2_ASAP7_75t_L g911 ( .A(n_829), .B(n_912), .Y(n_911) );
AOI21xp33_ASAP7_75t_SL g830 ( .A1(n_831), .A2(n_833), .B(n_835), .Y(n_830) );
INVx2_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
AOI221xp5_ASAP7_75t_L g836 ( .A1(n_837), .A2(n_838), .B1(n_840), .B2(n_841), .C(n_844), .Y(n_836) );
INVx1_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
INVx1_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
INVx2_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
OAI22xp33_ASAP7_75t_L g844 ( .A1(n_845), .A2(n_846), .B1(n_848), .B2(n_850), .Y(n_844) );
INVx2_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
INVx1_ASAP7_75t_L g858 ( .A(n_849), .Y(n_858) );
INVx2_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
INVx2_ASAP7_75t_L g893 ( .A(n_852), .Y(n_893) );
NOR4xp25_ASAP7_75t_L g853 ( .A(n_854), .B(n_876), .C(n_896), .D(n_910), .Y(n_853) );
OAI322xp33_ASAP7_75t_L g854 ( .A1(n_855), .A2(n_858), .A3(n_859), .B1(n_861), .B2(n_866), .C1(n_868), .C2(n_874), .Y(n_854) );
INVx1_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
INVx1_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
INVx1_ASAP7_75t_L g859 ( .A(n_860), .Y(n_859) );
INVx1_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
AND2x2_ASAP7_75t_L g862 ( .A(n_863), .B(n_864), .Y(n_862) );
INVx1_ASAP7_75t_L g873 ( .A(n_865), .Y(n_873) );
INVx1_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
INVx1_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
NAND2xp5_ASAP7_75t_L g869 ( .A(n_870), .B(n_871), .Y(n_869) );
INVxp67_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
HB1xp67_ASAP7_75t_L g874 ( .A(n_875), .Y(n_874) );
NAND3xp33_ASAP7_75t_SL g876 ( .A(n_877), .B(n_882), .C(n_886), .Y(n_876) );
INVx1_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
AND2x2_ASAP7_75t_L g888 ( .A(n_889), .B(n_890), .Y(n_888) );
INVx1_ASAP7_75t_L g891 ( .A(n_892), .Y(n_891) );
OR2x2_ASAP7_75t_L g892 ( .A(n_893), .B(n_894), .Y(n_892) );
INVx1_ASAP7_75t_L g894 ( .A(n_895), .Y(n_894) );
INVx1_ASAP7_75t_L g897 ( .A(n_898), .Y(n_897) );
INVx1_ASAP7_75t_L g900 ( .A(n_901), .Y(n_900) );
OAI21xp5_ASAP7_75t_L g903 ( .A1(n_904), .A2(n_905), .B(n_908), .Y(n_903) );
INVx1_ASAP7_75t_L g905 ( .A(n_906), .Y(n_905) );
AOI21x1_ASAP7_75t_L g939 ( .A1(n_914), .A2(n_940), .B(n_941), .Y(n_939) );
NOR2xp67_ASAP7_75t_SL g914 ( .A(n_915), .B(n_916), .Y(n_914) );
INVx2_ASAP7_75t_L g916 ( .A(n_917), .Y(n_916) );
INVx5_ASAP7_75t_SL g917 ( .A(n_918), .Y(n_917) );
BUFx6f_ASAP7_75t_L g918 ( .A(n_919), .Y(n_918) );
BUFx8_ASAP7_75t_SL g940 ( .A(n_919), .Y(n_940) );
BUFx6f_ASAP7_75t_L g919 ( .A(n_920), .Y(n_919) );
NOR2xp33_ASAP7_75t_L g922 ( .A(n_923), .B(n_924), .Y(n_922) );
CKINVDCx5p33_ASAP7_75t_R g924 ( .A(n_925), .Y(n_924) );
INVx1_ASAP7_75t_L g925 ( .A(n_926), .Y(n_925) );
OAI22xp5_ASAP7_75t_L g928 ( .A1(n_929), .A2(n_932), .B1(n_934), .B2(n_936), .Y(n_928) );
BUFx12f_ASAP7_75t_L g929 ( .A(n_930), .Y(n_929) );
CKINVDCx11_ASAP7_75t_R g930 ( .A(n_931), .Y(n_930) );
INVx1_ASAP7_75t_L g932 ( .A(n_933), .Y(n_932) );
INVx1_ASAP7_75t_L g934 ( .A(n_935), .Y(n_934) );
NOR2x1_ASAP7_75t_SL g937 ( .A(n_938), .B(n_939), .Y(n_937) );
INVx2_ASAP7_75t_SL g941 ( .A(n_942), .Y(n_941) );
INVx1_ASAP7_75t_SL g946 ( .A(n_947), .Y(n_946) );
BUFx3_ASAP7_75t_L g947 ( .A(n_948), .Y(n_947) );
BUFx3_ASAP7_75t_L g958 ( .A(n_948), .Y(n_958) );
OR2x2_ASAP7_75t_SL g948 ( .A(n_949), .B(n_955), .Y(n_948) );
NAND3xp33_ASAP7_75t_L g949 ( .A(n_950), .B(n_951), .C(n_953), .Y(n_949) );
CKINVDCx5p33_ASAP7_75t_R g951 ( .A(n_952), .Y(n_951) );
CKINVDCx5p33_ASAP7_75t_R g956 ( .A(n_957), .Y(n_956) );
INVx1_ASAP7_75t_L g957 ( .A(n_958), .Y(n_957) );
endmodule