module fake_jpeg_26392_n_202 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_202);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_202;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_9),
.B(n_12),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_6),
.B(n_14),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx6_ASAP7_75t_SL g30 ( 
.A(n_3),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_21),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_32),
.B(n_33),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_21),
.B(n_0),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_34),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_38),
.Y(n_60)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

BUFx4f_ASAP7_75t_SL g40 ( 
.A(n_30),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_40),
.Y(n_46)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_31),
.A2(n_20),
.B1(n_19),
.B2(n_16),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_43),
.A2(n_52),
.B1(n_56),
.B2(n_57),
.Y(n_69)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_25),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_47),
.B(n_54),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_32),
.B(n_33),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_22),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_31),
.A2(n_20),
.B1(n_19),
.B2(n_16),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_39),
.B(n_23),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_39),
.A2(n_20),
.B1(n_23),
.B2(n_18),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_41),
.A2(n_18),
.B1(n_28),
.B2(n_15),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_26),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_37),
.Y(n_73)
);

NAND2xp33_ASAP7_75t_SL g59 ( 
.A(n_37),
.B(n_26),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_59),
.B(n_25),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_61),
.A2(n_47),
.B1(n_59),
.B2(n_48),
.Y(n_84)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_66),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_56),
.A2(n_41),
.B1(n_38),
.B2(n_34),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_65),
.A2(n_72),
.B1(n_43),
.B2(n_52),
.Y(n_81)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_50),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_68),
.B(n_74),
.Y(n_96)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_71),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_R g71 ( 
.A(n_57),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_49),
.A2(n_41),
.B1(n_38),
.B2(n_34),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_73),
.B(n_75),
.Y(n_90)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_54),
.B(n_22),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_77),
.B(n_55),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_73),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_78),
.B(n_80),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_79),
.B(n_81),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_55),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_85),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_84),
.A2(n_45),
.B(n_67),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_68),
.B(n_46),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_47),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_89),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_64),
.B(n_47),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_69),
.A2(n_48),
.B1(n_53),
.B2(n_36),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_91),
.A2(n_93),
.B1(n_62),
.B2(n_45),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_69),
.A2(n_58),
.B1(n_46),
.B2(n_42),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_75),
.B(n_58),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_94),
.B(n_60),
.Y(n_102)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_95),
.B(n_74),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_94),
.B(n_61),
.C(n_70),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_98),
.B(n_99),
.C(n_109),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_44),
.C(n_60),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_102),
.B(n_112),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_103),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_96),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_104),
.B(n_108),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_105),
.A2(n_87),
.B1(n_36),
.B2(n_42),
.Y(n_127)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_106),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_96),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_107),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_86),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_63),
.C(n_66),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_63),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_110),
.B(n_95),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_28),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_111),
.B(n_29),
.Y(n_130)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_91),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_113),
.A2(n_104),
.B(n_115),
.Y(n_126)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_87),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_114),
.B(n_90),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_89),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_116),
.B(n_126),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_117),
.B(n_122),
.Y(n_135)
);

OAI32xp33_ASAP7_75t_L g118 ( 
.A1(n_101),
.A2(n_81),
.A3(n_79),
.B1(n_90),
.B2(n_92),
.Y(n_118)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_118),
.Y(n_134)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_97),
.Y(n_122)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_114),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_124),
.B(n_125),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_92),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_127),
.A2(n_42),
.B1(n_36),
.B2(n_15),
.Y(n_143)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_128),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_130),
.B(n_111),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_102),
.B(n_29),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_131),
.B(n_133),
.Y(n_144)
);

INVx1_ASAP7_75t_SL g133 ( 
.A(n_100),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_129),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_136),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_132),
.B(n_109),
.C(n_99),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_138),
.B(n_140),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_132),
.B(n_113),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_141),
.B(n_148),
.Y(n_150)
);

AOI22x1_ASAP7_75t_L g142 ( 
.A1(n_118),
.A2(n_105),
.B1(n_112),
.B2(n_100),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_142),
.A2(n_146),
.B1(n_128),
.B2(n_123),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g153 ( 
.A(n_143),
.Y(n_153)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_121),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_145),
.B(n_147),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_123),
.A2(n_17),
.B1(n_26),
.B2(n_25),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_116),
.B(n_40),
.C(n_51),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_120),
.B(n_17),
.Y(n_149)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_149),
.Y(n_158)
);

A2O1A1Ixp33_ASAP7_75t_SL g169 ( 
.A1(n_151),
.A2(n_40),
.B(n_51),
.C(n_2),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_139),
.B(n_133),
.Y(n_152)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_152),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_134),
.A2(n_119),
.B1(n_124),
.B2(n_126),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_155),
.A2(n_156),
.B1(n_161),
.B2(n_146),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_142),
.A2(n_119),
.B1(n_130),
.B2(n_27),
.Y(n_156)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_137),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_159),
.B(n_10),
.Y(n_172)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_135),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_160),
.B(n_140),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_144),
.A2(n_27),
.B1(n_14),
.B2(n_13),
.Y(n_161)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_162),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_163),
.B(n_166),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g164 ( 
.A(n_150),
.B(n_147),
.Y(n_164)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_164),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_155),
.A2(n_148),
.B(n_141),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_154),
.B(n_138),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_167),
.B(n_171),
.Y(n_177)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_168),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_169),
.A2(n_153),
.B(n_1),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_160),
.A2(n_157),
.B(n_152),
.Y(n_170)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_170),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_154),
.B(n_51),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_172),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_181)
);

O2A1O1Ixp33_ASAP7_75t_SL g187 ( 
.A1(n_178),
.A2(n_169),
.B(n_5),
.C(n_7),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_165),
.A2(n_156),
.B(n_158),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_179),
.B(n_169),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_168),
.A2(n_150),
.B1(n_10),
.B2(n_3),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_180),
.B(n_172),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_181),
.B(n_178),
.Y(n_188)
);

OR2x2_ASAP7_75t_L g193 ( 
.A(n_183),
.B(n_188),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_180),
.B(n_173),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_184),
.B(n_189),
.Y(n_194)
);

INVx11_ASAP7_75t_L g185 ( 
.A(n_176),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_185),
.B(n_186),
.Y(n_192)
);

OAI21x1_ASAP7_75t_SL g190 ( 
.A1(n_187),
.A2(n_4),
.B(n_7),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_175),
.B(n_4),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_190),
.B(n_191),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_187),
.A2(n_182),
.B(n_174),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_193),
.B(n_177),
.C(n_186),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_195),
.B(n_196),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_192),
.B(n_185),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_197),
.A2(n_194),
.B(n_40),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_199),
.A2(n_4),
.B(n_8),
.Y(n_200)
);

AO21x1_ASAP7_75t_L g201 ( 
.A1(n_200),
.A2(n_198),
.B(n_8),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_201),
.B(n_8),
.Y(n_202)
);


endmodule