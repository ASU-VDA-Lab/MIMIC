module real_aes_1435_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_794, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_794;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_766;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_769;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_288;
wire n_147;
wire n_150;
wire n_404;
wire n_713;
wire n_598;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_785;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_749;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_481;
wire n_148;
wire n_498;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_762;
wire n_210;
wire n_212;
wire n_325;
wire n_575;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_0), .B(n_145), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g175 ( .A1(n_1), .A2(n_154), .B(n_176), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_2), .B(n_110), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_3), .B(n_145), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_4), .B(n_161), .Y(n_534) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_5), .B(n_161), .Y(n_224) );
INVx1_ASAP7_75t_L g152 ( .A(n_6), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_7), .B(n_161), .Y(n_199) );
CKINVDCx16_ASAP7_75t_R g110 ( .A(n_8), .Y(n_110) );
NAND2xp33_ASAP7_75t_L g162 ( .A(n_9), .B(n_163), .Y(n_162) );
AND2x2_ASAP7_75t_L g476 ( .A(n_10), .B(n_171), .Y(n_476) );
AND2x2_ASAP7_75t_L g536 ( .A(n_11), .B(n_140), .Y(n_536) );
INVx2_ASAP7_75t_L g142 ( .A(n_12), .Y(n_142) );
AOI221x1_ASAP7_75t_L g240 ( .A1(n_13), .A2(n_24), .B1(n_145), .B2(n_154), .C(n_241), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_14), .B(n_161), .Y(n_510) );
CKINVDCx16_ASAP7_75t_R g111 ( .A(n_15), .Y(n_111) );
NAND2xp5_ASAP7_75t_SL g144 ( .A(n_16), .B(n_145), .Y(n_144) );
AO21x2_ASAP7_75t_L g139 ( .A1(n_17), .A2(n_140), .B(n_143), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_18), .B(n_179), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_19), .B(n_161), .Y(n_188) );
AO21x1_ASAP7_75t_L g219 ( .A1(n_20), .A2(n_145), .B(n_220), .Y(n_219) );
NAND2xp5_ASAP7_75t_SL g541 ( .A(n_21), .B(n_145), .Y(n_541) );
NOR2xp33_ASAP7_75t_SL g106 ( .A(n_22), .B(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g125 ( .A(n_22), .Y(n_125) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_23), .A2(n_91), .B1(n_145), .B2(n_481), .Y(n_480) );
NAND2x1_ASAP7_75t_L g210 ( .A(n_25), .B(n_161), .Y(n_210) );
NAND2x1_ASAP7_75t_L g198 ( .A(n_26), .B(n_163), .Y(n_198) );
OA21x2_ASAP7_75t_L g141 ( .A1(n_27), .A2(n_88), .B(n_142), .Y(n_141) );
OR2x2_ASAP7_75t_L g166 ( .A(n_27), .B(n_88), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_28), .B(n_163), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_29), .B(n_161), .Y(n_160) );
AO21x2_ASAP7_75t_L g505 ( .A1(n_30), .A2(n_171), .B(n_506), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_31), .B(n_163), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_32), .A2(n_154), .B(n_532), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_33), .B(n_161), .Y(n_517) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_34), .A2(n_154), .B(n_230), .Y(n_229) );
AND2x2_ASAP7_75t_L g151 ( .A(n_35), .B(n_152), .Y(n_151) );
AND2x2_ASAP7_75t_L g155 ( .A(n_35), .B(n_156), .Y(n_155) );
INVx1_ASAP7_75t_L g489 ( .A(n_35), .Y(n_489) );
NOR3xp33_ASAP7_75t_L g108 ( .A(n_36), .B(n_109), .C(n_111), .Y(n_108) );
OR2x6_ASAP7_75t_L g123 ( .A(n_36), .B(n_124), .Y(n_123) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_37), .B(n_145), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_38), .B(n_145), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_39), .B(n_161), .Y(n_501) );
CKINVDCx20_ASAP7_75t_R g192 ( .A(n_40), .Y(n_192) );
XNOR2xp5_ASAP7_75t_L g777 ( .A(n_40), .B(n_778), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_41), .B(n_163), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_42), .B(n_145), .Y(n_462) );
XNOR2xp5_ASAP7_75t_L g763 ( .A(n_43), .B(n_764), .Y(n_763) );
AOI21xp5_ASAP7_75t_L g471 ( .A1(n_44), .A2(n_154), .B(n_472), .Y(n_471) );
OAI22xp5_ASAP7_75t_SL g779 ( .A1(n_45), .A2(n_780), .B1(n_781), .B2(n_782), .Y(n_779) );
CKINVDCx20_ASAP7_75t_R g780 ( .A(n_45), .Y(n_780) );
AOI21xp5_ASAP7_75t_L g196 ( .A1(n_46), .A2(n_154), .B(n_197), .Y(n_196) );
XNOR2xp5_ASAP7_75t_L g762 ( .A(n_47), .B(n_763), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_48), .B(n_163), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_49), .B(n_163), .Y(n_211) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_50), .B(n_145), .Y(n_507) );
INVx1_ASAP7_75t_L g148 ( .A(n_51), .Y(n_148) );
INVx1_ASAP7_75t_L g158 ( .A(n_51), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_52), .B(n_161), .Y(n_474) );
AND2x2_ASAP7_75t_L g496 ( .A(n_53), .B(n_179), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_54), .B(n_163), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_55), .B(n_161), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_56), .B(n_163), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_57), .A2(n_154), .B(n_209), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g475 ( .A(n_58), .B(n_145), .Y(n_475) );
NAND2xp5_ASAP7_75t_SL g498 ( .A(n_59), .B(n_145), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_60), .A2(n_154), .B(n_515), .Y(n_514) );
AOI22xp5_ASAP7_75t_L g764 ( .A1(n_61), .A2(n_100), .B1(n_765), .B2(n_766), .Y(n_764) );
CKINVDCx20_ASAP7_75t_R g766 ( .A(n_61), .Y(n_766) );
AO21x1_ASAP7_75t_L g221 ( .A1(n_62), .A2(n_154), .B(n_222), .Y(n_221) );
AND2x2_ASAP7_75t_L g547 ( .A(n_63), .B(n_180), .Y(n_547) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_64), .B(n_145), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_65), .B(n_163), .Y(n_502) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_66), .B(n_145), .Y(n_200) );
AOI22xp5_ASAP7_75t_L g782 ( .A1(n_67), .A2(n_80), .B1(n_783), .B2(n_784), .Y(n_782) );
CKINVDCx20_ASAP7_75t_R g784 ( .A(n_67), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_68), .B(n_163), .Y(n_511) );
AOI22xp5_ASAP7_75t_L g486 ( .A1(n_69), .A2(n_95), .B1(n_154), .B2(n_487), .Y(n_486) );
AND2x2_ASAP7_75t_L g234 ( .A(n_70), .B(n_180), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_71), .B(n_161), .Y(n_544) );
INVx1_ASAP7_75t_L g150 ( .A(n_72), .Y(n_150) );
INVx1_ASAP7_75t_L g156 ( .A(n_72), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_73), .B(n_119), .Y(n_118) );
AND2x2_ASAP7_75t_L g202 ( .A(n_74), .B(n_171), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_75), .B(n_163), .Y(n_533) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_76), .A2(n_154), .B(n_500), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g463 ( .A1(n_77), .A2(n_154), .B(n_464), .Y(n_463) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_78), .A2(n_154), .B(n_509), .Y(n_508) );
AND2x2_ASAP7_75t_L g519 ( .A(n_79), .B(n_180), .Y(n_519) );
CKINVDCx20_ASAP7_75t_R g783 ( .A(n_80), .Y(n_783) );
NAND2xp5_ASAP7_75t_SL g478 ( .A(n_81), .B(n_179), .Y(n_478) );
INVx1_ASAP7_75t_L g107 ( .A(n_82), .Y(n_107) );
AND2x2_ASAP7_75t_L g170 ( .A(n_83), .B(n_171), .Y(n_170) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_84), .B(n_145), .Y(n_190) );
AND2x2_ASAP7_75t_L g467 ( .A(n_85), .B(n_140), .Y(n_467) );
AND2x2_ASAP7_75t_L g220 ( .A(n_86), .B(n_165), .Y(n_220) );
INVxp33_ASAP7_75t_L g789 ( .A(n_87), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_89), .B(n_163), .Y(n_189) );
AND2x2_ASAP7_75t_L g214 ( .A(n_90), .B(n_171), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_92), .B(n_161), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g186 ( .A1(n_93), .A2(n_154), .B(n_187), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_94), .B(n_163), .Y(n_242) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_96), .A2(n_154), .B(n_543), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_97), .B(n_161), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_98), .B(n_161), .Y(n_177) );
BUFx2_ASAP7_75t_L g546 ( .A(n_99), .Y(n_546) );
CKINVDCx20_ASAP7_75t_R g765 ( .A(n_100), .Y(n_765) );
BUFx2_ASAP7_75t_L g117 ( .A(n_101), .Y(n_117) );
AOI21xp5_ASAP7_75t_L g153 ( .A1(n_102), .A2(n_154), .B(n_159), .Y(n_153) );
CKINVDCx20_ASAP7_75t_R g773 ( .A(n_103), .Y(n_773) );
AOI21xp33_ASAP7_75t_SL g104 ( .A1(n_105), .A2(n_112), .B(n_788), .Y(n_104) );
INVx2_ASAP7_75t_L g792 ( .A(n_105), .Y(n_792) );
AND2x2_ASAP7_75t_SL g105 ( .A(n_106), .B(n_108), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_107), .B(n_125), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g121 ( .A(n_111), .B(n_122), .Y(n_121) );
OR2x6_ASAP7_75t_SL g132 ( .A(n_111), .B(n_122), .Y(n_132) );
AND2x6_ASAP7_75t_SL g761 ( .A(n_111), .B(n_123), .Y(n_761) );
OR2x2_ASAP7_75t_L g775 ( .A(n_111), .B(n_123), .Y(n_775) );
OA22x2_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_117), .B1(n_126), .B2(n_776), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_114), .B(n_118), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_116), .Y(n_115) );
HB1xp67_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
OAI21xp5_ASAP7_75t_L g776 ( .A1(n_118), .A2(n_777), .B(n_785), .Y(n_776) );
INVx1_ASAP7_75t_SL g119 ( .A(n_120), .Y(n_119) );
BUFx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
BUFx2_ASAP7_75t_L g787 ( .A(n_121), .Y(n_787) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_123), .Y(n_122) );
OAI21xp5_ASAP7_75t_SL g126 ( .A1(n_127), .A2(n_762), .B(n_767), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
OAI22xp5_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_133), .B1(n_455), .B2(n_758), .Y(n_128) );
BUFx4f_ASAP7_75t_SL g129 ( .A(n_130), .Y(n_129) );
OAI22x1_ASAP7_75t_L g768 ( .A1(n_130), .A2(n_769), .B1(n_770), .B2(n_771), .Y(n_768) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_131), .Y(n_130) );
CKINVDCx11_ASAP7_75t_R g131 ( .A(n_132), .Y(n_131) );
INVx1_ASAP7_75t_L g769 ( .A(n_133), .Y(n_769) );
AND2x4_ASAP7_75t_L g133 ( .A(n_134), .B(n_376), .Y(n_133) );
NOR3xp33_ASAP7_75t_SL g134 ( .A(n_135), .B(n_288), .C(n_328), .Y(n_134) );
OAI221xp5_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_203), .B1(n_252), .B2(n_267), .C(n_270), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
AND2x2_ASAP7_75t_L g137 ( .A(n_138), .B(n_167), .Y(n_137) );
INVx2_ASAP7_75t_L g285 ( .A(n_138), .Y(n_285) );
AND2x2_ASAP7_75t_L g315 ( .A(n_138), .B(n_316), .Y(n_315) );
BUFx3_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
AND2x2_ASAP7_75t_L g253 ( .A(n_139), .B(n_254), .Y(n_253) );
OR2x2_ASAP7_75t_L g260 ( .A(n_139), .B(n_193), .Y(n_260) );
INVx2_ASAP7_75t_L g266 ( .A(n_139), .Y(n_266) );
AND2x2_ASAP7_75t_L g275 ( .A(n_139), .B(n_169), .Y(n_275) );
INVx1_ASAP7_75t_L g291 ( .A(n_139), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_139), .B(n_337), .Y(n_336) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_140), .A2(n_541), .B(n_542), .Y(n_540) );
BUFx4f_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx3_ASAP7_75t_L g172 ( .A(n_141), .Y(n_172) );
AND2x4_ASAP7_75t_L g165 ( .A(n_142), .B(n_166), .Y(n_165) );
AND2x2_ASAP7_75t_SL g180 ( .A(n_142), .B(n_166), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_153), .B(n_165), .Y(n_143) );
AND2x4_ASAP7_75t_L g145 ( .A(n_146), .B(n_151), .Y(n_145) );
AND2x4_ASAP7_75t_L g146 ( .A(n_147), .B(n_149), .Y(n_146) );
AND2x6_ASAP7_75t_L g163 ( .A(n_147), .B(n_156), .Y(n_163) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
AND2x4_ASAP7_75t_L g161 ( .A(n_149), .B(n_158), .Y(n_161) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx5_ASAP7_75t_L g164 ( .A(n_151), .Y(n_164) );
AND2x2_ASAP7_75t_L g157 ( .A(n_152), .B(n_158), .Y(n_157) );
HB1xp67_ASAP7_75t_L g484 ( .A(n_152), .Y(n_484) );
AND2x6_ASAP7_75t_L g154 ( .A(n_155), .B(n_157), .Y(n_154) );
BUFx3_ASAP7_75t_L g485 ( .A(n_155), .Y(n_485) );
INVx2_ASAP7_75t_L g491 ( .A(n_156), .Y(n_491) );
AND2x4_ASAP7_75t_L g487 ( .A(n_157), .B(n_488), .Y(n_487) );
INVx2_ASAP7_75t_L g483 ( .A(n_158), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g159 ( .A1(n_160), .A2(n_162), .B(n_164), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_163), .B(n_546), .Y(n_545) );
AOI21xp5_ASAP7_75t_L g176 ( .A1(n_164), .A2(n_177), .B(n_178), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_164), .A2(n_188), .B(n_189), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g197 ( .A1(n_164), .A2(n_198), .B(n_199), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_164), .A2(n_210), .B(n_211), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_164), .A2(n_223), .B(n_224), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_164), .A2(n_231), .B(n_232), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_164), .A2(n_242), .B(n_243), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g464 ( .A1(n_164), .A2(n_465), .B(n_466), .Y(n_464) );
AOI21xp5_ASAP7_75t_L g472 ( .A1(n_164), .A2(n_473), .B(n_474), .Y(n_472) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_164), .A2(n_501), .B(n_502), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g509 ( .A1(n_164), .A2(n_510), .B(n_511), .Y(n_509) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_164), .A2(n_516), .B(n_517), .Y(n_515) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_164), .A2(n_533), .B(n_534), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_164), .A2(n_544), .B(n_545), .Y(n_543) );
INVx1_ASAP7_75t_SL g184 ( .A(n_165), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_165), .B(n_226), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_165), .A2(n_498), .B(n_499), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_165), .A2(n_507), .B(n_508), .Y(n_506) );
AND2x2_ASAP7_75t_SL g167 ( .A(n_168), .B(n_181), .Y(n_167) );
INVx4_ASAP7_75t_L g256 ( .A(n_168), .Y(n_256) );
AND2x2_ASAP7_75t_L g287 ( .A(n_168), .B(n_194), .Y(n_287) );
AND2x2_ASAP7_75t_L g363 ( .A(n_168), .B(n_337), .Y(n_363) );
NAND2x1p5_ASAP7_75t_L g405 ( .A(n_168), .B(n_193), .Y(n_405) );
INVx5_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_169), .B(n_193), .Y(n_292) );
AND2x2_ASAP7_75t_L g316 ( .A(n_169), .B(n_194), .Y(n_316) );
BUFx2_ASAP7_75t_L g332 ( .A(n_169), .Y(n_332) );
NOR2x1_ASAP7_75t_SL g435 ( .A(n_169), .B(n_337), .Y(n_435) );
OR2x6_ASAP7_75t_L g169 ( .A(n_170), .B(n_173), .Y(n_169) );
INVx3_ASAP7_75t_L g213 ( .A(n_171), .Y(n_213) );
INVx4_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
AO21x2_ASAP7_75t_L g469 ( .A1(n_172), .A2(n_470), .B(n_476), .Y(n_469) );
AOI21xp5_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_175), .B(n_179), .Y(n_173) );
CKINVDCx5p33_ASAP7_75t_R g201 ( .A(n_179), .Y(n_201) );
OA21x2_ASAP7_75t_L g239 ( .A1(n_179), .A2(n_240), .B(n_244), .Y(n_239) );
OA21x2_ASAP7_75t_L g302 ( .A1(n_179), .A2(n_240), .B(n_244), .Y(n_302) );
AOI21xp5_ASAP7_75t_L g461 ( .A1(n_179), .A2(n_462), .B(n_463), .Y(n_461) );
AO21x2_ASAP7_75t_L g479 ( .A1(n_179), .A2(n_480), .B(n_486), .Y(n_479) );
BUFx6f_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx2_ASAP7_75t_L g312 ( .A(n_181), .Y(n_312) );
AOI221xp5_ASAP7_75t_L g378 ( .A1(n_181), .A2(n_379), .B1(n_381), .B2(n_383), .C(n_388), .Y(n_378) );
AND2x2_ASAP7_75t_L g398 ( .A(n_181), .B(n_291), .Y(n_398) );
AND2x4_ASAP7_75t_L g181 ( .A(n_182), .B(n_193), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx2_ASAP7_75t_L g254 ( .A(n_183), .Y(n_254) );
INVx1_ASAP7_75t_L g307 ( .A(n_183), .Y(n_307) );
AO21x2_ASAP7_75t_L g183 ( .A1(n_184), .A2(n_185), .B(n_191), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g191 ( .A(n_184), .B(n_192), .Y(n_191) );
AO21x2_ASAP7_75t_L g337 ( .A1(n_184), .A2(n_185), .B(n_191), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_186), .B(n_190), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_193), .B(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g276 ( .A(n_193), .B(n_264), .Y(n_276) );
INVx2_ASAP7_75t_L g318 ( .A(n_193), .Y(n_318) );
AND2x2_ASAP7_75t_L g451 ( .A(n_193), .B(n_266), .Y(n_451) );
INVx4_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_194), .Y(n_308) );
AO21x2_ASAP7_75t_L g194 ( .A1(n_195), .A2(n_201), .B(n_202), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_196), .B(n_200), .Y(n_195) );
AOI21x1_ASAP7_75t_L g529 ( .A1(n_201), .A2(n_530), .B(n_536), .Y(n_529) );
NOR3xp33_ASAP7_75t_L g203 ( .A(n_204), .B(n_235), .C(n_250), .Y(n_203) );
AND2x2_ASAP7_75t_L g204 ( .A(n_205), .B(n_215), .Y(n_204) );
INVx2_ASAP7_75t_L g365 ( .A(n_205), .Y(n_365) );
AND2x2_ASAP7_75t_L g410 ( .A(n_205), .B(n_287), .Y(n_410) );
BUFx2_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
INVx1_ASAP7_75t_L g355 ( .A(n_206), .Y(n_355) );
AND2x4_ASAP7_75t_SL g370 ( .A(n_206), .B(n_282), .Y(n_370) );
AO21x2_ASAP7_75t_L g206 ( .A1(n_207), .A2(n_213), .B(n_214), .Y(n_206) );
AO21x2_ASAP7_75t_L g249 ( .A1(n_207), .A2(n_213), .B(n_214), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_208), .B(n_212), .Y(n_207) );
AO21x2_ASAP7_75t_L g227 ( .A1(n_213), .A2(n_228), .B(n_234), .Y(n_227) );
AO21x2_ASAP7_75t_L g247 ( .A1(n_213), .A2(n_228), .B(n_234), .Y(n_247) );
AO21x1_ASAP7_75t_SL g512 ( .A1(n_213), .A2(n_513), .B(n_519), .Y(n_512) );
AO21x2_ASAP7_75t_L g570 ( .A1(n_213), .A2(n_513), .B(n_519), .Y(n_570) );
INVx2_ASAP7_75t_L g324 ( .A(n_215), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_215), .B(n_354), .Y(n_380) );
AND2x4_ASAP7_75t_L g413 ( .A(n_215), .B(n_360), .Y(n_413) );
AND2x4_ASAP7_75t_L g215 ( .A(n_216), .B(n_227), .Y(n_215) );
AND2x2_ASAP7_75t_L g251 ( .A(n_216), .B(n_246), .Y(n_251) );
OR2x2_ASAP7_75t_L g281 ( .A(n_216), .B(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_SL g350 ( .A(n_216), .B(n_302), .Y(n_350) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
BUFx2_ASAP7_75t_L g295 ( .A(n_217), .Y(n_295) );
INVx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVx2_ASAP7_75t_L g269 ( .A(n_218), .Y(n_269) );
OAI21x1_ASAP7_75t_SL g218 ( .A1(n_219), .A2(n_221), .B(n_225), .Y(n_218) );
INVx1_ASAP7_75t_L g226 ( .A(n_220), .Y(n_226) );
INVx2_ASAP7_75t_L g282 ( .A(n_227), .Y(n_282) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_229), .B(n_233), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g444 ( .A(n_235), .B(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_237), .B(n_245), .Y(n_236) );
AND2x2_ASAP7_75t_L g250 ( .A(n_237), .B(n_251), .Y(n_250) );
OR2x2_ASAP7_75t_L g323 ( .A(n_237), .B(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g408 ( .A(n_237), .Y(n_408) );
BUFx2_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
AND2x4_ASAP7_75t_L g268 ( .A(n_238), .B(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g387 ( .A(n_238), .B(n_247), .Y(n_387) );
AND2x2_ASAP7_75t_L g391 ( .A(n_238), .B(n_257), .Y(n_391) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
INVx2_ASAP7_75t_L g360 ( .A(n_239), .Y(n_360) );
HB1xp67_ASAP7_75t_L g428 ( .A(n_239), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_245), .B(n_268), .Y(n_344) );
AND2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_248), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_246), .B(n_269), .Y(n_454) );
INVx2_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g258 ( .A(n_247), .B(n_249), .Y(n_258) );
AND2x2_ASAP7_75t_L g340 ( .A(n_247), .B(n_302), .Y(n_340) );
AND2x2_ASAP7_75t_L g359 ( .A(n_247), .B(n_248), .Y(n_359) );
BUFx2_ASAP7_75t_L g280 ( .A(n_248), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_248), .B(n_340), .Y(n_339) );
INVx2_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
BUFx3_ASAP7_75t_L g257 ( .A(n_249), .Y(n_257) );
INVxp67_ASAP7_75t_L g300 ( .A(n_249), .Y(n_300) );
INVx1_ASAP7_75t_L g273 ( .A(n_251), .Y(n_273) );
AND2x2_ASAP7_75t_L g309 ( .A(n_251), .B(n_280), .Y(n_309) );
NAND2xp33_ASAP7_75t_L g390 ( .A(n_251), .B(n_391), .Y(n_390) );
AND2x2_ASAP7_75t_L g427 ( .A(n_251), .B(n_428), .Y(n_427) );
AOI221xp5_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_255), .B1(n_258), .B2(n_259), .C(n_261), .Y(n_252) );
AND2x2_ASAP7_75t_L g356 ( .A(n_253), .B(n_256), .Y(n_356) );
AND2x2_ASAP7_75t_SL g375 ( .A(n_253), .B(n_316), .Y(n_375) );
AND2x2_ASAP7_75t_L g393 ( .A(n_253), .B(n_318), .Y(n_393) );
AND2x2_ASAP7_75t_L g448 ( .A(n_253), .B(n_287), .Y(n_448) );
INVx1_ASAP7_75t_L g264 ( .A(n_254), .Y(n_264) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_254), .Y(n_320) );
CKINVDCx16_ASAP7_75t_R g400 ( .A(n_255), .Y(n_400) );
AND2x4_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_256), .B(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_256), .B(n_307), .Y(n_382) );
AND2x2_ASAP7_75t_L g349 ( .A(n_257), .B(n_350), .Y(n_349) );
INVx1_ASAP7_75t_SL g385 ( .A(n_257), .Y(n_385) );
AND2x2_ASAP7_75t_L g294 ( .A(n_258), .B(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_258), .B(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g436 ( .A(n_258), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_258), .B(n_360), .Y(n_446) );
AND2x4_ASAP7_75t_L g362 ( .A(n_259), .B(n_363), .Y(n_362) );
INVx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
OR2x2_ASAP7_75t_L g433 ( .A(n_260), .B(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
OR2x2_ASAP7_75t_L g262 ( .A(n_263), .B(n_265), .Y(n_262) );
OR2x2_ASAP7_75t_L g304 ( .A(n_265), .B(n_305), .Y(n_304) );
OR2x2_ASAP7_75t_L g311 ( .A(n_266), .B(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g342 ( .A(n_266), .B(n_316), .Y(n_342) );
AND2x2_ASAP7_75t_L g416 ( .A(n_266), .B(n_337), .Y(n_416) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g364 ( .A(n_268), .B(n_365), .Y(n_364) );
OAI32xp33_ASAP7_75t_L g429 ( .A1(n_268), .A2(n_430), .A3(n_432), .B1(n_433), .B2(n_436), .Y(n_429) );
AND2x4_ASAP7_75t_L g301 ( .A(n_269), .B(n_302), .Y(n_301) );
OR2x2_ASAP7_75t_L g399 ( .A(n_269), .B(n_302), .Y(n_399) );
AOI22xp5_ASAP7_75t_L g270 ( .A1(n_271), .A2(n_274), .B1(n_277), .B2(n_283), .Y(n_270) );
INVxp67_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
O2A1O1Ixp33_ASAP7_75t_SL g388 ( .A1(n_272), .A2(n_286), .B(n_389), .C(n_390), .Y(n_388) );
HB1xp67_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
OR2x2_ASAP7_75t_L g372 ( .A(n_273), .B(n_300), .Y(n_372) );
INVx1_ASAP7_75t_SL g443 ( .A(n_274), .Y(n_443) );
AND2x4_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
AND2x4_ASAP7_75t_L g346 ( .A(n_276), .B(n_285), .Y(n_346) );
AOI221xp5_ASAP7_75t_L g424 ( .A1(n_276), .A2(n_425), .B1(n_426), .B2(n_427), .C(n_429), .Y(n_424) );
INVx1_ASAP7_75t_SL g277 ( .A(n_278), .Y(n_277) );
OR2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_281), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
NOR2xp33_ASAP7_75t_L g352 ( .A(n_281), .B(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
OAI22xp33_ASAP7_75t_L g366 ( .A1(n_284), .A2(n_314), .B1(n_367), .B2(n_368), .Y(n_366) );
OR2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
OAI211xp5_ASAP7_75t_SL g402 ( .A1(n_285), .A2(n_403), .B(n_411), .C(n_424), .Y(n_402) );
INVx2_ASAP7_75t_SL g286 ( .A(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g322 ( .A(n_287), .B(n_291), .Y(n_322) );
OAI211xp5_ASAP7_75t_SL g288 ( .A1(n_289), .A2(n_293), .B(n_296), .C(n_325), .Y(n_288) );
OR2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_292), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g319 ( .A(n_291), .B(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g439 ( .A(n_291), .B(n_435), .Y(n_439) );
OAI32xp33_ASAP7_75t_L g396 ( .A1(n_292), .A2(n_397), .A3(n_399), .B1(n_400), .B2(n_401), .Y(n_396) );
INVx1_ASAP7_75t_SL g293 ( .A(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_SL g386 ( .A(n_295), .B(n_387), .Y(n_386) );
AOI221xp5_ASAP7_75t_L g296 ( .A1(n_297), .A2(n_303), .B1(n_309), .B2(n_310), .C(n_313), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_SL g298 ( .A(n_299), .B(n_301), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
OR2x2_ASAP7_75t_L g453 ( .A(n_300), .B(n_454), .Y(n_453) );
NAND2xp5_ASAP7_75t_SL g367 ( .A(n_301), .B(n_365), .Y(n_367) );
A2O1A1O1Ixp25_ASAP7_75t_L g438 ( .A1(n_301), .A2(n_370), .B(n_386), .C(n_432), .D(n_439), .Y(n_438) );
AOI31xp33_ASAP7_75t_L g440 ( .A1(n_301), .A2(n_322), .A3(n_432), .B(n_439), .Y(n_440) );
AND2x2_ASAP7_75t_L g354 ( .A(n_302), .B(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_SL g442 ( .A(n_304), .B(n_443), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_306), .B(n_308), .Y(n_305) );
INVx2_ASAP7_75t_L g431 ( .A(n_306), .Y(n_431) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g426 ( .A(n_307), .B(n_318), .Y(n_426) );
INVx1_ASAP7_75t_L g341 ( .A(n_309), .Y(n_341) );
AND2x2_ASAP7_75t_L g326 ( .A(n_310), .B(n_327), .Y(n_326) );
INVx2_ASAP7_75t_SL g310 ( .A(n_311), .Y(n_310) );
AOI31xp33_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_317), .A3(n_321), .B(n_323), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_316), .B(n_431), .Y(n_430) );
AND2x2_ASAP7_75t_L g449 ( .A(n_316), .B(n_395), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
AND2x2_ASAP7_75t_L g394 ( .A(n_318), .B(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g420 ( .A(n_318), .Y(n_420) );
INVxp67_ASAP7_75t_L g389 ( .A(n_319), .Y(n_389) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx2_ASAP7_75t_L g327 ( .A(n_323), .Y(n_327) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
NAND3xp33_ASAP7_75t_SL g328 ( .A(n_329), .B(n_345), .C(n_361), .Y(n_328) );
AOI22xp5_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_338), .B1(n_342), .B2(n_343), .Y(n_329) );
INVxp67_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_332), .B(n_333), .Y(n_331) );
INVx2_ASAP7_75t_L g415 ( .A(n_332), .Y(n_415) );
INVx1_ASAP7_75t_SL g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVxp67_ASAP7_75t_SL g395 ( .A(n_336), .Y(n_395) );
INVxp67_ASAP7_75t_SL g421 ( .A(n_336), .Y(n_421) );
OR2x2_ASAP7_75t_L g422 ( .A(n_336), .B(n_405), .Y(n_422) );
NAND2xp33_ASAP7_75t_L g338 ( .A(n_339), .B(n_341), .Y(n_338) );
INVx1_ASAP7_75t_L g373 ( .A(n_340), .Y(n_373) );
INVx1_ASAP7_75t_SL g343 ( .A(n_344), .Y(n_343) );
AOI22xp33_ASAP7_75t_L g345 ( .A1(n_346), .A2(n_347), .B1(n_356), .B2(n_357), .Y(n_345) );
NAND2xp5_ASAP7_75t_SL g347 ( .A(n_348), .B(n_351), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_SL g353 ( .A(n_354), .Y(n_353) );
AOI221xp5_ASAP7_75t_L g392 ( .A1(n_354), .A2(n_359), .B1(n_393), .B2(n_394), .C(n_396), .Y(n_392) );
INVx2_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
NAND2x1_ASAP7_75t_L g358 ( .A(n_359), .B(n_360), .Y(n_358) );
INVx1_ASAP7_75t_L g432 ( .A(n_359), .Y(n_432) );
AND2x2_ASAP7_75t_L g369 ( .A(n_360), .B(n_370), .Y(n_369) );
O2A1O1Ixp33_ASAP7_75t_SL g417 ( .A1(n_360), .A2(n_418), .B(n_422), .C(n_423), .Y(n_417) );
AOI211xp5_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_364), .B(n_366), .C(n_371), .Y(n_361) );
AND2x2_ASAP7_75t_L g412 ( .A(n_365), .B(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g423 ( .A(n_370), .Y(n_423) );
AOI21xp33_ASAP7_75t_SL g371 ( .A1(n_372), .A2(n_373), .B(n_374), .Y(n_371) );
INVx2_ASAP7_75t_SL g374 ( .A(n_375), .Y(n_374) );
NOR3xp33_ASAP7_75t_L g376 ( .A(n_377), .B(n_402), .C(n_437), .Y(n_376) );
NAND2xp5_ASAP7_75t_SL g377 ( .A(n_378), .B(n_392), .Y(n_377) );
INVx1_ASAP7_75t_SL g379 ( .A(n_380), .Y(n_379) );
INVxp67_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
NAND2xp5_ASAP7_75t_SL g384 ( .A(n_385), .B(n_386), .Y(n_384) );
INVx1_ASAP7_75t_L g401 ( .A(n_386), .Y(n_401) );
INVxp67_ASAP7_75t_L g425 ( .A(n_390), .Y(n_425) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_SL g409 ( .A(n_399), .Y(n_409) );
AOI22xp5_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_406), .B1(n_409), .B2(n_410), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
AOI21xp5_ASAP7_75t_L g411 ( .A1(n_412), .A2(n_414), .B(n_417), .Y(n_411) );
AND2x2_ASAP7_75t_L g414 ( .A(n_415), .B(n_416), .Y(n_414) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_420), .B(n_421), .Y(n_419) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
AND2x2_ASAP7_75t_L g450 ( .A(n_435), .B(n_451), .Y(n_450) );
OAI221xp5_ASAP7_75t_L g437 ( .A1(n_438), .A2(n_440), .B1(n_441), .B2(n_444), .C(n_447), .Y(n_437) );
INVxp67_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
OAI31xp33_ASAP7_75t_SL g447 ( .A1(n_448), .A2(n_449), .A3(n_450), .B(n_452), .Y(n_447) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx3_ASAP7_75t_SL g770 ( .A(n_455), .Y(n_770) );
XNOR2xp5_ASAP7_75t_L g778 ( .A(n_455), .B(n_779), .Y(n_778) );
AND2x4_ASAP7_75t_SL g455 ( .A(n_456), .B(n_654), .Y(n_455) );
NOR3xp33_ASAP7_75t_SL g456 ( .A(n_457), .B(n_563), .C(n_595), .Y(n_456) );
OAI221xp5_ASAP7_75t_L g457 ( .A1(n_458), .A2(n_492), .B1(n_520), .B2(n_537), .C(n_548), .Y(n_457) );
OR2x2_ASAP7_75t_L g458 ( .A(n_459), .B(n_468), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
AND2x2_ASAP7_75t_L g526 ( .A(n_460), .B(n_469), .Y(n_526) );
INVx4_ASAP7_75t_L g554 ( .A(n_460), .Y(n_554) );
AND2x4_ASAP7_75t_SL g594 ( .A(n_460), .B(n_528), .Y(n_594) );
BUFx2_ASAP7_75t_L g604 ( .A(n_460), .Y(n_604) );
NOR2x1_ASAP7_75t_L g670 ( .A(n_460), .B(n_609), .Y(n_670) );
AND2x2_ASAP7_75t_L g679 ( .A(n_460), .B(n_607), .Y(n_679) );
OR2x2_ASAP7_75t_L g687 ( .A(n_460), .B(n_688), .Y(n_687) );
AND2x2_ASAP7_75t_L g713 ( .A(n_460), .B(n_552), .Y(n_713) );
AND2x4_ASAP7_75t_L g732 ( .A(n_460), .B(n_733), .Y(n_732) );
OR2x6_ASAP7_75t_L g460 ( .A(n_461), .B(n_467), .Y(n_460) );
INVx2_ASAP7_75t_SL g645 ( .A(n_468), .Y(n_645) );
OR2x2_ASAP7_75t_L g468 ( .A(n_469), .B(n_477), .Y(n_468) );
AND2x2_ASAP7_75t_L g552 ( .A(n_469), .B(n_529), .Y(n_552) );
INVx2_ASAP7_75t_L g579 ( .A(n_469), .Y(n_579) );
INVx2_ASAP7_75t_L g609 ( .A(n_469), .Y(n_609) );
AND2x2_ASAP7_75t_L g623 ( .A(n_469), .B(n_528), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_471), .B(n_475), .Y(n_470) );
AND2x2_ASAP7_75t_L g553 ( .A(n_477), .B(n_554), .Y(n_553) );
INVx2_ASAP7_75t_L g576 ( .A(n_477), .Y(n_576) );
BUFx3_ASAP7_75t_L g590 ( .A(n_477), .Y(n_590) );
AND2x2_ASAP7_75t_L g619 ( .A(n_477), .B(n_620), .Y(n_619) );
AND2x4_ASAP7_75t_L g477 ( .A(n_478), .B(n_479), .Y(n_477) );
AND2x4_ASAP7_75t_L g524 ( .A(n_478), .B(n_479), .Y(n_524) );
AND2x4_ASAP7_75t_L g481 ( .A(n_482), .B(n_485), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_483), .B(n_484), .Y(n_482) );
NOR2x1p5_ASAP7_75t_L g488 ( .A(n_489), .B(n_490), .Y(n_488) );
INVx3_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx1_ASAP7_75t_L g625 ( .A(n_492), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_493), .B(n_503), .Y(n_492) );
OR2x2_ASAP7_75t_L g736 ( .A(n_493), .B(n_537), .Y(n_736) );
INVx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
AND2x2_ASAP7_75t_L g592 ( .A(n_494), .B(n_593), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_494), .B(n_503), .Y(n_653) );
OR2x2_ASAP7_75t_L g751 ( .A(n_494), .B(n_673), .Y(n_751) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
AND2x2_ASAP7_75t_L g562 ( .A(n_495), .B(n_538), .Y(n_562) );
OR2x2_ASAP7_75t_SL g572 ( .A(n_495), .B(n_573), .Y(n_572) );
INVx4_ASAP7_75t_L g583 ( .A(n_495), .Y(n_583) );
HB1xp67_ASAP7_75t_L g634 ( .A(n_495), .Y(n_634) );
NAND2x1_ASAP7_75t_L g640 ( .A(n_495), .B(n_539), .Y(n_640) );
AND2x2_ASAP7_75t_L g665 ( .A(n_495), .B(n_505), .Y(n_665) );
OR2x2_ASAP7_75t_L g686 ( .A(n_495), .B(n_569), .Y(n_686) );
OR2x6_ASAP7_75t_L g495 ( .A(n_496), .B(n_497), .Y(n_495) );
INVx1_ASAP7_75t_L g581 ( .A(n_503), .Y(n_581) );
O2A1O1Ixp33_ASAP7_75t_L g674 ( .A1(n_503), .A2(n_675), .B(n_678), .C(n_680), .Y(n_674) );
AND2x2_ASAP7_75t_L g747 ( .A(n_503), .B(n_523), .Y(n_747) );
AND2x2_ASAP7_75t_L g503 ( .A(n_504), .B(n_512), .Y(n_503) );
INVx1_ASAP7_75t_L g614 ( .A(n_504), .Y(n_614) );
AND2x2_ASAP7_75t_L g684 ( .A(n_504), .B(n_539), .Y(n_684) );
INVx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g558 ( .A(n_505), .Y(n_558) );
OR2x2_ASAP7_75t_L g573 ( .A(n_505), .B(n_539), .Y(n_573) );
INVx1_ASAP7_75t_L g589 ( .A(n_505), .Y(n_589) );
AND2x2_ASAP7_75t_L g601 ( .A(n_505), .B(n_512), .Y(n_601) );
HB1xp67_ASAP7_75t_L g707 ( .A(n_505), .Y(n_707) );
NOR2x1_ASAP7_75t_SL g538 ( .A(n_512), .B(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_514), .B(n_518), .Y(n_513) );
INVxp67_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_522), .B(n_525), .Y(n_521) );
OR2x2_ASAP7_75t_L g671 ( .A(n_522), .B(n_606), .Y(n_671) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_523), .B(n_689), .Y(n_688) );
OR2x2_ASAP7_75t_L g753 ( .A(n_523), .B(n_650), .Y(n_753) );
INVx3_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
AND2x2_ASAP7_75t_L g598 ( .A(n_524), .B(n_579), .Y(n_598) );
AND2x2_ASAP7_75t_L g694 ( .A(n_524), .B(n_607), .Y(n_694) );
INVx1_ASAP7_75t_L g611 ( .A(n_525), .Y(n_611) );
AND2x2_ASAP7_75t_L g525 ( .A(n_526), .B(n_527), .Y(n_525) );
INVx1_ASAP7_75t_L g661 ( .A(n_526), .Y(n_661) );
INVx2_ASAP7_75t_L g628 ( .A(n_527), .Y(n_628) );
HB1xp67_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
AND2x2_ASAP7_75t_L g578 ( .A(n_528), .B(n_579), .Y(n_578) );
INVx2_ASAP7_75t_L g608 ( .A(n_528), .Y(n_608) );
INVx1_ASAP7_75t_L g733 ( .A(n_528), .Y(n_733) );
INVx3_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
HB1xp67_ASAP7_75t_L g690 ( .A(n_529), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_531), .B(n_535), .Y(n_530) );
OR2x2_ASAP7_75t_L g704 ( .A(n_537), .B(n_705), .Y(n_704) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx2_ASAP7_75t_SL g559 ( .A(n_539), .Y(n_559) );
OR2x2_ASAP7_75t_L g582 ( .A(n_539), .B(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g593 ( .A(n_539), .B(n_569), .Y(n_593) );
AND2x2_ASAP7_75t_L g667 ( .A(n_539), .B(n_583), .Y(n_667) );
BUFx2_ASAP7_75t_L g750 ( .A(n_539), .Y(n_750) );
OR2x6_ASAP7_75t_L g539 ( .A(n_540), .B(n_547), .Y(n_539) );
AOI21xp5_ASAP7_75t_L g548 ( .A1(n_549), .A2(n_555), .B(n_560), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_551), .B(n_553), .Y(n_550) );
AND2x2_ASAP7_75t_L g702 ( .A(n_551), .B(n_624), .Y(n_702) );
BUFx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g561 ( .A(n_552), .B(n_554), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_553), .B(n_623), .Y(n_724) );
INVx1_ASAP7_75t_L g754 ( .A(n_553), .Y(n_754) );
NAND2x1p5_ASAP7_75t_L g650 ( .A(n_554), .B(n_651), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_554), .B(n_690), .Y(n_727) );
INVxp67_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_557), .B(n_559), .Y(n_556) );
AND2x4_ASAP7_75t_SL g591 ( .A(n_557), .B(n_592), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_557), .B(n_585), .Y(n_738) );
INVx3_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
NOR2xp33_ASAP7_75t_L g696 ( .A(n_558), .B(n_640), .Y(n_696) );
AND2x2_ASAP7_75t_L g714 ( .A(n_558), .B(n_667), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_559), .B(n_601), .Y(n_617) );
A2O1A1Ixp33_ASAP7_75t_L g646 ( .A1(n_559), .A2(n_605), .B(n_647), .C(n_652), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_559), .B(n_677), .Y(n_676) );
AND2x2_ASAP7_75t_L g560 ( .A(n_561), .B(n_562), .Y(n_560) );
AOI221xp5_ASAP7_75t_L g741 ( .A1(n_561), .A2(n_634), .B1(n_742), .B2(n_748), .C(n_752), .Y(n_741) );
INVx1_ASAP7_75t_SL g729 ( .A(n_562), .Y(n_729) );
OAI221xp5_ASAP7_75t_L g563 ( .A1(n_564), .A2(n_574), .B1(n_580), .B2(n_584), .C(n_794), .Y(n_563) );
INVx2_ASAP7_75t_SL g564 ( .A(n_565), .Y(n_564) );
AND2x4_ASAP7_75t_L g565 ( .A(n_566), .B(n_571), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g639 ( .A(n_568), .Y(n_639) );
HB1xp67_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g613 ( .A(n_569), .B(n_614), .Y(n_613) );
AND2x2_ASAP7_75t_L g644 ( .A(n_569), .B(n_589), .Y(n_644) );
INVx2_ASAP7_75t_L g677 ( .A(n_569), .Y(n_677) );
INVx3_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
OAI32xp33_ASAP7_75t_L g728 ( .A1(n_572), .A2(n_619), .A3(n_650), .B1(n_729), .B2(n_730), .Y(n_728) );
OR2x2_ASAP7_75t_L g699 ( .A(n_573), .B(n_686), .Y(n_699) );
INVx1_ASAP7_75t_L g709 ( .A(n_574), .Y(n_709) );
OR2x2_ASAP7_75t_L g574 ( .A(n_575), .B(n_577), .Y(n_574) );
INVx2_ASAP7_75t_L g624 ( .A(n_575), .Y(n_624) );
AND2x2_ASAP7_75t_L g695 ( .A(n_575), .B(n_670), .Y(n_695) );
OR2x2_ASAP7_75t_L g726 ( .A(n_575), .B(n_727), .Y(n_726) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_576), .B(n_631), .Y(n_630) );
INVx1_ASAP7_75t_SL g577 ( .A(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g620 ( .A(n_579), .Y(n_620) );
OR2x2_ASAP7_75t_L g580 ( .A(n_581), .B(n_582), .Y(n_580) );
INVx2_ASAP7_75t_SL g585 ( .A(n_582), .Y(n_585) );
OR2x2_ASAP7_75t_L g672 ( .A(n_582), .B(n_673), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_583), .B(n_601), .Y(n_600) );
NOR2xp67_ASAP7_75t_L g706 ( .A(n_583), .B(n_707), .Y(n_706) );
BUFx2_ASAP7_75t_L g719 ( .A(n_583), .Y(n_719) );
A2O1A1Ixp33_ASAP7_75t_L g584 ( .A1(n_585), .A2(n_586), .B(n_591), .C(n_594), .Y(n_584) );
AND2x2_ASAP7_75t_L g734 ( .A(n_586), .B(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
OR2x2_ASAP7_75t_L g587 ( .A(n_588), .B(n_590), .Y(n_587) );
BUFx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
OR2x2_ASAP7_75t_L g660 ( .A(n_590), .B(n_661), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_590), .B(n_594), .Y(n_681) );
AND2x2_ASAP7_75t_L g712 ( .A(n_590), .B(n_713), .Y(n_712) );
O2A1O1Ixp33_ASAP7_75t_L g722 ( .A1(n_592), .A2(n_723), .B(n_725), .C(n_728), .Y(n_722) );
AOI222xp33_ASAP7_75t_L g596 ( .A1(n_593), .A2(n_597), .B1(n_599), .B2(n_602), .C1(n_610), .C2(n_612), .Y(n_596) );
AND2x2_ASAP7_75t_L g664 ( .A(n_593), .B(n_665), .Y(n_664) );
AND2x2_ASAP7_75t_L g597 ( .A(n_594), .B(n_598), .Y(n_597) );
INVx2_ASAP7_75t_SL g618 ( .A(n_594), .Y(n_618) );
NAND4xp25_ASAP7_75t_L g595 ( .A(n_596), .B(n_615), .C(n_636), .D(n_646), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_598), .B(n_604), .Y(n_658) );
INVx1_ASAP7_75t_SL g599 ( .A(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g666 ( .A(n_601), .B(n_667), .Y(n_666) );
INVx2_ASAP7_75t_SL g673 ( .A(n_601), .Y(n_673) );
AND2x2_ASAP7_75t_L g602 ( .A(n_603), .B(n_605), .Y(n_602) );
A2O1A1Ixp33_ASAP7_75t_L g636 ( .A1(n_603), .A2(n_637), .B(n_641), .C(n_645), .Y(n_636) );
INVx2_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_604), .B(n_619), .Y(n_740) );
OR2x2_ASAP7_75t_L g744 ( .A(n_604), .B(n_630), .Y(n_744) );
INVx1_ASAP7_75t_L g717 ( .A(n_605), .Y(n_717) );
INVx2_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .Y(n_607) );
INVx1_ASAP7_75t_SL g651 ( .A(n_608), .Y(n_651) );
INVx1_ASAP7_75t_L g631 ( .A(n_609), .Y(n_631) );
INVx2_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_611), .B(n_648), .Y(n_647) );
BUFx2_ASAP7_75t_SL g612 ( .A(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g635 ( .A(n_613), .Y(n_635) );
AOI322xp5_ASAP7_75t_L g615 ( .A1(n_616), .A2(n_618), .A3(n_619), .B1(n_621), .B2(n_625), .C1(n_626), .C2(n_632), .Y(n_615) );
INVxp67_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
O2A1O1Ixp33_ASAP7_75t_SL g697 ( .A1(n_618), .A2(n_698), .B(n_699), .C(n_700), .Y(n_697) );
INVx1_ASAP7_75t_L g720 ( .A(n_619), .Y(n_720) );
NOR2xp67_ASAP7_75t_L g621 ( .A(n_622), .B(n_624), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g678 ( .A(n_624), .B(n_679), .Y(n_678) );
AND2x2_ASAP7_75t_L g626 ( .A(n_627), .B(n_629), .Y(n_626) );
INVx2_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx2_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
HB1xp67_ASAP7_75t_L g700 ( .A(n_630), .Y(n_700) );
INVx2_ASAP7_75t_SL g632 ( .A(n_633), .Y(n_632) );
OR2x2_ASAP7_75t_L g633 ( .A(n_634), .B(n_635), .Y(n_633) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
OR2x2_ASAP7_75t_L g638 ( .A(n_639), .B(n_640), .Y(n_638) );
INVx3_ASAP7_75t_L g643 ( .A(n_640), .Y(n_643) );
OR2x2_ASAP7_75t_L g711 ( .A(n_640), .B(n_673), .Y(n_711) );
NOR2xp33_ASAP7_75t_L g756 ( .A(n_640), .B(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_643), .B(n_644), .Y(n_642) );
INVx1_ASAP7_75t_SL g743 ( .A(n_644), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_645), .B(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
NAND3xp33_ASAP7_75t_SL g748 ( .A(n_653), .B(n_749), .C(n_751), .Y(n_748) );
NOR3xp33_ASAP7_75t_SL g654 ( .A(n_655), .B(n_692), .C(n_721), .Y(n_654) );
NAND2xp5_ASAP7_75t_SL g655 ( .A(n_656), .B(n_674), .Y(n_655) );
O2A1O1Ixp33_ASAP7_75t_L g656 ( .A1(n_657), .A2(n_659), .B(n_662), .C(n_668), .Y(n_656) );
OAI31xp33_ASAP7_75t_L g701 ( .A1(n_657), .A2(n_679), .A3(n_702), .B(n_703), .Y(n_701) );
INVx1_ASAP7_75t_SL g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_SL g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
NOR2xp33_ASAP7_75t_L g663 ( .A(n_664), .B(n_666), .Y(n_663) );
INVx2_ASAP7_75t_L g716 ( .A(n_664), .Y(n_716) );
INVx1_ASAP7_75t_L g691 ( .A(n_666), .Y(n_691) );
AOI21xp5_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_671), .B(n_672), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
OR2x2_ASAP7_75t_L g718 ( .A(n_676), .B(n_719), .Y(n_718) );
INVxp67_ASAP7_75t_L g757 ( .A(n_677), .Y(n_757) );
OAI22xp33_ASAP7_75t_SL g680 ( .A1(n_681), .A2(n_682), .B1(n_687), .B2(n_691), .Y(n_680) );
INVx3_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
AND2x4_ASAP7_75t_L g683 ( .A(n_684), .B(n_685), .Y(n_683) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
HB1xp67_ASAP7_75t_L g698 ( .A(n_686), .Y(n_698) );
OR2x2_ASAP7_75t_L g749 ( .A(n_686), .B(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
NAND3xp33_ASAP7_75t_SL g692 ( .A(n_693), .B(n_701), .C(n_708), .Y(n_692) );
O2A1O1Ixp33_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_695), .B(n_696), .C(n_697), .Y(n_693) );
INVx2_ASAP7_75t_L g730 ( .A(n_694), .Y(n_730) );
INVx1_ASAP7_75t_SL g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
AOI221xp5_ASAP7_75t_L g708 ( .A1(n_709), .A2(n_710), .B1(n_712), .B2(n_714), .C(n_715), .Y(n_708) );
INVx2_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
OAI22xp33_ASAP7_75t_L g715 ( .A1(n_716), .A2(n_717), .B1(n_718), .B2(n_720), .Y(n_715) );
NAND3xp33_ASAP7_75t_SL g721 ( .A(n_722), .B(n_731), .C(n_741), .Y(n_721) );
INVxp33_ASAP7_75t_SL g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_SL g725 ( .A(n_726), .Y(n_725) );
AOI22xp5_ASAP7_75t_L g731 ( .A1(n_732), .A2(n_734), .B1(n_737), .B2(n_739), .Y(n_731) );
INVx2_ASAP7_75t_L g745 ( .A(n_732), .Y(n_745) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
OAI22xp5_ASAP7_75t_L g742 ( .A1(n_743), .A2(n_744), .B1(n_745), .B2(n_746), .Y(n_742) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
OAI22xp33_ASAP7_75t_SL g752 ( .A1(n_751), .A2(n_753), .B1(n_754), .B2(n_755), .Y(n_752) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx4_ASAP7_75t_SL g758 ( .A(n_759), .Y(n_758) );
CKINVDCx6p67_ASAP7_75t_R g771 ( .A(n_759), .Y(n_771) );
INVx3_ASAP7_75t_SL g759 ( .A(n_760), .Y(n_759) );
CKINVDCx5p33_ASAP7_75t_R g760 ( .A(n_761), .Y(n_760) );
AOI21xp5_ASAP7_75t_L g767 ( .A1(n_762), .A2(n_768), .B(n_772), .Y(n_767) );
NOR2xp33_ASAP7_75t_L g772 ( .A(n_773), .B(n_774), .Y(n_772) );
BUFx2_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
CKINVDCx16_ASAP7_75t_R g781 ( .A(n_782), .Y(n_781) );
INVx1_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
HB1xp67_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
NOR2xp33_ASAP7_75t_L g788 ( .A(n_789), .B(n_790), .Y(n_788) );
HB1xp67_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
INVx3_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
endmodule