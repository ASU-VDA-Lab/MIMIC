module fake_jpeg_8180_n_145 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_145);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_145;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx6_ASAP7_75t_SL g14 ( 
.A(n_13),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_3),
.B(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

INVx8_ASAP7_75t_SL g23 ( 
.A(n_12),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_7),
.B(n_13),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_30),
.B(n_32),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_24),
.B(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_37),
.B(n_38),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_24),
.B(n_1),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_24),
.B(n_1),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_39),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_34),
.A2(n_14),
.B1(n_18),
.B2(n_15),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_40),
.A2(n_49),
.B1(n_17),
.B2(n_20),
.Y(n_67)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_45),
.B(n_51),
.Y(n_66)
);

OR2x2_ASAP7_75t_SL g48 ( 
.A(n_35),
.B(n_28),
.Y(n_48)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_48),
.B(n_26),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_30),
.A2(n_18),
.B1(n_28),
.B2(n_15),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_51),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_53),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_38),
.C(n_28),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_54),
.B(n_16),
.C(n_58),
.Y(n_86)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_52),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_55),
.B(n_64),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_19),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_56),
.B(n_62),
.Y(n_83)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_63),
.Y(n_77)
);

OAI22x1_ASAP7_75t_SL g58 ( 
.A1(n_48),
.A2(n_29),
.B1(n_21),
.B2(n_33),
.Y(n_58)
);

AOI32xp33_ASAP7_75t_L g85 ( 
.A1(n_58),
.A2(n_69),
.A3(n_71),
.B1(n_29),
.B2(n_21),
.Y(n_85)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_18),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_61),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_33),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_50),
.B(n_15),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_43),
.A2(n_36),
.B1(n_37),
.B2(n_20),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_51),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_70),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_31),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_68),
.B(n_2),
.Y(n_90)
);

O2A1O1Ixp33_ASAP7_75t_SL g69 ( 
.A1(n_46),
.A2(n_29),
.B(n_21),
.C(n_17),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_44),
.Y(n_70)
);

OA22x2_ASAP7_75t_L g71 ( 
.A1(n_44),
.A2(n_29),
.B1(n_21),
.B2(n_26),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_41),
.B(n_19),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_73),
.Y(n_81)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_79),
.B(n_82),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_61),
.A2(n_16),
.B(n_27),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_80),
.A2(n_22),
.B(n_56),
.Y(n_100)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_85),
.A2(n_69),
.B1(n_71),
.B2(n_29),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_86),
.B(n_54),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_55),
.B(n_27),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_87),
.B(n_90),
.Y(n_92)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_4),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_91),
.B(n_93),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_86),
.B(n_73),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_89),
.A2(n_59),
.B(n_70),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_84),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_57),
.Y(n_95)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_95),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_64),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_96),
.B(n_102),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_97),
.B(n_99),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_89),
.A2(n_71),
.B(n_72),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_100),
.B(n_81),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_75),
.A2(n_71),
.B1(n_29),
.B2(n_21),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_101),
.A2(n_103),
.B1(n_90),
.B2(n_76),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_2),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_77),
.A2(n_22),
.B1(n_21),
.B2(n_53),
.Y(n_103)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_104),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_98),
.B(n_75),
.Y(n_106)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_106),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_110),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_96),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_96),
.B(n_91),
.Y(n_111)
);

FAx1_ASAP7_75t_SL g118 ( 
.A(n_111),
.B(n_100),
.CI(n_80),
.CON(n_118),
.SN(n_118)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_113),
.A2(n_115),
.B1(n_103),
.B2(n_74),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_114),
.B(n_93),
.C(n_101),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_116),
.B(n_118),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_105),
.Y(n_117)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_117),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_114),
.B(n_88),
.C(n_78),
.Y(n_120)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_120),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_107),
.B(n_102),
.Y(n_122)
);

OAI21xp33_ASAP7_75t_SL g126 ( 
.A1(n_122),
.A2(n_123),
.B(n_105),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_126),
.A2(n_129),
.B(n_121),
.Y(n_131)
);

AOI322xp5_ASAP7_75t_L g128 ( 
.A1(n_122),
.A2(n_108),
.A3(n_111),
.B1(n_115),
.B2(n_102),
.C1(n_106),
.C2(n_92),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_128),
.B(n_120),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_119),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_125),
.B(n_116),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_130),
.B(n_134),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_131),
.B(n_132),
.Y(n_138)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_127),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_126),
.Y(n_133)
);

OAI31xp33_ASAP7_75t_L g136 ( 
.A1(n_133),
.A2(n_118),
.A3(n_124),
.B(n_83),
.Y(n_136)
);

HAxp5_ASAP7_75t_SL g135 ( 
.A(n_130),
.B(n_117),
.CON(n_135),
.SN(n_135)
);

AO21x1_ASAP7_75t_L g141 ( 
.A1(n_135),
.A2(n_136),
.B(n_11),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_137),
.B(n_112),
.C(n_83),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_139),
.B(n_140),
.C(n_135),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_137),
.B(n_118),
.C(n_84),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_141),
.A2(n_138),
.B1(n_5),
.B2(n_9),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_142),
.Y(n_144)
);

AOI221xp5_ASAP7_75t_L g145 ( 
.A1(n_144),
.A2(n_143),
.B1(n_5),
.B2(n_10),
.C(n_11),
.Y(n_145)
);


endmodule