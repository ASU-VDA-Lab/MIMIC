module fake_jpeg_16678_n_67 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_67);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_67;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_50;
wire n_43;
wire n_12;
wire n_32;
wire n_15;
wire n_66;

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_6),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_0),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_0),
.B(n_5),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

AOI21xp33_ASAP7_75t_L g17 ( 
.A1(n_3),
.A2(n_4),
.B(n_2),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

HB1xp67_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_21),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_18),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_20),
.A2(n_18),
.B1(n_10),
.B2(n_17),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_12),
.B(n_1),
.Y(n_21)
);

BUFx2_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

INVx2_ASAP7_75t_SL g30 ( 
.A(n_22),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

OR2x2_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_24),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_12),
.B(n_2),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_25),
.A2(n_17),
.B1(n_10),
.B2(n_13),
.Y(n_36)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_21),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_31),
.B(n_32),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_29),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_29),
.B(n_26),
.Y(n_33)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_28),
.Y(n_34)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

AOI32xp33_ASAP7_75t_L g46 ( 
.A1(n_36),
.A2(n_16),
.A3(n_14),
.B1(n_15),
.B2(n_5),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

AO21x2_ASAP7_75t_SL g41 ( 
.A1(n_37),
.A2(n_30),
.B(n_28),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_30),
.A2(n_20),
.B1(n_13),
.B2(n_3),
.Y(n_39)
);

XOR2xp5_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_40),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_9),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_41),
.A2(n_35),
.B1(n_14),
.B2(n_15),
.Y(n_52)
);

NAND2xp33_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_9),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_45),
.B(n_38),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_46),
.A2(n_39),
.B1(n_16),
.B2(n_37),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_48),
.A2(n_50),
.B1(n_52),
.B2(n_42),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_38),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_SL g55 ( 
.A(n_49),
.B(n_47),
.Y(n_55)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_51),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_42),
.B(n_44),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_53),
.B(n_41),
.C(n_43),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_54),
.B(n_52),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_55),
.B(n_56),
.C(n_41),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_SL g61 ( 
.A1(n_58),
.A2(n_59),
.B(n_55),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_57),
.A2(n_49),
.B1(n_41),
.B2(n_35),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_60),
.B(n_14),
.C(n_15),
.Y(n_62)
);

AO21x1_ASAP7_75t_L g64 ( 
.A1(n_61),
.A2(n_4),
.B(n_8),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_62),
.B(n_60),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_63),
.Y(n_65)
);

INVxp33_ASAP7_75t_L g66 ( 
.A(n_65),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_66),
.B(n_64),
.Y(n_67)
);


endmodule