module fake_jpeg_14427_n_238 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_238);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_238;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_122;
wire n_75;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

CKINVDCx9p33_ASAP7_75t_R g38 ( 
.A(n_25),
.Y(n_38)
);

CKINVDCx6p67_ASAP7_75t_R g82 ( 
.A(n_38),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_19),
.B(n_14),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_39),
.B(n_42),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_26),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_41),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_26),
.B(n_0),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_25),
.B(n_1),
.C(n_2),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_20),
.B(n_14),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_48),
.B(n_53),
.Y(n_65)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_30),
.B(n_1),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_54),
.Y(n_97)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_1),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_59),
.Y(n_74)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_30),
.B(n_3),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_61),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_33),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_62),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_38),
.A2(n_21),
.B1(n_28),
.B2(n_22),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_63),
.A2(n_70),
.B1(n_90),
.B2(n_91),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_51),
.A2(n_28),
.B1(n_27),
.B2(n_36),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_40),
.B(n_27),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_71),
.B(n_73),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_41),
.B(n_42),
.Y(n_73)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_77),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_55),
.B(n_35),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_86),
.Y(n_99)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_84),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_56),
.B(n_35),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_85),
.B(n_88),
.Y(n_101)
);

NOR2x1_ASAP7_75t_L g86 ( 
.A(n_56),
.B(n_33),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_44),
.B(n_17),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_45),
.A2(n_36),
.B1(n_31),
.B2(n_24),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_47),
.A2(n_31),
.B1(n_24),
.B2(n_17),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_50),
.B(n_34),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_92),
.B(n_94),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_54),
.B(n_34),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_59),
.B(n_29),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_96),
.B(n_98),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_58),
.B(n_29),
.Y(n_98)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_100),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_73),
.A2(n_62),
.B1(n_52),
.B2(n_43),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_104),
.A2(n_128),
.B1(n_102),
.B2(n_125),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_67),
.B(n_49),
.C(n_4),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_105),
.B(n_8),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_66),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_110),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_67),
.B(n_71),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_108),
.B(n_122),
.Y(n_138)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_74),
.A2(n_3),
.B(n_5),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_111),
.A2(n_72),
.B(n_82),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_83),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_112),
.B(n_115),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_64),
.B(n_78),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_114),
.B(n_117),
.Y(n_149)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_69),
.Y(n_115)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_116),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_65),
.B(n_10),
.Y(n_117)
);

INVx2_ASAP7_75t_SL g118 ( 
.A(n_89),
.Y(n_118)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_118),
.Y(n_143)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_93),
.Y(n_119)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_119),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_74),
.B(n_5),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_121),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_86),
.B(n_7),
.Y(n_122)
);

BUFx2_ASAP7_75t_L g123 ( 
.A(n_76),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_123),
.Y(n_135)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_69),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_124),
.B(n_126),
.Y(n_141)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_80),
.Y(n_125)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_125),
.Y(n_153)
);

OAI32xp33_ASAP7_75t_L g126 ( 
.A1(n_74),
.A2(n_8),
.A3(n_9),
.B1(n_10),
.B2(n_87),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_95),
.B(n_79),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_127),
.B(n_102),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_95),
.A2(n_8),
.B1(n_9),
.B2(n_80),
.Y(n_128)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_76),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_129),
.B(n_82),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_112),
.A2(n_82),
.B1(n_68),
.B2(n_89),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_130),
.B(n_132),
.Y(n_160)
);

OAI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_104),
.A2(n_82),
.B1(n_79),
.B2(n_97),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_133),
.B(n_152),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_127),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_151),
.Y(n_158)
);

OAI21xp33_ASAP7_75t_L g167 ( 
.A1(n_139),
.A2(n_155),
.B(n_126),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_140),
.B(n_148),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_107),
.A2(n_75),
.B1(n_72),
.B2(n_97),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_144),
.A2(n_121),
.B(n_109),
.Y(n_165)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_145),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_101),
.B(n_81),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_121),
.B(n_81),
.Y(n_150)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_150),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_122),
.B(n_75),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_99),
.B(n_108),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_154),
.B(n_103),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_105),
.B(n_111),
.Y(n_155)
);

AOI221xp5_ASAP7_75t_L g192 ( 
.A1(n_157),
.A2(n_167),
.B1(n_176),
.B2(n_146),
.C(n_141),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_149),
.B(n_113),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_161),
.B(n_164),
.Y(n_182)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_143),
.Y(n_162)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_162),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_149),
.B(n_120),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_165),
.A2(n_150),
.B(n_151),
.Y(n_180)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_143),
.Y(n_166)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_166),
.Y(n_189)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_131),
.Y(n_168)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_168),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_148),
.B(n_120),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_169),
.B(n_134),
.Y(n_193)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_131),
.Y(n_170)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_170),
.Y(n_191)
);

OR2x2_ASAP7_75t_L g171 ( 
.A(n_154),
.B(n_129),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_171),
.A2(n_133),
.B(n_134),
.Y(n_179)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_137),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_172),
.B(n_173),
.Y(n_185)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_137),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_137),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_174),
.B(n_175),
.Y(n_187)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_145),
.Y(n_175)
);

OAI21xp33_ASAP7_75t_L g176 ( 
.A1(n_150),
.A2(n_128),
.B(n_100),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_158),
.B(n_159),
.Y(n_178)
);

OAI322xp33_ASAP7_75t_L g204 ( 
.A1(n_178),
.A2(n_193),
.A3(n_162),
.B1(n_174),
.B2(n_173),
.C1(n_172),
.C2(n_147),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_179),
.A2(n_194),
.B(n_180),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_180),
.B(n_192),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_177),
.B(n_140),
.C(n_155),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_181),
.B(n_178),
.C(n_171),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_158),
.A2(n_141),
.B1(n_136),
.B2(n_144),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_183),
.A2(n_188),
.B1(n_156),
.B2(n_166),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_171),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_186),
.B(n_168),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_159),
.A2(n_152),
.B1(n_160),
.B2(n_170),
.Y(n_188)
);

A2O1A1O1Ixp25_ASAP7_75t_L g194 ( 
.A1(n_177),
.A2(n_138),
.B(n_146),
.C(n_139),
.D(n_118),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_195),
.B(n_198),
.Y(n_214)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_187),
.Y(n_196)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_196),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_181),
.B(n_163),
.C(n_159),
.Y(n_198)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_199),
.Y(n_210)
);

AOI322xp5_ASAP7_75t_SL g200 ( 
.A1(n_182),
.A2(n_138),
.A3(n_139),
.B1(n_160),
.B2(n_163),
.C1(n_165),
.C2(n_175),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_200),
.B(n_201),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_190),
.B(n_156),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_202),
.B(n_204),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_190),
.B(n_147),
.Y(n_203)
);

AOI322xp5_ASAP7_75t_L g211 ( 
.A1(n_203),
.A2(n_191),
.A3(n_184),
.B1(n_189),
.B2(n_142),
.C1(n_187),
.C2(n_153),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_186),
.A2(n_153),
.B1(n_135),
.B2(n_142),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_205),
.A2(n_206),
.B(n_191),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_185),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_207),
.B(n_194),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_211),
.A2(n_202),
.B1(n_196),
.B2(n_206),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_207),
.A2(n_179),
.B(n_188),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_213),
.B(n_197),
.Y(n_219)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_215),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_216),
.B(n_205),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_217),
.B(n_212),
.C(n_208),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_219),
.B(n_222),
.Y(n_225)
);

INVxp67_ASAP7_75t_SL g220 ( 
.A(n_210),
.Y(n_220)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_220),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_209),
.A2(n_195),
.B1(n_198),
.B2(n_197),
.Y(n_221)
);

OR2x2_ASAP7_75t_L g228 ( 
.A(n_221),
.B(n_223),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_216),
.A2(n_184),
.B1(n_189),
.B2(n_185),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_226),
.B(n_227),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_221),
.B(n_214),
.C(n_222),
.Y(n_227)
);

O2A1O1Ixp33_ASAP7_75t_SL g229 ( 
.A1(n_228),
.A2(n_218),
.B(n_215),
.C(n_213),
.Y(n_229)
);

A2O1A1Ixp33_ASAP7_75t_SL g233 ( 
.A1(n_229),
.A2(n_232),
.B(n_212),
.C(n_225),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_224),
.B(n_214),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_231),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_228),
.A2(n_218),
.B(n_223),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_233),
.A2(n_230),
.B1(n_118),
.B2(n_123),
.Y(n_236)
);

BUFx24_ASAP7_75t_SL g235 ( 
.A(n_234),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_235),
.B(n_236),
.C(n_116),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_237),
.B(n_119),
.Y(n_238)
);


endmodule