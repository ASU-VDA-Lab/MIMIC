module real_jpeg_19767_n_16 (n_333, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_333;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_0),
.A2(n_26),
.B1(n_33),
.B2(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_0),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_0),
.A2(n_30),
.B1(n_31),
.B2(n_132),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_0),
.A2(n_44),
.B1(n_45),
.B2(n_132),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_0),
.A2(n_62),
.B1(n_63),
.B2(n_132),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g130 ( 
.A(n_1),
.Y(n_130)
);

AOI21xp33_ASAP7_75t_L g178 ( 
.A1(n_1),
.A2(n_14),
.B(n_63),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_1),
.A2(n_44),
.B1(n_45),
.B2(n_130),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_1),
.A2(n_105),
.B1(n_186),
.B2(n_187),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_1),
.B(n_87),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_1),
.B(n_31),
.Y(n_215)
);

AOI21xp33_ASAP7_75t_L g219 ( 
.A1(n_1),
.A2(n_31),
.B(n_215),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_3),
.A2(n_30),
.B1(n_31),
.B2(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_3),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_3),
.A2(n_26),
.B1(n_33),
.B2(n_125),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_3),
.A2(n_62),
.B1(n_63),
.B2(n_125),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_3),
.A2(n_44),
.B1(n_45),
.B2(n_125),
.Y(n_204)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_4),
.Y(n_106)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_4),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_4),
.A2(n_139),
.B(n_161),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_4),
.A2(n_170),
.B1(n_171),
.B2(n_173),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_5),
.A2(n_26),
.B1(n_33),
.B2(n_34),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_5),
.A2(n_34),
.B1(n_44),
.B2(n_45),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_5),
.A2(n_34),
.B1(n_62),
.B2(n_63),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_5),
.A2(n_30),
.B1(n_31),
.B2(n_34),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_6),
.A2(n_30),
.B1(n_31),
.B2(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_6),
.A2(n_44),
.B1(n_45),
.B2(n_50),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_6),
.A2(n_50),
.B1(n_62),
.B2(n_63),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_6),
.A2(n_26),
.B1(n_33),
.B2(n_50),
.Y(n_285)
);

BUFx8_ASAP7_75t_L g63 ( 
.A(n_7),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_8),
.A2(n_30),
.B1(n_31),
.B2(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_8),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_8),
.A2(n_26),
.B1(n_33),
.B2(n_57),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_8),
.A2(n_57),
.B1(n_62),
.B2(n_63),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_8),
.A2(n_44),
.B1(n_45),
.B2(n_57),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_9),
.A2(n_26),
.B1(n_33),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_9),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_9),
.A2(n_30),
.B1(n_31),
.B2(n_36),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_9),
.A2(n_36),
.B1(n_62),
.B2(n_63),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_9),
.A2(n_36),
.B1(n_44),
.B2(n_45),
.Y(n_257)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_11),
.A2(n_30),
.B1(n_31),
.B2(n_127),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_11),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_11),
.A2(n_62),
.B1(n_63),
.B2(n_127),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_11),
.A2(n_44),
.B1(n_45),
.B2(n_127),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_11),
.A2(n_26),
.B1(n_33),
.B2(n_127),
.Y(n_265)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_13),
.A2(n_25),
.B1(n_30),
.B2(n_31),
.Y(n_29)
);

A2O1A1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_14),
.A2(n_44),
.B(n_60),
.C(n_61),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_14),
.B(n_44),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_14),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_61)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_14),
.Y(n_64)
);

INVx11_ASAP7_75t_SL g46 ( 
.A(n_15),
.Y(n_46)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_94),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_92),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_78),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_19),
.B(n_78),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_70),
.C(n_73),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_20),
.A2(n_21),
.B1(n_70),
.B2(n_319),
.Y(n_325)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_38),
.B1(n_39),
.B2(n_69),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_22),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_32),
.B1(n_35),
.B2(n_37),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_23),
.A2(n_37),
.B1(n_144),
.B2(n_145),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_23),
.A2(n_37),
.B1(n_145),
.B2(n_265),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_23),
.A2(n_265),
.B(n_284),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_23),
.A2(n_84),
.B(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_24),
.B(n_72),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_24),
.A2(n_82),
.B(n_83),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_24),
.A2(n_29),
.B1(n_129),
.B2(n_131),
.Y(n_128)
);

O2A1O1Ixp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B(n_28),
.C(n_29),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_25),
.B(n_26),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_25),
.B(n_31),
.Y(n_136)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

HAxp5_ASAP7_75t_SL g129 ( 
.A(n_26),
.B(n_130),
.CON(n_129),
.SN(n_129)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_28),
.A2(n_30),
.B1(n_129),
.B2(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_29),
.B(n_72),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_29),
.B(n_285),
.Y(n_284)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_30),
.Y(n_31)
);

AOI32xp33_ASAP7_75t_L g214 ( 
.A1(n_30),
.A2(n_44),
.A3(n_48),
.B1(n_215),
.B2(n_216),
.Y(n_214)
);

A2O1A1Ixp33_ASAP7_75t_L g53 ( 
.A1(n_31),
.A2(n_43),
.B(n_47),
.C(n_54),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_31),
.B(n_47),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_32),
.A2(n_37),
.B(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_35),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_37),
.B(n_130),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_58),
.B1(n_67),
.B2(n_68),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_40),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_51),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_42),
.A2(n_52),
.B(n_148),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_49),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_43),
.B(n_56),
.Y(n_77)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_43),
.A2(n_53),
.B1(n_124),
.B2(n_126),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_43),
.A2(n_53),
.B1(n_124),
.B2(n_157),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_43),
.A2(n_53),
.B1(n_157),
.B2(n_219),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_43),
.A2(n_51),
.B(n_281),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_43),
.A2(n_53),
.B1(n_76),
.B2(n_281),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_44),
.A2(n_45),
.B1(n_47),
.B2(n_48),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

A2O1A1Ixp33_ASAP7_75t_L g177 ( 
.A1(n_45),
.A2(n_64),
.B(n_130),
.C(n_178),
.Y(n_177)
);

NAND2xp33_ASAP7_75t_SL g216 ( 
.A(n_45),
.B(n_47),
.Y(n_216)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_49),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_52),
.B(n_55),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_52),
.A2(n_75),
.B(n_77),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_52),
.A2(n_87),
.B(n_88),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_52),
.A2(n_77),
.B(n_88),
.Y(n_267)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_58),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_58),
.B(n_68),
.C(n_69),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_58),
.A2(n_67),
.B1(n_74),
.B2(n_322),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_61),
.B(n_65),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_59),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_59),
.A2(n_65),
.B(n_120),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_59),
.A2(n_61),
.B1(n_181),
.B2(n_182),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_59),
.A2(n_61),
.B1(n_182),
.B2(n_204),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_59),
.A2(n_61),
.B1(n_204),
.B2(n_222),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_59),
.A2(n_222),
.B(n_238),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_59),
.A2(n_61),
.B1(n_112),
.B2(n_257),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_59),
.A2(n_120),
.B(n_257),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_61),
.A2(n_112),
.B(n_113),
.Y(n_111)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_61),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_61),
.B(n_130),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_62),
.B(n_193),
.Y(n_192)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_63),
.B(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_66),
.B(n_121),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_67),
.B(n_70),
.C(n_74),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_70),
.A2(n_319),
.B1(n_320),
.B2(n_321),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_70),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_73),
.B(n_325),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_74),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_79),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_81),
.B1(n_85),
.B2(n_86),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

OAI321xp33_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_316),
.A3(n_326),
.B1(n_329),
.B2(n_330),
.C(n_333),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_296),
.B(n_315),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_272),
.B(n_295),
.Y(n_96)
);

O2A1O1Ixp33_ASAP7_75t_SL g97 ( 
.A1(n_98),
.A2(n_162),
.B(n_247),
.C(n_271),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_150),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_99),
.B(n_150),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_101),
.B1(n_133),
.B2(n_149),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_SL g101 ( 
.A(n_102),
.B(n_117),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_102),
.B(n_117),
.C(n_149),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_104),
.B1(n_111),
.B2(n_116),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_103),
.B(n_116),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_107),
.B(n_108),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_105),
.A2(n_107),
.B1(n_138),
.B2(n_140),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_105),
.B(n_110),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g170 ( 
.A(n_105),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_105),
.A2(n_172),
.B1(n_186),
.B2(n_187),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_105),
.A2(n_174),
.B(n_206),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_105),
.A2(n_106),
.B(n_291),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_106),
.B(n_110),
.Y(n_109)
);

INVx5_ASAP7_75t_L g188 ( 
.A(n_106),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_106),
.B(n_130),
.Y(n_193)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_109),
.A2(n_170),
.B(n_207),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_111),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_113),
.B(n_238),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_115),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_114),
.B(n_121),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_122),
.C(n_128),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_118),
.A2(n_119),
.B1(n_122),
.B2(n_123),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_126),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_SL g151 ( 
.A(n_128),
.B(n_152),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_131),
.Y(n_144)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_133),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_141),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_134),
.B(n_142),
.C(n_147),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_137),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_135),
.B(n_137),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_142),
.A2(n_143),
.B1(n_146),
.B2(n_147),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_153),
.C(n_155),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_151),
.B(n_243),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_153),
.A2(n_154),
.B1(n_155),
.B2(n_244),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_155),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_158),
.C(n_159),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_156),
.B(n_232),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_158),
.A2(n_159),
.B1(n_160),
.B2(n_233),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_158),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_161),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_163),
.B(n_246),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_240),
.B(n_245),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_227),
.B(n_239),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_209),
.B(n_226),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_196),
.B(n_208),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_183),
.B(n_195),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_175),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_169),
.B(n_175),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_177),
.B1(n_179),
.B2(n_180),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_177),
.B(n_179),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_180),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_184),
.A2(n_190),
.B(n_194),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_189),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_185),
.B(n_189),
.Y(n_194)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_188),
.B(n_207),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_197),
.B(n_198),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_205),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_201),
.B1(n_202),
.B2(n_203),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_200),
.B(n_203),
.C(n_205),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_203),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_206),
.B(n_255),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_207),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_210),
.B(n_211),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_217),
.B1(n_224),
.B2(n_225),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_212),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_213),
.B(n_214),
.Y(n_236)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_217),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_220),
.B1(n_221),
.B2(n_223),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_218),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_220),
.B(n_223),
.C(n_224),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_221),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_228),
.B(n_229),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_230),
.A2(n_231),
.B1(n_234),
.B2(n_235),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_230),
.B(n_236),
.C(n_237),
.Y(n_241)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_235),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_241),
.B(n_242),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_248),
.B(n_249),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_269),
.B2(n_270),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_253),
.B1(n_258),
.B2(n_259),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_252),
.B(n_259),
.C(n_270),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_253),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_256),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_254),
.B(n_256),
.Y(n_278)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_260),
.A2(n_261),
.B1(n_262),
.B2(n_268),
.Y(n_259)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_260),
.Y(n_268)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_266),
.B2(n_267),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_263),
.B(n_267),
.C(n_268),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_264),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_267),
.Y(n_266)
);

CKINVDCx14_ASAP7_75t_R g270 ( 
.A(n_269),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_273),
.B(n_274),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_294),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_276),
.A2(n_277),
.B1(n_287),
.B2(n_288),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_276),
.B(n_288),
.C(n_294),
.Y(n_297)
);

CKINVDCx14_ASAP7_75t_R g276 ( 
.A(n_277),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_278),
.B(n_282),
.C(n_286),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_280),
.A2(n_282),
.B1(n_283),
.B2(n_286),
.Y(n_279)
);

CKINVDCx14_ASAP7_75t_R g286 ( 
.A(n_280),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_283),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_285),
.Y(n_311)
);

CKINVDCx14_ASAP7_75t_R g287 ( 
.A(n_288),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_289),
.A2(n_290),
.B1(n_292),
.B2(n_293),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_289),
.A2(n_290),
.B1(n_310),
.B2(n_312),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_289),
.A2(n_306),
.B(n_310),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_290),
.B(n_292),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_292),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_297),
.B(n_298),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_299),
.A2(n_300),
.B1(n_313),
.B2(n_314),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_305),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_301),
.B(n_305),
.C(n_314),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_302),
.A2(n_303),
.B(n_304),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_302),
.B(n_303),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_304),
.B(n_318),
.C(n_323),
.Y(n_317)
);

FAx1_ASAP7_75t_SL g328 ( 
.A(n_304),
.B(n_318),
.CI(n_323),
.CON(n_328),
.SN(n_328)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_306),
.A2(n_307),
.B1(n_308),
.B2(n_309),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_310),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_313),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_324),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_317),
.B(n_324),
.Y(n_330)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_327),
.B(n_328),
.Y(n_329)
);

BUFx24_ASAP7_75t_SL g331 ( 
.A(n_328),
.Y(n_331)
);


endmodule