module real_jpeg_26735_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_131;
wire n_47;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_173;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_195;
wire n_61;
wire n_110;
wire n_258;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_278;
wire n_130;
wire n_144;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_277;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_187;
wire n_97;
wire n_75;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_202;
wire n_244;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_269;
wire n_96;
wire n_273;
wire n_253;
wire n_89;

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_0),
.Y(n_65)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_0),
.Y(n_66)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_0),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_1),
.A2(n_78),
.B1(n_79),
.B2(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_1),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_1),
.A2(n_49),
.B1(n_50),
.B2(n_151),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_1),
.A2(n_27),
.B1(n_30),
.B2(n_151),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_1),
.A2(n_33),
.B1(n_36),
.B2(n_151),
.Y(n_236)
);

OAI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_2),
.A2(n_27),
.B1(n_30),
.B2(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_2),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_2),
.A2(n_43),
.B1(n_78),
.B2(n_79),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_2),
.A2(n_33),
.B1(n_36),
.B2(n_43),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_2),
.A2(n_43),
.B1(n_49),
.B2(n_50),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_3),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_3),
.A2(n_29),
.B1(n_33),
.B2(n_36),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_3),
.A2(n_29),
.B1(n_78),
.B2(n_79),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_3),
.A2(n_29),
.B1(n_49),
.B2(n_50),
.Y(n_126)
);

BUFx12_ASAP7_75t_L g77 ( 
.A(n_4),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_6),
.A2(n_78),
.B1(n_79),
.B2(n_131),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_6),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_6),
.A2(n_49),
.B1(n_50),
.B2(n_131),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_6),
.A2(n_27),
.B1(n_30),
.B2(n_131),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_6),
.A2(n_33),
.B1(n_36),
.B2(n_131),
.Y(n_228)
);

INVx13_ASAP7_75t_L g79 ( 
.A(n_7),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_8),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_8),
.B(n_81),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_8),
.B(n_49),
.Y(n_188)
);

AOI21xp33_ASAP7_75t_L g192 ( 
.A1(n_8),
.A2(n_49),
.B(n_188),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_8),
.A2(n_27),
.B1(n_30),
.B2(n_149),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_8),
.A2(n_33),
.B(n_37),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_8),
.B(n_99),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_8),
.A2(n_63),
.B1(n_66),
.B2(n_236),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_9),
.A2(n_49),
.B1(n_50),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_9),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_9),
.A2(n_27),
.B1(n_30),
.B2(n_56),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_9),
.A2(n_33),
.B1(n_36),
.B2(n_56),
.Y(n_165)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_11),
.A2(n_49),
.B1(n_50),
.B2(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_11),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_11),
.A2(n_27),
.B1(n_30),
.B2(n_58),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_11),
.A2(n_33),
.B1(n_36),
.B2(n_58),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_12),
.A2(n_78),
.B1(n_79),
.B2(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_12),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_12),
.A2(n_49),
.B1(n_50),
.B2(n_106),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_12),
.A2(n_27),
.B1(n_30),
.B2(n_106),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_12),
.A2(n_33),
.B1(n_36),
.B2(n_106),
.Y(n_223)
);

BUFx24_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_14),
.A2(n_27),
.B1(n_30),
.B2(n_52),
.Y(n_53)
);

INVx11_ASAP7_75t_SL g34 ( 
.A(n_15),
.Y(n_34)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_133),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_132),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_109),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_20),
.B(n_109),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_87),
.B2(n_108),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_60),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_44),
.B(n_59),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_24),
.B(n_44),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_38),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_25),
.A2(n_40),
.B(n_196),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_31),
.Y(n_25)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_26),
.Y(n_142)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

OAI22xp33_ASAP7_75t_L g41 ( 
.A1(n_27),
.A2(n_30),
.B1(n_35),
.B2(n_37),
.Y(n_41)
);

NAND2xp33_ASAP7_75t_SL g189 ( 
.A(n_27),
.B(n_47),
.Y(n_189)
);

A2O1A1Ixp33_ASAP7_75t_L g214 ( 
.A1(n_27),
.A2(n_35),
.B(n_149),
.C(n_215),
.Y(n_214)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI32xp33_ASAP7_75t_L g186 ( 
.A1(n_30),
.A2(n_50),
.A3(n_187),
.B1(n_188),
.B2(n_189),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_31),
.B(n_42),
.Y(n_71)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_41),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_32),
.A2(n_40),
.B1(n_70),
.B2(n_97),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_32),
.A2(n_38),
.B(n_97),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_32),
.A2(n_40),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_32),
.A2(n_40),
.B1(n_212),
.B2(n_213),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_32),
.A2(n_40),
.B1(n_195),
.B2(n_213),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_32),
.B(n_149),
.Y(n_234)
);

OA22x2_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_32)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_36),
.B(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_36),
.B(n_240),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_39),
.B(n_42),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g69 ( 
.A1(n_40),
.A2(n_70),
.B(n_71),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_40),
.A2(n_71),
.B(n_142),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_45),
.A2(n_53),
.B1(n_54),
.B2(n_57),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_45),
.B(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_45),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_45),
.A2(n_53),
.B1(n_145),
.B2(n_146),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_45),
.A2(n_53),
.B1(n_145),
.B2(n_174),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_45),
.A2(n_53),
.B1(n_174),
.B2(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_53),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_49),
.B1(n_50),
.B2(n_52),
.Y(n_46)
);

INVx6_ASAP7_75t_L g187 ( 
.A(n_47),
.Y(n_187)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_49),
.A2(n_50),
.B1(n_76),
.B2(n_77),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_49),
.B(n_76),
.Y(n_163)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_50),
.A2(n_80),
.B1(n_148),
.B2(n_163),
.Y(n_162)
);

BUFx4f_ASAP7_75t_SL g50 ( 
.A(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_53),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_53),
.B(n_101),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_53),
.B(n_126),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_55),
.A2(n_99),
.B(n_100),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_72),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_69),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_62),
.A2(n_73),
.B1(n_74),
.B2(n_86),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_62),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_62),
.A2(n_69),
.B1(n_86),
.B2(n_115),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_66),
.B(n_67),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_63),
.A2(n_119),
.B(n_120),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_63),
.A2(n_95),
.B1(n_119),
.B2(n_165),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_63),
.A2(n_93),
.B(n_223),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_63),
.A2(n_66),
.B1(n_228),
.B2(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_64),
.B(n_91),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_64),
.A2(n_68),
.B(n_121),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_64),
.A2(n_94),
.B1(n_227),
.B2(n_229),
.Y(n_226)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_65),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_66),
.B(n_92),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_66),
.A2(n_90),
.B(n_165),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_68),
.B(n_94),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_69),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_82),
.B(n_83),
.Y(n_74)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_75),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_75),
.A2(n_81),
.B1(n_148),
.B2(n_150),
.Y(n_147)
);

O2A1O1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_78),
.B(n_80),
.C(n_81),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_76),
.B(n_78),
.Y(n_80)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

HAxp5_ASAP7_75t_SL g148 ( 
.A(n_78),
.B(n_149),
.CON(n_148),
.SN(n_148)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_81),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_81),
.B(n_82),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_85),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_84),
.A2(n_104),
.B1(n_105),
.B2(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_84),
.A2(n_104),
.B1(n_130),
.B2(n_156),
.Y(n_155)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_87),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_98),
.C(n_102),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_96),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_89),
.B(n_96),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_93),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_98),
.A2(n_102),
.B1(n_103),
.B2(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_98),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_104),
.A2(n_105),
.B(n_107),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_114),
.C(n_116),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_110),
.A2(n_111),
.B1(n_114),
.B2(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_114),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_116),
.B(n_277),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_123),
.C(n_128),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_117),
.B(n_269),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_122),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_122),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_123),
.A2(n_128),
.B1(n_129),
.B2(n_270),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_123),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_125),
.B(n_127),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_124),
.A2(n_159),
.B(n_160),
.Y(n_158)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_274),
.B(n_279),
.Y(n_133)
);

O2A1O1Ixp33_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_178),
.B(n_260),
.C(n_273),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_166),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_136),
.B(n_166),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_152),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_139),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_138),
.B(n_139),
.C(n_152),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_143),
.C(n_147),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_140),
.A2(n_141),
.B1(n_143),
.B2(n_144),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_146),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g168 ( 
.A(n_147),
.B(n_169),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_149),
.B(n_241),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_150),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_153),
.B(n_161),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_155),
.B1(n_157),
.B2(n_158),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_154),
.B(n_158),
.C(n_161),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_164),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_162),
.B(n_164),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_170),
.C(n_172),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_167),
.A2(n_168),
.B1(n_255),
.B2(n_257),
.Y(n_254)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_170),
.A2(n_171),
.B1(n_172),
.B2(n_256),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_172),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_175),
.C(n_177),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_173),
.B(n_200),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_175),
.A2(n_176),
.B1(n_177),
.B2(n_201),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_177),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_179),
.B(n_259),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_252),
.B(n_258),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_206),
.B(n_251),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_197),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_182),
.B(n_197),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_190),
.C(n_193),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_183),
.A2(n_184),
.B1(n_248),
.B2(n_249),
.Y(n_247)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_185),
.B(n_186),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_190),
.A2(n_191),
.B1(n_193),
.B2(n_194),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_198),
.A2(n_199),
.B1(n_202),
.B2(n_203),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_198),
.B(n_204),
.C(n_205),
.Y(n_253)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_245),
.B(n_250),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_224),
.B(n_244),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_216),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_209),
.B(n_216),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_210),
.B(n_214),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_210),
.A2(n_211),
.B1(n_214),
.B2(n_231),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_214),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_222),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_220),
.B2(n_221),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_218),
.B(n_221),
.C(n_222),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_219),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_221),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_223),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_232),
.B(n_243),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_230),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_226),
.B(n_230),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_237),
.B(n_242),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_234),
.B(n_235),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_246),
.B(n_247),
.Y(n_250)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_253),
.B(n_254),
.Y(n_258)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_255),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_261),
.B(n_262),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_271),
.B2(n_272),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_267),
.B2(n_268),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_265),
.B(n_268),
.C(n_272),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_271),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_275),
.B(n_276),
.Y(n_279)
);


endmodule