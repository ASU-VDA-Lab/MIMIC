module real_aes_12461_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_924, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_924;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_887;
wire n_187;
wire n_436;
wire n_599;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_905;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_919;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_666;
wire n_320;
wire n_537;
wire n_551;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_889;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_356;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_892;
wire n_528;
wire n_578;
wire n_202;
wire n_372;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_920;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_909;
wire n_298;
wire n_523;
wire n_860;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_913;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_917;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_898;
wire n_115;
wire n_604;
wire n_110;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_756;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_891;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_914;
wire n_707;
wire n_622;
wire n_915;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_907;
wire n_847;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_899;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_922;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_888;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_911;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
INVx2_ASAP7_75t_SL g633 ( .A(n_0), .Y(n_633) );
CKINVDCx5p33_ASAP7_75t_R g530 ( .A(n_1), .Y(n_530) );
OA21x2_ASAP7_75t_L g134 ( .A1(n_2), .A2(n_47), .B(n_135), .Y(n_134) );
INVx1_ASAP7_75t_L g233 ( .A(n_2), .Y(n_233) );
NAND2xp5_ASAP7_75t_SL g589 ( .A(n_3), .B(n_217), .Y(n_589) );
NAND2xp5_ASAP7_75t_SL g643 ( .A(n_4), .B(n_212), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_5), .B(n_252), .Y(n_251) );
NAND2xp33_ASAP7_75t_L g272 ( .A(n_6), .B(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g555 ( .A(n_7), .B(n_167), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_8), .B(n_143), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_9), .B(n_176), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_10), .B(n_179), .Y(n_584) );
CKINVDCx5p33_ASAP7_75t_R g288 ( .A(n_11), .Y(n_288) );
BUFx3_ASAP7_75t_L g141 ( .A(n_12), .Y(n_141) );
INVx1_ASAP7_75t_L g146 ( .A(n_12), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_13), .B(n_166), .Y(n_591) );
A2O1A1Ixp33_ASAP7_75t_L g239 ( .A1(n_14), .A2(n_156), .B(n_240), .C(n_242), .Y(n_239) );
AOI22xp33_ASAP7_75t_SL g906 ( .A1(n_15), .A2(n_907), .B1(n_908), .B2(n_909), .Y(n_906) );
INVx1_ASAP7_75t_L g909 ( .A(n_15), .Y(n_909) );
BUFx10_ASAP7_75t_L g896 ( .A(n_16), .Y(n_896) );
CKINVDCx5p33_ASAP7_75t_R g211 ( .A(n_17), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_18), .B(n_143), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_19), .B(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_20), .B(n_195), .Y(n_194) );
A2O1A1Ixp33_ASAP7_75t_L g224 ( .A1(n_21), .A2(n_225), .B(n_226), .C(n_228), .Y(n_224) );
CKINVDCx5p33_ASAP7_75t_R g578 ( .A(n_22), .Y(n_578) );
NAND3xp33_ASAP7_75t_L g648 ( .A(n_23), .B(n_139), .C(n_646), .Y(n_648) );
AND2x2_ASAP7_75t_L g208 ( .A(n_24), .B(n_133), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_25), .B(n_252), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_26), .B(n_166), .Y(n_185) );
AOI22xp33_ASAP7_75t_L g299 ( .A1(n_27), .A2(n_71), .B1(n_174), .B2(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g164 ( .A(n_28), .Y(n_164) );
INVx1_ASAP7_75t_L g255 ( .A(n_29), .Y(n_255) );
AOI22xp33_ASAP7_75t_L g99 ( .A1(n_30), .A2(n_100), .B1(n_112), .B2(n_921), .Y(n_99) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_31), .B(n_628), .Y(n_627) );
NAND2xp5_ASAP7_75t_SL g173 ( .A(n_32), .B(n_174), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_33), .B(n_166), .Y(n_274) );
INVx1_ASAP7_75t_L g107 ( .A(n_34), .Y(n_107) );
AND3x2_ASAP7_75t_L g920 ( .A(n_34), .B(n_891), .C(n_893), .Y(n_920) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_35), .B(n_193), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g614 ( .A(n_36), .B(n_156), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_37), .B(n_166), .Y(n_165) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_38), .B(n_217), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g533 ( .A(n_39), .B(n_214), .Y(n_533) );
AOI22xp5_ASAP7_75t_L g114 ( .A1(n_40), .A2(n_115), .B1(n_116), .B2(n_887), .Y(n_114) );
INVx1_ASAP7_75t_L g887 ( .A(n_40), .Y(n_887) );
CKINVDCx5p33_ASAP7_75t_R g241 ( .A(n_41), .Y(n_241) );
AND2x4_ASAP7_75t_L g163 ( .A(n_42), .B(n_164), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_43), .B(n_166), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_44), .B(n_133), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_45), .B(n_166), .Y(n_662) );
AOI22xp33_ASAP7_75t_L g297 ( .A1(n_46), .A2(n_83), .B1(n_174), .B2(n_176), .Y(n_297) );
INVx1_ASAP7_75t_L g232 ( .A(n_47), .Y(n_232) );
CKINVDCx5p33_ASAP7_75t_R g549 ( .A(n_48), .Y(n_549) );
A2O1A1Ixp33_ASAP7_75t_L g631 ( .A1(n_49), .A2(n_550), .B(n_632), .C(n_634), .Y(n_631) );
INVx1_ASAP7_75t_L g135 ( .A(n_50), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_51), .B(n_166), .Y(n_535) );
AND2x4_ASAP7_75t_L g104 ( .A(n_52), .B(n_105), .Y(n_104) );
INVx3_ASAP7_75t_L g576 ( .A(n_53), .Y(n_576) );
AOI22xp5_ASAP7_75t_L g897 ( .A1(n_54), .A2(n_898), .B1(n_915), .B2(n_917), .Y(n_897) );
HB1xp67_ASAP7_75t_L g109 ( .A(n_55), .Y(n_109) );
NOR2xp67_ASAP7_75t_L g892 ( .A(n_55), .B(n_73), .Y(n_892) );
AND2x2_ASAP7_75t_L g203 ( .A(n_56), .B(n_167), .Y(n_203) );
INVx1_ASAP7_75t_L g105 ( .A(n_57), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_58), .B(n_195), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g670 ( .A(n_59), .B(n_572), .Y(n_670) );
NAND2x1_ASAP7_75t_L g155 ( .A(n_60), .B(n_156), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_61), .B(n_271), .Y(n_270) );
INVx1_ASAP7_75t_L g587 ( .A(n_62), .Y(n_587) );
NAND2xp5_ASAP7_75t_SL g181 ( .A(n_63), .B(n_182), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_64), .B(n_153), .Y(n_248) );
NOR3xp33_ASAP7_75t_L g102 ( .A(n_65), .B(n_103), .C(n_106), .Y(n_102) );
INVx2_ASAP7_75t_L g894 ( .A(n_65), .Y(n_894) );
CKINVDCx5p33_ASAP7_75t_R g543 ( .A(n_66), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_67), .B(n_176), .Y(n_642) );
NAND2xp5_ASAP7_75t_SL g138 ( .A(n_68), .B(n_139), .Y(n_138) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_69), .B(n_139), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_70), .B(n_237), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g201 ( .A(n_72), .B(n_193), .Y(n_201) );
HB1xp67_ASAP7_75t_L g111 ( .A(n_73), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g151 ( .A(n_74), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_75), .B(n_618), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_76), .B(n_143), .Y(n_142) );
NAND2xp33_ASAP7_75t_SL g250 ( .A(n_77), .B(n_144), .Y(n_250) );
NAND2xp5_ASAP7_75t_SL g247 ( .A(n_78), .B(n_214), .Y(n_247) );
INVx1_ASAP7_75t_L g626 ( .A(n_79), .Y(n_626) );
CKINVDCx5p33_ASAP7_75t_R g551 ( .A(n_80), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_81), .B(n_153), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_82), .B(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g149 ( .A(n_84), .Y(n_149) );
INVx1_ASAP7_75t_L g160 ( .A(n_84), .Y(n_160) );
BUFx3_ASAP7_75t_L g179 ( .A(n_84), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_85), .B(n_200), .Y(n_199) );
CKINVDCx5p33_ASAP7_75t_R g227 ( .A(n_86), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_87), .B(n_176), .Y(n_528) );
INVx1_ASAP7_75t_L g574 ( .A(n_88), .Y(n_574) );
NAND2xp5_ASAP7_75t_SL g616 ( .A(n_89), .B(n_182), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_90), .B(n_167), .Y(n_619) );
NAND2xp33_ASAP7_75t_L g267 ( .A(n_91), .B(n_268), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_92), .B(n_669), .Y(n_668) );
CKINVDCx5p33_ASAP7_75t_R g569 ( .A(n_93), .Y(n_569) );
INVx1_ASAP7_75t_L g565 ( .A(n_94), .Y(n_565) );
CKINVDCx5p33_ASAP7_75t_R g545 ( .A(n_95), .Y(n_545) );
CKINVDCx5p33_ASAP7_75t_R g912 ( .A(n_96), .Y(n_912) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_97), .B(n_214), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_98), .B(n_572), .Y(n_665) );
BUFx6f_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
BUFx6f_ASAP7_75t_L g922 ( .A(n_101), .Y(n_922) );
AND2x4_ASAP7_75t_L g101 ( .A(n_102), .B(n_108), .Y(n_101) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_L g121 ( .A(n_106), .Y(n_121) );
BUFx2_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
NAND2xp5_ASAP7_75t_L g905 ( .A(n_107), .B(n_892), .Y(n_905) );
NOR2xp33_ASAP7_75t_L g108 ( .A(n_109), .B(n_110), .Y(n_108) );
INVx1_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
OR2x2_ASAP7_75t_L g112 ( .A(n_113), .B(n_911), .Y(n_112) );
OAI21xp5_ASAP7_75t_SL g113 ( .A1(n_114), .A2(n_888), .B(n_897), .Y(n_113) );
INVx1_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
HB1xp67_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
OAI22xp5_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_122), .B1(n_516), .B2(n_885), .Y(n_117) );
INVx2_ASAP7_75t_SL g118 ( .A(n_119), .Y(n_118) );
INVx11_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
BUFx8_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
BUFx6f_ASAP7_75t_SL g886 ( .A(n_121), .Y(n_886) );
INVx2_ASAP7_75t_L g908 ( .A(n_122), .Y(n_908) );
AND2x2_ASAP7_75t_L g122 ( .A(n_123), .B(n_455), .Y(n_122) );
NOR2xp33_ASAP7_75t_L g123 ( .A(n_124), .B(n_399), .Y(n_123) );
NAND4xp25_ASAP7_75t_L g124 ( .A(n_125), .B(n_315), .C(n_342), .D(n_367), .Y(n_124) );
AOI221x1_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_219), .B1(n_275), .B2(n_282), .C(n_303), .Y(n_125) );
AND2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_186), .Y(n_126) );
INVx1_ASAP7_75t_L g410 ( .A(n_127), .Y(n_410) );
INVx2_ASAP7_75t_SL g127 ( .A(n_128), .Y(n_127) );
INVx2_ASAP7_75t_L g308 ( .A(n_128), .Y(n_308) );
OR2x2_ASAP7_75t_L g489 ( .A(n_128), .B(n_490), .Y(n_489) );
OR2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_169), .Y(n_128) );
BUFx2_ASAP7_75t_L g324 ( .A(n_129), .Y(n_324) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx1_ASAP7_75t_L g279 ( .A(n_130), .Y(n_279) );
INVx1_ASAP7_75t_L g365 ( .A(n_130), .Y(n_365) );
OAI21x1_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_136), .B(n_165), .Y(n_130) );
OAI21x1_ASAP7_75t_L g170 ( .A1(n_131), .A2(n_171), .B(n_185), .Y(n_170) );
OAI21xp5_ASAP7_75t_L g339 ( .A1(n_131), .A2(n_171), .B(n_185), .Y(n_339) );
OAI21x1_ASAP7_75t_L g605 ( .A1(n_131), .A2(n_539), .B(n_606), .Y(n_605) );
OAI21x1_ASAP7_75t_L g610 ( .A1(n_131), .A2(n_611), .B(n_619), .Y(n_610) );
OAI21x1_ASAP7_75t_L g658 ( .A1(n_131), .A2(n_611), .B(n_619), .Y(n_658) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
NOR2x1_ASAP7_75t_SL g671 ( .A(n_132), .B(n_672), .Y(n_671) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
NOR2xp67_ASAP7_75t_SL g189 ( .A(n_133), .B(n_190), .Y(n_189) );
INVxp67_ASAP7_75t_SL g207 ( .A(n_133), .Y(n_207) );
INVx1_ASAP7_75t_L g690 ( .A(n_133), .Y(n_690) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g168 ( .A(n_134), .Y(n_168) );
INVxp33_ASAP7_75t_L g256 ( .A(n_134), .Y(n_256) );
BUFx2_ASAP7_75t_L g259 ( .A(n_134), .Y(n_259) );
INVx1_ASAP7_75t_L g234 ( .A(n_135), .Y(n_234) );
OAI21xp5_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_150), .B(n_161), .Y(n_136) );
AOI21xp5_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_142), .B(n_147), .Y(n_137) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx2_ASAP7_75t_L g174 ( .A(n_140), .Y(n_174) );
INVx2_ASAP7_75t_L g273 ( .A(n_140), .Y(n_273) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_141), .Y(n_154) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_141), .Y(n_177) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g214 ( .A(n_145), .Y(n_214) );
INVx2_ASAP7_75t_L g217 ( .A(n_145), .Y(n_217) );
INVx1_ASAP7_75t_L g268 ( .A(n_145), .Y(n_268) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g158 ( .A(n_146), .Y(n_158) );
AOI21xp5_ASAP7_75t_L g180 ( .A1(n_147), .A2(n_181), .B(n_183), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_147), .A2(n_216), .B(n_218), .Y(n_215) );
AO21x1_ASAP7_75t_L g246 ( .A1(n_147), .A2(n_247), .B(n_248), .Y(n_246) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_147), .A2(n_527), .B(n_528), .Y(n_526) );
AOI21xp5_ASAP7_75t_L g588 ( .A1(n_147), .A2(n_589), .B(n_590), .Y(n_588) );
AOI21xp5_ASAP7_75t_L g615 ( .A1(n_147), .A2(n_616), .B(n_617), .Y(n_615) );
BUFx10_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g646 ( .A(n_148), .Y(n_646) );
INVx1_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
BUFx3_ASAP7_75t_L g546 ( .A(n_149), .Y(n_546) );
O2A1O1Ixp5_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_152), .B(n_155), .C(n_159), .Y(n_150) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g200 ( .A(n_154), .Y(n_200) );
INVx2_ASAP7_75t_L g266 ( .A(n_154), .Y(n_266) );
INVx2_ASAP7_75t_L g300 ( .A(n_154), .Y(n_300) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx2_ASAP7_75t_L g182 ( .A(n_157), .Y(n_182) );
INVx2_ASAP7_75t_L g212 ( .A(n_157), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_157), .B(n_227), .Y(n_226) );
HB1xp67_ASAP7_75t_L g628 ( .A(n_157), .Y(n_628) );
INVx3_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
BUFx6f_ASAP7_75t_L g193 ( .A(n_158), .Y(n_193) );
INVx2_ASAP7_75t_L g196 ( .A(n_159), .Y(n_196) );
NAND3xp33_ASAP7_75t_L g298 ( .A(n_159), .B(n_291), .C(n_295), .Y(n_298) );
AOI21xp5_ASAP7_75t_L g612 ( .A1(n_159), .A2(n_613), .B(n_614), .Y(n_612) );
BUFx3_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx2_ASAP7_75t_L g243 ( .A(n_160), .Y(n_243) );
INVx1_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx2_ASAP7_75t_SL g235 ( .A(n_162), .Y(n_235) );
INVx1_ASAP7_75t_L g534 ( .A(n_162), .Y(n_534) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
BUFx6f_ASAP7_75t_SL g184 ( .A(n_163), .Y(n_184) );
INVx1_ASAP7_75t_L g190 ( .A(n_163), .Y(n_190) );
INVx1_ASAP7_75t_L g292 ( .A(n_163), .Y(n_292) );
INVx3_ASAP7_75t_L g567 ( .A(n_163), .Y(n_567) );
HB1xp67_ASAP7_75t_L g639 ( .A(n_166), .Y(n_639) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
AND2x2_ASAP7_75t_L g281 ( .A(n_169), .B(n_187), .Y(n_281) );
INVx1_ASAP7_75t_L g398 ( .A(n_169), .Y(n_398) );
AND2x2_ASAP7_75t_L g429 ( .A(n_169), .B(n_365), .Y(n_429) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
OR2x2_ASAP7_75t_L g331 ( .A(n_170), .B(n_187), .Y(n_331) );
OAI21x1_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_180), .B(n_184), .Y(n_171) );
AOI21xp5_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_175), .B(n_178), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_174), .B(n_586), .Y(n_585) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx2_ASAP7_75t_L g195 ( .A(n_177), .Y(n_195) );
INVx2_ASAP7_75t_L g252 ( .A(n_177), .Y(n_252) );
INVx2_ASAP7_75t_L g271 ( .A(n_177), .Y(n_271) );
INVx2_ASAP7_75t_L g532 ( .A(n_177), .Y(n_532) );
INVx3_ASAP7_75t_L g542 ( .A(n_177), .Y(n_542) );
INVx3_ASAP7_75t_L g625 ( .A(n_177), .Y(n_625) );
AO21x1_ASAP7_75t_L g249 ( .A1(n_178), .A2(n_250), .B(n_251), .Y(n_249) );
O2A1O1Ixp5_ASAP7_75t_L g529 ( .A1(n_178), .A2(n_530), .B(n_531), .C(n_533), .Y(n_529) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVx1_ASAP7_75t_L g202 ( .A(n_179), .Y(n_202) );
AOI211x1_ASAP7_75t_L g209 ( .A1(n_179), .A2(n_208), .B(n_210), .C(n_215), .Y(n_209) );
INVx2_ASAP7_75t_L g229 ( .A(n_179), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_179), .B(n_567), .Y(n_566) );
NOR3xp33_ASAP7_75t_L g573 ( .A(n_179), .B(n_567), .C(n_574), .Y(n_573) );
INVx2_ASAP7_75t_L g544 ( .A(n_182), .Y(n_544) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_184), .A2(n_207), .B(n_208), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_184), .A2(n_254), .B(n_258), .Y(n_257) );
OAI21x1_ASAP7_75t_L g263 ( .A1(n_184), .A2(n_264), .B(n_269), .Y(n_263) );
OAI21x1_ASAP7_75t_L g581 ( .A1(n_184), .A2(n_582), .B(n_588), .Y(n_581) );
OAI21x1_ASAP7_75t_L g611 ( .A1(n_184), .A2(n_612), .B(n_615), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_186), .B(n_446), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_186), .B(n_429), .Y(n_454) );
AND2x4_ASAP7_75t_L g186 ( .A(n_187), .B(n_204), .Y(n_186) );
INVx2_ASAP7_75t_L g338 ( .A(n_187), .Y(n_338) );
INVx1_ASAP7_75t_L g382 ( .A(n_187), .Y(n_382) );
AND2x4_ASAP7_75t_L g187 ( .A(n_188), .B(n_197), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_189), .B(n_191), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g197 ( .A1(n_189), .A2(n_198), .B(n_203), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g191 ( .A1(n_192), .A2(n_194), .B(n_196), .Y(n_191) );
INVx1_ASAP7_75t_L g225 ( .A(n_193), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_193), .B(n_241), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g564 ( .A(n_193), .B(n_565), .Y(n_564) );
INVx2_ASAP7_75t_L g618 ( .A(n_193), .Y(n_618) );
INVxp67_ASAP7_75t_L g548 ( .A(n_195), .Y(n_548) );
INVxp67_ASAP7_75t_L g583 ( .A(n_195), .Y(n_583) );
AOI21xp5_ASAP7_75t_L g667 ( .A1(n_196), .A2(n_668), .B(n_670), .Y(n_667) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_199), .A2(n_201), .B(n_202), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g632 ( .A(n_200), .B(n_633), .Y(n_632) );
AOI21xp5_ASAP7_75t_L g264 ( .A1(n_202), .A2(n_265), .B(n_267), .Y(n_264) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
INVx2_ASAP7_75t_L g307 ( .A(n_205), .Y(n_307) );
INVx1_ASAP7_75t_L g312 ( .A(n_205), .Y(n_312) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_205), .Y(n_323) );
BUFx2_ASAP7_75t_L g335 ( .A(n_205), .Y(n_335) );
AND2x2_ASAP7_75t_L g366 ( .A(n_205), .B(n_338), .Y(n_366) );
INVx2_ASAP7_75t_L g460 ( .A(n_205), .Y(n_460) );
AND2x2_ASAP7_75t_L g476 ( .A(n_205), .B(n_339), .Y(n_476) );
OR2x6_ASAP7_75t_L g205 ( .A(n_206), .B(n_209), .Y(n_205) );
OAI21xp5_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_212), .B(n_213), .Y(n_210) );
INVx2_ASAP7_75t_L g550 ( .A(n_217), .Y(n_550) );
AND2x2_ASAP7_75t_L g219 ( .A(n_220), .B(n_244), .Y(n_219) );
OR2x2_ASAP7_75t_L g378 ( .A(n_220), .B(n_341), .Y(n_378) );
NAND2x1p5_ASAP7_75t_L g439 ( .A(n_220), .B(n_440), .Y(n_439) );
INVx2_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVx1_ASAP7_75t_L g328 ( .A(n_222), .Y(n_328) );
AND2x2_ASAP7_75t_L g359 ( .A(n_222), .B(n_360), .Y(n_359) );
BUFx2_ASAP7_75t_L g386 ( .A(n_222), .Y(n_386) );
AND2x2_ASAP7_75t_L g434 ( .A(n_222), .B(n_307), .Y(n_434) );
HB1xp67_ASAP7_75t_L g470 ( .A(n_222), .Y(n_470) );
NAND2x1p5_ASAP7_75t_L g222 ( .A(n_223), .B(n_238), .Y(n_222) );
NAND2x1p5_ASAP7_75t_L g302 ( .A(n_223), .B(n_238), .Y(n_302) );
OA21x2_ASAP7_75t_L g223 ( .A1(n_224), .A2(n_230), .B(n_236), .Y(n_223) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_225), .A2(n_572), .B1(n_573), .B2(n_575), .Y(n_571) );
AOI21xp5_ASAP7_75t_L g269 ( .A1(n_228), .A2(n_270), .B(n_272), .Y(n_269) );
INVx1_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g586 ( .A(n_229), .B(n_587), .Y(n_586) );
OR2x2_ASAP7_75t_L g238 ( .A(n_230), .B(n_239), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_231), .B(n_235), .Y(n_230) );
INVx2_ASAP7_75t_L g237 ( .A(n_231), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g287 ( .A(n_231), .B(n_288), .Y(n_287) );
AO21x2_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_233), .B(n_234), .Y(n_231) );
AOI21x1_ASAP7_75t_L g296 ( .A1(n_232), .A2(n_233), .B(n_234), .Y(n_296) );
INVx1_ASAP7_75t_L g672 ( .A(n_235), .Y(n_672) );
INVxp67_ASAP7_75t_L g553 ( .A(n_237), .Y(n_553) );
OAI21xp33_ASAP7_75t_L g635 ( .A1(n_237), .A2(n_292), .B(n_630), .Y(n_635) );
INVx1_ASAP7_75t_L g552 ( .A(n_242), .Y(n_552) );
AOI21xp5_ASAP7_75t_L g664 ( .A1(n_242), .A2(n_665), .B(n_666), .Y(n_664) );
INVx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
INVx2_ASAP7_75t_L g294 ( .A(n_243), .Y(n_294) );
INVx3_ASAP7_75t_L g341 ( .A(n_244), .Y(n_341) );
AND2x2_ASAP7_75t_L g421 ( .A(n_244), .B(n_373), .Y(n_421) );
AND2x2_ASAP7_75t_L g511 ( .A(n_244), .B(n_385), .Y(n_511) );
AND2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_260), .Y(n_244) );
OR2x2_ASAP7_75t_L g301 ( .A(n_245), .B(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g314 ( .A(n_245), .B(n_261), .Y(n_314) );
AND2x2_ASAP7_75t_L g327 ( .A(n_245), .B(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g350 ( .A(n_245), .B(n_302), .Y(n_350) );
INVx2_ASAP7_75t_L g360 ( .A(n_245), .Y(n_360) );
INVx1_ASAP7_75t_L g407 ( .A(n_245), .Y(n_407) );
AO31x2_ASAP7_75t_L g245 ( .A1(n_246), .A2(n_249), .A3(n_253), .B(n_257), .Y(n_245) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
BUFx3_ASAP7_75t_L g262 ( .A(n_259), .Y(n_262) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVx1_ASAP7_75t_L g362 ( .A(n_261), .Y(n_362) );
AND2x2_ASAP7_75t_L g387 ( .A(n_261), .B(n_286), .Y(n_387) );
INVx1_ASAP7_75t_L g414 ( .A(n_261), .Y(n_414) );
AND2x2_ASAP7_75t_L g467 ( .A(n_261), .B(n_442), .Y(n_467) );
OAI21x1_ASAP7_75t_L g261 ( .A1(n_262), .A2(n_263), .B(n_274), .Y(n_261) );
OAI21x1_ASAP7_75t_L g524 ( .A1(n_262), .A2(n_525), .B(n_535), .Y(n_524) );
OAI21x1_ASAP7_75t_L g580 ( .A1(n_262), .A2(n_581), .B(n_591), .Y(n_580) );
NOR2xp33_ASAP7_75t_L g568 ( .A(n_266), .B(n_569), .Y(n_568) );
INVx2_ASAP7_75t_L g572 ( .A(n_266), .Y(n_572) );
INVx1_ASAP7_75t_L g669 ( .A(n_268), .Y(n_669) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
OR2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_280), .Y(n_276) );
HB1xp67_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g311 ( .A(n_278), .B(n_312), .Y(n_311) );
OR2x2_ASAP7_75t_L g332 ( .A(n_278), .B(n_312), .Y(n_332) );
INVx2_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g355 ( .A(n_279), .Y(n_355) );
OR2x2_ASAP7_75t_L g423 ( .A(n_280), .B(n_371), .Y(n_423) );
INVx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g310 ( .A(n_281), .B(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g506 ( .A(n_281), .B(n_306), .Y(n_506) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
OR2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_301), .Y(n_283) );
OR2x2_ASAP7_75t_L g340 ( .A(n_284), .B(n_341), .Y(n_340) );
OR2x2_ASAP7_75t_L g499 ( .A(n_284), .B(n_341), .Y(n_499) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
HB1xp67_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g318 ( .A(n_286), .Y(n_318) );
INVxp67_ASAP7_75t_L g349 ( .A(n_286), .Y(n_349) );
AND2x2_ASAP7_75t_L g361 ( .A(n_286), .B(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g373 ( .A(n_286), .Y(n_373) );
AND2x2_ASAP7_75t_L g395 ( .A(n_286), .B(n_302), .Y(n_395) );
INVx1_ASAP7_75t_L g442 ( .A(n_286), .Y(n_442) );
OR2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_289), .Y(n_286) );
OAI22xp5_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_297), .B1(n_298), .B2(n_299), .Y(n_289) );
NAND3xp33_ASAP7_75t_L g290 ( .A(n_291), .B(n_293), .C(n_295), .Y(n_290) );
BUFx2_ASAP7_75t_L g554 ( .A(n_291), .Y(n_554) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
NOR2xp33_ASAP7_75t_L g570 ( .A(n_294), .B(n_567), .Y(n_570) );
NOR3xp33_ASAP7_75t_L g575 ( .A(n_294), .B(n_567), .C(n_576), .Y(n_575) );
HB1xp67_ASAP7_75t_L g561 ( .A(n_295), .Y(n_561) );
NOR2xp33_ASAP7_75t_SL g577 ( .A(n_295), .B(n_578), .Y(n_577) );
INVx2_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
OR2x2_ASAP7_75t_L g322 ( .A(n_301), .B(n_323), .Y(n_322) );
INVx2_ASAP7_75t_L g374 ( .A(n_301), .Y(n_374) );
NOR2xp33_ASAP7_75t_L g419 ( .A(n_301), .B(n_420), .Y(n_419) );
OR2x2_ASAP7_75t_L g492 ( .A(n_301), .B(n_493), .Y(n_492) );
AND2x2_ASAP7_75t_L g357 ( .A(n_302), .B(n_318), .Y(n_357) );
INVx2_ASAP7_75t_L g488 ( .A(n_302), .Y(n_488) );
AOI21xp33_ASAP7_75t_L g303 ( .A1(n_304), .A2(n_309), .B(n_313), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_305), .B(n_308), .Y(n_304) );
NAND3xp33_ASAP7_75t_L g495 ( .A(n_305), .B(n_369), .C(n_370), .Y(n_495) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_306), .B(n_397), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_306), .B(n_353), .Y(n_462) );
BUFx3_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
OR2x2_ASAP7_75t_L g490 ( .A(n_307), .B(n_338), .Y(n_490) );
AND2x4_ASAP7_75t_SL g380 ( .A(n_308), .B(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g432 ( .A(n_308), .Y(n_432) );
OAI22xp5_ASAP7_75t_L g409 ( .A1(n_309), .A2(n_410), .B1(n_411), .B2(n_415), .Y(n_409) );
INVx2_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g356 ( .A(n_314), .B(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g394 ( .A(n_314), .B(n_395), .Y(n_394) );
AOI21xp5_ASAP7_75t_L g315 ( .A1(n_316), .A2(n_319), .B(n_325), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_316), .B(n_327), .Y(n_326) );
INVx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_321), .B(n_324), .Y(n_320) );
INVx2_ASAP7_75t_SL g321 ( .A(n_322), .Y(n_321) );
OAI32xp33_ASAP7_75t_L g424 ( .A1(n_322), .A2(n_359), .A3(n_425), .B1(n_426), .B2(n_427), .Y(n_424) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_324), .B(n_491), .Y(n_513) );
OAI22xp33_ASAP7_75t_L g325 ( .A1(n_326), .A2(n_329), .B1(n_333), .B2(n_340), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_327), .B(n_428), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_327), .B(n_467), .Y(n_501) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
NOR2x1_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
INVx4_ASAP7_75t_L g369 ( .A(n_331), .Y(n_369) );
HB1xp67_ASAP7_75t_L g408 ( .A(n_331), .Y(n_408) );
OR2x2_ASAP7_75t_L g448 ( .A(n_331), .B(n_364), .Y(n_448) );
INVx1_ASAP7_75t_L g346 ( .A(n_332), .Y(n_346) );
OR2x2_ASAP7_75t_L g425 ( .A(n_332), .B(n_381), .Y(n_425) );
OR2x2_ASAP7_75t_L g333 ( .A(n_334), .B(n_336), .Y(n_333) );
AND2x2_ASAP7_75t_L g453 ( .A(n_334), .B(n_337), .Y(n_453) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_335), .B(n_353), .Y(n_418) );
INVx1_ASAP7_75t_L g437 ( .A(n_335), .Y(n_437) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
HB1xp67_ASAP7_75t_L g345 ( .A(n_337), .Y(n_345) );
AND2x2_ASAP7_75t_L g377 ( .A(n_337), .B(n_364), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_337), .B(n_437), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_337), .B(n_371), .Y(n_473) );
AND2x2_ASAP7_75t_L g337 ( .A(n_338), .B(n_339), .Y(n_337) );
AND2x4_ASAP7_75t_SL g459 ( .A(n_338), .B(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g354 ( .A(n_339), .Y(n_354) );
AOI222xp33_ASAP7_75t_L g342 ( .A1(n_343), .A2(n_347), .B1(n_351), .B2(n_356), .C1(n_358), .C2(n_363), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_345), .B(n_346), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_346), .B(n_403), .Y(n_402) );
NOR4xp25_ASAP7_75t_L g505 ( .A(n_346), .B(n_429), .C(n_506), .D(n_507), .Y(n_505) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_349), .B(n_350), .Y(n_348) );
INVx2_ASAP7_75t_L g515 ( .A(n_350), .Y(n_515) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_354), .B(n_355), .Y(n_353) );
INVx1_ASAP7_75t_L g446 ( .A(n_354), .Y(n_446) );
INVx2_ASAP7_75t_L g371 ( .A(n_355), .Y(n_371) );
INVx2_ASAP7_75t_L g415 ( .A(n_357), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g457 ( .A1(n_358), .A2(n_458), .B1(n_461), .B2(n_463), .Y(n_457) );
AND2x4_ASAP7_75t_SL g358 ( .A(n_359), .B(n_361), .Y(n_358) );
AND2x2_ASAP7_75t_L g463 ( .A(n_359), .B(n_387), .Y(n_463) );
INVx1_ASAP7_75t_L g466 ( .A(n_359), .Y(n_466) );
AND2x2_ASAP7_75t_L g441 ( .A(n_360), .B(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g478 ( .A(n_360), .Y(n_478) );
INVx1_ASAP7_75t_L g426 ( .A(n_361), .Y(n_426) );
AND2x2_ASAP7_75t_L g469 ( .A(n_361), .B(n_470), .Y(n_469) );
AND2x2_ASAP7_75t_L g487 ( .A(n_362), .B(n_488), .Y(n_487) );
AND2x2_ASAP7_75t_L g363 ( .A(n_364), .B(n_366), .Y(n_363) );
HB1xp67_ASAP7_75t_L g503 ( .A(n_364), .Y(n_503) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
AND2x2_ASAP7_75t_L g397 ( .A(n_365), .B(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g508 ( .A(n_366), .Y(n_508) );
AOI211xp5_ASAP7_75t_L g367 ( .A1(n_368), .A2(n_372), .B(n_375), .C(n_388), .Y(n_367) );
NOR2x1_ASAP7_75t_L g481 ( .A(n_368), .B(n_482), .Y(n_481) );
AOI322xp5_ASAP7_75t_L g497 ( .A1(n_368), .A2(n_369), .A3(n_434), .B1(n_498), .B2(n_500), .C1(n_502), .C2(n_924), .Y(n_497) );
AND2x4_ASAP7_75t_L g368 ( .A(n_369), .B(n_370), .Y(n_368) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g458 ( .A(n_371), .B(n_459), .Y(n_458) );
OR2x2_ASAP7_75t_L g483 ( .A(n_371), .B(n_484), .Y(n_483) );
AND2x2_ASAP7_75t_L g372 ( .A(n_373), .B(n_374), .Y(n_372) );
HB1xp67_ASAP7_75t_L g391 ( .A(n_373), .Y(n_391) );
INVx2_ASAP7_75t_L g510 ( .A(n_373), .Y(n_510) );
INVx1_ASAP7_75t_L g451 ( .A(n_374), .Y(n_451) );
OAI22xp5_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_378), .B1(n_379), .B2(n_383), .Y(n_375) );
OAI22xp33_ASAP7_75t_L g474 ( .A1(n_376), .A2(n_393), .B1(n_475), .B2(n_477), .Y(n_474) );
INVx2_ASAP7_75t_SL g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g491 ( .A(n_381), .Y(n_491) );
INVx4_ASAP7_75t_R g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_385), .B(n_387), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g392 ( .A(n_386), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_387), .B(n_405), .Y(n_404) );
INVx2_ASAP7_75t_L g493 ( .A(n_387), .Y(n_493) );
AOI21xp5_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_393), .B(n_396), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
AND2x4_ASAP7_75t_L g390 ( .A(n_391), .B(n_392), .Y(n_390) );
INVx2_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
NAND4xp25_ASAP7_75t_L g399 ( .A(n_400), .B(n_416), .C(n_430), .D(n_443), .Y(n_399) );
AOI21xp5_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_408), .B(n_409), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_407), .B(n_413), .Y(n_412) );
INVx2_ASAP7_75t_L g449 ( .A(n_411), .Y(n_449) );
OR2x2_ASAP7_75t_L g411 ( .A(n_412), .B(n_415), .Y(n_411) );
INVxp67_ASAP7_75t_SL g413 ( .A(n_414), .Y(n_413) );
BUFx3_ASAP7_75t_L g420 ( .A(n_414), .Y(n_420) );
AOI221xp5_ASAP7_75t_L g416 ( .A1(n_417), .A2(n_419), .B1(n_421), .B2(n_422), .C(n_424), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx2_ASAP7_75t_L g428 ( .A(n_420), .Y(n_428) );
AND2x2_ASAP7_75t_L g440 ( .A(n_420), .B(n_441), .Y(n_440) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_420), .B(n_515), .Y(n_514) );
AND2x2_ASAP7_75t_L g433 ( .A(n_421), .B(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
O2A1O1Ixp33_ASAP7_75t_L g450 ( .A1(n_426), .A2(n_451), .B(n_452), .C(n_454), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_428), .B(n_429), .Y(n_427) );
AOI22xp5_ASAP7_75t_L g430 ( .A1(n_431), .A2(n_433), .B1(n_435), .B2(n_438), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g496 ( .A(n_441), .Y(n_496) );
O2A1O1Ixp33_ASAP7_75t_L g443 ( .A1(n_444), .A2(n_447), .B(n_449), .C(n_450), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
AOI22xp5_ASAP7_75t_L g512 ( .A1(n_449), .A2(n_458), .B1(n_513), .B2(n_514), .Y(n_512) );
INVxp67_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
NOR3xp33_ASAP7_75t_L g455 ( .A(n_456), .B(n_494), .C(n_504), .Y(n_455) );
NAND3xp33_ASAP7_75t_SL g456 ( .A(n_457), .B(n_464), .C(n_479), .Y(n_456) );
INVx1_ASAP7_75t_L g484 ( .A(n_459), .Y(n_484) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
AOI21xp5_ASAP7_75t_L g479 ( .A1(n_463), .A2(n_480), .B(n_485), .Y(n_479) );
AOI21xp5_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_472), .B(n_474), .Y(n_464) );
OAI211xp5_ASAP7_75t_L g465 ( .A1(n_466), .A2(n_467), .B(n_468), .C(n_471), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_467), .B(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx2_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
OAI22xp5_ASAP7_75t_L g485 ( .A1(n_486), .A2(n_489), .B1(n_491), .B2(n_492), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
OAI21xp33_ASAP7_75t_SL g494 ( .A1(n_495), .A2(n_496), .B(n_497), .Y(n_494) );
INVx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
OAI21xp33_ASAP7_75t_L g504 ( .A1(n_505), .A2(n_509), .B(n_512), .Y(n_504) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_510), .B(n_511), .Y(n_509) );
AND2x4_ASAP7_75t_L g516 ( .A(n_517), .B(n_783), .Y(n_516) );
NOR3xp33_ASAP7_75t_L g517 ( .A(n_518), .B(n_705), .C(n_756), .Y(n_517) );
OAI221xp5_ASAP7_75t_SL g518 ( .A1(n_519), .A2(n_607), .B1(n_650), .B2(n_655), .C(n_674), .Y(n_518) );
AOI211xp5_ASAP7_75t_L g519 ( .A1(n_520), .A2(n_556), .B(n_592), .C(n_600), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
AND2x4_ASAP7_75t_L g880 ( .A(n_521), .B(n_596), .Y(n_880) );
AND2x2_ASAP7_75t_L g521 ( .A(n_522), .B(n_536), .Y(n_521) );
INVx1_ASAP7_75t_L g594 ( .A(n_522), .Y(n_594) );
AND2x2_ASAP7_75t_L g735 ( .A(n_522), .B(n_681), .Y(n_735) );
HB1xp67_ASAP7_75t_L g780 ( .A(n_522), .Y(n_780) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx2_ASAP7_75t_L g603 ( .A(n_523), .Y(n_603) );
INVx3_ASAP7_75t_L g683 ( .A(n_523), .Y(n_683) );
AND2x2_ASAP7_75t_L g711 ( .A(n_523), .B(n_605), .Y(n_711) );
AND2x2_ASAP7_75t_L g718 ( .A(n_523), .B(n_719), .Y(n_718) );
INVx3_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
OAI21xp5_ASAP7_75t_L g525 ( .A1(n_526), .A2(n_529), .B(n_534), .Y(n_525) );
INVx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
OAI21x1_ASAP7_75t_L g640 ( .A1(n_534), .A2(n_641), .B(n_644), .Y(n_640) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
OR2x2_ASAP7_75t_L g692 ( .A(n_537), .B(n_654), .Y(n_692) );
AO31x2_ASAP7_75t_L g537 ( .A1(n_538), .A2(n_553), .A3(n_554), .B(n_555), .Y(n_537) );
AO31x2_ASAP7_75t_L g703 ( .A1(n_538), .A2(n_553), .A3(n_554), .B(n_555), .Y(n_703) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
AOI22x1_ASAP7_75t_L g539 ( .A1(n_540), .A2(n_546), .B1(n_547), .B2(n_552), .Y(n_539) );
OAI22x1_ASAP7_75t_L g540 ( .A1(n_541), .A2(n_543), .B1(n_544), .B2(n_545), .Y(n_540) );
INVxp67_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx1_ASAP7_75t_L g634 ( .A(n_546), .Y(n_634) );
AOI21x1_ASAP7_75t_L g641 ( .A1(n_546), .A2(n_642), .B(n_643), .Y(n_641) );
OAI22xp5_ASAP7_75t_L g547 ( .A1(n_548), .A2(n_549), .B1(n_550), .B2(n_551), .Y(n_547) );
AOI21x1_ASAP7_75t_SL g623 ( .A1(n_552), .A2(n_624), .B(n_627), .Y(n_623) );
INVx1_ASAP7_75t_L g606 ( .A(n_555), .Y(n_606) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
AOI322xp5_ASAP7_75t_L g706 ( .A1(n_557), .A2(n_707), .A3(n_711), .B1(n_712), .B2(n_715), .C1(n_722), .C2(n_730), .Y(n_706) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
HB1xp67_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g730 ( .A(n_559), .B(n_682), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_559), .B(n_682), .Y(n_745) );
AND2x2_ASAP7_75t_L g798 ( .A(n_559), .B(n_711), .Y(n_798) );
AND2x2_ASAP7_75t_L g559 ( .A(n_560), .B(n_579), .Y(n_559) );
INVx3_ASAP7_75t_L g598 ( .A(n_560), .Y(n_598) );
AO21x2_ASAP7_75t_L g560 ( .A1(n_561), .A2(n_562), .B(n_577), .Y(n_560) );
AO21x1_ASAP7_75t_L g720 ( .A1(n_561), .A2(n_562), .B(n_577), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_563), .B(n_571), .Y(n_562) );
AOI22xp5_ASAP7_75t_L g563 ( .A1(n_564), .A2(n_566), .B1(n_568), .B2(n_570), .Y(n_563) );
INVx1_ASAP7_75t_L g599 ( .A(n_579), .Y(n_599) );
AND2x2_ASAP7_75t_L g604 ( .A(n_579), .B(n_605), .Y(n_604) );
INVx3_ASAP7_75t_L g654 ( .A(n_579), .Y(n_654) );
HB1xp67_ASAP7_75t_L g740 ( .A(n_579), .Y(n_740) );
INVx2_ASAP7_75t_L g753 ( .A(n_579), .Y(n_753) );
AND2x2_ASAP7_75t_L g763 ( .A(n_579), .B(n_598), .Y(n_763) );
INVx1_ASAP7_75t_L g824 ( .A(n_579), .Y(n_824) );
BUFx6f_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
OAI21xp5_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_584), .B(n_585), .Y(n_582) );
NOR2xp67_ASAP7_75t_L g592 ( .A(n_593), .B(n_595), .Y(n_592) );
HB1xp67_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx2_ASAP7_75t_L g841 ( .A(n_594), .Y(n_841) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
OR2x2_ASAP7_75t_L g867 ( .A(n_597), .B(n_702), .Y(n_867) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_598), .B(n_599), .Y(n_597) );
INVx1_ASAP7_75t_L g681 ( .A(n_598), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_598), .B(n_683), .Y(n_704) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_SL g601 ( .A(n_602), .B(n_604), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g813 ( .A(n_602), .B(n_789), .Y(n_813) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
NOR2xp67_ASAP7_75t_L g652 ( .A(n_603), .B(n_653), .Y(n_652) );
AND2x4_ASAP7_75t_L g772 ( .A(n_604), .B(n_773), .Y(n_772) );
AND2x4_ASAP7_75t_L g682 ( .A(n_605), .B(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g791 ( .A(n_605), .Y(n_791) );
OR2x2_ASAP7_75t_L g607 ( .A(n_608), .B(n_620), .Y(n_607) );
AND2x2_ASAP7_75t_L g697 ( .A(n_608), .B(n_660), .Y(n_697) );
OR2x2_ASAP7_75t_L g864 ( .A(n_608), .B(n_695), .Y(n_864) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g677 ( .A(n_609), .B(n_678), .Y(n_677) );
BUFx3_ASAP7_75t_L g709 ( .A(n_609), .Y(n_709) );
AND2x2_ASAP7_75t_L g836 ( .A(n_609), .B(n_621), .Y(n_836) );
AND2x4_ASAP7_75t_L g852 ( .A(n_609), .B(n_749), .Y(n_852) );
INVx2_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
HB1xp67_ASAP7_75t_L g796 ( .A(n_610), .Y(n_796) );
INVxp67_ASAP7_75t_L g647 ( .A(n_618), .Y(n_647) );
OR2x2_ASAP7_75t_L g713 ( .A(n_620), .B(n_714), .Y(n_713) );
INVx2_ASAP7_75t_L g760 ( .A(n_620), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_621), .B(n_636), .Y(n_620) );
AND2x4_ASAP7_75t_L g657 ( .A(n_621), .B(n_658), .Y(n_657) );
HB1xp67_ASAP7_75t_L g699 ( .A(n_621), .Y(n_699) );
INVx1_ASAP7_75t_L g725 ( .A(n_621), .Y(n_725) );
AND2x2_ASAP7_75t_L g768 ( .A(n_621), .B(n_688), .Y(n_768) );
INVx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx2_ASAP7_75t_L g687 ( .A(n_622), .Y(n_687) );
OAI21x1_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_629), .B(n_635), .Y(n_622) );
OR2x2_ASAP7_75t_L g624 ( .A(n_625), .B(n_626), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_630), .B(n_631), .Y(n_629) );
AND2x4_ASAP7_75t_L g729 ( .A(n_636), .B(n_660), .Y(n_729) );
INVx1_ASAP7_75t_L g743 ( .A(n_636), .Y(n_743) );
INVx2_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVxp67_ASAP7_75t_SL g673 ( .A(n_637), .Y(n_673) );
INVx2_ASAP7_75t_L g696 ( .A(n_637), .Y(n_696) );
INVx2_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
OAI21x1_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_640), .B(n_649), .Y(n_638) );
OA21x2_ASAP7_75t_L g688 ( .A1(n_640), .A2(n_649), .B(n_689), .Y(n_688) );
OAI21xp5_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_647), .B(n_648), .Y(n_644) );
INVxp67_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
HB1xp67_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
OR2x2_ASAP7_75t_L g810 ( .A(n_653), .B(n_811), .Y(n_810) );
BUFx2_ASAP7_75t_L g831 ( .A(n_653), .Y(n_831) );
INVx2_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g834 ( .A(n_654), .B(n_820), .Y(n_834) );
OR2x2_ASAP7_75t_L g655 ( .A(n_656), .B(n_659), .Y(n_655) );
INVx2_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
AND2x2_ASAP7_75t_L g741 ( .A(n_657), .B(n_742), .Y(n_741) );
AND2x2_ASAP7_75t_L g804 ( .A(n_657), .B(n_805), .Y(n_804) );
AND2x2_ASAP7_75t_L g829 ( .A(n_657), .B(n_830), .Y(n_829) );
INVx1_ASAP7_75t_L g873 ( .A(n_657), .Y(n_873) );
AND2x2_ASAP7_75t_L g726 ( .A(n_658), .B(n_696), .Y(n_726) );
AND2x4_ASAP7_75t_L g728 ( .A(n_658), .B(n_729), .Y(n_728) );
OR2x2_ASAP7_75t_L g733 ( .A(n_658), .B(n_686), .Y(n_733) );
AND2x4_ASAP7_75t_L g748 ( .A(n_658), .B(n_749), .Y(n_748) );
OR2x2_ASAP7_75t_L g659 ( .A(n_660), .B(n_673), .Y(n_659) );
INVx2_ASAP7_75t_L g678 ( .A(n_660), .Y(n_678) );
INVx2_ASAP7_75t_L g700 ( .A(n_660), .Y(n_700) );
BUFx2_ASAP7_75t_L g714 ( .A(n_660), .Y(n_714) );
INVx1_ASAP7_75t_L g770 ( .A(n_660), .Y(n_770) );
AND2x2_ASAP7_75t_L g830 ( .A(n_660), .B(n_688), .Y(n_830) );
BUFx6f_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
NAND2x1_ASAP7_75t_L g661 ( .A(n_662), .B(n_663), .Y(n_661) );
OAI21x1_ASAP7_75t_SL g663 ( .A1(n_664), .A2(n_667), .B(n_671), .Y(n_663) );
AND2x2_ASAP7_75t_L g710 ( .A(n_673), .B(n_678), .Y(n_710) );
AOI21xp5_ASAP7_75t_L g674 ( .A1(n_675), .A2(n_684), .B(n_691), .Y(n_674) );
INVxp67_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_677), .B(n_679), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_677), .B(n_760), .Y(n_759) );
INVx1_ASAP7_75t_L g853 ( .A(n_677), .Y(n_853) );
AND2x2_ASAP7_75t_L g865 ( .A(n_677), .B(n_685), .Y(n_865) );
BUFx2_ASAP7_75t_L g805 ( .A(n_678), .Y(n_805) );
INVx1_ASAP7_75t_L g879 ( .A(n_678), .Y(n_879) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_681), .B(n_682), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_682), .B(n_739), .Y(n_738) );
INVx2_ASAP7_75t_L g754 ( .A(n_682), .Y(n_754) );
INVx2_ASAP7_75t_SL g684 ( .A(n_685), .Y(n_684) );
AOI22xp33_ASAP7_75t_L g875 ( .A1(n_685), .A2(n_876), .B1(n_878), .B2(n_880), .Y(n_875) );
INVx2_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
OR2x2_ASAP7_75t_SL g686 ( .A(n_687), .B(n_688), .Y(n_686) );
OR2x6_ASAP7_75t_L g695 ( .A(n_687), .B(n_696), .Y(n_695) );
INVx2_ASAP7_75t_L g749 ( .A(n_687), .Y(n_749) );
INVx1_ASAP7_75t_SL g689 ( .A(n_690), .Y(n_689) );
OAI22xp5_ASAP7_75t_L g691 ( .A1(n_692), .A2(n_693), .B1(n_698), .B2(n_701), .Y(n_691) );
INVx2_ASAP7_75t_SL g736 ( .A(n_692), .Y(n_736) );
OR2x2_ASAP7_75t_L g765 ( .A(n_692), .B(n_704), .Y(n_765) );
INVx2_ASAP7_75t_L g802 ( .A(n_693), .Y(n_802) );
NAND2x1p5_ASAP7_75t_L g693 ( .A(n_694), .B(n_697), .Y(n_693) );
INVx2_ASAP7_75t_SL g694 ( .A(n_695), .Y(n_694) );
OR2x2_ASAP7_75t_L g850 ( .A(n_695), .B(n_700), .Y(n_850) );
OR2x2_ASAP7_75t_L g883 ( .A(n_695), .B(n_709), .Y(n_883) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_699), .B(n_700), .Y(n_698) );
AND2x2_ASAP7_75t_L g771 ( .A(n_699), .B(n_726), .Y(n_771) );
INVx1_ASAP7_75t_L g747 ( .A(n_700), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g787 ( .A(n_700), .B(n_724), .Y(n_787) );
OR2x2_ASAP7_75t_L g823 ( .A(n_700), .B(n_824), .Y(n_823) );
OR2x2_ASAP7_75t_L g701 ( .A(n_702), .B(n_704), .Y(n_701) );
INVx1_ASAP7_75t_L g820 ( .A(n_702), .Y(n_820) );
BUFx3_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx2_ASAP7_75t_L g721 ( .A(n_703), .Y(n_721) );
INVx1_ASAP7_75t_L g773 ( .A(n_704), .Y(n_773) );
HB1xp67_ASAP7_75t_L g807 ( .A(n_704), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_706), .B(n_731), .Y(n_705) );
INVx2_ASAP7_75t_SL g707 ( .A(n_708), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_709), .B(n_710), .Y(n_708) );
INVx2_ASAP7_75t_L g777 ( .A(n_709), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_709), .B(n_729), .Y(n_782) );
AND2x2_ASAP7_75t_L g795 ( .A(n_710), .B(n_796), .Y(n_795) );
BUFx3_ASAP7_75t_L g855 ( .A(n_710), .Y(n_855) );
INVx1_ASAP7_75t_L g857 ( .A(n_711), .Y(n_857) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
AND2x2_ASAP7_75t_L g835 ( .A(n_714), .B(n_836), .Y(n_835) );
NAND2x1_ASAP7_75t_L g821 ( .A(n_715), .B(n_822), .Y(n_821) );
INVx3_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx2_ASAP7_75t_L g848 ( .A(n_716), .Y(n_848) );
OR2x6_ASAP7_75t_L g716 ( .A(n_717), .B(n_721), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g811 ( .A(n_718), .Y(n_811) );
AND2x2_ASAP7_75t_L g871 ( .A(n_718), .B(n_721), .Y(n_871) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
AND2x2_ASAP7_75t_L g752 ( .A(n_720), .B(n_753), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_720), .B(n_791), .Y(n_790) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_721), .B(n_763), .Y(n_762) );
INVx2_ASAP7_75t_L g862 ( .A(n_721), .Y(n_862) );
NAND2x1_ASAP7_75t_L g722 ( .A(n_723), .B(n_727), .Y(n_722) );
INVx2_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
HB1xp67_ASAP7_75t_L g825 ( .A(n_724), .Y(n_825) );
AND2x2_ASAP7_75t_L g724 ( .A(n_725), .B(n_726), .Y(n_724) );
INVx2_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
AOI221x1_ASAP7_75t_L g731 ( .A1(n_732), .A2(n_734), .B1(n_737), .B2(n_741), .C(n_744), .Y(n_731) );
INVx3_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
AOI22xp5_ASAP7_75t_L g766 ( .A1(n_734), .A2(n_767), .B1(n_771), .B2(n_772), .Y(n_766) );
AOI22xp5_ASAP7_75t_L g774 ( .A1(n_734), .A2(n_775), .B1(n_778), .B2(n_781), .Y(n_774) );
INVxp67_ASAP7_75t_SL g872 ( .A(n_734), .Y(n_872) );
AND2x4_ASAP7_75t_L g734 ( .A(n_735), .B(n_736), .Y(n_734) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
OR2x2_ASAP7_75t_L g812 ( .A(n_739), .B(n_813), .Y(n_812) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVxp67_ASAP7_75t_SL g755 ( .A(n_742), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_742), .B(n_777), .Y(n_776) );
HB1xp67_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
OAI22xp5_ASAP7_75t_L g744 ( .A1(n_745), .A2(n_746), .B1(n_750), .B2(n_755), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_747), .B(n_748), .Y(n_746) );
AND2x4_ASAP7_75t_L g815 ( .A(n_747), .B(n_760), .Y(n_815) );
AOI22xp5_ASAP7_75t_L g757 ( .A1(n_748), .A2(n_758), .B1(n_761), .B2(n_764), .Y(n_757) );
AND2x2_ASAP7_75t_L g838 ( .A(n_748), .B(n_805), .Y(n_838) );
OR2x2_ASAP7_75t_L g750 ( .A(n_751), .B(n_754), .Y(n_750) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
AND2x2_ASAP7_75t_L g819 ( .A(n_752), .B(n_820), .Y(n_819) );
INVx1_ASAP7_75t_L g840 ( .A(n_752), .Y(n_840) );
AND2x2_ASAP7_75t_L g861 ( .A(n_752), .B(n_862), .Y(n_861) );
AND2x2_ASAP7_75t_L g878 ( .A(n_752), .B(n_879), .Y(n_878) );
NAND3xp33_ASAP7_75t_SL g756 ( .A(n_757), .B(n_766), .C(n_774), .Y(n_756) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx1_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_763), .B(n_780), .Y(n_779) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
AND2x2_ASAP7_75t_L g767 ( .A(n_768), .B(n_769), .Y(n_767) );
INVx2_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
INVxp67_ASAP7_75t_L g809 ( .A(n_771), .Y(n_809) );
OAI21xp5_ASAP7_75t_L g832 ( .A1(n_772), .A2(n_833), .B(n_835), .Y(n_832) );
INVx1_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
INVxp67_ASAP7_75t_SL g778 ( .A(n_779), .Y(n_778) );
INVx1_ASAP7_75t_L g877 ( .A(n_780), .Y(n_877) );
INVx1_ASAP7_75t_L g793 ( .A(n_781), .Y(n_793) );
INVx2_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
NOR2x1_ASAP7_75t_L g783 ( .A(n_784), .B(n_842), .Y(n_783) );
NAND3xp33_ASAP7_75t_SL g784 ( .A(n_785), .B(n_799), .C(n_816), .Y(n_784) );
AOI21xp5_ASAP7_75t_L g785 ( .A1(n_786), .A2(n_788), .B(n_792), .Y(n_785) );
INVx1_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
HB1xp67_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
INVx2_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
AOI21xp5_ASAP7_75t_L g792 ( .A1(n_793), .A2(n_794), .B(n_797), .Y(n_792) );
INVx1_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
OAI22xp5_ASAP7_75t_SL g876 ( .A1(n_796), .A2(n_851), .B1(n_862), .B2(n_877), .Y(n_876) );
INVx1_ASAP7_75t_L g884 ( .A(n_796), .Y(n_884) );
INVx2_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
AOI21xp5_ASAP7_75t_L g799 ( .A1(n_800), .A2(n_806), .B(n_808), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_801), .B(n_803), .Y(n_800) );
INVx2_ASAP7_75t_SL g801 ( .A(n_802), .Y(n_801) );
INVx1_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
INVx1_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
OAI22xp5_ASAP7_75t_L g808 ( .A1(n_809), .A2(n_810), .B1(n_812), .B2(n_814), .Y(n_808) );
INVx1_ASAP7_75t_L g828 ( .A(n_811), .Y(n_828) );
INVx2_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
AOI21xp5_ASAP7_75t_L g858 ( .A1(n_815), .A2(n_839), .B(n_859), .Y(n_858) );
AOI21xp5_ASAP7_75t_L g816 ( .A1(n_817), .A2(n_825), .B(n_826), .Y(n_816) );
NAND2xp5_ASAP7_75t_L g817 ( .A(n_818), .B(n_821), .Y(n_817) );
INVx1_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g870 ( .A(n_822), .B(n_871), .Y(n_870) );
INVx2_ASAP7_75t_SL g822 ( .A(n_823), .Y(n_822) );
INVx2_ASAP7_75t_L g847 ( .A(n_824), .Y(n_847) );
NAND3xp33_ASAP7_75t_SL g826 ( .A(n_827), .B(n_832), .C(n_837), .Y(n_826) );
NAND3xp33_ASAP7_75t_SL g827 ( .A(n_828), .B(n_829), .C(n_831), .Y(n_827) );
AND2x2_ASAP7_75t_L g859 ( .A(n_830), .B(n_852), .Y(n_859) );
INVx1_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
NAND3xp33_ASAP7_75t_L g837 ( .A(n_838), .B(n_839), .C(n_841), .Y(n_837) );
INVx1_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
NAND2xp5_ASAP7_75t_L g842 ( .A(n_843), .B(n_868), .Y(n_842) );
AOI21xp5_ASAP7_75t_L g843 ( .A1(n_844), .A2(n_849), .B(n_856), .Y(n_843) );
INVx1_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
NAND2x1p5_ASAP7_75t_L g845 ( .A(n_846), .B(n_848), .Y(n_845) );
INVx1_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
NAND4xp25_ASAP7_75t_SL g849 ( .A(n_850), .B(n_851), .C(n_853), .D(n_854), .Y(n_849) );
INVx3_ASAP7_75t_R g851 ( .A(n_852), .Y(n_851) );
INVx1_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
OAI21xp5_ASAP7_75t_SL g856 ( .A1(n_857), .A2(n_858), .B(n_860), .Y(n_856) );
AOI22xp5_ASAP7_75t_L g860 ( .A1(n_861), .A2(n_863), .B1(n_865), .B2(n_866), .Y(n_860) );
INVx2_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
INVx2_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
NOR2xp33_ASAP7_75t_L g868 ( .A(n_869), .B(n_874), .Y(n_868) );
AOI21xp5_ASAP7_75t_SL g869 ( .A1(n_870), .A2(n_872), .B(n_873), .Y(n_869) );
AOI22xp5_ASAP7_75t_L g881 ( .A1(n_871), .A2(n_880), .B1(n_882), .B2(n_884), .Y(n_881) );
NAND2xp5_ASAP7_75t_SL g874 ( .A(n_875), .B(n_881), .Y(n_874) );
INVx2_ASAP7_75t_SL g882 ( .A(n_883), .Y(n_882) );
CKINVDCx10_ASAP7_75t_R g885 ( .A(n_886), .Y(n_885) );
BUFx4f_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
OR2x6_ASAP7_75t_L g889 ( .A(n_890), .B(n_895), .Y(n_889) );
AND2x2_ASAP7_75t_L g890 ( .A(n_891), .B(n_893), .Y(n_890) );
HB1xp67_ASAP7_75t_L g891 ( .A(n_892), .Y(n_891) );
BUFx2_ASAP7_75t_L g893 ( .A(n_894), .Y(n_893) );
INVx1_ASAP7_75t_L g904 ( .A(n_894), .Y(n_904) );
INVx3_ASAP7_75t_L g895 ( .A(n_896), .Y(n_895) );
BUFx6f_ASAP7_75t_L g916 ( .A(n_896), .Y(n_916) );
NAND2xp5_ASAP7_75t_L g919 ( .A(n_896), .B(n_920), .Y(n_919) );
OAI21xp5_ASAP7_75t_SL g898 ( .A1(n_899), .A2(n_906), .B(n_910), .Y(n_898) );
CKINVDCx5p33_ASAP7_75t_R g899 ( .A(n_900), .Y(n_899) );
INVx1_ASAP7_75t_L g900 ( .A(n_901), .Y(n_900) );
INVxp67_ASAP7_75t_L g901 ( .A(n_902), .Y(n_901) );
BUFx3_ASAP7_75t_L g914 ( .A(n_902), .Y(n_914) );
INVx2_ASAP7_75t_L g902 ( .A(n_903), .Y(n_902) );
NOR2x1p5_ASAP7_75t_L g903 ( .A(n_904), .B(n_905), .Y(n_903) );
INVx2_ASAP7_75t_SL g907 ( .A(n_908), .Y(n_907) );
INVxp67_ASAP7_75t_L g910 ( .A(n_911), .Y(n_910) );
NOR2xp33_ASAP7_75t_L g911 ( .A(n_912), .B(n_913), .Y(n_911) );
BUFx6f_ASAP7_75t_L g913 ( .A(n_914), .Y(n_913) );
CKINVDCx5p33_ASAP7_75t_R g915 ( .A(n_916), .Y(n_915) );
INVx2_ASAP7_75t_SL g917 ( .A(n_918), .Y(n_917) );
BUFx3_ASAP7_75t_L g918 ( .A(n_919), .Y(n_918) );
INVx4_ASAP7_75t_SL g921 ( .A(n_922), .Y(n_921) );
endmodule