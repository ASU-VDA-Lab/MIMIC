module real_aes_7608_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_666;
wire n_537;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_746;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_754;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_527;
wire n_434;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_349;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g551 ( .A1(n_0), .A2(n_176), .B(n_552), .C(n_555), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_1), .B(n_502), .Y(n_556) );
INVx1_ASAP7_75t_L g110 ( .A(n_2), .Y(n_110) );
INVx1_ASAP7_75t_L g188 ( .A(n_3), .Y(n_188) );
NAND2xp5_ASAP7_75t_SL g542 ( .A(n_4), .B(n_148), .Y(n_542) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_5), .A2(n_475), .B(n_496), .Y(n_495) );
AO21x2_ASAP7_75t_L g504 ( .A1(n_6), .A2(n_168), .B(n_505), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g196 ( .A1(n_7), .A2(n_38), .B1(n_142), .B2(n_197), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_8), .B(n_168), .Y(n_177) );
AND2x6_ASAP7_75t_L g160 ( .A(n_9), .B(n_161), .Y(n_160) );
A2O1A1Ixp33_ASAP7_75t_L g564 ( .A1(n_10), .A2(n_160), .B(n_480), .C(n_565), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_11), .B(n_116), .Y(n_115) );
NOR2xp33_ASAP7_75t_L g436 ( .A(n_11), .B(n_39), .Y(n_436) );
INVx1_ASAP7_75t_L g138 ( .A(n_12), .Y(n_138) );
INVx1_ASAP7_75t_L g181 ( .A(n_13), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_14), .B(n_146), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g510 ( .A(n_15), .B(n_148), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_16), .B(n_134), .Y(n_252) );
AO32x2_ASAP7_75t_L g194 ( .A1(n_17), .A2(n_133), .A3(n_159), .B1(n_168), .B2(n_195), .Y(n_194) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_18), .B(n_142), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_19), .B(n_134), .Y(n_190) );
AOI22xp33_ASAP7_75t_L g198 ( .A1(n_20), .A2(n_54), .B1(n_142), .B2(n_197), .Y(n_198) );
AOI22xp33_ASAP7_75t_SL g236 ( .A1(n_21), .A2(n_81), .B1(n_142), .B2(n_146), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_22), .B(n_142), .Y(n_209) );
A2O1A1Ixp33_ASAP7_75t_L g528 ( .A1(n_23), .A2(n_159), .B(n_480), .C(n_529), .Y(n_528) );
OAI22xp5_ASAP7_75t_SL g123 ( .A1(n_24), .A2(n_60), .B1(n_124), .B2(n_125), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_24), .Y(n_124) );
A2O1A1Ixp33_ASAP7_75t_L g507 ( .A1(n_25), .A2(n_159), .B(n_480), .C(n_508), .Y(n_507) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_26), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_27), .B(n_163), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_28), .B(n_441), .Y(n_440) );
AOI21xp5_ASAP7_75t_L g548 ( .A1(n_29), .A2(n_475), .B(n_549), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_30), .B(n_163), .Y(n_211) );
INVx2_ASAP7_75t_L g144 ( .A(n_31), .Y(n_144) );
A2O1A1Ixp33_ASAP7_75t_L g517 ( .A1(n_32), .A2(n_478), .B(n_488), .C(n_518), .Y(n_517) );
NAND2xp5_ASAP7_75t_SL g141 ( .A(n_33), .B(n_142), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_34), .B(n_163), .Y(n_222) );
XNOR2x2_ASAP7_75t_SL g121 ( .A(n_35), .B(n_122), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_36), .B(n_218), .Y(n_509) );
OAI22xp5_ASAP7_75t_L g456 ( .A1(n_37), .A2(n_85), .B1(n_457), .B2(n_458), .Y(n_456) );
CKINVDCx20_ASAP7_75t_R g457 ( .A(n_37), .Y(n_457) );
INVx1_ASAP7_75t_L g116 ( .A(n_39), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_40), .B(n_527), .Y(n_526) );
CKINVDCx20_ASAP7_75t_R g569 ( .A(n_41), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_42), .B(n_148), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_43), .B(n_475), .Y(n_506) );
A2O1A1Ixp33_ASAP7_75t_L g477 ( .A1(n_44), .A2(n_478), .B(n_482), .C(n_488), .Y(n_477) );
OAI321xp33_ASAP7_75t_L g120 ( .A1(n_45), .A2(n_121), .A3(n_430), .B1(n_437), .B2(n_438), .C(n_440), .Y(n_120) );
INVx1_ASAP7_75t_L g437 ( .A(n_45), .Y(n_437) );
NAND2xp5_ASAP7_75t_SL g171 ( .A(n_46), .B(n_142), .Y(n_171) );
INVx1_ASAP7_75t_L g553 ( .A(n_47), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g234 ( .A1(n_48), .A2(n_91), .B1(n_197), .B2(n_235), .Y(n_234) );
INVx1_ASAP7_75t_L g483 ( .A(n_49), .Y(n_483) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_50), .B(n_142), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_51), .B(n_142), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_52), .B(n_475), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_53), .B(n_154), .Y(n_175) );
AOI22xp33_ASAP7_75t_SL g250 ( .A1(n_55), .A2(n_61), .B1(n_142), .B2(n_146), .Y(n_250) );
CKINVDCx20_ASAP7_75t_R g534 ( .A(n_56), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_57), .B(n_447), .Y(n_446) );
NAND2xp5_ASAP7_75t_SL g156 ( .A(n_58), .B(n_142), .Y(n_156) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_59), .B(n_142), .Y(n_215) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_60), .Y(n_125) );
OAI22xp5_ASAP7_75t_SL g463 ( .A1(n_60), .A2(n_125), .B1(n_126), .B2(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g161 ( .A(n_62), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_63), .B(n_475), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_64), .B(n_502), .Y(n_501) );
A2O1A1Ixp33_ASAP7_75t_L g498 ( .A1(n_65), .A2(n_154), .B(n_184), .C(n_499), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_66), .B(n_142), .Y(n_189) );
INVx1_ASAP7_75t_L g137 ( .A(n_67), .Y(n_137) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_68), .Y(n_119) );
NAND2xp5_ASAP7_75t_SL g520 ( .A(n_69), .B(n_148), .Y(n_520) );
AO32x2_ASAP7_75t_L g232 ( .A1(n_70), .A2(n_159), .A3(n_168), .B1(n_233), .B2(n_237), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_71), .B(n_149), .Y(n_566) );
INVx1_ASAP7_75t_L g152 ( .A(n_72), .Y(n_152) );
INVx1_ASAP7_75t_L g206 ( .A(n_73), .Y(n_206) );
CKINVDCx16_ASAP7_75t_R g550 ( .A(n_74), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_75), .B(n_485), .Y(n_530) );
A2O1A1Ixp33_ASAP7_75t_L g539 ( .A1(n_76), .A2(n_480), .B(n_488), .C(n_540), .Y(n_539) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_77), .B(n_146), .Y(n_207) );
CKINVDCx16_ASAP7_75t_R g497 ( .A(n_78), .Y(n_497) );
INVx1_ASAP7_75t_L g113 ( .A(n_79), .Y(n_113) );
NAND2xp5_ASAP7_75t_SL g531 ( .A(n_80), .B(n_484), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_82), .B(n_197), .Y(n_221) );
CKINVDCx20_ASAP7_75t_R g522 ( .A(n_83), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_84), .B(n_146), .Y(n_210) );
INVx1_ASAP7_75t_L g458 ( .A(n_85), .Y(n_458) );
INVx2_ASAP7_75t_L g135 ( .A(n_86), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g546 ( .A(n_87), .Y(n_546) );
NAND2xp5_ASAP7_75t_SL g567 ( .A(n_88), .B(n_158), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_89), .B(n_146), .Y(n_172) );
NAND3xp33_ASAP7_75t_SL g109 ( .A(n_90), .B(n_110), .C(n_111), .Y(n_109) );
OR2x2_ASAP7_75t_L g433 ( .A(n_90), .B(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g450 ( .A(n_90), .Y(n_450) );
OR2x2_ASAP7_75t_L g462 ( .A(n_90), .B(n_435), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g249 ( .A1(n_92), .A2(n_103), .B1(n_146), .B2(n_147), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_93), .B(n_475), .Y(n_516) );
INVx1_ASAP7_75t_L g519 ( .A(n_94), .Y(n_519) );
INVxp67_ASAP7_75t_L g500 ( .A(n_95), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_96), .B(n_146), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_97), .B(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g541 ( .A(n_98), .Y(n_541) );
INVx1_ASAP7_75t_L g562 ( .A(n_99), .Y(n_562) );
AOI22xp5_ASAP7_75t_L g104 ( .A1(n_100), .A2(n_105), .B1(n_117), .B2(n_771), .Y(n_104) );
AOI22xp5_ASAP7_75t_L g453 ( .A1(n_101), .A2(n_454), .B1(n_455), .B2(n_456), .Y(n_453) );
CKINVDCx20_ASAP7_75t_R g454 ( .A(n_101), .Y(n_454) );
AND2x2_ASAP7_75t_L g490 ( .A(n_102), .B(n_163), .Y(n_490) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx2_ASAP7_75t_SL g773 ( .A(n_107), .Y(n_773) );
AND2x2_ASAP7_75t_SL g107 ( .A(n_108), .B(n_114), .Y(n_107) );
CKINVDCx16_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
AND2x2_ASAP7_75t_L g435 ( .A(n_110), .B(n_436), .Y(n_435) );
OA211x2_ASAP7_75t_L g117 ( .A1(n_111), .A2(n_118), .B(n_120), .C(n_444), .Y(n_117) );
INVx1_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
INVxp67_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_L g445 ( .A(n_119), .Y(n_445) );
NAND2x1p5_ASAP7_75t_L g438 ( .A(n_121), .B(n_439), .Y(n_438) );
XNOR2xp5_ASAP7_75t_L g122 ( .A(n_123), .B(n_126), .Y(n_122) );
INVx1_ASAP7_75t_SL g464 ( .A(n_126), .Y(n_464) );
OR3x1_ASAP7_75t_L g126 ( .A(n_127), .B(n_358), .C(n_407), .Y(n_126) );
NAND5xp2_ASAP7_75t_L g127 ( .A(n_128), .B(n_273), .C(n_301), .D(n_331), .E(n_345), .Y(n_127) );
AOI221xp5_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_191), .B1(n_223), .B2(n_228), .C(n_239), .Y(n_128) );
NOR2xp33_ASAP7_75t_L g129 ( .A(n_130), .B(n_164), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_130), .B(n_225), .Y(n_224) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx2_ASAP7_75t_L g253 ( .A(n_131), .Y(n_253) );
AND2x2_ASAP7_75t_L g261 ( .A(n_131), .B(n_167), .Y(n_261) );
AND2x2_ASAP7_75t_L g284 ( .A(n_131), .B(n_166), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_131), .B(n_178), .Y(n_299) );
OR2x2_ASAP7_75t_L g308 ( .A(n_131), .B(n_246), .Y(n_308) );
HB1xp67_ASAP7_75t_L g311 ( .A(n_131), .Y(n_311) );
AND2x2_ASAP7_75t_L g419 ( .A(n_131), .B(n_246), .Y(n_419) );
OA21x2_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_139), .B(n_162), .Y(n_131) );
OA21x2_ASAP7_75t_L g178 ( .A1(n_132), .A2(n_179), .B(n_190), .Y(n_178) );
INVx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
NOR2xp33_ASAP7_75t_L g568 ( .A(n_133), .B(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_134), .Y(n_168) );
AND2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_136), .Y(n_134) );
AND2x2_ASAP7_75t_SL g163 ( .A(n_135), .B(n_136), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_137), .B(n_138), .Y(n_136) );
OAI21xp5_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_151), .B(n_159), .Y(n_139) );
AOI21xp5_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_145), .B(n_148), .Y(n_140) );
INVx3_ASAP7_75t_L g205 ( .A(n_142), .Y(n_205) );
HB1xp67_ASAP7_75t_L g543 ( .A(n_142), .Y(n_543) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx1_ASAP7_75t_L g197 ( .A(n_143), .Y(n_197) );
BUFx3_ASAP7_75t_L g235 ( .A(n_143), .Y(n_235) );
AND2x6_ASAP7_75t_L g480 ( .A(n_143), .B(n_481), .Y(n_480) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx1_ASAP7_75t_L g147 ( .A(n_144), .Y(n_147) );
INVx1_ASAP7_75t_L g155 ( .A(n_144), .Y(n_155) );
INVx2_ASAP7_75t_L g182 ( .A(n_146), .Y(n_182) );
INVx3_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_148), .A2(n_171), .B(n_172), .Y(n_170) );
INVx2_ASAP7_75t_L g176 ( .A(n_148), .Y(n_176) );
O2A1O1Ixp5_ASAP7_75t_SL g204 ( .A1(n_148), .A2(n_205), .B(n_206), .C(n_207), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_148), .B(n_500), .Y(n_499) );
INVx5_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
OAI22xp5_ASAP7_75t_SL g233 ( .A1(n_149), .A2(n_158), .B1(n_234), .B2(n_236), .Y(n_233) );
INVx3_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_150), .Y(n_158) );
BUFx6f_ASAP7_75t_L g186 ( .A(n_150), .Y(n_186) );
INVx1_ASAP7_75t_L g218 ( .A(n_150), .Y(n_218) );
AND2x2_ASAP7_75t_L g476 ( .A(n_150), .B(n_155), .Y(n_476) );
INVx1_ASAP7_75t_L g481 ( .A(n_150), .Y(n_481) );
O2A1O1Ixp5_ASAP7_75t_L g151 ( .A1(n_152), .A2(n_153), .B(n_156), .C(n_157), .Y(n_151) );
O2A1O1Ixp33_ASAP7_75t_L g187 ( .A1(n_153), .A2(n_176), .B(n_188), .C(n_189), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_153), .A2(n_530), .B(n_531), .Y(n_529) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_157), .A2(n_220), .B(n_221), .Y(n_219) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
OAI22xp5_ASAP7_75t_L g195 ( .A1(n_158), .A2(n_176), .B1(n_196), .B2(n_198), .Y(n_195) );
OAI22xp5_ASAP7_75t_L g248 ( .A1(n_158), .A2(n_176), .B1(n_249), .B2(n_250), .Y(n_248) );
INVx4_ASAP7_75t_L g554 ( .A(n_158), .Y(n_554) );
NAND3xp33_ASAP7_75t_L g272 ( .A(n_159), .B(n_247), .C(n_248), .Y(n_272) );
BUFx3_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
OAI21xp5_ASAP7_75t_L g169 ( .A1(n_160), .A2(n_170), .B(n_173), .Y(n_169) );
OAI21xp5_ASAP7_75t_L g179 ( .A1(n_160), .A2(n_180), .B(n_187), .Y(n_179) );
OAI21xp5_ASAP7_75t_L g203 ( .A1(n_160), .A2(n_204), .B(n_208), .Y(n_203) );
OAI21xp5_ASAP7_75t_L g213 ( .A1(n_160), .A2(n_214), .B(n_219), .Y(n_213) );
AND2x4_ASAP7_75t_L g475 ( .A(n_160), .B(n_476), .Y(n_475) );
INVx4_ASAP7_75t_SL g489 ( .A(n_160), .Y(n_489) );
NAND2x1p5_ASAP7_75t_L g563 ( .A(n_160), .B(n_476), .Y(n_563) );
OA21x2_ASAP7_75t_L g202 ( .A1(n_163), .A2(n_203), .B(n_211), .Y(n_202) );
OA21x2_ASAP7_75t_L g212 ( .A1(n_163), .A2(n_213), .B(n_222), .Y(n_212) );
INVx2_ASAP7_75t_L g237 ( .A(n_163), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g473 ( .A1(n_163), .A2(n_474), .B(n_477), .Y(n_473) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_163), .A2(n_516), .B(n_517), .Y(n_515) );
INVx1_ASAP7_75t_L g535 ( .A(n_163), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g367 ( .A(n_164), .B(n_311), .Y(n_367) );
INVx2_ASAP7_75t_SL g164 ( .A(n_165), .Y(n_164) );
OAI311xp33_ASAP7_75t_L g309 ( .A1(n_165), .A2(n_310), .A3(n_311), .B1(n_312), .C1(n_327), .Y(n_309) );
AND2x2_ASAP7_75t_L g165 ( .A(n_166), .B(n_178), .Y(n_165) );
AND2x2_ASAP7_75t_L g270 ( .A(n_166), .B(n_271), .Y(n_270) );
INVx2_ASAP7_75t_L g277 ( .A(n_166), .Y(n_277) );
AND2x2_ASAP7_75t_L g398 ( .A(n_166), .B(n_227), .Y(n_398) );
INVx3_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_167), .B(n_227), .Y(n_226) );
AND2x2_ASAP7_75t_L g254 ( .A(n_167), .B(n_178), .Y(n_254) );
AND2x2_ASAP7_75t_L g306 ( .A(n_167), .B(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g320 ( .A(n_167), .B(n_253), .Y(n_320) );
OA21x2_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_169), .B(n_177), .Y(n_167) );
INVx4_ASAP7_75t_L g247 ( .A(n_168), .Y(n_247) );
HB1xp67_ASAP7_75t_L g494 ( .A(n_168), .Y(n_494) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_168), .A2(n_506), .B(n_507), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_175), .B(n_176), .Y(n_173) );
INVx2_ASAP7_75t_L g227 ( .A(n_178), .Y(n_227) );
AND2x2_ASAP7_75t_L g269 ( .A(n_178), .B(n_253), .Y(n_269) );
O2A1O1Ixp33_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_182), .B(n_183), .C(n_184), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_182), .A2(n_509), .B(n_510), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g565 ( .A1(n_182), .A2(n_566), .B(n_567), .Y(n_565) );
O2A1O1Ixp33_ASAP7_75t_L g540 ( .A1(n_184), .A2(n_541), .B(n_542), .C(n_543), .Y(n_540) );
INVx1_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_185), .A2(n_209), .B(n_210), .Y(n_208) );
INVx4_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
INVx2_ASAP7_75t_L g485 ( .A(n_186), .Y(n_485) );
AND2x2_ASAP7_75t_L g191 ( .A(n_192), .B(n_199), .Y(n_191) );
OR2x2_ASAP7_75t_L g364 ( .A(n_192), .B(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_192), .B(n_370), .Y(n_381) );
INVx2_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g376 ( .A(n_193), .B(n_377), .Y(n_376) );
BUFx2_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
INVx2_ASAP7_75t_L g238 ( .A(n_194), .Y(n_238) );
AND2x2_ASAP7_75t_L g305 ( .A(n_194), .B(n_232), .Y(n_305) );
AND2x2_ASAP7_75t_L g316 ( .A(n_194), .B(n_212), .Y(n_316) );
AND2x2_ASAP7_75t_L g325 ( .A(n_194), .B(n_326), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_199), .B(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_199), .B(n_266), .Y(n_310) );
INVx2_ASAP7_75t_SL g199 ( .A(n_200), .Y(n_199) );
OR2x2_ASAP7_75t_L g297 ( .A(n_200), .B(n_256), .Y(n_297) );
OR2x2_ASAP7_75t_L g200 ( .A(n_201), .B(n_212), .Y(n_200) );
INVx2_ASAP7_75t_L g230 ( .A(n_201), .Y(n_230) );
AND2x2_ASAP7_75t_L g324 ( .A(n_201), .B(n_325), .Y(n_324) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx2_ASAP7_75t_L g242 ( .A(n_202), .Y(n_242) );
OR2x2_ASAP7_75t_L g341 ( .A(n_202), .B(n_342), .Y(n_341) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_202), .Y(n_404) );
AND2x2_ASAP7_75t_L g243 ( .A(n_212), .B(n_238), .Y(n_243) );
INVx1_ASAP7_75t_L g264 ( .A(n_212), .Y(n_264) );
AND2x2_ASAP7_75t_L g285 ( .A(n_212), .B(n_286), .Y(n_285) );
INVx2_ASAP7_75t_L g326 ( .A(n_212), .Y(n_326) );
INVx1_ASAP7_75t_L g342 ( .A(n_212), .Y(n_342) );
HB1xp67_ASAP7_75t_L g417 ( .A(n_212), .Y(n_417) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_215), .A2(n_216), .B(n_217), .Y(n_214) );
INVx1_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVxp67_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_225), .B(n_330), .Y(n_371) );
OAI22xp5_ASAP7_75t_L g373 ( .A1(n_225), .A2(n_315), .B1(n_364), .B2(n_374), .Y(n_373) );
INVx1_ASAP7_75t_SL g225 ( .A(n_226), .Y(n_225) );
OAI211xp5_ASAP7_75t_SL g407 ( .A1(n_226), .A2(n_408), .B(n_410), .C(n_428), .Y(n_407) );
INVx2_ASAP7_75t_L g260 ( .A(n_227), .Y(n_260) );
AND2x2_ASAP7_75t_L g318 ( .A(n_227), .B(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g329 ( .A(n_227), .B(n_330), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_228), .B(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g228 ( .A(n_229), .B(n_231), .Y(n_228) );
AND2x2_ASAP7_75t_L g302 ( .A(n_229), .B(n_266), .Y(n_302) );
BUFx2_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
AND2x2_ASAP7_75t_L g334 ( .A(n_230), .B(n_325), .Y(n_334) );
AND2x2_ASAP7_75t_L g353 ( .A(n_230), .B(n_267), .Y(n_353) );
AND2x4_ASAP7_75t_L g289 ( .A(n_231), .B(n_263), .Y(n_289) );
AND2x2_ASAP7_75t_L g427 ( .A(n_231), .B(n_403), .Y(n_427) );
AND2x2_ASAP7_75t_L g231 ( .A(n_232), .B(n_238), .Y(n_231) );
BUFx6f_ASAP7_75t_L g256 ( .A(n_232), .Y(n_256) );
INVx1_ASAP7_75t_L g267 ( .A(n_232), .Y(n_267) );
INVx1_ASAP7_75t_L g366 ( .A(n_232), .Y(n_366) );
HB1xp67_ASAP7_75t_L g487 ( .A(n_235), .Y(n_487) );
INVx2_ASAP7_75t_L g555 ( .A(n_235), .Y(n_555) );
INVx1_ASAP7_75t_L g532 ( .A(n_237), .Y(n_532) );
OR2x2_ASAP7_75t_L g257 ( .A(n_238), .B(n_242), .Y(n_257) );
AND2x2_ASAP7_75t_L g266 ( .A(n_238), .B(n_267), .Y(n_266) );
NOR2xp67_ASAP7_75t_L g286 ( .A(n_238), .B(n_287), .Y(n_286) );
OAI221xp5_ASAP7_75t_L g239 ( .A1(n_240), .A2(n_244), .B1(n_255), .B2(n_258), .C(n_262), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
A2O1A1Ixp33_ASAP7_75t_L g262 ( .A1(n_241), .A2(n_263), .B(n_265), .C(n_268), .Y(n_262) );
AND2x2_ASAP7_75t_L g241 ( .A(n_242), .B(n_243), .Y(n_241) );
INVx1_ASAP7_75t_L g287 ( .A(n_242), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_242), .B(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_SL g370 ( .A(n_242), .B(n_264), .Y(n_370) );
HB1xp67_ASAP7_75t_L g377 ( .A(n_242), .Y(n_377) );
AND2x2_ASAP7_75t_L g295 ( .A(n_243), .B(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g332 ( .A(n_243), .B(n_333), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_245), .B(n_254), .Y(n_244) );
INVx2_ASAP7_75t_L g323 ( .A(n_245), .Y(n_323) );
AOI222xp33_ASAP7_75t_L g372 ( .A1(n_245), .A2(n_256), .B1(n_373), .B2(n_375), .C1(n_376), .C2(n_378), .Y(n_372) );
AND2x2_ASAP7_75t_L g429 ( .A(n_245), .B(n_398), .Y(n_429) );
AND2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_253), .Y(n_245) );
INVx1_ASAP7_75t_L g319 ( .A(n_246), .Y(n_319) );
AO21x1_ASAP7_75t_L g246 ( .A1(n_247), .A2(n_248), .B(n_251), .Y(n_246) );
INVx3_ASAP7_75t_L g502 ( .A(n_247), .Y(n_502) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_247), .B(n_522), .Y(n_521) );
AO21x2_ASAP7_75t_L g537 ( .A1(n_247), .A2(n_538), .B(n_545), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g545 ( .A(n_247), .B(n_546), .Y(n_545) );
AO21x2_ASAP7_75t_L g560 ( .A1(n_247), .A2(n_561), .B(n_568), .Y(n_560) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
AND2x4_ASAP7_75t_L g271 ( .A(n_252), .B(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g357 ( .A(n_254), .B(n_291), .Y(n_357) );
AOI21xp33_ASAP7_75t_L g368 ( .A1(n_255), .A2(n_369), .B(n_371), .Y(n_368) );
OR2x2_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .Y(n_255) );
INVx2_ASAP7_75t_L g296 ( .A(n_256), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_256), .B(n_263), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_256), .B(n_409), .Y(n_408) );
INVx1_ASAP7_75t_SL g258 ( .A(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_261), .Y(n_259) );
INVx3_ASAP7_75t_L g322 ( .A(n_260), .Y(n_322) );
OR2x2_ASAP7_75t_L g374 ( .A(n_260), .B(n_296), .Y(n_374) );
AND2x2_ASAP7_75t_L g290 ( .A(n_261), .B(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g328 ( .A(n_261), .B(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_261), .B(n_322), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_261), .B(n_318), .Y(n_344) );
AND2x2_ASAP7_75t_L g348 ( .A(n_261), .B(n_330), .Y(n_348) );
INVxp67_ASAP7_75t_L g280 ( .A(n_263), .Y(n_280) );
BUFx3_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
OAI22xp5_ASAP7_75t_L g337 ( .A1(n_265), .A2(n_338), .B1(n_343), .B2(n_344), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_265), .B(n_370), .Y(n_400) );
INVx1_ASAP7_75t_SL g265 ( .A(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g386 ( .A(n_266), .B(n_377), .Y(n_386) );
AND2x2_ASAP7_75t_L g415 ( .A(n_266), .B(n_416), .Y(n_415) );
AND2x2_ASAP7_75t_L g420 ( .A(n_266), .B(n_370), .Y(n_420) );
INVx1_ASAP7_75t_L g333 ( .A(n_267), .Y(n_333) );
BUFx2_ASAP7_75t_L g339 ( .A(n_267), .Y(n_339) );
INVx1_ASAP7_75t_L g424 ( .A(n_268), .Y(n_424) );
AND2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
NAND2x1p5_ASAP7_75t_L g275 ( .A(n_269), .B(n_276), .Y(n_275) );
INVx1_ASAP7_75t_L g300 ( .A(n_270), .Y(n_300) );
NOR2x1_ASAP7_75t_L g276 ( .A(n_271), .B(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g283 ( .A(n_271), .B(n_284), .Y(n_283) );
INVx2_ASAP7_75t_L g292 ( .A(n_271), .Y(n_292) );
INVx3_ASAP7_75t_L g330 ( .A(n_271), .Y(n_330) );
OR2x2_ASAP7_75t_L g396 ( .A(n_271), .B(n_397), .Y(n_396) );
AOI211xp5_ASAP7_75t_L g273 ( .A1(n_274), .A2(n_278), .B(n_281), .C(n_293), .Y(n_273) );
AOI221xp5_ASAP7_75t_L g410 ( .A1(n_274), .A2(n_411), .B1(n_418), .B2(n_420), .C(n_421), .Y(n_410) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
NAND2xp5_ASAP7_75t_SL g281 ( .A(n_282), .B(n_288), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_283), .B(n_285), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_284), .B(n_322), .Y(n_336) );
AND2x2_ASAP7_75t_L g378 ( .A(n_284), .B(n_318), .Y(n_378) );
INVx1_ASAP7_75t_SL g391 ( .A(n_285), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_285), .B(n_339), .Y(n_394) );
INVx1_ASAP7_75t_L g412 ( .A(n_286), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
AOI221xp5_ASAP7_75t_L g379 ( .A1(n_290), .A2(n_380), .B1(n_382), .B2(n_386), .C(n_387), .Y(n_379) );
AND2x2_ASAP7_75t_L g406 ( .A(n_291), .B(n_398), .Y(n_406) );
INVx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
INVx1_ASAP7_75t_L g390 ( .A(n_292), .Y(n_390) );
AOI21xp33_ASAP7_75t_SL g293 ( .A1(n_294), .A2(n_297), .B(n_298), .Y(n_293) );
INVx1_ASAP7_75t_SL g294 ( .A(n_295), .Y(n_294) );
OR2x2_ASAP7_75t_L g361 ( .A(n_296), .B(n_362), .Y(n_361) );
INVx2_ASAP7_75t_L g347 ( .A(n_297), .Y(n_347) );
INVx1_ASAP7_75t_L g375 ( .A(n_298), .Y(n_375) );
OR2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
O2A1O1Ixp33_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_303), .B(n_306), .C(n_309), .Y(n_301) );
OAI31xp33_ASAP7_75t_L g428 ( .A1(n_302), .A2(n_340), .A3(n_427), .B(n_429), .Y(n_428) );
INVxp67_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g402 ( .A(n_305), .B(n_403), .Y(n_402) );
INVx1_ASAP7_75t_SL g423 ( .A(n_305), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_307), .B(n_322), .Y(n_350) );
INVx1_ASAP7_75t_SL g307 ( .A(n_308), .Y(n_307) );
OR2x2_ASAP7_75t_L g425 ( .A(n_308), .B(n_322), .Y(n_425) );
AOI22xp5_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_317), .B1(n_321), .B2(n_324), .Y(n_312) );
NAND2xp33_ASAP7_75t_L g313 ( .A(n_314), .B(n_315), .Y(n_313) );
INVx2_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_316), .B(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g352 ( .A(n_316), .B(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g355 ( .A(n_316), .B(n_339), .Y(n_355) );
AND2x2_ASAP7_75t_L g409 ( .A(n_316), .B(n_404), .Y(n_409) );
AND2x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_320), .Y(n_317) );
INVx1_ASAP7_75t_L g384 ( .A(n_320), .Y(n_384) );
NOR2xp67_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
OAI32xp33_ASAP7_75t_L g387 ( .A1(n_322), .A2(n_356), .A3(n_388), .B1(n_390), .B2(n_391), .Y(n_387) );
INVx1_ASAP7_75t_L g362 ( .A(n_325), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_325), .B(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g385 ( .A(n_329), .Y(n_385) );
O2A1O1Ixp33_ASAP7_75t_L g331 ( .A1(n_332), .A2(n_334), .B(n_335), .C(n_337), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_333), .B(n_370), .Y(n_369) );
AOI221xp5_ASAP7_75t_L g345 ( .A1(n_334), .A2(n_346), .B1(n_347), .B2(n_348), .C(n_349), .Y(n_345) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
INVx2_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g346 ( .A(n_344), .Y(n_346) );
OAI22xp5_ASAP7_75t_L g349 ( .A1(n_350), .A2(n_351), .B1(n_354), .B2(n_356), .Y(n_349) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
NAND4xp25_ASAP7_75t_SL g411 ( .A(n_354), .B(n_412), .C(n_413), .D(n_414), .Y(n_411) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx1_ASAP7_75t_SL g356 ( .A(n_357), .Y(n_356) );
NAND4xp25_ASAP7_75t_SL g358 ( .A(n_359), .B(n_372), .C(n_379), .D(n_392), .Y(n_358) );
O2A1O1Ixp33_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_363), .B(n_367), .C(n_368), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_SL g389 ( .A(n_365), .Y(n_389) );
INVx2_ASAP7_75t_L g413 ( .A(n_370), .Y(n_413) );
OR2x2_ASAP7_75t_L g422 ( .A(n_377), .B(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
OR2x2_ASAP7_75t_L g383 ( .A(n_384), .B(n_385), .Y(n_383) );
AOI21xp5_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_395), .B(n_399), .Y(n_392) );
INVxp67_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
AND2x2_ASAP7_75t_L g418 ( .A(n_398), .B(n_419), .Y(n_418) );
AOI21xp33_ASAP7_75t_SL g399 ( .A1(n_400), .A2(n_401), .B(n_405), .Y(n_399) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
CKINVDCx16_ASAP7_75t_R g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
OAI22xp5_ASAP7_75t_L g421 ( .A1(n_422), .A2(n_424), .B1(n_425), .B2(n_426), .Y(n_421) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g439 ( .A(n_432), .Y(n_439) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_SL g443 ( .A(n_433), .Y(n_443) );
NOR2x2_ASAP7_75t_L g449 ( .A(n_434), .B(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
OR2x2_ASAP7_75t_L g467 ( .A(n_435), .B(n_450), .Y(n_467) );
NAND4xp25_ASAP7_75t_SL g444 ( .A(n_440), .B(n_445), .C(n_446), .D(n_451), .Y(n_444) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_SL g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_SL g447 ( .A(n_448), .Y(n_447) );
INVx3_ASAP7_75t_SL g448 ( .A(n_449), .Y(n_448) );
AOI22xp5_ASAP7_75t_L g451 ( .A1(n_452), .A2(n_453), .B1(n_459), .B2(n_766), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
OAI22xp5_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_463), .B1(n_465), .B2(n_468), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g767 ( .A(n_461), .Y(n_767) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g768 ( .A(n_463), .Y(n_768) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g769 ( .A(n_466), .Y(n_769) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx4_ASAP7_75t_L g770 ( .A(n_468), .Y(n_770) );
BUFx6f_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
OR5x1_ASAP7_75t_L g469 ( .A(n_470), .B(n_639), .C(n_717), .D(n_741), .E(n_758), .Y(n_469) );
OAI211xp5_ASAP7_75t_SL g470 ( .A1(n_471), .A2(n_511), .B(n_557), .C(n_616), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_472), .B(n_491), .Y(n_471) );
AND2x2_ASAP7_75t_L g570 ( .A(n_472), .B(n_493), .Y(n_570) );
INVx5_ASAP7_75t_SL g598 ( .A(n_472), .Y(n_598) );
AND2x2_ASAP7_75t_L g634 ( .A(n_472), .B(n_619), .Y(n_634) );
OR2x2_ASAP7_75t_L g673 ( .A(n_472), .B(n_492), .Y(n_673) );
OR2x2_ASAP7_75t_L g704 ( .A(n_472), .B(n_595), .Y(n_704) );
NOR2xp33_ASAP7_75t_L g740 ( .A(n_472), .B(n_608), .Y(n_740) );
AND2x2_ASAP7_75t_L g752 ( .A(n_472), .B(n_595), .Y(n_752) );
OR2x6_ASAP7_75t_L g472 ( .A(n_473), .B(n_490), .Y(n_472) );
BUFx2_ASAP7_75t_L g527 ( .A(n_475), .Y(n_527) );
INVx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
O2A1O1Ixp33_ASAP7_75t_L g496 ( .A1(n_479), .A2(n_489), .B(n_497), .C(n_498), .Y(n_496) );
O2A1O1Ixp33_ASAP7_75t_SL g549 ( .A1(n_479), .A2(n_489), .B(n_550), .C(n_551), .Y(n_549) );
INVx5_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
O2A1O1Ixp33_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_484), .B(n_486), .C(n_487), .Y(n_482) );
O2A1O1Ixp33_ASAP7_75t_L g518 ( .A1(n_484), .A2(n_487), .B(n_519), .C(n_520), .Y(n_518) );
INVx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
AND2x2_ASAP7_75t_L g751 ( .A(n_491), .B(n_752), .Y(n_751) );
INVx1_ASAP7_75t_SL g491 ( .A(n_492), .Y(n_491) );
OR2x2_ASAP7_75t_L g614 ( .A(n_492), .B(n_615), .Y(n_614) );
OR2x2_ASAP7_75t_L g492 ( .A(n_493), .B(n_503), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_493), .B(n_595), .Y(n_594) );
HB1xp67_ASAP7_75t_L g607 ( .A(n_493), .Y(n_607) );
INVx3_ASAP7_75t_L g622 ( .A(n_493), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_493), .B(n_503), .Y(n_646) );
OR2x2_ASAP7_75t_L g655 ( .A(n_493), .B(n_598), .Y(n_655) );
AND2x2_ASAP7_75t_L g659 ( .A(n_493), .B(n_619), .Y(n_659) );
AND2x2_ASAP7_75t_L g665 ( .A(n_493), .B(n_666), .Y(n_665) );
INVxp67_ASAP7_75t_L g702 ( .A(n_493), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_493), .B(n_560), .Y(n_716) );
OA21x2_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_495), .B(n_501), .Y(n_493) );
OA21x2_ASAP7_75t_L g547 ( .A1(n_502), .A2(n_548), .B(n_556), .Y(n_547) );
OR2x2_ASAP7_75t_L g608 ( .A(n_503), .B(n_560), .Y(n_608) );
AND2x2_ASAP7_75t_L g619 ( .A(n_503), .B(n_595), .Y(n_619) );
AND2x2_ASAP7_75t_L g631 ( .A(n_503), .B(n_622), .Y(n_631) );
NAND2xp5_ASAP7_75t_SL g654 ( .A(n_503), .B(n_560), .Y(n_654) );
INVx1_ASAP7_75t_SL g666 ( .A(n_503), .Y(n_666) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
AND2x2_ASAP7_75t_L g559 ( .A(n_504), .B(n_560), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_504), .B(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_513), .B(n_523), .Y(n_512) );
AND2x2_ASAP7_75t_L g579 ( .A(n_513), .B(n_580), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_513), .B(n_536), .Y(n_583) );
AND2x2_ASAP7_75t_L g586 ( .A(n_513), .B(n_587), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_513), .B(n_589), .Y(n_588) );
OR2x2_ASAP7_75t_L g611 ( .A(n_513), .B(n_602), .Y(n_611) );
HB1xp67_ASAP7_75t_L g630 ( .A(n_513), .Y(n_630) );
AND2x2_ASAP7_75t_L g651 ( .A(n_513), .B(n_652), .Y(n_651) );
OR2x2_ASAP7_75t_L g661 ( .A(n_513), .B(n_662), .Y(n_661) );
AND2x2_ASAP7_75t_L g707 ( .A(n_513), .B(n_590), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_513), .B(n_613), .Y(n_734) );
INVx5_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
BUFx2_ASAP7_75t_L g604 ( .A(n_514), .Y(n_604) );
AND2x2_ASAP7_75t_L g670 ( .A(n_514), .B(n_602), .Y(n_670) );
AND2x2_ASAP7_75t_L g754 ( .A(n_514), .B(n_622), .Y(n_754) );
OR2x6_ASAP7_75t_L g514 ( .A(n_515), .B(n_521), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_523), .B(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g743 ( .A(n_523), .Y(n_743) );
AND2x2_ASAP7_75t_L g523 ( .A(n_524), .B(n_536), .Y(n_523) );
AND2x2_ASAP7_75t_L g573 ( .A(n_524), .B(n_574), .Y(n_573) );
AND2x4_ASAP7_75t_L g582 ( .A(n_524), .B(n_580), .Y(n_582) );
INVx5_ASAP7_75t_L g590 ( .A(n_524), .Y(n_590) );
AND2x2_ASAP7_75t_L g613 ( .A(n_524), .B(n_547), .Y(n_613) );
HB1xp67_ASAP7_75t_L g650 ( .A(n_524), .Y(n_650) );
OR2x6_ASAP7_75t_L g524 ( .A(n_525), .B(n_533), .Y(n_524) );
AOI21xp5_ASAP7_75t_SL g525 ( .A1(n_526), .A2(n_528), .B(n_532), .Y(n_525) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_534), .B(n_535), .Y(n_533) );
INVx1_ASAP7_75t_L g691 ( .A(n_536), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_536), .B(n_707), .Y(n_706) );
AND2x2_ASAP7_75t_L g724 ( .A(n_536), .B(n_590), .Y(n_724) );
A2O1A1Ixp33_ASAP7_75t_L g753 ( .A1(n_536), .A2(n_647), .B(n_754), .C(n_755), .Y(n_753) );
AND2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_547), .Y(n_536) );
BUFx2_ASAP7_75t_L g574 ( .A(n_537), .Y(n_574) );
INVx2_ASAP7_75t_L g578 ( .A(n_537), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_539), .B(n_544), .Y(n_538) );
INVx2_ASAP7_75t_L g580 ( .A(n_547), .Y(n_580) );
AND2x2_ASAP7_75t_L g587 ( .A(n_547), .B(n_578), .Y(n_587) );
AND2x2_ASAP7_75t_L g678 ( .A(n_547), .B(n_590), .Y(n_678) );
NOR2xp33_ASAP7_75t_L g552 ( .A(n_553), .B(n_554), .Y(n_552) );
AOI211x1_ASAP7_75t_SL g557 ( .A1(n_558), .A2(n_571), .B(n_584), .C(n_609), .Y(n_557) );
INVx1_ASAP7_75t_L g675 ( .A(n_558), .Y(n_675) );
AND2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_570), .Y(n_558) );
INVx5_ASAP7_75t_SL g595 ( .A(n_560), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_560), .B(n_665), .Y(n_664) );
AOI311xp33_ASAP7_75t_L g683 ( .A1(n_560), .A2(n_684), .A3(n_686), .B(n_687), .C(n_693), .Y(n_683) );
A2O1A1Ixp33_ASAP7_75t_L g718 ( .A1(n_560), .A2(n_631), .B(n_719), .C(n_722), .Y(n_718) );
OAI21xp5_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_563), .B(n_564), .Y(n_561) );
INVxp67_ASAP7_75t_L g638 ( .A(n_570), .Y(n_638) );
NAND4xp25_ASAP7_75t_SL g571 ( .A(n_572), .B(n_575), .C(n_581), .D(n_583), .Y(n_571) );
NOR2xp33_ASAP7_75t_L g636 ( .A(n_572), .B(n_637), .Y(n_636) );
INVx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g629 ( .A(n_573), .B(n_630), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_576), .B(n_579), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_576), .B(n_582), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_576), .B(n_589), .Y(n_709) );
BUFx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_577), .B(n_590), .Y(n_727) );
HB1xp67_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx2_ASAP7_75t_L g602 ( .A(n_578), .Y(n_602) );
INVxp67_ASAP7_75t_L g637 ( .A(n_579), .Y(n_637) );
AND2x4_ASAP7_75t_L g589 ( .A(n_580), .B(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g663 ( .A(n_580), .B(n_602), .Y(n_663) );
INVx1_ASAP7_75t_L g690 ( .A(n_580), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_580), .B(n_677), .Y(n_737) );
NOR2xp33_ASAP7_75t_L g671 ( .A(n_581), .B(n_651), .Y(n_671) );
INVx1_ASAP7_75t_SL g581 ( .A(n_582), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_582), .B(n_604), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_582), .B(n_651), .Y(n_750) );
INVx1_ASAP7_75t_L g761 ( .A(n_583), .Y(n_761) );
A2O1A1Ixp33_ASAP7_75t_L g584 ( .A1(n_585), .A2(n_588), .B(n_591), .C(n_599), .Y(n_584) );
INVx1_ASAP7_75t_SL g585 ( .A(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g603 ( .A(n_587), .B(n_604), .Y(n_603) );
AND2x2_ASAP7_75t_L g641 ( .A(n_587), .B(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g623 ( .A(n_588), .Y(n_623) );
AND2x2_ASAP7_75t_L g600 ( .A(n_589), .B(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_589), .B(n_651), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_589), .B(n_670), .Y(n_694) );
OR2x2_ASAP7_75t_L g610 ( .A(n_590), .B(n_611), .Y(n_610) );
INVx2_ASAP7_75t_L g642 ( .A(n_590), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_590), .B(n_602), .Y(n_657) );
AND2x2_ASAP7_75t_L g714 ( .A(n_590), .B(n_670), .Y(n_714) );
HB1xp67_ASAP7_75t_L g721 ( .A(n_590), .Y(n_721) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AOI221xp5_ASAP7_75t_L g725 ( .A1(n_592), .A2(n_604), .B1(n_726), .B2(n_728), .C(n_731), .Y(n_725) );
AND2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_596), .Y(n_592) );
INVx1_ASAP7_75t_SL g593 ( .A(n_594), .Y(n_593) );
OR2x2_ASAP7_75t_L g615 ( .A(n_595), .B(n_598), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_595), .B(n_665), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_595), .B(n_622), .Y(n_730) );
INVx1_ASAP7_75t_SL g596 ( .A(n_597), .Y(n_596) );
OR2x2_ASAP7_75t_L g715 ( .A(n_597), .B(n_716), .Y(n_715) );
OR2x2_ASAP7_75t_L g729 ( .A(n_597), .B(n_730), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_598), .B(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g626 ( .A(n_598), .B(n_619), .Y(n_626) );
AND2x2_ASAP7_75t_L g696 ( .A(n_598), .B(n_697), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_598), .B(n_645), .Y(n_742) );
NOR2xp33_ASAP7_75t_L g745 ( .A(n_598), .B(n_746), .Y(n_745) );
OAI21xp5_ASAP7_75t_SL g599 ( .A1(n_600), .A2(n_603), .B(n_605), .Y(n_599) );
INVx2_ASAP7_75t_L g632 ( .A(n_600), .Y(n_632) );
HB1xp67_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g652 ( .A(n_602), .Y(n_652) );
OR2x2_ASAP7_75t_L g656 ( .A(n_604), .B(n_657), .Y(n_656) );
OR2x2_ASAP7_75t_L g759 ( .A(n_604), .B(n_727), .Y(n_759) );
INVx1_ASAP7_75t_SL g605 ( .A(n_606), .Y(n_605) );
OR2x2_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
AOI21xp33_ASAP7_75t_SL g609 ( .A1(n_610), .A2(n_612), .B(n_614), .Y(n_609) );
INVx1_ASAP7_75t_L g763 ( .A(n_610), .Y(n_763) );
INVx2_ASAP7_75t_SL g677 ( .A(n_611), .Y(n_677) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
A2O1A1Ixp33_ASAP7_75t_L g758 ( .A1(n_614), .A2(n_695), .B(n_759), .C(n_760), .Y(n_758) );
OAI322xp33_ASAP7_75t_SL g627 ( .A1(n_615), .A2(n_628), .A3(n_631), .B1(n_632), .B2(n_633), .C1(n_635), .C2(n_638), .Y(n_627) );
INVx2_ASAP7_75t_L g647 ( .A(n_615), .Y(n_647) );
AOI221xp5_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_623), .B1(n_624), .B2(n_626), .C(n_627), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
OAI22xp33_ASAP7_75t_SL g693 ( .A1(n_618), .A2(n_694), .B1(n_695), .B2(n_698), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_619), .B(n_620), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_619), .B(n_622), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_619), .B(n_757), .Y(n_756) );
INVx2_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
OR2x2_ASAP7_75t_L g692 ( .A(n_621), .B(n_654), .Y(n_692) );
INVx1_ASAP7_75t_L g682 ( .A(n_622), .Y(n_682) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
AOI21xp5_ASAP7_75t_L g735 ( .A1(n_626), .A2(n_736), .B(n_738), .Y(n_735) );
AOI21xp33_ASAP7_75t_L g660 ( .A1(n_628), .A2(n_661), .B(n_664), .Y(n_660) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
NOR2xp67_ASAP7_75t_SL g689 ( .A(n_630), .B(n_690), .Y(n_689) );
NOR2xp33_ASAP7_75t_L g722 ( .A(n_630), .B(n_723), .Y(n_722) );
INVx1_ASAP7_75t_SL g746 ( .A(n_631), .Y(n_746) );
INVx1_ASAP7_75t_SL g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
NAND4xp25_ASAP7_75t_L g639 ( .A(n_640), .B(n_667), .C(n_683), .D(n_699), .Y(n_639) );
AOI211xp5_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_643), .B(n_648), .C(n_660), .Y(n_640) );
INVx1_ASAP7_75t_L g732 ( .A(n_641), .Y(n_732) );
AND2x2_ASAP7_75t_L g680 ( .A(n_642), .B(n_663), .Y(n_680) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_645), .B(n_647), .Y(n_644) );
INVx1_ASAP7_75t_SL g645 ( .A(n_646), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_647), .B(n_682), .Y(n_681) );
OAI22xp33_ASAP7_75t_L g648 ( .A1(n_649), .A2(n_653), .B1(n_656), .B2(n_658), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_650), .B(n_651), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_650), .B(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g698 ( .A(n_651), .Y(n_698) );
O2A1O1Ixp33_ASAP7_75t_L g712 ( .A1(n_651), .A2(n_690), .B(n_713), .C(n_715), .Y(n_712) );
OR2x2_ASAP7_75t_L g653 ( .A(n_654), .B(n_655), .Y(n_653) );
INVx1_ASAP7_75t_L g697 ( .A(n_654), .Y(n_697) );
INVx1_ASAP7_75t_L g757 ( .A(n_655), .Y(n_757) );
NAND2xp33_ASAP7_75t_SL g747 ( .A(n_656), .B(n_748), .Y(n_747) );
INVx1_ASAP7_75t_SL g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx2_ASAP7_75t_L g686 ( .A(n_665), .Y(n_686) );
O2A1O1Ixp33_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_671), .B(n_672), .C(n_674), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
OAI22xp5_ASAP7_75t_L g674 ( .A1(n_675), .A2(n_676), .B1(n_679), .B2(n_681), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_677), .B(n_678), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_677), .B(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_682), .B(n_703), .Y(n_765) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
AOI21xp33_ASAP7_75t_SL g687 ( .A1(n_688), .A2(n_691), .B(n_692), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_SL g695 ( .A(n_696), .Y(n_695) );
AOI221xp5_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_705), .B1(n_708), .B2(n_710), .C(n_712), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_702), .B(n_703), .Y(n_701) );
INVx1_ASAP7_75t_SL g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVxp67_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
OAI22xp5_ASAP7_75t_L g731 ( .A1(n_715), .A2(n_732), .B1(n_733), .B2(n_734), .Y(n_731) );
NAND3xp33_ASAP7_75t_SL g717 ( .A(n_718), .B(n_725), .C(n_735), .Y(n_717) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_SL g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
CKINVDCx16_ASAP7_75t_R g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVxp67_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
OAI211xp5_ASAP7_75t_L g741 ( .A1(n_742), .A2(n_743), .B(n_744), .C(n_753), .Y(n_741) );
INVx1_ASAP7_75t_L g762 ( .A(n_742), .Y(n_762) );
AOI22xp33_ASAP7_75t_L g744 ( .A1(n_745), .A2(n_747), .B1(n_749), .B2(n_751), .Y(n_744) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
AOI22xp5_ASAP7_75t_L g760 ( .A1(n_761), .A2(n_762), .B1(n_763), .B2(n_764), .Y(n_760) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
OAI22x1_ASAP7_75t_SL g766 ( .A1(n_767), .A2(n_768), .B1(n_769), .B2(n_770), .Y(n_766) );
INVx1_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
INVx1_ASAP7_75t_SL g772 ( .A(n_773), .Y(n_772) );
endmodule