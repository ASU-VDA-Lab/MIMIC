module fake_jpeg_11194_n_120 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_120);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_120;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_29),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_36),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_5),
.B(n_9),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_11),
.B(n_3),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_12),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_25),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_28),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_10),
.Y(n_51)
);

BUFx16f_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_49),
.Y(n_53)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_52),
.Y(n_55)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

AND2x2_ASAP7_75t_SL g56 ( 
.A(n_42),
.B(n_0),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_57),
.Y(n_74)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_58),
.B(n_59),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_0),
.Y(n_59)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_60),
.B(n_61),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_1),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_19),
.C(n_31),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_62),
.B(n_39),
.C(n_44),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_70),
.Y(n_81)
);

INVx6_ASAP7_75t_SL g65 ( 
.A(n_55),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_65),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_41),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_67),
.B(n_69),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_51),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_57),
.Y(n_70)
);

NOR2x1_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_50),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_71),
.B(n_45),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_72),
.A2(n_60),
.B1(n_53),
.B2(n_39),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_75),
.A2(n_79),
.B(n_16),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_74),
.A2(n_47),
.B1(n_46),
.B2(n_40),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_76),
.A2(n_84),
.B1(n_20),
.B2(n_22),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_83),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_74),
.A2(n_38),
.B1(n_2),
.B2(n_4),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_1),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_88),
.Y(n_93)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_63),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_73),
.A2(n_2),
.B1(n_4),
.B2(n_6),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_85),
.Y(n_90)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_86),
.Y(n_92)
);

OR2x2_ASAP7_75t_SL g88 ( 
.A(n_66),
.B(n_6),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_64),
.A2(n_7),
.B1(n_8),
.B2(n_13),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_89),
.A2(n_32),
.B1(n_24),
.B2(n_26),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_75),
.A2(n_21),
.B1(n_30),
.B2(n_14),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_91),
.A2(n_102),
.B1(n_83),
.B2(n_27),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_81),
.A2(n_7),
.B(n_8),
.Y(n_94)
);

NOR3xp33_ASAP7_75t_L g104 ( 
.A(n_94),
.B(n_98),
.C(n_23),
.Y(n_104)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_95),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_80),
.Y(n_97)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_97),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_17),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_100),
.B(n_101),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_87),
.B(n_18),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_103),
.B(n_91),
.C(n_94),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_104),
.B(n_105),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_107),
.A2(n_96),
.B1(n_92),
.B2(n_99),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_93),
.C(n_90),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_109),
.B(n_99),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_111),
.B(n_113),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_113),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_115),
.A2(n_110),
.B(n_108),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_116),
.B(n_114),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_112),
.C(n_106),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_118),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_104),
.Y(n_120)
);


endmodule