module fake_jpeg_11034_n_412 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_412);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_412;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx8_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx4f_ASAP7_75t_SL g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_14),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_11),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_4),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_8),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_12),
.Y(n_48)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

BUFx16f_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_55),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_24),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_56),
.B(n_76),
.Y(n_115)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_57),
.Y(n_111)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_58),
.Y(n_122)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

BUFx10_ASAP7_75t_L g120 ( 
.A(n_59),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_60),
.Y(n_131)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_61),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_62),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_37),
.B(n_7),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_63),
.B(n_93),
.Y(n_158)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_64),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_65),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

INVx8_ASAP7_75t_L g138 ( 
.A(n_66),
.Y(n_138)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_67),
.Y(n_126)
);

INVx2_ASAP7_75t_SL g68 ( 
.A(n_20),
.Y(n_68)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_68),
.Y(n_166)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_69),
.Y(n_128)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_20),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_70),
.B(n_79),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

INVx8_ASAP7_75t_L g144 ( 
.A(n_71),
.Y(n_144)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_19),
.Y(n_72)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_72),
.Y(n_143)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_18),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g145 ( 
.A(n_73),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_44),
.B(n_7),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_74),
.B(n_96),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_23),
.Y(n_75)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_75),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_45),
.B(n_9),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_77),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_26),
.Y(n_78)
);

INVx8_ASAP7_75t_L g171 ( 
.A(n_78),
.Y(n_171)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

BUFx10_ASAP7_75t_L g152 ( 
.A(n_80),
.Y(n_152)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_81),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_26),
.Y(n_82)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_82),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_39),
.Y(n_83)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_83),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_39),
.Y(n_84)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_84),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_85),
.Y(n_136)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_21),
.Y(n_86)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_86),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_87),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_20),
.Y(n_88)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_88),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_47),
.B(n_9),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_89),
.B(n_92),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_33),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_90),
.Y(n_169)
);

BUFx8_ASAP7_75t_L g91 ( 
.A(n_24),
.Y(n_91)
);

INVx6_ASAP7_75t_SL g118 ( 
.A(n_91),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_24),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_48),
.B(n_4),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_27),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_94),
.B(n_104),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_30),
.B(n_10),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_95),
.B(n_98),
.Y(n_123)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_17),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_17),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_97),
.B(n_100),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_32),
.B(n_12),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_32),
.B(n_15),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_99),
.B(n_40),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_33),
.Y(n_100)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_35),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_101),
.B(n_102),
.Y(n_173)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_35),
.Y(n_102)
);

INVx11_ASAP7_75t_L g103 ( 
.A(n_24),
.Y(n_103)
);

BUFx2_ASAP7_75t_R g157 ( 
.A(n_103),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_49),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_27),
.B(n_15),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_105),
.B(n_108),
.Y(n_161)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_23),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_106),
.A2(n_40),
.B1(n_52),
.B2(n_49),
.Y(n_119)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_35),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_107),
.B(n_3),
.Y(n_150)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_21),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_34),
.B(n_16),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_51),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_40),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_110),
.B(n_91),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_58),
.A2(n_38),
.B1(n_42),
.B2(n_46),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_112),
.A2(n_163),
.B(n_169),
.Y(n_188)
);

OAI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_65),
.A2(n_38),
.B1(n_42),
.B2(n_46),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_116),
.A2(n_132),
.B1(n_134),
.B2(n_147),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_119),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_124),
.B(n_168),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_109),
.A2(n_34),
.B1(n_50),
.B2(n_52),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_133),
.B(n_139),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_66),
.A2(n_50),
.B1(n_52),
.B2(n_51),
.Y(n_134)
);

OA22x2_ASAP7_75t_L g135 ( 
.A1(n_71),
.A2(n_28),
.B1(n_53),
.B2(n_54),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_135),
.A2(n_119),
.B1(n_112),
.B2(n_163),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_106),
.A2(n_28),
.B1(n_53),
.B2(n_54),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_137),
.A2(n_151),
.B1(n_131),
.B2(n_159),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_90),
.B(n_0),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_107),
.B(n_1),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_142),
.B(n_149),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_78),
.A2(n_2),
.B1(n_3),
.B2(n_83),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_55),
.B(n_2),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_150),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_61),
.A2(n_3),
.B1(n_75),
.B2(n_96),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_60),
.B(n_62),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_153),
.B(n_162),
.Y(n_196)
);

AND2x2_ASAP7_75t_SL g160 ( 
.A(n_68),
.B(n_70),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_160),
.B(n_146),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_75),
.B(n_110),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_103),
.A2(n_87),
.B1(n_82),
.B2(n_84),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_100),
.B(n_88),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_164),
.B(n_165),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_97),
.B(n_85),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_59),
.B(n_80),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_172),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_161),
.B(n_129),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_175),
.B(n_207),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_135),
.A2(n_141),
.B1(n_137),
.B2(n_118),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_177),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_178),
.A2(n_179),
.B1(n_199),
.B2(n_180),
.Y(n_259)
);

OAI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_150),
.A2(n_116),
.B1(n_135),
.B2(n_151),
.Y(n_179)
);

OAI21xp33_ASAP7_75t_L g255 ( 
.A1(n_180),
.A2(n_183),
.B(n_192),
.Y(n_255)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_118),
.Y(n_181)
);

BUFx2_ASAP7_75t_L g236 ( 
.A(n_181),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_115),
.A2(n_125),
.B(n_123),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_182),
.A2(n_205),
.B(n_185),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_160),
.B(n_146),
.Y(n_183)
);

A2O1A1Ixp33_ASAP7_75t_L g184 ( 
.A1(n_160),
.A2(n_130),
.B(n_166),
.C(n_158),
.Y(n_184)
);

A2O1A1Ixp33_ASAP7_75t_L g239 ( 
.A1(n_184),
.A2(n_180),
.B(n_183),
.C(n_187),
.Y(n_239)
);

BUFx10_ASAP7_75t_L g186 ( 
.A(n_120),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_186),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_188),
.B(n_224),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_141),
.A2(n_148),
.B1(n_145),
.B2(n_155),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_190),
.Y(n_269)
);

INVx11_ASAP7_75t_L g191 ( 
.A(n_120),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_191),
.Y(n_254)
);

HAxp5_ASAP7_75t_SL g192 ( 
.A(n_157),
.B(n_120),
.CON(n_192),
.SN(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_128),
.Y(n_193)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_193),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_173),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_194),
.B(n_201),
.Y(n_261)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_143),
.Y(n_197)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_197),
.Y(n_244)
);

OAI22xp33_ASAP7_75t_L g199 ( 
.A1(n_140),
.A2(n_170),
.B1(n_117),
.B2(n_167),
.Y(n_199)
);

CKINVDCx14_ASAP7_75t_R g200 ( 
.A(n_157),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_200),
.B(n_206),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_113),
.B(n_121),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_148),
.A2(n_145),
.B1(n_155),
.B2(n_156),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_202),
.A2(n_221),
.B1(n_229),
.B2(n_176),
.Y(n_246)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_126),
.Y(n_203)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_203),
.Y(n_233)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_114),
.Y(n_204)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_204),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_113),
.B(n_111),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_138),
.B(n_144),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_138),
.B(n_144),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_208),
.B(n_216),
.Y(n_268)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_114),
.Y(n_209)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_209),
.Y(n_242)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_127),
.Y(n_210)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_210),
.Y(n_245)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_127),
.Y(n_211)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_211),
.Y(n_249)
);

CKINVDCx14_ASAP7_75t_R g212 ( 
.A(n_156),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_212),
.B(n_213),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_152),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_136),
.Y(n_214)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_214),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_171),
.B(n_170),
.Y(n_216)
);

AOI21xp33_ASAP7_75t_L g217 ( 
.A1(n_152),
.A2(n_145),
.B(n_111),
.Y(n_217)
);

OR2x2_ASAP7_75t_L g240 ( 
.A(n_217),
.B(n_181),
.Y(n_240)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_131),
.Y(n_218)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_218),
.Y(n_256)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_136),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_219),
.B(n_222),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_171),
.B(n_117),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_220),
.B(n_216),
.Y(n_234)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_154),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_159),
.B(n_122),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_223),
.B(n_225),
.Y(n_253)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_154),
.Y(n_224)
);

OR2x2_ASAP7_75t_L g225 ( 
.A(n_152),
.B(n_122),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_174),
.B(n_115),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_226),
.B(n_228),
.Y(n_257)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_174),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_227),
.B(n_209),
.Y(n_250)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_166),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_174),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_189),
.A2(n_175),
.B1(n_176),
.B2(n_198),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_231),
.A2(n_248),
.B1(n_258),
.B2(n_263),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_234),
.B(n_260),
.Y(n_279)
);

OAI21xp33_ASAP7_75t_L g291 ( 
.A1(n_239),
.A2(n_247),
.B(n_266),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_240),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_246),
.A2(n_267),
.B1(n_236),
.B2(n_264),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_207),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_189),
.A2(n_187),
.B1(n_178),
.B2(n_215),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_250),
.B(n_271),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_252),
.B(n_260),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_188),
.A2(n_195),
.B1(n_225),
.B2(n_208),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_259),
.A2(n_270),
.B1(n_237),
.B2(n_269),
.Y(n_275)
);

OR2x2_ASAP7_75t_L g262 ( 
.A(n_196),
.B(n_184),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_262),
.B(n_272),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_195),
.A2(n_220),
.B1(n_199),
.B2(n_183),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_203),
.B(n_182),
.C(n_210),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_265),
.B(n_238),
.C(n_271),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_186),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_227),
.A2(n_229),
.B1(n_224),
.B2(n_204),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_192),
.A2(n_218),
.B1(n_191),
.B2(n_186),
.Y(n_270)
);

AND2x2_ASAP7_75t_SL g271 ( 
.A(n_186),
.B(n_175),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_205),
.B(n_124),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_240),
.A2(n_238),
.B(n_237),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_273),
.A2(n_283),
.B(n_284),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_261),
.B(n_257),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_274),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_275),
.A2(n_289),
.B1(n_296),
.B2(n_299),
.Y(n_320)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_243),
.Y(n_276)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_276),
.Y(n_316)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_243),
.Y(n_278)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_278),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_279),
.B(n_281),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_280),
.B(n_282),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_247),
.B(n_268),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_244),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_234),
.B(n_271),
.C(n_265),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_284),
.B(n_293),
.Y(n_306)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_244),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_285),
.B(n_288),
.Y(n_312)
);

BUFx12_ASAP7_75t_L g287 ( 
.A(n_236),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_252),
.B(n_262),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_259),
.A2(n_231),
.B1(n_248),
.B2(n_253),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_230),
.B(n_232),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_290),
.B(n_292),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_235),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_268),
.B(n_258),
.C(n_239),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_250),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_294),
.B(n_295),
.Y(n_326)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_256),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_263),
.A2(n_270),
.B1(n_269),
.B2(n_238),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_249),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_297),
.B(n_302),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_255),
.A2(n_266),
.B1(n_256),
.B2(n_249),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_L g313 ( 
.A1(n_301),
.A2(n_267),
.B1(n_250),
.B2(n_264),
.Y(n_313)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_251),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_245),
.Y(n_303)
);

INVx5_ASAP7_75t_L g304 ( 
.A(n_241),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_251),
.B(n_236),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_305),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_300),
.A2(n_254),
.B1(n_241),
.B2(n_242),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_307),
.A2(n_310),
.B1(n_315),
.B2(n_297),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_300),
.A2(n_242),
.B1(n_233),
.B2(n_245),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_313),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_281),
.A2(n_233),
.B1(n_286),
.B2(n_293),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_287),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_317),
.B(n_294),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_277),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_319),
.B(n_322),
.Y(n_331)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_277),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_273),
.A2(n_286),
.B(n_283),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_323),
.A2(n_278),
.B(n_282),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_324),
.B(n_291),
.Y(n_330)
);

CKINVDCx16_ASAP7_75t_R g327 ( 
.A(n_277),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_327),
.B(n_285),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_328),
.B(n_332),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_308),
.B(n_279),
.Y(n_329)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_329),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_330),
.B(n_335),
.C(n_341),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_309),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_320),
.A2(n_280),
.B1(n_298),
.B2(n_292),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_333),
.A2(n_344),
.B1(n_307),
.B2(n_310),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_SL g334 ( 
.A(n_325),
.B(n_302),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_SL g348 ( 
.A(n_334),
.B(n_339),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_324),
.B(n_276),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_SL g357 ( 
.A1(n_336),
.A2(n_342),
.B(n_326),
.Y(n_357)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_316),
.Y(n_337)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_337),
.Y(n_351)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_338),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_311),
.B(n_325),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g353 ( 
.A(n_340),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_306),
.B(n_295),
.C(n_303),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_326),
.B(n_304),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_309),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_343),
.B(n_314),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_320),
.A2(n_287),
.B1(n_311),
.B2(n_313),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_312),
.B(n_287),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_SL g361 ( 
.A(n_346),
.B(n_312),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_306),
.B(n_323),
.C(n_327),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_347),
.B(n_323),
.C(n_315),
.Y(n_356)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_350),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_342),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_355),
.B(n_360),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_356),
.B(n_363),
.C(n_343),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_357),
.A2(n_361),
.B(n_331),
.Y(n_365)
);

AND2x6_ASAP7_75t_L g359 ( 
.A(n_330),
.B(n_320),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_SL g364 ( 
.A1(n_359),
.A2(n_345),
.B(n_336),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_342),
.Y(n_360)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_362),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_335),
.B(n_322),
.C(n_319),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_364),
.A2(n_374),
.B(n_357),
.Y(n_377)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_365),
.Y(n_384)
);

INVx3_ASAP7_75t_L g366 ( 
.A(n_358),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_366),
.B(n_369),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_358),
.A2(n_344),
.B1(n_333),
.B2(n_345),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_368),
.A2(n_376),
.B1(n_362),
.B2(n_353),
.Y(n_382)
);

INVx1_ASAP7_75t_SL g369 ( 
.A(n_351),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_SL g370 ( 
.A(n_363),
.B(n_347),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_SL g378 ( 
.A(n_370),
.B(n_352),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_352),
.B(n_341),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_371),
.B(n_373),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_354),
.A2(n_338),
.B(n_332),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_355),
.A2(n_360),
.B1(n_354),
.B2(n_349),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g387 ( 
.A1(n_377),
.A2(n_375),
.B(n_368),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_378),
.B(n_348),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_376),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_379),
.A2(n_381),
.B1(n_386),
.B2(n_337),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_371),
.B(n_373),
.C(n_370),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_380),
.B(n_329),
.C(n_308),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_367),
.A2(n_366),
.B1(n_349),
.B2(n_372),
.Y(n_381)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_382),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_369),
.A2(n_359),
.B1(n_356),
.B2(n_310),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_387),
.A2(n_381),
.B(n_384),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_389),
.B(n_392),
.Y(n_397)
);

OAI21xp33_ASAP7_75t_L g390 ( 
.A1(n_377),
.A2(n_314),
.B(n_351),
.Y(n_390)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_390),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_391),
.A2(n_316),
.B1(n_318),
.B2(n_317),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_383),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_393),
.B(n_321),
.Y(n_398)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_394),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_SL g396 ( 
.A1(n_389),
.A2(n_380),
.B(n_386),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_396),
.A2(n_392),
.B(n_385),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_398),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_399),
.B(n_388),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_400),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_403),
.B(n_394),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_405),
.B(n_406),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_402),
.B(n_397),
.C(n_385),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g408 ( 
.A1(n_404),
.A2(n_401),
.B(n_395),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_408),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_409),
.B(n_407),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_410),
.B(n_405),
.C(n_399),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_411),
.B(n_378),
.Y(n_412)
);


endmodule