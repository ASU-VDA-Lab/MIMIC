module fake_jpeg_9366_n_115 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_115);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_115;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_9),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

BUFx4f_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx4f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_26),
.B(n_28),
.Y(n_48)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_0),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_32),
.Y(n_41)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_20),
.B(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_19),
.B(n_1),
.Y(n_34)
);

OAI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_34),
.A2(n_19),
.B1(n_24),
.B2(n_12),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_40),
.B(n_33),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

OA22x2_ASAP7_75t_L g44 ( 
.A1(n_30),
.A2(n_18),
.B1(n_13),
.B2(n_23),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_23),
.C(n_18),
.Y(n_64)
);

NOR2x1_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_12),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_49),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_27),
.A2(n_22),
.B1(n_25),
.B2(n_17),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_31),
.A2(n_22),
.B1(n_25),
.B2(n_17),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_51),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_36),
.A2(n_24),
.B1(n_15),
.B2(n_23),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_52),
.B(n_53),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_45),
.B(n_26),
.Y(n_53)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

AND2x6_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_1),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_57),
.A2(n_46),
.B1(n_47),
.B2(n_42),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_29),
.Y(n_59)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_15),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_65),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_64),
.A2(n_46),
.B1(n_47),
.B2(n_44),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_66),
.B(n_13),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_68),
.A2(n_73),
.B1(n_58),
.B2(n_56),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_64),
.B(n_41),
.C(n_42),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_75),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_62),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_1),
.Y(n_75)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

INVxp67_ASAP7_75t_SL g94 ( 
.A(n_80),
.Y(n_94)
);

CKINVDCx5p33_ASAP7_75t_R g81 ( 
.A(n_67),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_81),
.Y(n_96)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

INVxp33_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_83),
.B(n_84),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_54),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_62),
.Y(n_85)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_85),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_86),
.Y(n_93)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_87),
.A2(n_88),
.B1(n_57),
.B2(n_77),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_79),
.B(n_72),
.C(n_76),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_89),
.B(n_84),
.C(n_79),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_95),
.A2(n_55),
.B1(n_58),
.B2(n_71),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_96),
.B(n_81),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_97),
.A2(n_98),
.B(n_67),
.Y(n_105)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_92),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_99),
.B(n_92),
.Y(n_102)
);

A2O1A1Ixp33_ASAP7_75t_SL g100 ( 
.A1(n_93),
.A2(n_83),
.B(n_85),
.C(n_74),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_100),
.A2(n_93),
.B1(n_95),
.B2(n_91),
.Y(n_103)
);

AOI321xp33_ASAP7_75t_L g104 ( 
.A1(n_101),
.A2(n_91),
.A3(n_96),
.B1(n_90),
.B2(n_94),
.C(n_89),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_102),
.B(n_2),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_103),
.A2(n_104),
.B1(n_105),
.B2(n_38),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_102),
.A2(n_100),
.B1(n_78),
.B2(n_65),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_106),
.A2(n_38),
.B1(n_3),
.B2(n_5),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_107),
.B(n_108),
.Y(n_109)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_110),
.Y(n_112)
);

AOI322xp5_ASAP7_75t_L g111 ( 
.A1(n_109),
.A2(n_106),
.A3(n_7),
.B1(n_8),
.B2(n_11),
.C1(n_4),
.C2(n_38),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_111),
.B(n_110),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_113),
.A2(n_112),
.B1(n_8),
.B2(n_4),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_38),
.Y(n_115)
);


endmodule