module fake_jpeg_10815_n_33 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_33);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_33;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx3_ASAP7_75t_L g7 ( 
.A(n_6),
.Y(n_7)
);

INVx2_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

BUFx3_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

NOR2x1_ASAP7_75t_L g13 ( 
.A(n_12),
.B(n_0),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_13),
.B(n_15),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_8),
.B(n_0),
.Y(n_14)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_14),
.B(n_5),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_9),
.B(n_0),
.Y(n_15)
);

INVx4_ASAP7_75t_SL g16 ( 
.A(n_8),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_SL g22 ( 
.A1(n_16),
.A2(n_18),
.B(n_5),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_SL g17 ( 
.A1(n_7),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_17),
.A2(n_10),
.B1(n_11),
.B2(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_19),
.A2(n_18),
.B1(n_13),
.B2(n_16),
.Y(n_26)
);

MAJx2_ASAP7_75t_L g20 ( 
.A(n_14),
.B(n_10),
.C(n_4),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_20),
.B(n_21),
.C(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_22),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_21),
.B(n_23),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_26),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_27),
.B(n_20),
.Y(n_28)
);

AO21x1_ASAP7_75t_L g31 ( 
.A1(n_28),
.A2(n_25),
.B(n_27),
.Y(n_31)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_29),
.B(n_16),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_31),
.A2(n_32),
.B1(n_30),
.B2(n_24),
.Y(n_33)
);


endmodule