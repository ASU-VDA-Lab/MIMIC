module fake_jpeg_12627_n_563 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_563);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_563;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVxp33_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_18),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_14),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_6),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_18),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_7),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

INVxp33_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_53),
.Y(n_109)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_54),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_55),
.Y(n_108)
);

INVx6_ASAP7_75t_SL g56 ( 
.A(n_24),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_56),
.Y(n_159)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_57),
.Y(n_133)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_58),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_59),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_60),
.Y(n_114)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_61),
.Y(n_157)
);

INVx3_ASAP7_75t_SL g62 ( 
.A(n_24),
.Y(n_62)
);

BUFx8_ASAP7_75t_L g125 ( 
.A(n_62),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_63),
.Y(n_118)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_64),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_29),
.B(n_0),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_65),
.B(n_91),
.Y(n_112)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_66),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_67),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_68),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_69),
.Y(n_107)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_70),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_71),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_27),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g168 ( 
.A(n_72),
.Y(n_168)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_19),
.Y(n_73)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_73),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_27),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_74),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_75),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_19),
.B(n_0),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_76),
.B(n_97),
.Y(n_129)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_77),
.Y(n_167)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_24),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_78),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

INVx8_ASAP7_75t_L g170 ( 
.A(n_79),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_80),
.Y(n_141)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_24),
.Y(n_81)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_81),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_28),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_82),
.B(n_83),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_28),
.B(n_0),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_84),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_85),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_86),
.Y(n_128)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_87),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_88),
.Y(n_130)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_19),
.Y(n_89)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_89),
.Y(n_131)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_35),
.Y(n_90)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_90),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_20),
.B(n_17),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_44),
.Y(n_92)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_92),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_30),
.Y(n_93)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_52),
.B(n_0),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_94),
.B(n_105),
.Y(n_149)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_35),
.Y(n_95)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_95),
.Y(n_124)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_30),
.Y(n_96)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_96),
.Y(n_169)
);

INVx5_ASAP7_75t_SL g97 ( 
.A(n_26),
.Y(n_97)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_35),
.Y(n_98)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_98),
.Y(n_166)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_35),
.Y(n_99)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_99),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_47),
.Y(n_100)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_100),
.Y(n_145)
);

INVx6_ASAP7_75t_SL g101 ( 
.A(n_22),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_101),
.B(n_104),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_47),
.Y(n_102)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_102),
.Y(n_150)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_21),
.Y(n_103)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_103),
.Y(n_154)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_47),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_29),
.B(n_1),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_21),
.Y(n_106)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_106),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_41),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_117),
.B(n_122),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_83),
.B(n_41),
.Y(n_122)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_82),
.Y(n_136)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_136),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_76),
.B(n_46),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_138),
.B(n_139),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_61),
.B(n_31),
.Y(n_139)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_66),
.Y(n_142)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_142),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_54),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_144),
.B(n_148),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_70),
.B(n_46),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_146),
.B(n_153),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_58),
.A2(n_21),
.B1(n_25),
.B2(n_51),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_147),
.A2(n_161),
.B1(n_93),
.B2(n_77),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_62),
.B(n_31),
.C(n_50),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_55),
.B(n_50),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_64),
.A2(n_25),
.B1(n_51),
.B2(n_47),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_104),
.Y(n_163)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_163),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_60),
.B(n_39),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_164),
.B(n_48),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_59),
.A2(n_25),
.B1(n_49),
.B2(n_38),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_165),
.A2(n_39),
.B1(n_38),
.B2(n_49),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_134),
.A2(n_72),
.B1(n_74),
.B2(n_28),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_171),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_129),
.A2(n_79),
.B1(n_80),
.B2(n_84),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_173),
.A2(n_191),
.B1(n_221),
.B2(n_222),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_111),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_174),
.B(n_194),
.Y(n_236)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_130),
.Y(n_175)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_175),
.Y(n_234)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_137),
.Y(n_176)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_176),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_108),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_177),
.Y(n_274)
);

NAND2xp33_ASAP7_75t_SL g178 ( 
.A(n_129),
.B(n_78),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_178),
.A2(n_184),
.B(n_219),
.Y(n_248)
);

INVx6_ASAP7_75t_L g180 ( 
.A(n_108),
.Y(n_180)
);

INVx6_ASAP7_75t_L g246 ( 
.A(n_180),
.Y(n_246)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_145),
.Y(n_181)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_181),
.Y(n_268)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_125),
.Y(n_183)
);

INVx4_ASAP7_75t_L g271 ( 
.A(n_183),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_110),
.B(n_60),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_111),
.Y(n_185)
);

NAND3xp33_ASAP7_75t_L g281 ( 
.A(n_185),
.B(n_213),
.C(n_3),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_124),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_187),
.Y(n_284)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_150),
.Y(n_188)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_188),
.Y(n_277)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_113),
.Y(n_189)
);

INVx6_ASAP7_75t_L g247 ( 
.A(n_189),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_190),
.A2(n_230),
.B1(n_109),
.B2(n_143),
.Y(n_275)
);

INVx5_ASAP7_75t_L g192 ( 
.A(n_168),
.Y(n_192)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_192),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_112),
.A2(n_71),
.B1(n_102),
.B2(n_100),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_193),
.A2(n_198),
.B1(n_228),
.B2(n_126),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_115),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_156),
.Y(n_195)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_195),
.Y(n_286)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_135),
.Y(n_197)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_197),
.Y(n_233)
);

O2A1O1Ixp33_ASAP7_75t_L g198 ( 
.A1(n_152),
.A2(n_34),
.B(n_48),
.C(n_45),
.Y(n_198)
);

OAI32xp33_ASAP7_75t_L g199 ( 
.A1(n_149),
.A2(n_81),
.A3(n_92),
.B1(n_88),
.B2(n_86),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_199),
.B(n_223),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_159),
.B(n_104),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_200),
.B(n_217),
.Y(n_287)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_154),
.Y(n_201)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_201),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_113),
.Y(n_202)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_202),
.Y(n_262)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_132),
.Y(n_204)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_204),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_169),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_205),
.Y(n_257)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_125),
.Y(n_206)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_206),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_140),
.A2(n_48),
.B1(n_34),
.B2(n_36),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_207),
.Y(n_260)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_127),
.Y(n_208)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_208),
.Y(n_261)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_168),
.Y(n_209)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_209),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_121),
.A2(n_85),
.B1(n_75),
.B2(n_69),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_210),
.A2(n_123),
.B1(n_118),
.B2(n_143),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_140),
.A2(n_43),
.B1(n_34),
.B2(n_36),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_211),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_168),
.Y(n_212)
);

BUFx4f_ASAP7_75t_SL g250 ( 
.A(n_212),
.Y(n_250)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_121),
.Y(n_215)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_215),
.Y(n_269)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_131),
.Y(n_216)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_216),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_133),
.B(n_45),
.Y(n_217)
);

INVx8_ASAP7_75t_L g218 ( 
.A(n_167),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_218),
.Y(n_283)
);

AO22x1_ASAP7_75t_L g219 ( 
.A1(n_152),
.A2(n_45),
.B1(n_43),
.B2(n_36),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_114),
.Y(n_220)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_220),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_116),
.A2(n_43),
.B1(n_51),
.B2(n_63),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_L g222 ( 
.A1(n_170),
.A2(n_68),
.B1(n_67),
.B2(n_51),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g223 ( 
.A(n_120),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_157),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_224),
.B(n_225),
.Y(n_259)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_160),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_166),
.B(n_1),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_226),
.B(n_3),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_125),
.B(n_1),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_227),
.B(n_178),
.Y(n_245)
);

OAI22xp33_ASAP7_75t_L g228 ( 
.A1(n_147),
.A2(n_42),
.B1(n_33),
.B2(n_22),
.Y(n_228)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_167),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_229),
.B(n_231),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_109),
.A2(n_42),
.B1(n_33),
.B2(n_22),
.Y(n_230)
);

AOI32xp33_ASAP7_75t_L g231 ( 
.A1(n_109),
.A2(n_42),
.A3(n_33),
.B1(n_22),
.B2(n_6),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_119),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_232),
.B(n_155),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_214),
.B(n_119),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_239),
.B(n_241),
.Y(n_313)
);

AOI22x1_ASAP7_75t_SL g240 ( 
.A1(n_199),
.A2(n_161),
.B1(n_114),
.B2(n_141),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_240),
.A2(n_220),
.B(n_42),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_196),
.B(n_128),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_L g243 ( 
.A1(n_191),
.A2(n_170),
.B1(n_128),
.B2(n_158),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_243),
.A2(n_266),
.B1(n_273),
.B2(n_275),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_227),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_244),
.B(n_270),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_245),
.B(n_42),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_251),
.A2(n_258),
.B1(n_198),
.B2(n_202),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_253),
.B(n_228),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_203),
.B(n_162),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_256),
.B(n_185),
.C(n_183),
.Y(n_291)
);

OAI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_210),
.A2(n_155),
.B1(n_141),
.B2(n_123),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_264),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_265),
.B(n_279),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_L g266 ( 
.A1(n_184),
.A2(n_158),
.B1(n_151),
.B2(n_107),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_227),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_179),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_272),
.B(n_276),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_L g273 ( 
.A1(n_184),
.A2(n_151),
.B1(n_107),
.B2(n_118),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_204),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_186),
.B(n_3),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_281),
.B(n_206),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_195),
.B(n_201),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_282),
.B(n_232),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g363 ( 
.A1(n_288),
.A2(n_321),
.B(n_277),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_274),
.Y(n_290)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_290),
.Y(n_352)
);

XNOR2x1_ASAP7_75t_L g357 ( 
.A(n_291),
.B(n_298),
.Y(n_357)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_282),
.Y(n_292)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_292),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_238),
.A2(n_215),
.B1(n_229),
.B2(n_218),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_293),
.A2(n_294),
.B1(n_299),
.B2(n_308),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_263),
.A2(n_175),
.B1(n_176),
.B2(n_181),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_236),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_295),
.B(n_304),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_256),
.B(n_172),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_240),
.A2(n_188),
.B1(n_180),
.B2(n_189),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_261),
.Y(n_300)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_300),
.Y(n_355)
);

OAI21xp33_ASAP7_75t_SL g301 ( 
.A1(n_260),
.A2(n_223),
.B(n_219),
.Y(n_301)
);

NOR2x1_ASAP7_75t_R g370 ( 
.A(n_301),
.B(n_234),
.Y(n_370)
);

HB1xp67_ASAP7_75t_L g302 ( 
.A(n_254),
.Y(n_302)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_302),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_303),
.B(n_306),
.Y(n_344)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_269),
.Y(n_305)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_305),
.Y(n_371)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_259),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_239),
.B(n_182),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_307),
.B(n_311),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_253),
.A2(n_275),
.B1(n_244),
.B2(n_270),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_261),
.Y(n_309)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_309),
.Y(n_374)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_278),
.Y(n_310)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_310),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_287),
.B(n_225),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_312),
.A2(n_317),
.B1(n_289),
.B2(n_292),
.Y(n_346)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_278),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_314),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_241),
.A2(n_280),
.B1(n_260),
.B2(n_237),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_315),
.A2(n_332),
.B1(n_335),
.B2(n_251),
.Y(n_356)
);

AO22x2_ASAP7_75t_L g318 ( 
.A1(n_242),
.A2(n_177),
.B1(n_209),
.B2(n_192),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_318),
.B(n_320),
.Y(n_343)
);

AND2x4_ASAP7_75t_L g319 ( 
.A(n_248),
.B(n_212),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g378 ( 
.A1(n_319),
.A2(n_333),
.B(n_9),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_254),
.Y(n_320)
);

INVx3_ASAP7_75t_L g322 ( 
.A(n_262),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_SL g342 ( 
.A1(n_322),
.A2(n_271),
.B1(n_262),
.B2(n_252),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_272),
.B(n_4),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_323),
.B(n_324),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_285),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_325),
.B(n_8),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_233),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_326),
.B(n_328),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_245),
.B(n_33),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_327),
.B(n_336),
.C(n_257),
.Y(n_351)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_269),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_249),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_329),
.B(n_331),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_233),
.B(n_4),
.Y(n_330)
);

INVxp33_ASAP7_75t_L g349 ( 
.A(n_330),
.Y(n_349)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_249),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_280),
.A2(n_33),
.B1(n_22),
.B2(n_7),
.Y(n_332)
);

O2A1O1Ixp33_ASAP7_75t_L g333 ( 
.A1(n_237),
.A2(n_5),
.B(n_6),
.C(n_8),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_284),
.B(n_5),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_334),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_248),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_235),
.B(n_5),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_235),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_337),
.B(n_286),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_298),
.B(n_267),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_338),
.B(n_339),
.C(n_362),
.Y(n_405)
);

MAJx2_ASAP7_75t_L g339 ( 
.A(n_313),
.B(n_267),
.C(n_285),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_342),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_346),
.A2(n_376),
.B1(n_322),
.B2(n_324),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_321),
.A2(n_271),
.B(n_252),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_SL g394 ( 
.A1(n_347),
.A2(n_353),
.B(n_370),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_351),
.B(n_368),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_288),
.A2(n_283),
.B(n_257),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_356),
.A2(n_364),
.B1(n_377),
.B2(n_296),
.Y(n_388)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_359),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_313),
.B(n_283),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_360),
.B(n_379),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_325),
.B(n_286),
.C(n_277),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_363),
.B(n_378),
.Y(n_404)
);

AOI22xp33_ASAP7_75t_SL g364 ( 
.A1(n_315),
.A2(n_247),
.B1(n_246),
.B2(n_274),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_327),
.B(n_250),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_SL g408 ( 
.A(n_365),
.B(n_373),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_SL g367 ( 
.A1(n_288),
.A2(n_268),
.B(n_255),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_L g412 ( 
.A1(n_367),
.A2(n_380),
.B(n_337),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_291),
.B(n_268),
.C(n_255),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_308),
.B(n_234),
.C(n_250),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_372),
.B(n_375),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_294),
.B(n_250),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_312),
.A2(n_247),
.B1(n_246),
.B2(n_11),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_299),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_377)
);

OAI32xp33_ASAP7_75t_L g379 ( 
.A1(n_293),
.A2(n_12),
.A3(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_L g380 ( 
.A1(n_319),
.A2(n_13),
.B(n_15),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_343),
.A2(n_318),
.B1(n_317),
.B2(n_295),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_383),
.A2(n_388),
.B1(n_397),
.B2(n_398),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_357),
.B(n_338),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_384),
.B(n_389),
.C(n_362),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_341),
.B(n_326),
.Y(n_386)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_386),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_357),
.B(n_319),
.Y(n_389)
);

CKINVDCx14_ASAP7_75t_R g390 ( 
.A(n_341),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_390),
.B(n_402),
.Y(n_446)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_354),
.Y(n_391)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_391),
.Y(n_421)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_358),
.Y(n_392)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_392),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_372),
.A2(n_316),
.B1(n_319),
.B2(n_318),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_393),
.A2(n_409),
.B1(n_410),
.B2(n_345),
.Y(n_428)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_354),
.Y(n_395)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_395),
.Y(n_432)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_358),
.Y(n_396)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_396),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_343),
.A2(n_318),
.B1(n_309),
.B2(n_314),
.Y(n_397)
);

OAI22xp33_ASAP7_75t_SL g398 ( 
.A1(n_345),
.A2(n_318),
.B1(n_333),
.B2(n_320),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_360),
.B(n_310),
.Y(n_399)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_399),
.Y(n_435)
);

INVx1_ASAP7_75t_SL g400 ( 
.A(n_374),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_400),
.B(n_406),
.Y(n_426)
);

INVx8_ASAP7_75t_L g401 ( 
.A(n_349),
.Y(n_401)
);

BUFx2_ASAP7_75t_L g439 ( 
.A(n_401),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_359),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_374),
.Y(n_403)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_403),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_340),
.B(n_300),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_376),
.A2(n_328),
.B1(n_331),
.B2(n_329),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_SL g411 ( 
.A(n_348),
.B(n_297),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_SL g443 ( 
.A(n_411),
.B(n_415),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_412),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_378),
.A2(n_305),
.B(n_290),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_413),
.B(n_417),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_366),
.B(n_336),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_381),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_416),
.B(n_418),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_350),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_381),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_387),
.B(n_365),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_420),
.B(n_427),
.Y(n_463)
);

INVx3_ASAP7_75t_L g422 ( 
.A(n_401),
.Y(n_422)
);

INVx3_ASAP7_75t_L g467 ( 
.A(n_422),
.Y(n_467)
);

XOR2x2_ASAP7_75t_L g423 ( 
.A(n_408),
.B(n_368),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_423),
.B(n_394),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_SL g424 ( 
.A(n_384),
.B(n_351),
.Y(n_424)
);

XNOR2x1_ASAP7_75t_L g465 ( 
.A(n_424),
.B(n_425),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_387),
.B(n_405),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_428),
.A2(n_404),
.B1(n_382),
.B2(n_385),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_383),
.A2(n_370),
.B1(n_363),
.B2(n_347),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_429),
.A2(n_442),
.B1(n_413),
.B2(n_410),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_L g431 ( 
.A1(n_409),
.A2(n_356),
.B1(n_344),
.B2(n_377),
.Y(n_431)
);

BUFx2_ASAP7_75t_L g461 ( 
.A(n_431),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_408),
.B(n_339),
.C(n_375),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_434),
.B(n_436),
.C(n_438),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_405),
.B(n_373),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_389),
.B(n_361),
.C(n_353),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_397),
.A2(n_369),
.B1(n_355),
.B2(n_350),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_386),
.B(n_369),
.Y(n_444)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_444),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_SL g445 ( 
.A(n_407),
.B(n_361),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_445),
.B(n_449),
.Y(n_454)
);

MAJx2_ASAP7_75t_L g449 ( 
.A(n_407),
.B(n_367),
.C(n_371),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_396),
.B(n_371),
.C(n_380),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_450),
.B(n_412),
.C(n_404),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_444),
.B(n_399),
.Y(n_452)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_452),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_455),
.B(n_457),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_427),
.B(n_395),
.C(n_391),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_456),
.B(n_458),
.C(n_475),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_436),
.B(n_382),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_420),
.B(n_385),
.C(n_393),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_426),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_459),
.B(n_460),
.Y(n_484)
);

HB1xp67_ASAP7_75t_L g460 ( 
.A(n_422),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_462),
.A2(n_477),
.B1(n_429),
.B2(n_442),
.Y(n_480)
);

BUFx2_ASAP7_75t_L g464 ( 
.A(n_441),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_464),
.B(n_466),
.Y(n_485)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_426),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_443),
.B(n_406),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_468),
.B(n_470),
.Y(n_498)
);

OAI21xp5_ASAP7_75t_SL g479 ( 
.A1(n_469),
.A2(n_473),
.B(n_434),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_446),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_440),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g486 ( 
.A(n_471),
.Y(n_486)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_440),
.Y(n_472)
);

AOI21x1_ASAP7_75t_L g482 ( 
.A1(n_472),
.A2(n_478),
.B(n_421),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_448),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_L g474 ( 
.A1(n_447),
.A2(n_394),
.B(n_404),
.Y(n_474)
);

AO21x1_ASAP7_75t_L g490 ( 
.A1(n_474),
.A2(n_449),
.B(n_445),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_425),
.B(n_400),
.C(n_418),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_476),
.A2(n_438),
.B1(n_450),
.B2(n_414),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_419),
.A2(n_414),
.B1(n_416),
.B2(n_403),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_437),
.Y(n_478)
);

HB1xp67_ASAP7_75t_L g506 ( 
.A(n_479),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_480),
.A2(n_493),
.B1(n_496),
.B2(n_461),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_464),
.A2(n_435),
.B1(n_447),
.B2(n_432),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_SL g507 ( 
.A1(n_481),
.A2(n_488),
.B1(n_499),
.B2(n_477),
.Y(n_507)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_482),
.Y(n_503)
);

O2A1O1Ixp33_ASAP7_75t_L g487 ( 
.A1(n_451),
.A2(n_433),
.B(n_441),
.C(n_430),
.Y(n_487)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_487),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_475),
.B(n_423),
.C(n_424),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_489),
.B(n_501),
.C(n_465),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_490),
.B(n_491),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_463),
.B(n_439),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_462),
.A2(n_439),
.B1(n_379),
.B2(n_352),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_456),
.B(n_352),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_495),
.B(n_497),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_461),
.A2(n_290),
.B1(n_16),
.B2(n_17),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_457),
.B(n_15),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_476),
.A2(n_16),
.B1(n_17),
.B2(n_455),
.Y(n_499)
);

AOI21xp5_ASAP7_75t_L g500 ( 
.A1(n_474),
.A2(n_16),
.B(n_17),
.Y(n_500)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_500),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_458),
.B(n_463),
.Y(n_501)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_487),
.Y(n_504)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_504),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_507),
.A2(n_519),
.B1(n_480),
.B2(n_493),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g525 ( 
.A(n_508),
.B(n_489),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_486),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_509),
.B(n_511),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_495),
.B(n_453),
.C(n_465),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_491),
.B(n_453),
.C(n_454),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_512),
.B(n_514),
.Y(n_523)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_513),
.Y(n_527)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_484),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_485),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_515),
.B(n_496),
.Y(n_534)
);

CKINVDCx14_ASAP7_75t_R g517 ( 
.A(n_498),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_517),
.B(n_518),
.Y(n_528)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_481),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_SL g519 ( 
.A1(n_488),
.A2(n_452),
.B1(n_467),
.B2(n_454),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_SL g540 ( 
.A1(n_520),
.A2(n_499),
.B1(n_503),
.B2(n_505),
.Y(n_540)
);

XOR2xp5_ASAP7_75t_L g521 ( 
.A(n_516),
.B(n_501),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_521),
.B(n_525),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_502),
.Y(n_524)
);

INVx11_ASAP7_75t_L g545 ( 
.A(n_524),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_514),
.B(n_467),
.Y(n_529)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_529),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_519),
.B(n_494),
.Y(n_530)
);

MAJx2_ASAP7_75t_L g536 ( 
.A(n_530),
.B(n_507),
.C(n_512),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_511),
.B(n_483),
.C(n_494),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_531),
.B(n_533),
.C(n_508),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_506),
.B(n_492),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_532),
.A2(n_534),
.B1(n_515),
.B2(n_502),
.Y(n_535)
);

XOR2xp5_ASAP7_75t_L g533 ( 
.A(n_516),
.B(n_483),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_535),
.B(n_537),
.Y(n_552)
);

OAI21x1_ASAP7_75t_L g548 ( 
.A1(n_536),
.A2(n_524),
.B(n_520),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_531),
.B(n_533),
.C(n_522),
.Y(n_538)
);

AOI21xp5_ASAP7_75t_L g547 ( 
.A1(n_538),
.A2(n_539),
.B(n_542),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_530),
.B(n_513),
.C(n_490),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_540),
.B(n_527),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_521),
.B(n_510),
.C(n_497),
.Y(n_542)
);

INVxp67_ASAP7_75t_L g544 ( 
.A(n_523),
.Y(n_544)
);

NAND2xp33_ASAP7_75t_SL g546 ( 
.A(n_544),
.B(n_528),
.Y(n_546)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_546),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_548),
.Y(n_554)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_549),
.Y(n_556)
);

OAI22xp5_ASAP7_75t_SL g550 ( 
.A1(n_544),
.A2(n_526),
.B1(n_505),
.B2(n_500),
.Y(n_550)
);

HB1xp67_ASAP7_75t_L g555 ( 
.A(n_550),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_538),
.B(n_543),
.Y(n_551)
);

OAI21xp33_ASAP7_75t_SL g557 ( 
.A1(n_554),
.A2(n_545),
.B(n_552),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_557),
.B(n_558),
.C(n_555),
.Y(n_559)
);

O2A1O1Ixp33_ASAP7_75t_SL g558 ( 
.A1(n_553),
.A2(n_545),
.B(n_546),
.C(n_551),
.Y(n_558)
);

OA21x2_ASAP7_75t_L g560 ( 
.A1(n_559),
.A2(n_556),
.B(n_541),
.Y(n_560)
);

XNOR2xp5_ASAP7_75t_L g561 ( 
.A(n_560),
.B(n_547),
.Y(n_561)
);

OAI31xp33_ASAP7_75t_SL g562 ( 
.A1(n_561),
.A2(n_537),
.A3(n_536),
.B(n_525),
.Y(n_562)
);

OAI21xp5_ASAP7_75t_L g563 ( 
.A1(n_562),
.A2(n_539),
.B(n_542),
.Y(n_563)
);


endmodule