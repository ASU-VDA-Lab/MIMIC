module fake_jpeg_5110_n_331 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_331);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_331;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx2_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx4f_ASAP7_75t_SL g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_22),
.B(n_16),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_35),
.B(n_43),
.Y(n_62)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

HB1xp67_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_22),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_44),
.Y(n_50)
);

INVx6_ASAP7_75t_SL g38 ( 
.A(n_21),
.Y(n_38)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_42),
.A2(n_19),
.B1(n_33),
.B2(n_27),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_22),
.B(n_19),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_22),
.B(n_0),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_42),
.A2(n_22),
.B1(n_19),
.B2(n_18),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_35),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_47),
.B(n_69),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_33),
.C(n_21),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_48),
.B(n_51),
.C(n_56),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_33),
.C(n_21),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_37),
.B(n_17),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_52),
.B(n_54),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_53),
.A2(n_60),
.B1(n_66),
.B2(n_70),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_37),
.B(n_17),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_37),
.A2(n_19),
.B1(n_27),
.B2(n_30),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_55),
.A2(n_64),
.B1(n_34),
.B2(n_31),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_33),
.C(n_21),
.Y(n_56)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_42),
.A2(n_36),
.B1(n_32),
.B2(n_28),
.Y(n_60)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_63),
.B(n_68),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_40),
.A2(n_27),
.B1(n_21),
.B2(n_32),
.Y(n_64)
);

OR2x4_ASAP7_75t_SL g65 ( 
.A(n_38),
.B(n_27),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_65),
.A2(n_61),
.B1(n_67),
.B2(n_59),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_42),
.A2(n_28),
.B1(n_32),
.B2(n_17),
.Y(n_66)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_44),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_42),
.A2(n_28),
.B1(n_17),
.B2(n_34),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_36),
.A2(n_34),
.B1(n_18),
.B2(n_30),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_71),
.A2(n_23),
.B1(n_31),
.B2(n_30),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_69),
.A2(n_41),
.B1(n_40),
.B2(n_36),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_73),
.A2(n_83),
.B1(n_84),
.B2(n_72),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_41),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_74),
.B(n_45),
.Y(n_120)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_75),
.B(n_86),
.Y(n_113)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_76),
.B(n_90),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_54),
.B(n_34),
.Y(n_78)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_78),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_79),
.A2(n_82),
.B1(n_91),
.B2(n_67),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_47),
.B(n_24),
.Y(n_80)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_80),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_55),
.A2(n_41),
.B1(n_40),
.B2(n_38),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_68),
.A2(n_20),
.B1(n_29),
.B2(n_24),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_63),
.B(n_62),
.Y(n_85)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_85),
.Y(n_114)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

INVx2_ASAP7_75t_SL g87 ( 
.A(n_65),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_87),
.B(n_39),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_62),
.B(n_24),
.Y(n_89)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_89),
.Y(n_116)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_46),
.A2(n_31),
.B1(n_29),
.B2(n_20),
.Y(n_91)
);

A2O1A1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_94),
.A2(n_53),
.B(n_58),
.C(n_51),
.Y(n_110)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_95),
.B(n_67),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_65),
.A2(n_18),
.B1(n_29),
.B2(n_23),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_96),
.A2(n_99),
.B1(n_25),
.B2(n_16),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_50),
.B(n_23),
.Y(n_98)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_61),
.A2(n_20),
.B1(n_25),
.B2(n_39),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_73),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_101),
.B(n_128),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_97),
.B(n_74),
.C(n_56),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_103),
.B(n_115),
.C(n_94),
.Y(n_155)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_105),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_106),
.A2(n_111),
.B1(n_112),
.B2(n_118),
.Y(n_138)
);

AO32x1_ASAP7_75t_L g107 ( 
.A1(n_87),
.A2(n_96),
.A3(n_85),
.B1(n_86),
.B2(n_75),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_107),
.B(n_117),
.Y(n_151)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_77),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_109),
.A2(n_122),
.B1(n_75),
.B2(n_87),
.Y(n_152)
);

AOI221xp5_ASAP7_75t_L g132 ( 
.A1(n_110),
.A2(n_107),
.B1(n_121),
.B2(n_112),
.C(n_113),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_95),
.A2(n_48),
.B1(n_72),
.B2(n_60),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_88),
.A2(n_71),
.B1(n_70),
.B2(n_72),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_97),
.B(n_61),
.C(n_58),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_74),
.B(n_39),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_119),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_120),
.B(n_124),
.Y(n_130)
);

AND2x6_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_86),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_121),
.B(n_92),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_95),
.A2(n_39),
.B1(n_16),
.B2(n_15),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_98),
.B(n_100),
.Y(n_124)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_77),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_125),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_45),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_126),
.B(n_92),
.Y(n_135)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_127),
.Y(n_133)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_77),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_77),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_129),
.B(n_57),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_SL g181 ( 
.A(n_132),
.B(n_135),
.C(n_158),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_125),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_137),
.Y(n_162)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_124),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_140),
.B(n_141),
.Y(n_171)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_128),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_118),
.A2(n_101),
.B1(n_117),
.B2(n_106),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_142),
.A2(n_154),
.B1(n_109),
.B2(n_129),
.Y(n_185)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_102),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_143),
.B(n_145),
.Y(n_168)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_144),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_120),
.B(n_76),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_117),
.B(n_76),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_146),
.B(n_148),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_108),
.B(n_73),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_147),
.Y(n_184)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_102),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_103),
.B(n_93),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_149),
.B(n_153),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_126),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_150),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_152),
.Y(n_180)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_105),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_115),
.A2(n_79),
.B1(n_82),
.B2(n_87),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_155),
.B(n_149),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_156),
.B(n_91),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_114),
.B(n_89),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_157),
.B(n_159),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_123),
.B(n_104),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_114),
.B(n_78),
.Y(n_159)
);

A2O1A1O1Ixp25_ASAP7_75t_L g160 ( 
.A1(n_107),
.A2(n_94),
.B(n_81),
.C(n_91),
.D(n_93),
.Y(n_160)
);

NAND3xp33_ASAP7_75t_L g165 ( 
.A(n_160),
.B(n_110),
.C(n_84),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_131),
.A2(n_111),
.B1(n_90),
.B2(n_81),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_163),
.A2(n_172),
.B1(n_183),
.B2(n_185),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_164),
.B(n_179),
.Y(n_207)
);

OAI21xp33_ASAP7_75t_SL g205 ( 
.A1(n_165),
.A2(n_160),
.B(n_151),
.Y(n_205)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_141),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_166),
.B(n_177),
.Y(n_198)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_134),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_167),
.B(n_170),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_169),
.B(n_186),
.C(n_150),
.Y(n_195)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_134),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_131),
.A2(n_90),
.B1(n_123),
.B2(n_104),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_144),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_175),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_146),
.B(n_116),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_176),
.A2(n_159),
.B(n_142),
.Y(n_215)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_130),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_130),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_178),
.B(n_187),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_143),
.A2(n_116),
.B(n_108),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_153),
.A2(n_99),
.B1(n_83),
.B2(n_80),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_155),
.B(n_45),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_145),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_147),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_188),
.B(n_190),
.Y(n_220)
);

OAI32xp33_ASAP7_75t_L g189 ( 
.A1(n_132),
.A2(n_39),
.A3(n_25),
.B1(n_57),
.B2(n_109),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_189),
.B(n_192),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_148),
.A2(n_57),
.B1(n_25),
.B2(n_26),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_137),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_166),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_193),
.B(n_194),
.Y(n_235)
);

INVx8_ASAP7_75t_L g194 ( 
.A(n_189),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_195),
.B(n_197),
.C(n_219),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_191),
.B(n_135),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_162),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_199),
.B(n_203),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_168),
.B(n_187),
.Y(n_200)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_200),
.Y(n_237)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_171),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_168),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_204),
.B(n_206),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_205),
.A2(n_209),
.B(n_216),
.Y(n_239)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_174),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_177),
.B(n_140),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_208),
.Y(n_236)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_174),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_172),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_210),
.B(n_179),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_178),
.B(n_158),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_212),
.A2(n_215),
.B(n_184),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_185),
.A2(n_151),
.B1(n_160),
.B2(n_136),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_214),
.A2(n_217),
.B1(n_154),
.B2(n_163),
.Y(n_225)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_191),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_176),
.A2(n_151),
.B1(n_188),
.B2(n_180),
.Y(n_217)
);

BUFx12f_ASAP7_75t_SL g218 ( 
.A(n_181),
.Y(n_218)
);

OA22x2_ASAP7_75t_L g233 ( 
.A1(n_218),
.A2(n_157),
.B1(n_182),
.B2(n_161),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_169),
.B(n_156),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_194),
.A2(n_215),
.B1(n_196),
.B2(n_218),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_221),
.A2(n_224),
.B1(n_229),
.B2(n_231),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_219),
.B(n_186),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_222),
.B(n_241),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_L g263 ( 
.A1(n_223),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_196),
.A2(n_180),
.B1(n_176),
.B2(n_170),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_225),
.A2(n_202),
.B1(n_216),
.B2(n_200),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_198),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_227),
.B(n_245),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_206),
.A2(n_167),
.B1(n_173),
.B2(n_181),
.Y(n_229)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_230),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_209),
.A2(n_138),
.B1(n_164),
.B2(n_133),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_204),
.A2(n_138),
.B1(n_133),
.B2(n_175),
.Y(n_232)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_232),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_233),
.A2(n_238),
.B(n_217),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_202),
.A2(n_161),
.B1(n_139),
.B2(n_25),
.Y(n_234)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_234),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_213),
.A2(n_139),
.B1(n_49),
.B2(n_26),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_195),
.B(n_49),
.C(n_45),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_240),
.B(n_244),
.C(n_246),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_207),
.B(n_49),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_207),
.B(n_49),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_242),
.B(n_220),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_197),
.B(n_49),
.C(n_45),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_203),
.B(n_15),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_214),
.B(n_45),
.C(n_1),
.Y(n_246)
);

AO221x1_ASAP7_75t_L g247 ( 
.A1(n_233),
.A2(n_193),
.B1(n_201),
.B2(n_45),
.C(n_212),
.Y(n_247)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_247),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_248),
.A2(n_263),
.B(n_224),
.Y(n_275)
);

INVxp33_ASAP7_75t_SL g249 ( 
.A(n_233),
.Y(n_249)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_249),
.Y(n_273)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_251),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_222),
.B(n_208),
.C(n_211),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_254),
.B(n_258),
.C(n_264),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_255),
.B(n_241),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_226),
.B(n_0),
.C(n_1),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_236),
.B(n_223),
.Y(n_259)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_259),
.Y(n_283)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_233),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_261),
.Y(n_270)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_243),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_262),
.B(n_266),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_226),
.B(n_2),
.C(n_3),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_238),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_240),
.B(n_3),
.C(n_4),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_267),
.B(n_244),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_271),
.B(n_278),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_250),
.B(n_242),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_272),
.B(n_280),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_256),
.B(n_229),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_274),
.B(n_257),
.Y(n_287)
);

AO21x1_ASAP7_75t_L g284 ( 
.A1(n_275),
.A2(n_248),
.B(n_270),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_276),
.B(n_255),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_SL g278 ( 
.A(n_265),
.B(n_221),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_266),
.A2(n_237),
.B1(n_246),
.B2(n_225),
.Y(n_279)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_279),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_250),
.B(n_254),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_265),
.B(n_239),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_281),
.B(n_251),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_284),
.A2(n_271),
.B(n_282),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_283),
.B(n_231),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_285),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_286),
.B(n_297),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_287),
.B(n_3),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_269),
.B(n_253),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_288),
.A2(n_294),
.B(n_295),
.Y(n_308)
);

INVx1_ASAP7_75t_SL g290 ( 
.A(n_273),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_290),
.B(n_292),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_268),
.B(n_232),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_277),
.A2(n_261),
.B(n_239),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_279),
.B(n_228),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_278),
.A2(n_260),
.B1(n_281),
.B2(n_252),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_296),
.B(n_282),
.Y(n_304)
);

AOI21xp33_ASAP7_75t_L g298 ( 
.A1(n_284),
.A2(n_235),
.B(n_228),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_298),
.A2(n_307),
.B(n_14),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_296),
.B(n_280),
.C(n_272),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_300),
.B(n_289),
.C(n_293),
.Y(n_314)
);

OAI321xp33_ASAP7_75t_L g301 ( 
.A1(n_290),
.A2(n_275),
.A3(n_234),
.B1(n_276),
.B2(n_267),
.C(n_252),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_301),
.A2(n_303),
.B(n_304),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_293),
.B(n_264),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_305),
.B(n_4),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_291),
.A2(n_258),
.B1(n_15),
.B2(n_14),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_309),
.B(n_4),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_308),
.B(n_297),
.Y(n_310)
);

OAI21xp33_ASAP7_75t_L g319 ( 
.A1(n_310),
.A2(n_317),
.B(n_318),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_311),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_313),
.A2(n_5),
.B(n_6),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_314),
.A2(n_315),
.B(n_300),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_303),
.A2(n_286),
.B(n_14),
.Y(n_315)
);

NOR2xp67_ASAP7_75t_L g316 ( 
.A(n_299),
.B(n_13),
.Y(n_316)
);

AOI322xp5_ASAP7_75t_L g320 ( 
.A1(n_316),
.A2(n_307),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_4),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_302),
.B(n_299),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_L g328 ( 
.A1(n_320),
.A2(n_317),
.B1(n_10),
.B2(n_11),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_321),
.A2(n_322),
.B(n_323),
.Y(n_327)
);

AOI322xp5_ASAP7_75t_L g322 ( 
.A1(n_315),
.A2(n_306),
.A3(n_6),
.B1(n_8),
.B2(n_9),
.C1(n_10),
.C2(n_11),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_312),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_325),
.A2(n_8),
.B(n_9),
.Y(n_326)
);

OAI21x1_ASAP7_75t_L g329 ( 
.A1(n_326),
.A2(n_328),
.B(n_9),
.Y(n_329)
);

AOI322xp5_ASAP7_75t_SL g330 ( 
.A1(n_329),
.A2(n_324),
.A3(n_327),
.B1(n_11),
.B2(n_9),
.C1(n_10),
.C2(n_319),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_10),
.Y(n_331)
);


endmodule