module fake_jpeg_2915_n_159 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_159);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_159;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_4),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_22),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_0),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_13),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_0),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_59),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_40),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_61),
.Y(n_64)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_62),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_63),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_49),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_69),
.B(n_48),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_57),
.A2(n_43),
.B1(n_52),
.B2(n_47),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_71),
.A2(n_73),
.B1(n_74),
.B2(n_75),
.Y(n_82)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_72),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_63),
.A2(n_43),
.B1(n_47),
.B2(n_49),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_60),
.A2(n_45),
.B1(n_55),
.B2(n_56),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_61),
.A2(n_53),
.B1(n_48),
.B2(n_44),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_66),
.B(n_41),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_76),
.B(n_78),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_54),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_70),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_79),
.B(n_80),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_51),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_70),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_83),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_51),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_46),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_88),
.Y(n_95)
);

A2O1A1Ixp33_ASAP7_75t_L g87 ( 
.A1(n_65),
.A2(n_1),
.B(n_2),
.C(n_4),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_87),
.B(n_5),
.Y(n_101)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_89),
.Y(n_99)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_36),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_91),
.B(n_39),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_82),
.A2(n_46),
.B1(n_72),
.B2(n_6),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_101),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_90),
.A2(n_1),
.B1(n_5),
.B2(n_6),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_97),
.A2(n_104),
.B1(n_101),
.B2(n_102),
.Y(n_109)
);

OA22x2_ASAP7_75t_L g98 ( 
.A1(n_88),
.A2(n_21),
.B1(n_38),
.B2(n_37),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_100),
.B(n_103),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_105),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_7),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_87),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_77),
.B(n_35),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_77),
.B(n_33),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_107),
.B(n_11),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_113),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_95),
.A2(n_104),
.B1(n_108),
.B2(n_93),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_111),
.A2(n_117),
.B1(n_118),
.B2(n_119),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_106),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_106),
.A2(n_80),
.B(n_81),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_114),
.A2(n_110),
.B(n_122),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_105),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_116),
.B(n_120),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_99),
.A2(n_79),
.B1(n_89),
.B2(n_85),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_107),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_98),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_94),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_121),
.B(n_123),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_SL g124 ( 
.A(n_98),
.B(n_92),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_124),
.B(n_125),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_95),
.B(n_23),
.C(n_31),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_126),
.B(n_25),
.Y(n_136)
);

AOI221xp5_ASAP7_75t_L g127 ( 
.A1(n_111),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.C(n_16),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_127),
.B(n_128),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_117),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_15),
.Y(n_129)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_129),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_115),
.A2(n_26),
.B(n_30),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_130),
.B(n_133),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_123),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_133)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_136),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_138),
.B(n_139),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_124),
.A2(n_32),
.B(n_27),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_135),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_145),
.B(n_129),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_143),
.B(n_138),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_146),
.B(n_147),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_141),
.A2(n_134),
.B1(n_131),
.B2(n_129),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_148),
.B(n_149),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_141),
.A2(n_137),
.B1(n_142),
.B2(n_140),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_151),
.B(n_112),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_144),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_150),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_154),
.A2(n_147),
.B1(n_137),
.B2(n_143),
.Y(n_155)
);

A2O1A1Ixp33_ASAP7_75t_L g156 ( 
.A1(n_155),
.A2(n_130),
.B(n_133),
.C(n_109),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_156),
.A2(n_146),
.B(n_119),
.Y(n_157)
);

NOR3xp33_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_132),
.C(n_118),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_125),
.Y(n_159)
);


endmodule