module fake_netlist_6_445_n_1695 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_149, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1695);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_149;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1695;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_544;
wire n_250;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_153;
wire n_842;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_154;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_152;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_133),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_117),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_31),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_73),
.Y(n_155)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_89),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_26),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_41),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_29),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_36),
.Y(n_160)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_12),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_85),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_72),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_14),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_119),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_74),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_124),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_137),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_123),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_80),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_93),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_135),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_57),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_41),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_6),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_6),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_134),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_31),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_139),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_150),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_33),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_76),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_44),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_59),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_44),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_5),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_18),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_37),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_97),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_61),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_63),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_28),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_136),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_69),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_34),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_87),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_12),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_84),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_48),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_20),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_42),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_130),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_95),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_128),
.Y(n_204)
);

BUFx2_ASAP7_75t_L g205 ( 
.A(n_28),
.Y(n_205)
);

INVx2_ASAP7_75t_SL g206 ( 
.A(n_83),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_64),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_70),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_79),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_143),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_77),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_98),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_78),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_108),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_20),
.Y(n_215)
);

CKINVDCx14_ASAP7_75t_R g216 ( 
.A(n_122),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_51),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_109),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_99),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_103),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_7),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_27),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_62),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_102),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_125),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_112),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_144),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_0),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_5),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_126),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_129),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_131),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_1),
.Y(n_233)
);

BUFx8_ASAP7_75t_SL g234 ( 
.A(n_40),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_42),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_18),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_110),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_53),
.Y(n_238)
);

BUFx10_ASAP7_75t_L g239 ( 
.A(n_107),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_88),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_56),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_100),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_58),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_43),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_15),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_94),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_60),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_22),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_14),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_151),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_35),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_45),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_10),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_101),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_116),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_15),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_33),
.Y(n_257)
);

INVx2_ASAP7_75t_SL g258 ( 
.A(n_26),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_50),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_29),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_140),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_16),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_67),
.Y(n_263)
);

INVx2_ASAP7_75t_SL g264 ( 
.A(n_147),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g265 ( 
.A(n_3),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_92),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_120),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_40),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_52),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_71),
.Y(n_270)
);

BUFx8_ASAP7_75t_SL g271 ( 
.A(n_86),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_105),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_45),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_48),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_0),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_113),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_121),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_1),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_25),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_114),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_2),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_132),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_7),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_146),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_50),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_75),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_111),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_104),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_8),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_24),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_23),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_118),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_66),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_149),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_43),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_32),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_37),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_115),
.Y(n_298)
);

INVx2_ASAP7_75t_SL g299 ( 
.A(n_49),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_145),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_23),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_65),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_81),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_180),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_236),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_271),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_236),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_236),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_236),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_189),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_236),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_236),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_191),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_247),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_267),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_289),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_289),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_216),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_289),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_174),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_174),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_234),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_178),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_178),
.Y(n_324)
);

INVxp67_ASAP7_75t_SL g325 ( 
.A(n_237),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_161),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_228),
.Y(n_327)
);

INVxp33_ASAP7_75t_L g328 ( 
.A(n_161),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_228),
.Y(n_329)
);

HB1xp67_ASAP7_75t_L g330 ( 
.A(n_205),
.Y(n_330)
);

INVxp33_ASAP7_75t_SL g331 ( 
.A(n_205),
.Y(n_331)
);

INVx1_ASAP7_75t_SL g332 ( 
.A(n_186),
.Y(n_332)
);

INVxp33_ASAP7_75t_SL g333 ( 
.A(n_157),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_260),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g335 ( 
.A(n_239),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_152),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_269),
.Y(n_337)
);

CKINVDCx16_ASAP7_75t_R g338 ( 
.A(n_239),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_260),
.Y(n_339)
);

INVxp33_ASAP7_75t_L g340 ( 
.A(n_154),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_265),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_265),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_265),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_153),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_154),
.Y(n_345)
);

HB1xp67_ASAP7_75t_L g346 ( 
.A(n_158),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_164),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_164),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_165),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_166),
.Y(n_350)
);

CKINVDCx14_ASAP7_75t_R g351 ( 
.A(n_239),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_181),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_163),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_167),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_181),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_221),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_168),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_221),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_169),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_252),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_252),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_256),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_256),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_172),
.Y(n_364)
);

BUFx3_ASAP7_75t_L g365 ( 
.A(n_237),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_173),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_259),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_184),
.Y(n_368)
);

INVxp67_ASAP7_75t_SL g369 ( 
.A(n_237),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_259),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_273),
.Y(n_371)
);

BUFx3_ASAP7_75t_L g372 ( 
.A(n_240),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_190),
.Y(n_373)
);

INVxp67_ASAP7_75t_SL g374 ( 
.A(n_240),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_273),
.Y(n_375)
);

INVxp67_ASAP7_75t_SL g376 ( 
.A(n_240),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_285),
.Y(n_377)
);

BUFx3_ASAP7_75t_L g378 ( 
.A(n_239),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_305),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_305),
.Y(n_380)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_325),
.B(n_258),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_304),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_307),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_353),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_307),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_369),
.B(n_206),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_374),
.B(n_376),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_308),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_341),
.B(n_342),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_336),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_308),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_309),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_309),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_311),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_331),
.A2(n_192),
.B1(n_195),
.B2(n_283),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_350),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_311),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_353),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_332),
.A2(n_262),
.B1(n_197),
.B2(n_249),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_341),
.B(n_342),
.Y(n_400)
);

INVx3_ASAP7_75t_L g401 ( 
.A(n_312),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_312),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_346),
.Y(n_403)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_323),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_354),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_323),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_343),
.B(n_206),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_345),
.Y(n_408)
);

HB1xp67_ASAP7_75t_L g409 ( 
.A(n_326),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_345),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_347),
.Y(n_411)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_316),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_316),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_343),
.B(n_264),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_347),
.Y(n_415)
);

NOR2x1_ASAP7_75t_L g416 ( 
.A(n_378),
.B(n_163),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_348),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_359),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_317),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_348),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_365),
.B(n_264),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_365),
.B(n_163),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_368),
.Y(n_423)
);

BUFx2_ASAP7_75t_L g424 ( 
.A(n_378),
.Y(n_424)
);

AND2x4_ASAP7_75t_L g425 ( 
.A(n_372),
.B(n_193),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_310),
.B(n_251),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_352),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_352),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_355),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_330),
.A2(n_257),
.B1(n_275),
.B2(n_183),
.Y(n_430)
);

INVx3_ASAP7_75t_L g431 ( 
.A(n_317),
.Y(n_431)
);

AO22x1_ASAP7_75t_L g432 ( 
.A1(n_328),
.A2(n_258),
.B1(n_299),
.B2(n_285),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_319),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_372),
.B(n_194),
.Y(n_434)
);

AND2x4_ASAP7_75t_L g435 ( 
.A(n_319),
.B(n_193),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_355),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_356),
.Y(n_437)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_371),
.Y(n_438)
);

AND2x4_ASAP7_75t_L g439 ( 
.A(n_356),
.B(n_220),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_358),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_358),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_360),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_360),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_320),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_361),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_361),
.B(n_196),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_320),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_384),
.Y(n_448)
);

INVx2_ASAP7_75t_SL g449 ( 
.A(n_387),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_389),
.Y(n_450)
);

NAND3xp33_ASAP7_75t_L g451 ( 
.A(n_438),
.B(n_351),
.C(n_338),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_406),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_389),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_406),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_406),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_406),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_424),
.B(n_335),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_406),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_389),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_SL g460 ( 
.A(n_390),
.B(n_306),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_382),
.Y(n_461)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_384),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_408),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_406),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_379),
.Y(n_465)
);

AO21x2_ASAP7_75t_L g466 ( 
.A1(n_434),
.A2(n_162),
.B(n_155),
.Y(n_466)
);

INVx8_ASAP7_75t_L g467 ( 
.A(n_387),
.Y(n_467)
);

AOI22xp33_ASAP7_75t_L g468 ( 
.A1(n_387),
.A2(n_299),
.B1(n_291),
.B2(n_301),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_384),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_384),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_424),
.B(n_335),
.Y(n_471)
);

AND2x6_ASAP7_75t_L g472 ( 
.A(n_422),
.B(n_208),
.Y(n_472)
);

NAND2xp33_ASAP7_75t_SL g473 ( 
.A(n_386),
.B(n_159),
.Y(n_473)
);

BUFx10_ASAP7_75t_L g474 ( 
.A(n_396),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_384),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_384),
.Y(n_476)
);

AOI22x1_ASAP7_75t_L g477 ( 
.A1(n_422),
.A2(n_338),
.B1(n_292),
.B2(n_284),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_405),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_434),
.B(n_318),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_395),
.B(n_313),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_379),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_380),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_418),
.B(n_333),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_380),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_398),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_381),
.B(n_156),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_426),
.Y(n_487)
);

INVx4_ASAP7_75t_L g488 ( 
.A(n_402),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_408),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_410),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_398),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_381),
.B(n_232),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_410),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_398),
.Y(n_494)
);

INVx4_ASAP7_75t_L g495 ( 
.A(n_402),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_411),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_398),
.Y(n_497)
);

AND3x2_ASAP7_75t_L g498 ( 
.A(n_409),
.B(n_179),
.C(n_220),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_422),
.B(n_198),
.Y(n_499)
);

OR2x6_ASAP7_75t_L g500 ( 
.A(n_432),
.B(n_290),
.Y(n_500)
);

NAND2xp33_ASAP7_75t_R g501 ( 
.A(n_423),
.B(n_322),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_403),
.A2(n_357),
.B1(n_373),
.B2(n_366),
.Y(n_502)
);

INVx8_ASAP7_75t_L g503 ( 
.A(n_425),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_446),
.B(n_344),
.Y(n_504)
);

NAND2xp33_ASAP7_75t_SL g505 ( 
.A(n_438),
.B(n_160),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_411),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_403),
.B(n_349),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_398),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_415),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_398),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_425),
.B(n_321),
.Y(n_511)
);

INVx2_ASAP7_75t_SL g512 ( 
.A(n_425),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_446),
.B(n_364),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_385),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_413),
.Y(n_515)
);

OAI22xp33_ASAP7_75t_SL g516 ( 
.A1(n_421),
.A2(n_155),
.B1(n_303),
.B2(n_171),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_413),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_421),
.B(n_340),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_413),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_399),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_413),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_425),
.B(n_202),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_416),
.B(n_207),
.Y(n_523)
);

CKINVDCx16_ASAP7_75t_R g524 ( 
.A(n_426),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_415),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_417),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_413),
.Y(n_527)
);

BUFx4f_ASAP7_75t_L g528 ( 
.A(n_402),
.Y(n_528)
);

OAI21xp33_ASAP7_75t_SL g529 ( 
.A1(n_407),
.A2(n_170),
.B(n_162),
.Y(n_529)
);

NOR2x1p5_ASAP7_75t_L g530 ( 
.A(n_400),
.B(n_175),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_417),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_420),
.B(n_321),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_420),
.Y(n_533)
);

BUFx3_ASAP7_75t_L g534 ( 
.A(n_435),
.Y(n_534)
);

INVx1_ASAP7_75t_SL g535 ( 
.A(n_409),
.Y(n_535)
);

AOI21x1_ASAP7_75t_L g536 ( 
.A1(n_385),
.A2(n_171),
.B(n_170),
.Y(n_536)
);

INVx4_ASAP7_75t_L g537 ( 
.A(n_402),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_416),
.B(n_314),
.Y(n_538)
);

NAND2xp33_ASAP7_75t_L g539 ( 
.A(n_407),
.B(n_208),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_388),
.B(n_209),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_413),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_414),
.B(n_315),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_L g543 ( 
.A1(n_430),
.A2(n_253),
.B1(n_245),
.B2(n_244),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_427),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_383),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_383),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_427),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_388),
.Y(n_548)
);

INVx3_ASAP7_75t_L g549 ( 
.A(n_402),
.Y(n_549)
);

AOI22xp33_ASAP7_75t_L g550 ( 
.A1(n_439),
.A2(n_291),
.B1(n_290),
.B2(n_301),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_414),
.B(n_337),
.Y(n_551)
);

BUFx6f_ASAP7_75t_L g552 ( 
.A(n_402),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_391),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_391),
.B(n_210),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_383),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_393),
.Y(n_556)
);

INVx3_ASAP7_75t_L g557 ( 
.A(n_401),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_393),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_SL g559 ( 
.A(n_395),
.B(n_212),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_393),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_430),
.B(n_213),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g562 ( 
.A(n_435),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_392),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_392),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_397),
.Y(n_565)
);

NOR3xp33_ASAP7_75t_L g566 ( 
.A(n_399),
.B(n_248),
.C(n_176),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_394),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_394),
.Y(n_568)
);

OAI21xp33_ASAP7_75t_SL g569 ( 
.A1(n_428),
.A2(n_177),
.B(n_182),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_394),
.Y(n_570)
);

OAI22xp33_ASAP7_75t_L g571 ( 
.A1(n_400),
.A2(n_235),
.B1(n_233),
.B2(n_185),
.Y(n_571)
);

OR2x6_ASAP7_75t_L g572 ( 
.A(n_432),
.B(n_177),
.Y(n_572)
);

INVx4_ASAP7_75t_L g573 ( 
.A(n_435),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_428),
.B(n_324),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_397),
.B(n_214),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_447),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_447),
.Y(n_577)
);

INVx1_ASAP7_75t_SL g578 ( 
.A(n_439),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_447),
.Y(n_579)
);

BUFx6f_ASAP7_75t_L g580 ( 
.A(n_435),
.Y(n_580)
);

OR2x6_ASAP7_75t_L g581 ( 
.A(n_439),
.B(n_182),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_429),
.Y(n_582)
);

OA22x2_ASAP7_75t_L g583 ( 
.A1(n_439),
.A2(n_377),
.B1(n_375),
.B2(n_370),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_429),
.B(n_217),
.Y(n_584)
);

INVx3_ASAP7_75t_L g585 ( 
.A(n_401),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_436),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_436),
.B(n_187),
.Y(n_587)
);

INVxp33_ASAP7_75t_SL g588 ( 
.A(n_437),
.Y(n_588)
);

INVxp33_ASAP7_75t_L g589 ( 
.A(n_437),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_440),
.Y(n_590)
);

AOI22xp33_ASAP7_75t_L g591 ( 
.A1(n_440),
.A2(n_284),
.B1(n_292),
.B2(n_266),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_441),
.B(n_324),
.Y(n_592)
);

INVx3_ASAP7_75t_L g593 ( 
.A(n_401),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_441),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_404),
.B(n_219),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_518),
.B(n_442),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_512),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_512),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_465),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_545),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_578),
.B(n_412),
.Y(n_601)
);

OAI22x1_ASAP7_75t_SL g602 ( 
.A1(n_520),
.A2(n_229),
.B1(n_278),
.B2(n_279),
.Y(n_602)
);

OAI221xp5_ASAP7_75t_L g603 ( 
.A1(n_468),
.A2(n_442),
.B1(n_445),
.B2(n_443),
.C(n_277),
.Y(n_603)
);

AOI22xp33_ASAP7_75t_L g604 ( 
.A1(n_449),
.A2(n_226),
.B1(n_277),
.B2(n_203),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_545),
.Y(n_605)
);

AOI22xp5_ASAP7_75t_SL g606 ( 
.A1(n_520),
.A2(n_222),
.B1(n_215),
.B2(n_201),
.Y(n_606)
);

OAI21xp5_ASAP7_75t_L g607 ( 
.A1(n_450),
.A2(n_453),
.B(n_449),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_573),
.B(n_467),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_467),
.B(n_412),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_588),
.B(n_188),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_503),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_467),
.B(n_412),
.Y(n_612)
);

INVx2_ASAP7_75t_SL g613 ( 
.A(n_530),
.Y(n_613)
);

NAND2x1_ASAP7_75t_L g614 ( 
.A(n_573),
.B(n_412),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_546),
.Y(n_615)
);

NAND3xp33_ASAP7_75t_L g616 ( 
.A(n_542),
.B(n_297),
.C(n_296),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_546),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_450),
.B(n_431),
.Y(n_618)
);

HB1xp67_ASAP7_75t_L g619 ( 
.A(n_535),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_588),
.B(n_199),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_589),
.B(n_443),
.Y(n_621)
);

INVx2_ASAP7_75t_SL g622 ( 
.A(n_511),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_453),
.B(n_431),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_573),
.B(n_208),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_511),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_459),
.B(n_447),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_463),
.B(n_447),
.Y(n_627)
);

A2O1A1Ixp33_ASAP7_75t_L g628 ( 
.A1(n_569),
.A2(n_241),
.B(n_266),
.C(n_282),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_589),
.B(n_200),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_504),
.B(n_268),
.Y(n_630)
);

INVx2_ASAP7_75t_SL g631 ( 
.A(n_498),
.Y(n_631)
);

INVx2_ASAP7_75t_SL g632 ( 
.A(n_532),
.Y(n_632)
);

AO221x1_ASAP7_75t_L g633 ( 
.A1(n_571),
.A2(n_208),
.B1(n_203),
.B2(n_204),
.C(n_226),
.Y(n_633)
);

BUFx4f_ASAP7_75t_L g634 ( 
.A(n_572),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_534),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_489),
.B(n_447),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_479),
.B(n_274),
.Y(n_637)
);

NAND2xp33_ASAP7_75t_L g638 ( 
.A(n_503),
.B(n_224),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_562),
.B(n_208),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_490),
.B(n_204),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_493),
.B(n_211),
.Y(n_641)
);

NOR3xp33_ASAP7_75t_L g642 ( 
.A(n_507),
.B(n_281),
.C(n_295),
.Y(n_642)
);

AOI22xp5_ASAP7_75t_L g643 ( 
.A1(n_551),
.A2(n_263),
.B1(n_225),
.B2(n_302),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_496),
.B(n_211),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_562),
.B(n_208),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_486),
.B(n_218),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_506),
.B(n_218),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_509),
.B(n_223),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_525),
.B(n_223),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_526),
.B(n_241),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_534),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_531),
.B(n_282),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_492),
.B(n_300),
.Y(n_653)
);

INVx3_ASAP7_75t_L g654 ( 
.A(n_562),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_465),
.Y(n_655)
);

INVxp67_ASAP7_75t_L g656 ( 
.A(n_505),
.Y(n_656)
);

NAND2xp33_ASAP7_75t_SL g657 ( 
.A(n_457),
.B(n_227),
.Y(n_657)
);

AOI22xp33_ASAP7_75t_L g658 ( 
.A1(n_466),
.A2(n_300),
.B1(n_303),
.B2(n_445),
.Y(n_658)
);

OAI22xp5_ASAP7_75t_L g659 ( 
.A1(n_499),
.A2(n_288),
.B1(n_231),
.B2(n_238),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_562),
.B(n_230),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_533),
.B(n_404),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_544),
.B(n_404),
.Y(n_662)
);

OAI22xp5_ASAP7_75t_SL g663 ( 
.A1(n_480),
.A2(n_362),
.B1(n_377),
.B2(n_375),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_532),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_574),
.Y(n_665)
);

INVx1_ASAP7_75t_SL g666 ( 
.A(n_461),
.Y(n_666)
);

INVx3_ASAP7_75t_L g667 ( 
.A(n_562),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_561),
.B(n_242),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_513),
.B(n_243),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_SL g670 ( 
.A(n_478),
.B(n_246),
.Y(n_670)
);

NAND2x1p5_ASAP7_75t_L g671 ( 
.A(n_580),
.B(n_404),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_538),
.B(n_250),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_547),
.B(n_254),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_481),
.Y(n_674)
);

NOR2xp67_ASAP7_75t_L g675 ( 
.A(n_451),
.B(n_280),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_580),
.B(n_557),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_474),
.B(n_367),
.Y(n_677)
);

AOI22xp5_ASAP7_75t_L g678 ( 
.A1(n_473),
.A2(n_255),
.B1(n_261),
.B2(n_270),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_580),
.B(n_272),
.Y(n_679)
);

AND2x4_ASAP7_75t_L g680 ( 
.A(n_582),
.B(n_367),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_586),
.B(n_590),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_580),
.B(n_276),
.Y(n_682)
);

INVxp67_ASAP7_75t_L g683 ( 
.A(n_505),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_580),
.B(n_286),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_574),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_594),
.B(n_444),
.Y(n_686)
);

OR2x2_ASAP7_75t_L g687 ( 
.A(n_471),
.B(n_362),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_481),
.B(n_444),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_482),
.B(n_444),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_592),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_557),
.B(n_585),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_555),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_592),
.Y(n_693)
);

OR2x2_ASAP7_75t_L g694 ( 
.A(n_524),
.B(n_363),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_540),
.B(n_287),
.Y(n_695)
);

NOR3xp33_ASAP7_75t_L g696 ( 
.A(n_543),
.B(n_370),
.C(n_363),
.Y(n_696)
);

AOI21xp5_ASAP7_75t_L g697 ( 
.A1(n_503),
.A2(n_433),
.B(n_419),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_484),
.B(n_514),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_514),
.B(n_433),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_555),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_548),
.B(n_433),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_553),
.Y(n_702)
);

AOI22xp5_ASAP7_75t_L g703 ( 
.A1(n_473),
.A2(n_293),
.B1(n_294),
.B2(n_298),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_553),
.B(n_419),
.Y(n_704)
);

BUFx6f_ASAP7_75t_L g705 ( 
.A(n_503),
.Y(n_705)
);

O2A1O1Ixp33_ASAP7_75t_L g706 ( 
.A1(n_516),
.A2(n_339),
.B(n_334),
.C(n_329),
.Y(n_706)
);

INVx2_ASAP7_75t_SL g707 ( 
.A(n_522),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_563),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_557),
.B(n_339),
.Y(n_709)
);

INVx3_ASAP7_75t_L g710 ( 
.A(n_585),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_556),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_563),
.B(n_334),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_478),
.Y(n_713)
);

INVx5_ASAP7_75t_L g714 ( 
.A(n_472),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_564),
.B(n_329),
.Y(n_715)
);

O2A1O1Ixp33_ASAP7_75t_L g716 ( 
.A1(n_539),
.A2(n_327),
.B(n_3),
.C(n_4),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_585),
.B(n_327),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_556),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_564),
.B(n_148),
.Y(n_719)
);

INVx2_ASAP7_75t_SL g720 ( 
.A(n_583),
.Y(n_720)
);

OAI22xp5_ASAP7_75t_L g721 ( 
.A1(n_477),
.A2(n_142),
.B1(n_141),
.B2(n_138),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_565),
.B(n_127),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_565),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_593),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_554),
.B(n_2),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_593),
.B(n_106),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_593),
.B(n_96),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_583),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_558),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_575),
.B(n_91),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_558),
.Y(n_731)
);

OR2x2_ASAP7_75t_L g732 ( 
.A(n_502),
.B(n_500),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_466),
.B(n_90),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_560),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_560),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_583),
.Y(n_736)
);

A2O1A1Ixp33_ASAP7_75t_L g737 ( 
.A1(n_529),
.A2(n_4),
.B(n_8),
.C(n_9),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_466),
.B(n_82),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_477),
.B(n_68),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_567),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_587),
.B(n_55),
.Y(n_741)
);

OAI221xp5_ASAP7_75t_L g742 ( 
.A1(n_550),
.A2(n_591),
.B1(n_559),
.B2(n_500),
.C(n_572),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_523),
.B(n_54),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_567),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_568),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_595),
.B(n_9),
.Y(n_746)
);

BUFx6f_ASAP7_75t_L g747 ( 
.A(n_448),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_568),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_474),
.B(n_10),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_549),
.B(n_11),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_584),
.B(n_11),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_570),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_515),
.B(n_13),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_549),
.B(n_49),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_515),
.B(n_13),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_570),
.Y(n_756)
);

OAI221xp5_ASAP7_75t_L g757 ( 
.A1(n_500),
.A2(n_16),
.B1(n_17),
.B2(n_19),
.C(n_21),
.Y(n_757)
);

BUFx3_ASAP7_75t_L g758 ( 
.A(n_474),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_581),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_517),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_549),
.B(n_17),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_517),
.B(n_19),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_599),
.Y(n_763)
);

OAI21xp33_ASAP7_75t_L g764 ( 
.A1(n_630),
.A2(n_566),
.B(n_460),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_596),
.B(n_581),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_672),
.B(n_581),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_607),
.B(n_519),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_672),
.B(n_581),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_630),
.B(n_462),
.Y(n_769)
);

OR2x2_ASAP7_75t_L g770 ( 
.A(n_619),
.B(n_461),
.Y(n_770)
);

BUFx3_ASAP7_75t_L g771 ( 
.A(n_758),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_655),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_621),
.B(n_462),
.Y(n_773)
);

OR2x6_ASAP7_75t_L g774 ( 
.A(n_758),
.B(n_572),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_674),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_674),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_702),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_677),
.B(n_483),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_708),
.Y(n_779)
);

BUFx6f_ASAP7_75t_L g780 ( 
.A(n_611),
.Y(n_780)
);

NOR3xp33_ASAP7_75t_SL g781 ( 
.A(n_663),
.B(n_480),
.C(n_501),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_723),
.Y(n_782)
);

INVx5_ASAP7_75t_L g783 ( 
.A(n_611),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_714),
.B(n_519),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_729),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_729),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_724),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_625),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_597),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_734),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_734),
.Y(n_791)
);

INVx2_ASAP7_75t_SL g792 ( 
.A(n_694),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_598),
.Y(n_793)
);

INVx8_ASAP7_75t_L g794 ( 
.A(n_713),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_SL g795 ( 
.A(n_666),
.B(n_487),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_710),
.Y(n_796)
);

BUFx3_ASAP7_75t_L g797 ( 
.A(n_759),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_735),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_710),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_646),
.B(n_521),
.Y(n_800)
);

NAND2xp33_ASAP7_75t_R g801 ( 
.A(n_732),
.B(n_572),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_714),
.B(n_521),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_735),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_635),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_653),
.B(n_527),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_653),
.B(n_527),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_707),
.B(n_695),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_651),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_695),
.B(n_541),
.Y(n_809)
);

INVxp67_ASAP7_75t_SL g810 ( 
.A(n_747),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_622),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_626),
.Y(n_812)
);

INVx3_ASAP7_75t_L g813 ( 
.A(n_654),
.Y(n_813)
);

AO21x1_ASAP7_75t_L g814 ( 
.A1(n_739),
.A2(n_536),
.B(n_539),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_632),
.B(n_541),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_609),
.A2(n_528),
.B(n_488),
.Y(n_816)
);

AOI22xp33_ASAP7_75t_L g817 ( 
.A1(n_728),
.A2(n_472),
.B1(n_577),
.B2(n_576),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_740),
.Y(n_818)
);

INVx5_ASAP7_75t_L g819 ( 
.A(n_611),
.Y(n_819)
);

BUFx6f_ASAP7_75t_L g820 ( 
.A(n_611),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_637),
.B(n_469),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_610),
.B(n_620),
.Y(n_822)
);

INVx2_ASAP7_75t_SL g823 ( 
.A(n_687),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_714),
.B(n_705),
.Y(n_824)
);

AOI22xp5_ASAP7_75t_L g825 ( 
.A1(n_637),
.A2(n_472),
.B1(n_577),
.B2(n_576),
.Y(n_825)
);

INVxp67_ASAP7_75t_L g826 ( 
.A(n_629),
.Y(n_826)
);

INVxp67_ASAP7_75t_SL g827 ( 
.A(n_747),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_744),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_698),
.B(n_470),
.Y(n_829)
);

BUFx3_ASAP7_75t_L g830 ( 
.A(n_720),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_744),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_745),
.Y(n_832)
);

AOI22xp33_ASAP7_75t_L g833 ( 
.A1(n_736),
.A2(n_472),
.B1(n_579),
.B2(n_458),
.Y(n_833)
);

O2A1O1Ixp5_ASAP7_75t_L g834 ( 
.A1(n_739),
.A2(n_536),
.B(n_458),
.C(n_454),
.Y(n_834)
);

BUFx8_ASAP7_75t_L g835 ( 
.A(n_749),
.Y(n_835)
);

AOI21xp5_ASAP7_75t_L g836 ( 
.A1(n_612),
.A2(n_528),
.B(n_495),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_601),
.B(n_475),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_664),
.B(n_485),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_656),
.B(n_537),
.Y(n_839)
);

INVxp67_ASAP7_75t_SL g840 ( 
.A(n_747),
.Y(n_840)
);

AOI22xp33_ASAP7_75t_L g841 ( 
.A1(n_658),
.A2(n_472),
.B1(n_579),
.B2(n_456),
.Y(n_841)
);

NAND2xp33_ASAP7_75t_L g842 ( 
.A(n_705),
.B(n_476),
.Y(n_842)
);

BUFx3_ASAP7_75t_L g843 ( 
.A(n_665),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_745),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_685),
.Y(n_845)
);

AOI22xp5_ASAP7_75t_L g846 ( 
.A1(n_683),
.A2(n_469),
.B1(n_485),
.B2(n_510),
.Y(n_846)
);

NAND2xp33_ASAP7_75t_L g847 ( 
.A(n_705),
.B(n_476),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_610),
.B(n_487),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_714),
.B(n_741),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_620),
.B(n_452),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_690),
.Y(n_851)
);

BUFx6f_ASAP7_75t_L g852 ( 
.A(n_747),
.Y(n_852)
);

OR2x2_ASAP7_75t_SL g853 ( 
.A(n_616),
.B(n_452),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_600),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_605),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_693),
.B(n_681),
.Y(n_856)
);

BUFx6f_ASAP7_75t_L g857 ( 
.A(n_654),
.Y(n_857)
);

AOI22xp5_ASAP7_75t_L g858 ( 
.A1(n_668),
.A2(n_494),
.B1(n_491),
.B2(n_510),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_742),
.B(n_537),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_618),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_725),
.B(n_658),
.Y(n_861)
);

BUFx6f_ASAP7_75t_L g862 ( 
.A(n_667),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_725),
.B(n_491),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_623),
.Y(n_864)
);

INVx3_ASAP7_75t_L g865 ( 
.A(n_667),
.Y(n_865)
);

HB1xp67_ASAP7_75t_L g866 ( 
.A(n_680),
.Y(n_866)
);

AOI22xp33_ASAP7_75t_L g867 ( 
.A1(n_633),
.A2(n_604),
.B1(n_757),
.B2(n_751),
.Y(n_867)
);

BUFx6f_ASAP7_75t_L g868 ( 
.A(n_671),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_SL g869 ( 
.A(n_730),
.B(n_454),
.Y(n_869)
);

INVx2_ASAP7_75t_SL g870 ( 
.A(n_680),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_670),
.B(n_488),
.Y(n_871)
);

OR2x2_ASAP7_75t_L g872 ( 
.A(n_613),
.B(n_497),
.Y(n_872)
);

AOI22xp5_ASAP7_75t_L g873 ( 
.A1(n_668),
.A2(n_497),
.B1(n_455),
.B2(n_456),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_604),
.B(n_455),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_669),
.B(n_488),
.Y(n_875)
);

NAND2x1p5_ASAP7_75t_L g876 ( 
.A(n_608),
.B(n_495),
.Y(n_876)
);

AOI22xp5_ASAP7_75t_L g877 ( 
.A1(n_669),
.A2(n_464),
.B1(n_495),
.B2(n_537),
.Y(n_877)
);

AND2x4_ASAP7_75t_L g878 ( 
.A(n_631),
.B(n_464),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_688),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_689),
.Y(n_880)
);

BUFx3_ASAP7_75t_L g881 ( 
.A(n_634),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_748),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_615),
.Y(n_883)
);

AOI22xp33_ASAP7_75t_SL g884 ( 
.A1(n_751),
.A2(n_21),
.B1(n_22),
.B2(n_24),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_673),
.B(n_508),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_673),
.B(n_508),
.Y(n_886)
);

NOR2xp67_ASAP7_75t_L g887 ( 
.A(n_643),
.B(n_552),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_617),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_752),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_712),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_606),
.B(n_25),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_640),
.B(n_508),
.Y(n_892)
);

INVxp67_ASAP7_75t_L g893 ( 
.A(n_641),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_715),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_644),
.B(n_647),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_648),
.B(n_508),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_686),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_696),
.B(n_27),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_692),
.Y(n_899)
);

AND2x4_ASAP7_75t_L g900 ( 
.A(n_675),
.B(n_608),
.Y(n_900)
);

AOI22xp33_ASAP7_75t_L g901 ( 
.A1(n_721),
.A2(n_508),
.B1(n_476),
.B2(n_448),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_699),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_SL g903 ( 
.A(n_634),
.B(n_476),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_700),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_711),
.Y(n_905)
);

INVx2_ASAP7_75t_SL g906 ( 
.A(n_649),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_650),
.B(n_448),
.Y(n_907)
);

BUFx2_ASAP7_75t_L g908 ( 
.A(n_746),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_652),
.B(n_448),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_718),
.Y(n_910)
);

AOI22xp33_ASAP7_75t_SL g911 ( 
.A1(n_603),
.A2(n_733),
.B1(n_738),
.B2(n_737),
.Y(n_911)
);

BUFx2_ASAP7_75t_L g912 ( 
.A(n_657),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_701),
.Y(n_913)
);

OR2x6_ASAP7_75t_L g914 ( 
.A(n_753),
.B(n_552),
.Y(n_914)
);

AND2x6_ASAP7_75t_L g915 ( 
.A(n_726),
.B(n_552),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_691),
.B(n_552),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_SL g917 ( 
.A(n_719),
.B(n_552),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_704),
.B(n_30),
.Y(n_918)
);

INVx2_ASAP7_75t_SL g919 ( 
.A(n_709),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_676),
.A2(n_30),
.B(n_32),
.Y(n_920)
);

OAI22xp5_ASAP7_75t_L g921 ( 
.A1(n_676),
.A2(n_47),
.B1(n_35),
.B2(n_36),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_722),
.B(n_34),
.Y(n_922)
);

INVx4_ASAP7_75t_L g923 ( 
.A(n_671),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_SL g924 ( 
.A(n_727),
.B(n_38),
.Y(n_924)
);

INVx2_ASAP7_75t_SL g925 ( 
.A(n_709),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_731),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_756),
.Y(n_927)
);

NOR3xp33_ASAP7_75t_SL g928 ( 
.A(n_737),
.B(n_38),
.C(n_39),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_717),
.B(n_39),
.Y(n_929)
);

INVxp67_ASAP7_75t_SL g930 ( 
.A(n_717),
.Y(n_930)
);

BUFx6f_ASAP7_75t_L g931 ( 
.A(n_614),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_661),
.Y(n_932)
);

BUFx4f_ASAP7_75t_L g933 ( 
.A(n_760),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_662),
.Y(n_934)
);

INVx2_ASAP7_75t_SL g935 ( 
.A(n_750),
.Y(n_935)
);

NOR3xp33_ASAP7_75t_L g936 ( 
.A(n_642),
.B(n_46),
.C(n_47),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_660),
.B(n_46),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_678),
.B(n_703),
.Y(n_938)
);

OR2x6_ASAP7_75t_L g939 ( 
.A(n_762),
.B(n_755),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_697),
.A2(n_682),
.B(n_679),
.Y(n_940)
);

AOI22xp5_ASAP7_75t_L g941 ( 
.A1(n_660),
.A2(n_682),
.B1(n_679),
.B2(n_684),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_627),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_822),
.B(n_684),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_885),
.A2(n_638),
.B(n_743),
.Y(n_944)
);

INVx3_ASAP7_75t_L g945 ( 
.A(n_780),
.Y(n_945)
);

NAND2x1p5_ASAP7_75t_L g946 ( 
.A(n_783),
.B(n_743),
.Y(n_946)
);

AND2x4_ASAP7_75t_L g947 ( 
.A(n_797),
.B(n_843),
.Y(n_947)
);

A2O1A1Ixp33_ASAP7_75t_L g948 ( 
.A1(n_861),
.A2(n_938),
.B(n_764),
.C(n_826),
.Y(n_948)
);

OR2x6_ASAP7_75t_L g949 ( 
.A(n_794),
.B(n_762),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_778),
.B(n_755),
.Y(n_950)
);

OR2x2_ASAP7_75t_L g951 ( 
.A(n_770),
.B(n_659),
.Y(n_951)
);

CKINVDCx20_ASAP7_75t_R g952 ( 
.A(n_794),
.Y(n_952)
);

AND2x2_ASAP7_75t_L g953 ( 
.A(n_823),
.B(n_753),
.Y(n_953)
);

A2O1A1Ixp33_ASAP7_75t_L g954 ( 
.A1(n_938),
.A2(n_716),
.B(n_754),
.C(n_761),
.Y(n_954)
);

BUFx3_ASAP7_75t_L g955 ( 
.A(n_794),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_826),
.B(n_628),
.Y(n_956)
);

AOI22xp5_ASAP7_75t_L g957 ( 
.A1(n_801),
.A2(n_624),
.B1(n_636),
.B2(n_602),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_807),
.B(n_624),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_R g959 ( 
.A(n_801),
.B(n_639),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_L g960 ( 
.A(n_893),
.B(n_639),
.Y(n_960)
);

OAI22xp5_ASAP7_75t_L g961 ( 
.A1(n_911),
.A2(n_628),
.B1(n_645),
.B2(n_706),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_763),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_893),
.B(n_856),
.Y(n_963)
);

AOI22xp33_ASAP7_75t_L g964 ( 
.A1(n_922),
.A2(n_924),
.B1(n_898),
.B2(n_937),
.Y(n_964)
);

BUFx8_ASAP7_75t_SL g965 ( 
.A(n_848),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_775),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_842),
.A2(n_847),
.B(n_809),
.Y(n_967)
);

NOR2xp33_ASAP7_75t_L g968 ( 
.A(n_908),
.B(n_792),
.Y(n_968)
);

INVx3_ASAP7_75t_SL g969 ( 
.A(n_774),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_890),
.B(n_894),
.Y(n_970)
);

HB1xp67_ASAP7_75t_L g971 ( 
.A(n_866),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_842),
.A2(n_847),
.B(n_875),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_897),
.B(n_879),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_880),
.B(n_902),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_R g975 ( 
.A(n_795),
.B(n_771),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_776),
.Y(n_976)
);

OAI22xp5_ASAP7_75t_SL g977 ( 
.A1(n_884),
.A2(n_867),
.B1(n_774),
.B2(n_781),
.Y(n_977)
);

OAI21xp5_ASAP7_75t_L g978 ( 
.A1(n_859),
.A2(n_911),
.B(n_834),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_785),
.Y(n_979)
);

OAI22xp5_ASAP7_75t_L g980 ( 
.A1(n_867),
.A2(n_901),
.B1(n_841),
.B2(n_817),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_913),
.B(n_860),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_SL g982 ( 
.A(n_765),
.B(n_870),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_SL g983 ( 
.A(n_766),
.B(n_768),
.Y(n_983)
);

INVx4_ASAP7_75t_L g984 ( 
.A(n_783),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_L g985 ( 
.A(n_906),
.B(n_843),
.Y(n_985)
);

O2A1O1Ixp5_ASAP7_75t_L g986 ( 
.A1(n_875),
.A2(n_849),
.B(n_814),
.C(n_869),
.Y(n_986)
);

AND3x1_ASAP7_75t_SL g987 ( 
.A(n_811),
.B(n_851),
.C(n_845),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_940),
.A2(n_849),
.B(n_769),
.Y(n_988)
);

A2O1A1Ixp33_ASAP7_75t_L g989 ( 
.A1(n_859),
.A2(n_941),
.B(n_864),
.C(n_922),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_850),
.B(n_812),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_816),
.A2(n_836),
.B(n_819),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_783),
.A2(n_819),
.B(n_821),
.Y(n_992)
);

O2A1O1Ixp33_ASAP7_75t_L g993 ( 
.A1(n_924),
.A2(n_921),
.B(n_936),
.C(n_918),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_SL g994 ( 
.A(n_866),
.B(n_783),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_788),
.B(n_781),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_772),
.Y(n_996)
);

BUFx2_ASAP7_75t_L g997 ( 
.A(n_771),
.Y(n_997)
);

BUFx6f_ASAP7_75t_L g998 ( 
.A(n_780),
.Y(n_998)
);

A2O1A1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_895),
.A2(n_777),
.B(n_779),
.C(n_782),
.Y(n_999)
);

BUFx6f_ASAP7_75t_L g1000 ( 
.A(n_780),
.Y(n_1000)
);

HB1xp67_ASAP7_75t_L g1001 ( 
.A(n_830),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_830),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_R g1003 ( 
.A(n_780),
.B(n_820),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_818),
.Y(n_1004)
);

AOI22x1_ASAP7_75t_L g1005 ( 
.A1(n_935),
.A2(n_934),
.B1(n_932),
.B2(n_942),
.Y(n_1005)
);

OAI22xp5_ASAP7_75t_L g1006 ( 
.A1(n_901),
.A2(n_841),
.B1(n_817),
.B2(n_833),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_789),
.B(n_793),
.Y(n_1007)
);

A2O1A1Ixp33_ASAP7_75t_L g1008 ( 
.A1(n_839),
.A2(n_871),
.B(n_925),
.C(n_919),
.Y(n_1008)
);

O2A1O1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_936),
.A2(n_929),
.B(n_808),
.C(n_804),
.Y(n_1009)
);

OAI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_834),
.A2(n_767),
.B(n_874),
.Y(n_1010)
);

BUFx2_ASAP7_75t_L g1011 ( 
.A(n_774),
.Y(n_1011)
);

OR2x6_ASAP7_75t_L g1012 ( 
.A(n_881),
.B(n_820),
.Y(n_1012)
);

OAI22x1_ASAP7_75t_L g1013 ( 
.A1(n_891),
.A2(n_912),
.B1(n_903),
.B2(n_878),
.Y(n_1013)
);

BUFx4f_ASAP7_75t_L g1014 ( 
.A(n_820),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_786),
.Y(n_1015)
);

A2O1A1Ixp33_ASAP7_75t_L g1016 ( 
.A1(n_839),
.A2(n_871),
.B(n_887),
.C(n_900),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_790),
.Y(n_1017)
);

NOR2x1_ASAP7_75t_R g1018 ( 
.A(n_881),
.B(n_900),
.Y(n_1018)
);

NOR2x1_ASAP7_75t_L g1019 ( 
.A(n_923),
.B(n_903),
.Y(n_1019)
);

A2O1A1Ixp33_ASAP7_75t_L g1020 ( 
.A1(n_773),
.A2(n_930),
.B(n_787),
.C(n_920),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_930),
.B(n_800),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_805),
.B(n_806),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_829),
.A2(n_892),
.B(n_896),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_907),
.A2(n_909),
.B(n_837),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_933),
.B(n_820),
.Y(n_1025)
);

BUFx2_ASAP7_75t_L g1026 ( 
.A(n_835),
.Y(n_1026)
);

AO21x1_ASAP7_75t_L g1027 ( 
.A1(n_863),
.A2(n_917),
.B(n_767),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_882),
.B(n_889),
.Y(n_1028)
);

INVxp67_ASAP7_75t_L g1029 ( 
.A(n_835),
.Y(n_1029)
);

BUFx6f_ASAP7_75t_L g1030 ( 
.A(n_852),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_872),
.Y(n_1031)
);

AOI221xp5_ASAP7_75t_L g1032 ( 
.A1(n_884),
.A2(n_928),
.B1(n_838),
.B2(n_815),
.C(n_799),
.Y(n_1032)
);

OAI22xp5_ASAP7_75t_SL g1033 ( 
.A1(n_939),
.A2(n_914),
.B1(n_853),
.B2(n_833),
.Y(n_1033)
);

INVx3_ASAP7_75t_SL g1034 ( 
.A(n_939),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_810),
.A2(n_827),
.B(n_840),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_791),
.Y(n_1036)
);

INVx4_ASAP7_75t_L g1037 ( 
.A(n_852),
.Y(n_1037)
);

BUFx6f_ASAP7_75t_L g1038 ( 
.A(n_852),
.Y(n_1038)
);

INVx3_ASAP7_75t_L g1039 ( 
.A(n_868),
.Y(n_1039)
);

INVx5_ASAP7_75t_L g1040 ( 
.A(n_852),
.Y(n_1040)
);

NOR3xp33_ASAP7_75t_SL g1041 ( 
.A(n_784),
.B(n_802),
.C(n_796),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_798),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_L g1043 ( 
.A(n_939),
.B(n_865),
.Y(n_1043)
);

AND2x2_ASAP7_75t_L g1044 ( 
.A(n_928),
.B(n_905),
.Y(n_1044)
);

A2O1A1Ixp33_ASAP7_75t_L g1045 ( 
.A1(n_825),
.A2(n_854),
.B(n_927),
.C(n_883),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_L g1046 ( 
.A(n_813),
.B(n_865),
.Y(n_1046)
);

OR2x6_ASAP7_75t_L g1047 ( 
.A(n_868),
.B(n_923),
.Y(n_1047)
);

A2O1A1Ixp33_ASAP7_75t_L g1048 ( 
.A1(n_855),
.A2(n_904),
.B(n_899),
.C(n_888),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_SL g1049 ( 
.A(n_868),
.B(n_857),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_803),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_844),
.Y(n_1051)
);

BUFx6f_ASAP7_75t_L g1052 ( 
.A(n_857),
.Y(n_1052)
);

NOR2xp67_ASAP7_75t_SL g1053 ( 
.A(n_868),
.B(n_862),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_828),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_831),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_SL g1056 ( 
.A(n_857),
.B(n_862),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_832),
.B(n_813),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_SL g1058 ( 
.A(n_862),
.B(n_926),
.Y(n_1058)
);

OAI22xp5_ASAP7_75t_L g1059 ( 
.A1(n_914),
.A2(n_876),
.B1(n_862),
.B2(n_846),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_910),
.B(n_916),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_858),
.Y(n_1061)
);

NOR2xp33_ASAP7_75t_L g1062 ( 
.A(n_914),
.B(n_784),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_873),
.B(n_877),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_L g1064 ( 
.A(n_802),
.B(n_824),
.Y(n_1064)
);

INVxp67_ASAP7_75t_L g1065 ( 
.A(n_824),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_R g1066 ( 
.A(n_931),
.B(n_915),
.Y(n_1066)
);

OR2x6_ASAP7_75t_L g1067 ( 
.A(n_876),
.B(n_931),
.Y(n_1067)
);

A2O1A1Ixp33_ASAP7_75t_L g1068 ( 
.A1(n_931),
.A2(n_822),
.B(n_630),
.C(n_861),
.Y(n_1068)
);

INVx6_ASAP7_75t_L g1069 ( 
.A(n_931),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_915),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_915),
.B(n_822),
.Y(n_1071)
);

BUFx6f_ASAP7_75t_L g1072 ( 
.A(n_915),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_915),
.B(n_822),
.Y(n_1073)
);

INVx3_ASAP7_75t_L g1074 ( 
.A(n_780),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_885),
.A2(n_503),
.B(n_886),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_885),
.A2(n_503),
.B(n_886),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_794),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_763),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_822),
.B(n_826),
.Y(n_1079)
);

O2A1O1Ixp33_ASAP7_75t_L g1080 ( 
.A1(n_861),
.A2(n_630),
.B(n_822),
.C(n_826),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_1028),
.Y(n_1081)
);

AO31x2_ASAP7_75t_L g1082 ( 
.A1(n_1027),
.A2(n_954),
.A3(n_989),
.B(n_961),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_963),
.B(n_1079),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_970),
.B(n_973),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_974),
.B(n_981),
.Y(n_1085)
);

INVxp67_ASAP7_75t_SL g1086 ( 
.A(n_1053),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_981),
.B(n_948),
.Y(n_1087)
);

AND2x4_ASAP7_75t_L g1088 ( 
.A(n_947),
.B(n_1011),
.Y(n_1088)
);

OAI21xp33_ASAP7_75t_SL g1089 ( 
.A1(n_980),
.A2(n_1006),
.B(n_978),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_972),
.A2(n_944),
.B(n_1076),
.Y(n_1090)
);

AND2x4_ASAP7_75t_L g1091 ( 
.A(n_1012),
.B(n_955),
.Y(n_1091)
);

A2O1A1Ixp33_ASAP7_75t_L g1092 ( 
.A1(n_1080),
.A2(n_993),
.B(n_1068),
.C(n_978),
.Y(n_1092)
);

OR2x2_ASAP7_75t_L g1093 ( 
.A(n_971),
.B(n_951),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_1023),
.A2(n_1024),
.B(n_967),
.Y(n_1094)
);

NOR4xp25_ASAP7_75t_L g1095 ( 
.A(n_964),
.B(n_1009),
.C(n_980),
.D(n_961),
.Y(n_1095)
);

OA21x2_ASAP7_75t_L g1096 ( 
.A1(n_986),
.A2(n_1010),
.B(n_1063),
.Y(n_1096)
);

AOI21x1_ASAP7_75t_L g1097 ( 
.A1(n_983),
.A2(n_1063),
.B(n_1021),
.Y(n_1097)
);

AOI21xp33_ASAP7_75t_L g1098 ( 
.A1(n_943),
.A2(n_977),
.B(n_958),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_SL g1099 ( 
.A1(n_1016),
.A2(n_1006),
.B(n_1067),
.Y(n_1099)
);

INVx4_ASAP7_75t_L g1100 ( 
.A(n_1014),
.Y(n_1100)
);

A2O1A1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_960),
.A2(n_999),
.B(n_1043),
.C(n_1008),
.Y(n_1101)
);

AOI22xp5_ASAP7_75t_L g1102 ( 
.A1(n_950),
.A2(n_995),
.B1(n_1033),
.B2(n_956),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_990),
.B(n_985),
.Y(n_1103)
);

AOI221xp5_ASAP7_75t_SL g1104 ( 
.A1(n_1032),
.A2(n_1013),
.B1(n_1044),
.B2(n_1061),
.C(n_1071),
.Y(n_1104)
);

OAI21x1_ASAP7_75t_SL g1105 ( 
.A1(n_1073),
.A2(n_1005),
.B(n_1059),
.Y(n_1105)
);

A2O1A1Ixp33_ASAP7_75t_L g1106 ( 
.A1(n_957),
.A2(n_1073),
.B(n_1062),
.C(n_1064),
.Y(n_1106)
);

AOI211x1_ASAP7_75t_L g1107 ( 
.A1(n_1007),
.A2(n_982),
.B(n_953),
.C(n_1002),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_L g1108 ( 
.A(n_1031),
.B(n_968),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_1004),
.Y(n_1109)
);

AOI221x1_ASAP7_75t_L g1110 ( 
.A1(n_1059),
.A2(n_1010),
.B1(n_1020),
.B2(n_1022),
.C(n_1070),
.Y(n_1110)
);

AO21x1_ASAP7_75t_L g1111 ( 
.A1(n_946),
.A2(n_1035),
.B(n_1060),
.Y(n_1111)
);

BUFx4_ASAP7_75t_SL g1112 ( 
.A(n_952),
.Y(n_1112)
);

BUFx6f_ASAP7_75t_L g1113 ( 
.A(n_998),
.Y(n_1113)
);

INVx4_ASAP7_75t_L g1114 ( 
.A(n_1014),
.Y(n_1114)
);

OAI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_1045),
.A2(n_1048),
.B(n_992),
.Y(n_1115)
);

A2O1A1Ixp33_ASAP7_75t_L g1116 ( 
.A1(n_1065),
.A2(n_1041),
.B(n_1019),
.C(n_1046),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_1034),
.B(n_1001),
.Y(n_1117)
);

OAI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_946),
.A2(n_1057),
.B(n_1054),
.Y(n_1118)
);

OAI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_1057),
.A2(n_1055),
.B(n_996),
.Y(n_1119)
);

INVx3_ASAP7_75t_L g1120 ( 
.A(n_984),
.Y(n_1120)
);

BUFx2_ASAP7_75t_L g1121 ( 
.A(n_975),
.Y(n_1121)
);

AND2x2_ASAP7_75t_L g1122 ( 
.A(n_949),
.B(n_969),
.Y(n_1122)
);

OAI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_1051),
.A2(n_1078),
.B(n_976),
.Y(n_1123)
);

AO21x2_ASAP7_75t_L g1124 ( 
.A1(n_959),
.A2(n_1066),
.B(n_1058),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_962),
.B(n_966),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1015),
.Y(n_1126)
);

AOI31xp33_ASAP7_75t_L g1127 ( 
.A1(n_1018),
.A2(n_1029),
.A3(n_1077),
.B(n_994),
.Y(n_1127)
);

OAI21x1_ASAP7_75t_L g1128 ( 
.A1(n_1056),
.A2(n_1049),
.B(n_1050),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1017),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_1067),
.A2(n_984),
.B(n_1040),
.Y(n_1130)
);

AND2x4_ASAP7_75t_L g1131 ( 
.A(n_949),
.B(n_1047),
.Y(n_1131)
);

BUFx6f_ASAP7_75t_L g1132 ( 
.A(n_998),
.Y(n_1132)
);

A2O1A1Ixp33_ASAP7_75t_L g1133 ( 
.A1(n_1036),
.A2(n_1042),
.B(n_1025),
.C(n_1039),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_1047),
.B(n_945),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_945),
.B(n_1074),
.Y(n_1135)
);

BUFx6f_ASAP7_75t_L g1136 ( 
.A(n_998),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1074),
.B(n_1052),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1030),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1030),
.Y(n_1139)
);

A2O1A1Ixp33_ASAP7_75t_L g1140 ( 
.A1(n_1072),
.A2(n_987),
.B(n_1040),
.C(n_1052),
.Y(n_1140)
);

NAND2x1_ASAP7_75t_L g1141 ( 
.A(n_1069),
.B(n_1067),
.Y(n_1141)
);

A2O1A1Ixp33_ASAP7_75t_L g1142 ( 
.A1(n_1072),
.A2(n_1040),
.B(n_1052),
.C(n_1000),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_1040),
.A2(n_1072),
.B(n_1037),
.Y(n_1143)
);

A2O1A1Ixp33_ASAP7_75t_L g1144 ( 
.A1(n_1000),
.A2(n_1030),
.B(n_1038),
.C(n_1026),
.Y(n_1144)
);

O2A1O1Ixp5_ASAP7_75t_SL g1145 ( 
.A1(n_965),
.A2(n_1003),
.B(n_1069),
.C(n_1038),
.Y(n_1145)
);

AO31x2_ASAP7_75t_L g1146 ( 
.A1(n_1037),
.A2(n_1000),
.A3(n_1038),
.B(n_1027),
.Y(n_1146)
);

AOI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_977),
.A2(n_822),
.B1(n_630),
.B2(n_826),
.Y(n_1147)
);

OA21x2_ASAP7_75t_L g1148 ( 
.A1(n_978),
.A2(n_986),
.B(n_1010),
.Y(n_1148)
);

BUFx2_ASAP7_75t_L g1149 ( 
.A(n_975),
.Y(n_1149)
);

OAI21x1_ASAP7_75t_L g1150 ( 
.A1(n_991),
.A2(n_834),
.B(n_988),
.Y(n_1150)
);

O2A1O1Ixp5_ASAP7_75t_SL g1151 ( 
.A1(n_983),
.A2(n_739),
.B(n_924),
.C(n_922),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_963),
.B(n_822),
.Y(n_1152)
);

CKINVDCx8_ASAP7_75t_R g1153 ( 
.A(n_1077),
.Y(n_1153)
);

OA21x2_ASAP7_75t_L g1154 ( 
.A1(n_978),
.A2(n_986),
.B(n_1010),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_963),
.B(n_822),
.Y(n_1155)
);

OA21x2_ASAP7_75t_L g1156 ( 
.A1(n_978),
.A2(n_986),
.B(n_1010),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_963),
.B(n_822),
.Y(n_1157)
);

OAI21x1_ASAP7_75t_L g1158 ( 
.A1(n_991),
.A2(n_834),
.B(n_988),
.Y(n_1158)
);

AOI21x1_ASAP7_75t_L g1159 ( 
.A1(n_983),
.A2(n_972),
.B(n_944),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_972),
.A2(n_944),
.B(n_1075),
.Y(n_1160)
);

INVx2_ASAP7_75t_SL g1161 ( 
.A(n_997),
.Y(n_1161)
);

OAI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_978),
.A2(n_989),
.B(n_948),
.Y(n_1162)
);

NOR2xp33_ASAP7_75t_L g1163 ( 
.A(n_1079),
.B(n_822),
.Y(n_1163)
);

OR2x6_ASAP7_75t_L g1164 ( 
.A(n_1012),
.B(n_794),
.Y(n_1164)
);

A2O1A1Ixp33_ASAP7_75t_L g1165 ( 
.A1(n_1080),
.A2(n_822),
.B(n_764),
.C(n_993),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_963),
.B(n_822),
.Y(n_1166)
);

INVx4_ASAP7_75t_L g1167 ( 
.A(n_1014),
.Y(n_1167)
);

A2O1A1Ixp33_ASAP7_75t_L g1168 ( 
.A1(n_1080),
.A2(n_822),
.B(n_764),
.C(n_993),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_972),
.A2(n_944),
.B(n_1075),
.Y(n_1169)
);

AOI21x1_ASAP7_75t_SL g1170 ( 
.A1(n_1073),
.A2(n_861),
.B(n_822),
.Y(n_1170)
);

BUFx6f_ASAP7_75t_L g1171 ( 
.A(n_998),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1028),
.Y(n_1172)
);

AOI21x1_ASAP7_75t_L g1173 ( 
.A1(n_983),
.A2(n_972),
.B(n_944),
.Y(n_1173)
);

AO31x2_ASAP7_75t_L g1174 ( 
.A1(n_1027),
.A2(n_954),
.A3(n_814),
.B(n_989),
.Y(n_1174)
);

OAI21x1_ASAP7_75t_L g1175 ( 
.A1(n_991),
.A2(n_834),
.B(n_988),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_979),
.Y(n_1176)
);

NOR2xp33_ASAP7_75t_L g1177 ( 
.A(n_1079),
.B(n_822),
.Y(n_1177)
);

INVx2_ASAP7_75t_SL g1178 ( 
.A(n_997),
.Y(n_1178)
);

INVx2_ASAP7_75t_SL g1179 ( 
.A(n_997),
.Y(n_1179)
);

HB1xp67_ASAP7_75t_L g1180 ( 
.A(n_971),
.Y(n_1180)
);

OAI21x1_ASAP7_75t_L g1181 ( 
.A1(n_991),
.A2(n_834),
.B(n_988),
.Y(n_1181)
);

BUFx3_ASAP7_75t_L g1182 ( 
.A(n_955),
.Y(n_1182)
);

HB1xp67_ASAP7_75t_L g1183 ( 
.A(n_971),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1028),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_972),
.A2(n_944),
.B(n_1075),
.Y(n_1185)
);

NAND3xp33_ASAP7_75t_L g1186 ( 
.A(n_1080),
.B(n_630),
.C(n_822),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1028),
.Y(n_1187)
);

OAI21x1_ASAP7_75t_L g1188 ( 
.A1(n_991),
.A2(n_834),
.B(n_988),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1028),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1028),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_972),
.A2(n_944),
.B(n_1075),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_SL g1192 ( 
.A(n_1031),
.B(n_822),
.Y(n_1192)
);

BUFx10_ASAP7_75t_L g1193 ( 
.A(n_968),
.Y(n_1193)
);

INVx1_ASAP7_75t_SL g1194 ( 
.A(n_975),
.Y(n_1194)
);

OAI21x1_ASAP7_75t_L g1195 ( 
.A1(n_991),
.A2(n_834),
.B(n_988),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_963),
.B(n_822),
.Y(n_1196)
);

BUFx6f_ASAP7_75t_L g1197 ( 
.A(n_998),
.Y(n_1197)
);

OAI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_978),
.A2(n_989),
.B(n_948),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_972),
.A2(n_944),
.B(n_1075),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1028),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_948),
.B(n_981),
.Y(n_1201)
);

AND2x2_ASAP7_75t_L g1202 ( 
.A(n_950),
.B(n_778),
.Y(n_1202)
);

BUFx2_ASAP7_75t_L g1203 ( 
.A(n_975),
.Y(n_1203)
);

AND2x4_ASAP7_75t_L g1204 ( 
.A(n_947),
.B(n_881),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_972),
.A2(n_944),
.B(n_1075),
.Y(n_1205)
);

BUFx2_ASAP7_75t_L g1206 ( 
.A(n_975),
.Y(n_1206)
);

OAI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_978),
.A2(n_989),
.B(n_948),
.Y(n_1207)
);

NOR2xp33_ASAP7_75t_L g1208 ( 
.A(n_1079),
.B(n_822),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_963),
.B(n_822),
.Y(n_1209)
);

OAI22xp5_ASAP7_75t_SL g1210 ( 
.A1(n_977),
.A2(n_520),
.B1(n_884),
.B2(n_395),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1028),
.Y(n_1211)
);

AOI21x1_ASAP7_75t_L g1212 ( 
.A1(n_983),
.A2(n_972),
.B(n_944),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_963),
.B(n_822),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_972),
.A2(n_944),
.B(n_1075),
.Y(n_1214)
);

OAI22xp5_ASAP7_75t_L g1215 ( 
.A1(n_1147),
.A2(n_1085),
.B1(n_1084),
.B2(n_1210),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_L g1216 ( 
.A1(n_1150),
.A2(n_1175),
.B(n_1158),
.Y(n_1216)
);

OAI21x1_ASAP7_75t_L g1217 ( 
.A1(n_1181),
.A2(n_1195),
.B(n_1188),
.Y(n_1217)
);

INVxp67_ASAP7_75t_L g1218 ( 
.A(n_1108),
.Y(n_1218)
);

OA21x2_ASAP7_75t_L g1219 ( 
.A1(n_1110),
.A2(n_1198),
.B(n_1162),
.Y(n_1219)
);

OAI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1186),
.A2(n_1168),
.B(n_1165),
.Y(n_1220)
);

AND2x2_ASAP7_75t_L g1221 ( 
.A(n_1202),
.B(n_1163),
.Y(n_1221)
);

AOI21x1_ASAP7_75t_L g1222 ( 
.A1(n_1097),
.A2(n_1173),
.B(n_1159),
.Y(n_1222)
);

OAI21x1_ASAP7_75t_L g1223 ( 
.A1(n_1094),
.A2(n_1214),
.B(n_1169),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_1112),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_1153),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1152),
.B(n_1155),
.Y(n_1226)
);

AOI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1090),
.A2(n_1160),
.B(n_1191),
.Y(n_1227)
);

HB1xp67_ASAP7_75t_L g1228 ( 
.A(n_1082),
.Y(n_1228)
);

NAND2x1p5_ASAP7_75t_L g1229 ( 
.A(n_1141),
.B(n_1131),
.Y(n_1229)
);

BUFx3_ASAP7_75t_L g1230 ( 
.A(n_1204),
.Y(n_1230)
);

OAI21x1_ASAP7_75t_L g1231 ( 
.A1(n_1185),
.A2(n_1199),
.B(n_1205),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1126),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1207),
.A2(n_1087),
.B(n_1201),
.Y(n_1233)
);

AOI21xp33_ASAP7_75t_L g1234 ( 
.A1(n_1186),
.A2(n_1147),
.B(n_1177),
.Y(n_1234)
);

OAI21x1_ASAP7_75t_L g1235 ( 
.A1(n_1212),
.A2(n_1115),
.B(n_1170),
.Y(n_1235)
);

A2O1A1Ixp33_ASAP7_75t_L g1236 ( 
.A1(n_1089),
.A2(n_1092),
.B(n_1098),
.C(n_1208),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1157),
.B(n_1166),
.Y(n_1237)
);

BUFx2_ASAP7_75t_L g1238 ( 
.A(n_1121),
.Y(n_1238)
);

NOR2x1_ASAP7_75t_L g1239 ( 
.A(n_1100),
.B(n_1114),
.Y(n_1239)
);

OAI21x1_ASAP7_75t_L g1240 ( 
.A1(n_1115),
.A2(n_1105),
.B(n_1151),
.Y(n_1240)
);

OAI21x1_ASAP7_75t_L g1241 ( 
.A1(n_1128),
.A2(n_1118),
.B(n_1111),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1129),
.Y(n_1242)
);

OAI21x1_ASAP7_75t_L g1243 ( 
.A1(n_1118),
.A2(n_1119),
.B(n_1096),
.Y(n_1243)
);

AOI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1201),
.A2(n_1099),
.B(n_1101),
.Y(n_1244)
);

CKINVDCx12_ASAP7_75t_R g1245 ( 
.A(n_1164),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1196),
.B(n_1209),
.Y(n_1246)
);

OAI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1106),
.A2(n_1098),
.B(n_1213),
.Y(n_1247)
);

AO32x2_ASAP7_75t_L g1248 ( 
.A1(n_1210),
.A2(n_1095),
.A3(n_1148),
.B1(n_1154),
.B2(n_1156),
.Y(n_1248)
);

INVx1_ASAP7_75t_SL g1249 ( 
.A(n_1194),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_1176),
.Y(n_1250)
);

OAI22xp5_ASAP7_75t_L g1251 ( 
.A1(n_1083),
.A2(n_1103),
.B1(n_1102),
.B2(n_1211),
.Y(n_1251)
);

OA21x2_ASAP7_75t_L g1252 ( 
.A1(n_1104),
.A2(n_1119),
.B(n_1102),
.Y(n_1252)
);

OA21x2_ASAP7_75t_L g1253 ( 
.A1(n_1104),
.A2(n_1123),
.B(n_1116),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_1088),
.B(n_1081),
.Y(n_1254)
);

OAI222xp33_ASAP7_75t_L g1255 ( 
.A1(n_1192),
.A2(n_1093),
.B1(n_1172),
.B2(n_1184),
.C1(n_1187),
.C2(n_1200),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1189),
.Y(n_1256)
);

OAI21x1_ASAP7_75t_L g1257 ( 
.A1(n_1096),
.A2(n_1130),
.B(n_1123),
.Y(n_1257)
);

CKINVDCx16_ASAP7_75t_R g1258 ( 
.A(n_1182),
.Y(n_1258)
);

AND2x2_ASAP7_75t_L g1259 ( 
.A(n_1190),
.B(n_1194),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1125),
.Y(n_1260)
);

OAI21x1_ASAP7_75t_L g1261 ( 
.A1(n_1148),
.A2(n_1154),
.B(n_1156),
.Y(n_1261)
);

INVx1_ASAP7_75t_SL g1262 ( 
.A(n_1149),
.Y(n_1262)
);

OAI21x1_ASAP7_75t_L g1263 ( 
.A1(n_1143),
.A2(n_1134),
.B(n_1135),
.Y(n_1263)
);

AOI22xp33_ASAP7_75t_SL g1264 ( 
.A1(n_1203),
.A2(n_1206),
.B1(n_1122),
.B2(n_1193),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1095),
.B(n_1183),
.Y(n_1265)
);

OA21x2_ASAP7_75t_L g1266 ( 
.A1(n_1133),
.A2(n_1140),
.B(n_1082),
.Y(n_1266)
);

A2O1A1Ixp33_ASAP7_75t_L g1267 ( 
.A1(n_1144),
.A2(n_1127),
.B(n_1142),
.C(n_1086),
.Y(n_1267)
);

AOI21x1_ASAP7_75t_L g1268 ( 
.A1(n_1137),
.A2(n_1138),
.B(n_1139),
.Y(n_1268)
);

OAI22xp5_ASAP7_75t_L g1269 ( 
.A1(n_1107),
.A2(n_1127),
.B1(n_1164),
.B2(n_1117),
.Y(n_1269)
);

AND2x2_ASAP7_75t_L g1270 ( 
.A(n_1180),
.B(n_1178),
.Y(n_1270)
);

AOI22xp33_ASAP7_75t_L g1271 ( 
.A1(n_1124),
.A2(n_1193),
.B1(n_1091),
.B2(n_1161),
.Y(n_1271)
);

NOR2xp33_ASAP7_75t_L g1272 ( 
.A(n_1179),
.B(n_1167),
.Y(n_1272)
);

AO21x2_ASAP7_75t_L g1273 ( 
.A1(n_1174),
.A2(n_1082),
.B(n_1146),
.Y(n_1273)
);

OAI21x1_ASAP7_75t_SL g1274 ( 
.A1(n_1167),
.A2(n_1145),
.B(n_1146),
.Y(n_1274)
);

CKINVDCx11_ASAP7_75t_R g1275 ( 
.A(n_1113),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1146),
.Y(n_1276)
);

OAI22x1_ASAP7_75t_L g1277 ( 
.A1(n_1120),
.A2(n_1174),
.B1(n_1132),
.B2(n_1136),
.Y(n_1277)
);

OAI22xp5_ASAP7_75t_L g1278 ( 
.A1(n_1113),
.A2(n_1132),
.B1(n_1136),
.B2(n_1171),
.Y(n_1278)
);

AO21x2_ASAP7_75t_L g1279 ( 
.A1(n_1174),
.A2(n_1113),
.B(n_1132),
.Y(n_1279)
);

AOI21xp33_ASAP7_75t_L g1280 ( 
.A1(n_1136),
.A2(n_1171),
.B(n_1197),
.Y(n_1280)
);

INVx2_ASAP7_75t_L g1281 ( 
.A(n_1171),
.Y(n_1281)
);

OA21x2_ASAP7_75t_L g1282 ( 
.A1(n_1197),
.A2(n_1110),
.B(n_1162),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_1197),
.A2(n_1210),
.B1(n_822),
.B2(n_884),
.Y(n_1283)
);

OAI22xp5_ASAP7_75t_SL g1284 ( 
.A1(n_1210),
.A2(n_487),
.B1(n_480),
.B2(n_884),
.Y(n_1284)
);

AOI22xp33_ASAP7_75t_L g1285 ( 
.A1(n_1210),
.A2(n_822),
.B1(n_884),
.B2(n_977),
.Y(n_1285)
);

AOI21x1_ASAP7_75t_L g1286 ( 
.A1(n_1097),
.A2(n_972),
.B(n_983),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1109),
.Y(n_1287)
);

NAND3xp33_ASAP7_75t_L g1288 ( 
.A(n_1186),
.B(n_630),
.C(n_822),
.Y(n_1288)
);

A2O1A1Ixp33_ASAP7_75t_L g1289 ( 
.A1(n_1162),
.A2(n_980),
.B(n_1207),
.C(n_1198),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1202),
.B(n_1163),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1152),
.B(n_1157),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1109),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1109),
.Y(n_1293)
);

OA21x2_ASAP7_75t_L g1294 ( 
.A1(n_1110),
.A2(n_1198),
.B(n_1162),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_1112),
.Y(n_1295)
);

NAND2x1p5_ASAP7_75t_L g1296 ( 
.A(n_1141),
.B(n_1053),
.Y(n_1296)
);

NOR2xp67_ASAP7_75t_L g1297 ( 
.A(n_1108),
.B(n_619),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1109),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1109),
.Y(n_1299)
);

NAND2x1p5_ASAP7_75t_L g1300 ( 
.A(n_1141),
.B(n_1053),
.Y(n_1300)
);

NOR2xp33_ASAP7_75t_L g1301 ( 
.A(n_1210),
.B(n_822),
.Y(n_1301)
);

A2O1A1Ixp33_ASAP7_75t_L g1302 ( 
.A1(n_1162),
.A2(n_980),
.B(n_1207),
.C(n_1198),
.Y(n_1302)
);

NAND2x1p5_ASAP7_75t_L g1303 ( 
.A(n_1141),
.B(n_1053),
.Y(n_1303)
);

NOR2xp33_ASAP7_75t_SL g1304 ( 
.A(n_1153),
.B(n_713),
.Y(n_1304)
);

OR2x2_ASAP7_75t_L g1305 ( 
.A(n_1152),
.B(n_1155),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1202),
.B(n_1163),
.Y(n_1306)
);

OR2x6_ASAP7_75t_L g1307 ( 
.A(n_1099),
.B(n_1164),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1109),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1109),
.Y(n_1309)
);

OAI21x1_ASAP7_75t_L g1310 ( 
.A1(n_1150),
.A2(n_1175),
.B(n_1158),
.Y(n_1310)
);

AO21x2_ASAP7_75t_L g1311 ( 
.A1(n_1094),
.A2(n_978),
.B(n_1090),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1152),
.B(n_1157),
.Y(n_1312)
);

OR2x6_ASAP7_75t_L g1313 ( 
.A(n_1099),
.B(n_1164),
.Y(n_1313)
);

BUFx3_ASAP7_75t_L g1314 ( 
.A(n_1204),
.Y(n_1314)
);

BUFx2_ASAP7_75t_L g1315 ( 
.A(n_1121),
.Y(n_1315)
);

INVx2_ASAP7_75t_L g1316 ( 
.A(n_1109),
.Y(n_1316)
);

OR2x6_ASAP7_75t_L g1317 ( 
.A(n_1099),
.B(n_1164),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1109),
.Y(n_1318)
);

OAI21x1_ASAP7_75t_SL g1319 ( 
.A1(n_1201),
.A2(n_1009),
.B(n_1087),
.Y(n_1319)
);

OR2x6_ASAP7_75t_L g1320 ( 
.A(n_1099),
.B(n_1164),
.Y(n_1320)
);

BUFx2_ASAP7_75t_R g1321 ( 
.A(n_1153),
.Y(n_1321)
);

INVx2_ASAP7_75t_L g1322 ( 
.A(n_1109),
.Y(n_1322)
);

AOI21x1_ASAP7_75t_L g1323 ( 
.A1(n_1097),
.A2(n_972),
.B(n_983),
.Y(n_1323)
);

OAI21x1_ASAP7_75t_L g1324 ( 
.A1(n_1150),
.A2(n_1175),
.B(n_1158),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1152),
.B(n_1157),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1109),
.Y(n_1326)
);

AOI22xp33_ASAP7_75t_L g1327 ( 
.A1(n_1210),
.A2(n_822),
.B1(n_884),
.B2(n_977),
.Y(n_1327)
);

O2A1O1Ixp33_ASAP7_75t_L g1328 ( 
.A1(n_1301),
.A2(n_1236),
.B(n_1215),
.C(n_1220),
.Y(n_1328)
);

OAI22xp5_ASAP7_75t_L g1329 ( 
.A1(n_1285),
.A2(n_1327),
.B1(n_1283),
.B2(n_1301),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1226),
.B(n_1237),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1246),
.B(n_1291),
.Y(n_1331)
);

O2A1O1Ixp5_ASAP7_75t_L g1332 ( 
.A1(n_1244),
.A2(n_1302),
.B(n_1289),
.C(n_1247),
.Y(n_1332)
);

AOI21xp5_ASAP7_75t_SL g1333 ( 
.A1(n_1289),
.A2(n_1302),
.B(n_1236),
.Y(n_1333)
);

OA21x2_ASAP7_75t_L g1334 ( 
.A1(n_1240),
.A2(n_1227),
.B(n_1231),
.Y(n_1334)
);

NOR2xp67_ASAP7_75t_L g1335 ( 
.A(n_1218),
.B(n_1297),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_1224),
.Y(n_1336)
);

OR2x2_ASAP7_75t_L g1337 ( 
.A(n_1265),
.B(n_1221),
.Y(n_1337)
);

AND2x2_ASAP7_75t_L g1338 ( 
.A(n_1290),
.B(n_1306),
.Y(n_1338)
);

OAI22xp5_ASAP7_75t_L g1339 ( 
.A1(n_1285),
.A2(n_1327),
.B1(n_1283),
.B2(n_1284),
.Y(n_1339)
);

OA21x2_ASAP7_75t_L g1340 ( 
.A1(n_1240),
.A2(n_1231),
.B(n_1223),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1309),
.Y(n_1341)
);

AND2x4_ASAP7_75t_L g1342 ( 
.A(n_1307),
.B(n_1313),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1316),
.Y(n_1343)
);

CKINVDCx16_ASAP7_75t_R g1344 ( 
.A(n_1304),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1316),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1254),
.B(n_1259),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1312),
.B(n_1325),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1305),
.B(n_1251),
.Y(n_1348)
);

AND2x4_ASAP7_75t_L g1349 ( 
.A(n_1307),
.B(n_1313),
.Y(n_1349)
);

HB1xp67_ASAP7_75t_L g1350 ( 
.A(n_1273),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1260),
.B(n_1256),
.Y(n_1351)
);

OR2x2_ASAP7_75t_L g1352 ( 
.A(n_1322),
.B(n_1326),
.Y(n_1352)
);

AOI221x1_ASAP7_75t_SL g1353 ( 
.A1(n_1234),
.A2(n_1288),
.B1(n_1269),
.B2(n_1299),
.C(n_1318),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1270),
.B(n_1233),
.Y(n_1354)
);

AOI21xp5_ASAP7_75t_SL g1355 ( 
.A1(n_1267),
.A2(n_1320),
.B(n_1307),
.Y(n_1355)
);

AOI221x1_ASAP7_75t_SL g1356 ( 
.A1(n_1287),
.A2(n_1308),
.B1(n_1298),
.B2(n_1293),
.C(n_1292),
.Y(n_1356)
);

HB1xp67_ASAP7_75t_L g1357 ( 
.A(n_1276),
.Y(n_1357)
);

OR2x2_ASAP7_75t_L g1358 ( 
.A(n_1249),
.B(n_1232),
.Y(n_1358)
);

OAI22xp5_ASAP7_75t_L g1359 ( 
.A1(n_1264),
.A2(n_1267),
.B1(n_1262),
.B2(n_1271),
.Y(n_1359)
);

OR2x2_ASAP7_75t_L g1360 ( 
.A(n_1242),
.B(n_1238),
.Y(n_1360)
);

OA21x2_ASAP7_75t_L g1361 ( 
.A1(n_1223),
.A2(n_1261),
.B(n_1243),
.Y(n_1361)
);

AND2x4_ASAP7_75t_L g1362 ( 
.A(n_1313),
.B(n_1320),
.Y(n_1362)
);

OR2x2_ASAP7_75t_L g1363 ( 
.A(n_1315),
.B(n_1252),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1250),
.B(n_1319),
.Y(n_1364)
);

AOI21xp5_ASAP7_75t_SL g1365 ( 
.A1(n_1317),
.A2(n_1320),
.B(n_1300),
.Y(n_1365)
);

AOI21xp5_ASAP7_75t_SL g1366 ( 
.A1(n_1317),
.A2(n_1300),
.B(n_1303),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1268),
.Y(n_1367)
);

OAI22xp5_ASAP7_75t_L g1368 ( 
.A1(n_1271),
.A2(n_1229),
.B1(n_1272),
.B2(n_1303),
.Y(n_1368)
);

NOR2xp33_ASAP7_75t_R g1369 ( 
.A(n_1224),
.B(n_1295),
.Y(n_1369)
);

BUFx6f_ASAP7_75t_L g1370 ( 
.A(n_1275),
.Y(n_1370)
);

OAI22xp5_ASAP7_75t_L g1371 ( 
.A1(n_1229),
.A2(n_1272),
.B1(n_1296),
.B2(n_1317),
.Y(n_1371)
);

OA21x2_ASAP7_75t_L g1372 ( 
.A1(n_1235),
.A2(n_1216),
.B(n_1217),
.Y(n_1372)
);

HB1xp67_ASAP7_75t_L g1373 ( 
.A(n_1282),
.Y(n_1373)
);

AOI21xp5_ASAP7_75t_L g1374 ( 
.A1(n_1311),
.A2(n_1294),
.B(n_1219),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1230),
.B(n_1314),
.Y(n_1375)
);

INVx1_ASAP7_75t_SL g1376 ( 
.A(n_1321),
.Y(n_1376)
);

AND2x4_ASAP7_75t_L g1377 ( 
.A(n_1263),
.B(n_1279),
.Y(n_1377)
);

O2A1O1Ixp5_ASAP7_75t_L g1378 ( 
.A1(n_1255),
.A2(n_1323),
.B(n_1286),
.C(n_1222),
.Y(n_1378)
);

INVx1_ASAP7_75t_SL g1379 ( 
.A(n_1225),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1281),
.B(n_1252),
.Y(n_1380)
);

OAI22xp5_ASAP7_75t_L g1381 ( 
.A1(n_1258),
.A2(n_1239),
.B1(n_1252),
.B2(n_1253),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1281),
.B(n_1280),
.Y(n_1382)
);

OAI22xp5_ASAP7_75t_L g1383 ( 
.A1(n_1253),
.A2(n_1225),
.B1(n_1295),
.B2(n_1282),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1228),
.B(n_1278),
.Y(n_1384)
);

AND2x4_ASAP7_75t_L g1385 ( 
.A(n_1257),
.B(n_1241),
.Y(n_1385)
);

INVx2_ASAP7_75t_SL g1386 ( 
.A(n_1277),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1248),
.B(n_1275),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1248),
.B(n_1266),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1248),
.B(n_1266),
.Y(n_1389)
);

OA22x2_ASAP7_75t_L g1390 ( 
.A1(n_1274),
.A2(n_1245),
.B1(n_1257),
.B2(n_1248),
.Y(n_1390)
);

OAI22xp5_ASAP7_75t_L g1391 ( 
.A1(n_1310),
.A2(n_1327),
.B1(n_1285),
.B2(n_1210),
.Y(n_1391)
);

AND2x2_ASAP7_75t_SL g1392 ( 
.A(n_1324),
.B(n_1219),
.Y(n_1392)
);

OAI22xp5_ASAP7_75t_L g1393 ( 
.A1(n_1285),
.A2(n_1327),
.B1(n_1210),
.B2(n_1283),
.Y(n_1393)
);

OR2x2_ASAP7_75t_L g1394 ( 
.A(n_1265),
.B(n_1221),
.Y(n_1394)
);

O2A1O1Ixp5_ASAP7_75t_L g1395 ( 
.A1(n_1220),
.A2(n_1162),
.B(n_1207),
.C(n_1198),
.Y(n_1395)
);

NOR2xp67_ASAP7_75t_L g1396 ( 
.A(n_1218),
.B(n_1077),
.Y(n_1396)
);

CKINVDCx5p33_ASAP7_75t_R g1397 ( 
.A(n_1224),
.Y(n_1397)
);

BUFx3_ASAP7_75t_L g1398 ( 
.A(n_1238),
.Y(n_1398)
);

AOI21xp5_ASAP7_75t_L g1399 ( 
.A1(n_1244),
.A2(n_972),
.B(n_1094),
.Y(n_1399)
);

NOR2xp67_ASAP7_75t_L g1400 ( 
.A(n_1218),
.B(n_1077),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1221),
.B(n_1290),
.Y(n_1401)
);

BUFx3_ASAP7_75t_L g1402 ( 
.A(n_1238),
.Y(n_1402)
);

OR2x2_ASAP7_75t_L g1403 ( 
.A(n_1265),
.B(n_1221),
.Y(n_1403)
);

BUFx3_ASAP7_75t_L g1404 ( 
.A(n_1238),
.Y(n_1404)
);

NOR2xp67_ASAP7_75t_L g1405 ( 
.A(n_1218),
.B(n_1077),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1357),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1357),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1388),
.B(n_1389),
.Y(n_1408)
);

HB1xp67_ASAP7_75t_L g1409 ( 
.A(n_1373),
.Y(n_1409)
);

BUFx2_ASAP7_75t_L g1410 ( 
.A(n_1373),
.Y(n_1410)
);

AOI22xp33_ASAP7_75t_L g1411 ( 
.A1(n_1339),
.A2(n_1393),
.B1(n_1329),
.B2(n_1391),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1380),
.B(n_1392),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1392),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1387),
.B(n_1374),
.Y(n_1414)
);

OR2x6_ASAP7_75t_L g1415 ( 
.A(n_1399),
.B(n_1355),
.Y(n_1415)
);

INVx3_ASAP7_75t_L g1416 ( 
.A(n_1385),
.Y(n_1416)
);

INVxp67_ASAP7_75t_R g1417 ( 
.A(n_1381),
.Y(n_1417)
);

INVx3_ASAP7_75t_L g1418 ( 
.A(n_1385),
.Y(n_1418)
);

OR2x6_ASAP7_75t_L g1419 ( 
.A(n_1365),
.B(n_1342),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1367),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1377),
.B(n_1385),
.Y(n_1421)
);

AOI22xp33_ASAP7_75t_SL g1422 ( 
.A1(n_1359),
.A2(n_1333),
.B1(n_1328),
.B2(n_1348),
.Y(n_1422)
);

CKINVDCx6p67_ASAP7_75t_R g1423 ( 
.A(n_1370),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1390),
.B(n_1386),
.Y(n_1424)
);

OR2x6_ASAP7_75t_L g1425 ( 
.A(n_1349),
.B(n_1362),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1390),
.B(n_1386),
.Y(n_1426)
);

AND2x4_ASAP7_75t_L g1427 ( 
.A(n_1349),
.B(n_1362),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1341),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1343),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1345),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1350),
.B(n_1363),
.Y(n_1431)
);

OR2x2_ASAP7_75t_L g1432 ( 
.A(n_1350),
.B(n_1354),
.Y(n_1432)
);

OR2x2_ASAP7_75t_L g1433 ( 
.A(n_1383),
.B(n_1334),
.Y(n_1433)
);

NOR2xp67_ASAP7_75t_L g1434 ( 
.A(n_1364),
.B(n_1371),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1332),
.B(n_1361),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1330),
.B(n_1331),
.Y(n_1436)
);

HB1xp67_ASAP7_75t_L g1437 ( 
.A(n_1352),
.Y(n_1437)
);

OR2x6_ASAP7_75t_L g1438 ( 
.A(n_1366),
.B(n_1340),
.Y(n_1438)
);

AO21x2_ASAP7_75t_L g1439 ( 
.A1(n_1384),
.A2(n_1351),
.B(n_1368),
.Y(n_1439)
);

OR2x2_ASAP7_75t_L g1440 ( 
.A(n_1334),
.B(n_1340),
.Y(n_1440)
);

OR2x2_ASAP7_75t_L g1441 ( 
.A(n_1334),
.B(n_1340),
.Y(n_1441)
);

HB1xp67_ASAP7_75t_L g1442 ( 
.A(n_1409),
.Y(n_1442)
);

BUFx6f_ASAP7_75t_L g1443 ( 
.A(n_1438),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1420),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1420),
.Y(n_1445)
);

HB1xp67_ASAP7_75t_L g1446 ( 
.A(n_1409),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1432),
.B(n_1394),
.Y(n_1447)
);

OR2x2_ASAP7_75t_L g1448 ( 
.A(n_1410),
.B(n_1372),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1432),
.B(n_1437),
.Y(n_1449)
);

OR2x2_ASAP7_75t_L g1450 ( 
.A(n_1410),
.B(n_1372),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1408),
.B(n_1332),
.Y(n_1451)
);

BUFx2_ASAP7_75t_L g1452 ( 
.A(n_1410),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_1423),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1412),
.B(n_1395),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1412),
.B(n_1395),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1412),
.B(n_1378),
.Y(n_1456)
);

INVx2_ASAP7_75t_R g1457 ( 
.A(n_1435),
.Y(n_1457)
);

AND2x4_ASAP7_75t_L g1458 ( 
.A(n_1416),
.B(n_1418),
.Y(n_1458)
);

AND2x4_ASAP7_75t_SL g1459 ( 
.A(n_1419),
.B(n_1370),
.Y(n_1459)
);

AOI22xp33_ASAP7_75t_L g1460 ( 
.A1(n_1411),
.A2(n_1347),
.B1(n_1337),
.B2(n_1403),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1421),
.B(n_1401),
.Y(n_1461)
);

OR2x2_ASAP7_75t_L g1462 ( 
.A(n_1432),
.B(n_1360),
.Y(n_1462)
);

OR2x2_ASAP7_75t_L g1463 ( 
.A(n_1431),
.B(n_1413),
.Y(n_1463)
);

AND2x4_ASAP7_75t_L g1464 ( 
.A(n_1418),
.B(n_1382),
.Y(n_1464)
);

NOR2xp33_ASAP7_75t_L g1465 ( 
.A(n_1422),
.B(n_1402),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1442),
.Y(n_1466)
);

INVx3_ASAP7_75t_L g1467 ( 
.A(n_1458),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1464),
.B(n_1414),
.Y(n_1468)
);

OAI21xp5_ASAP7_75t_L g1469 ( 
.A1(n_1465),
.A2(n_1422),
.B(n_1411),
.Y(n_1469)
);

BUFx3_ASAP7_75t_L g1470 ( 
.A(n_1459),
.Y(n_1470)
);

A2O1A1Ixp33_ASAP7_75t_L g1471 ( 
.A1(n_1465),
.A2(n_1353),
.B(n_1434),
.C(n_1335),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1442),
.Y(n_1472)
);

AOI221xp5_ASAP7_75t_L g1473 ( 
.A1(n_1460),
.A2(n_1436),
.B1(n_1356),
.B2(n_1424),
.C(n_1426),
.Y(n_1473)
);

NAND4xp25_ASAP7_75t_L g1474 ( 
.A(n_1460),
.B(n_1436),
.C(n_1434),
.D(n_1358),
.Y(n_1474)
);

BUFx4f_ASAP7_75t_SL g1475 ( 
.A(n_1462),
.Y(n_1475)
);

AND2x4_ASAP7_75t_L g1476 ( 
.A(n_1458),
.B(n_1418),
.Y(n_1476)
);

BUFx2_ASAP7_75t_L g1477 ( 
.A(n_1452),
.Y(n_1477)
);

NOR2xp33_ASAP7_75t_R g1478 ( 
.A(n_1453),
.B(n_1336),
.Y(n_1478)
);

OAI22xp5_ASAP7_75t_L g1479 ( 
.A1(n_1453),
.A2(n_1423),
.B1(n_1415),
.B2(n_1419),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1446),
.Y(n_1480)
);

AOI22xp33_ASAP7_75t_L g1481 ( 
.A1(n_1459),
.A2(n_1415),
.B1(n_1439),
.B2(n_1419),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_L g1482 ( 
.A1(n_1459),
.A2(n_1415),
.B1(n_1439),
.B2(n_1419),
.Y(n_1482)
);

AOI22xp33_ASAP7_75t_L g1483 ( 
.A1(n_1459),
.A2(n_1415),
.B1(n_1439),
.B2(n_1419),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1447),
.B(n_1439),
.Y(n_1484)
);

OAI22xp33_ASAP7_75t_L g1485 ( 
.A1(n_1447),
.A2(n_1415),
.B1(n_1417),
.B2(n_1419),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1446),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1464),
.B(n_1454),
.Y(n_1487)
);

OAI221xp5_ASAP7_75t_L g1488 ( 
.A1(n_1462),
.A2(n_1415),
.B1(n_1405),
.B2(n_1396),
.C(n_1400),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1454),
.B(n_1437),
.Y(n_1489)
);

OR2x2_ASAP7_75t_L g1490 ( 
.A(n_1463),
.B(n_1431),
.Y(n_1490)
);

AOI222xp33_ASAP7_75t_L g1491 ( 
.A1(n_1451),
.A2(n_1338),
.B1(n_1376),
.B2(n_1370),
.C1(n_1379),
.C2(n_1346),
.Y(n_1491)
);

OAI22xp33_ASAP7_75t_L g1492 ( 
.A1(n_1463),
.A2(n_1417),
.B1(n_1425),
.B2(n_1423),
.Y(n_1492)
);

INVx3_ASAP7_75t_L g1493 ( 
.A(n_1458),
.Y(n_1493)
);

OAI33xp33_ASAP7_75t_L g1494 ( 
.A1(n_1449),
.A2(n_1406),
.A3(n_1407),
.B1(n_1430),
.B2(n_1429),
.B3(n_1428),
.Y(n_1494)
);

AOI33xp33_ASAP7_75t_L g1495 ( 
.A1(n_1456),
.A2(n_1424),
.A3(n_1426),
.B1(n_1435),
.B2(n_1431),
.B3(n_1428),
.Y(n_1495)
);

BUFx2_ASAP7_75t_L g1496 ( 
.A(n_1452),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1464),
.B(n_1424),
.Y(n_1497)
);

OAI221xp5_ASAP7_75t_SL g1498 ( 
.A1(n_1456),
.A2(n_1433),
.B1(n_1426),
.B2(n_1435),
.C(n_1425),
.Y(n_1498)
);

INVx3_ASAP7_75t_L g1499 ( 
.A(n_1476),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1466),
.Y(n_1500)
);

INVx4_ASAP7_75t_L g1501 ( 
.A(n_1470),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1466),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1472),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1480),
.Y(n_1504)
);

INVx1_ASAP7_75t_SL g1505 ( 
.A(n_1475),
.Y(n_1505)
);

OAI21x1_ASAP7_75t_L g1506 ( 
.A1(n_1467),
.A2(n_1441),
.B(n_1440),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1487),
.B(n_1457),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1490),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1480),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1486),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_SL g1511 ( 
.A(n_1491),
.B(n_1427),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1490),
.Y(n_1512)
);

OR2x6_ASAP7_75t_L g1513 ( 
.A(n_1479),
.B(n_1443),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1477),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1477),
.Y(n_1515)
);

HB1xp67_ASAP7_75t_L g1516 ( 
.A(n_1496),
.Y(n_1516)
);

HB1xp67_ASAP7_75t_L g1517 ( 
.A(n_1496),
.Y(n_1517)
);

AND2x4_ASAP7_75t_L g1518 ( 
.A(n_1467),
.B(n_1443),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1489),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1487),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1484),
.B(n_1454),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1468),
.B(n_1457),
.Y(n_1522)
);

HB1xp67_ASAP7_75t_L g1523 ( 
.A(n_1497),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1500),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1501),
.B(n_1523),
.Y(n_1525)
);

NAND2x1p5_ASAP7_75t_L g1526 ( 
.A(n_1501),
.B(n_1470),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1500),
.Y(n_1527)
);

NOR2xp33_ASAP7_75t_L g1528 ( 
.A(n_1505),
.B(n_1336),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1501),
.B(n_1468),
.Y(n_1529)
);

AOI22xp33_ASAP7_75t_L g1530 ( 
.A1(n_1511),
.A2(n_1469),
.B1(n_1474),
.B2(n_1485),
.Y(n_1530)
);

BUFx2_ASAP7_75t_L g1531 ( 
.A(n_1501),
.Y(n_1531)
);

OR2x2_ASAP7_75t_L g1532 ( 
.A(n_1519),
.B(n_1455),
.Y(n_1532)
);

CKINVDCx20_ASAP7_75t_R g1533 ( 
.A(n_1505),
.Y(n_1533)
);

AOI31xp33_ASAP7_75t_L g1534 ( 
.A1(n_1511),
.A2(n_1471),
.A3(n_1491),
.B(n_1473),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1507),
.B(n_1457),
.Y(n_1535)
);

OAI31xp33_ASAP7_75t_L g1536 ( 
.A1(n_1516),
.A2(n_1474),
.A3(n_1488),
.B(n_1498),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1500),
.Y(n_1537)
);

OR2x2_ASAP7_75t_L g1538 ( 
.A(n_1519),
.B(n_1455),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1506),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1502),
.B(n_1495),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1504),
.Y(n_1541)
);

BUFx3_ASAP7_75t_L g1542 ( 
.A(n_1501),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1504),
.Y(n_1543)
);

INVx3_ASAP7_75t_L g1544 ( 
.A(n_1518),
.Y(n_1544)
);

OAI33xp33_ASAP7_75t_L g1545 ( 
.A1(n_1515),
.A2(n_1492),
.A3(n_1450),
.B1(n_1448),
.B2(n_1445),
.B3(n_1444),
.Y(n_1545)
);

AOI22x1_ASAP7_75t_L g1546 ( 
.A1(n_1516),
.A2(n_1344),
.B1(n_1370),
.B2(n_1397),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1507),
.B(n_1523),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1506),
.Y(n_1548)
);

OR2x2_ASAP7_75t_L g1549 ( 
.A(n_1508),
.B(n_1455),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1507),
.B(n_1493),
.Y(n_1550)
);

NOR2xp33_ASAP7_75t_R g1551 ( 
.A(n_1514),
.B(n_1397),
.Y(n_1551)
);

BUFx3_ASAP7_75t_L g1552 ( 
.A(n_1515),
.Y(n_1552)
);

NOR3xp33_ASAP7_75t_L g1553 ( 
.A(n_1521),
.B(n_1494),
.C(n_1398),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1504),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1522),
.B(n_1493),
.Y(n_1555)
);

INVx2_ASAP7_75t_L g1556 ( 
.A(n_1506),
.Y(n_1556)
);

CKINVDCx20_ASAP7_75t_R g1557 ( 
.A(n_1513),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1522),
.B(n_1520),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1522),
.B(n_1520),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1509),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1502),
.B(n_1451),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1547),
.Y(n_1562)
);

AO21x1_ASAP7_75t_L g1563 ( 
.A1(n_1534),
.A2(n_1515),
.B(n_1514),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1524),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1547),
.Y(n_1565)
);

OR2x2_ASAP7_75t_L g1566 ( 
.A(n_1540),
.B(n_1521),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1524),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1527),
.Y(n_1568)
);

OR2x2_ASAP7_75t_L g1569 ( 
.A(n_1540),
.B(n_1508),
.Y(n_1569)
);

OR2x2_ASAP7_75t_L g1570 ( 
.A(n_1561),
.B(n_1508),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1547),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1534),
.B(n_1461),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1527),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1530),
.B(n_1461),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1526),
.B(n_1529),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1526),
.B(n_1499),
.Y(n_1576)
);

OR2x6_ASAP7_75t_L g1577 ( 
.A(n_1531),
.B(n_1542),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1537),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1553),
.B(n_1461),
.Y(n_1579)
);

OAI21xp5_ASAP7_75t_SL g1580 ( 
.A1(n_1536),
.A2(n_1481),
.B(n_1482),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1537),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1552),
.Y(n_1582)
);

OR2x2_ASAP7_75t_L g1583 ( 
.A(n_1561),
.B(n_1512),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1541),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1541),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1543),
.Y(n_1586)
);

INVx1_ASAP7_75t_SL g1587 ( 
.A(n_1533),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1543),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1554),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1554),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1560),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1560),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1526),
.B(n_1499),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1552),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1553),
.B(n_1512),
.Y(n_1595)
);

OR2x2_ASAP7_75t_L g1596 ( 
.A(n_1532),
.B(n_1512),
.Y(n_1596)
);

AND2x4_ASAP7_75t_L g1597 ( 
.A(n_1577),
.B(n_1542),
.Y(n_1597)
);

OR2x2_ASAP7_75t_L g1598 ( 
.A(n_1562),
.B(n_1532),
.Y(n_1598)
);

OAI21xp5_ASAP7_75t_L g1599 ( 
.A1(n_1580),
.A2(n_1536),
.B(n_1546),
.Y(n_1599)
);

HB1xp67_ASAP7_75t_L g1600 ( 
.A(n_1577),
.Y(n_1600)
);

INVx3_ASAP7_75t_L g1601 ( 
.A(n_1577),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1564),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1567),
.Y(n_1603)
);

OR2x2_ASAP7_75t_L g1604 ( 
.A(n_1562),
.B(n_1538),
.Y(n_1604)
);

INVx1_ASAP7_75t_SL g1605 ( 
.A(n_1587),
.Y(n_1605)
);

INVx1_ASAP7_75t_SL g1606 ( 
.A(n_1575),
.Y(n_1606)
);

HB1xp67_ASAP7_75t_L g1607 ( 
.A(n_1577),
.Y(n_1607)
);

INVx1_ASAP7_75t_SL g1608 ( 
.A(n_1575),
.Y(n_1608)
);

OR2x2_ASAP7_75t_L g1609 ( 
.A(n_1565),
.B(n_1538),
.Y(n_1609)
);

AOI22xp33_ASAP7_75t_L g1610 ( 
.A1(n_1563),
.A2(n_1557),
.B1(n_1545),
.B2(n_1513),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1565),
.B(n_1526),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1568),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1572),
.B(n_1525),
.Y(n_1613)
);

OR2x2_ASAP7_75t_L g1614 ( 
.A(n_1571),
.B(n_1552),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1573),
.Y(n_1615)
);

NOR2xp33_ASAP7_75t_L g1616 ( 
.A(n_1574),
.B(n_1528),
.Y(n_1616)
);

NOR2x1_ASAP7_75t_L g1617 ( 
.A(n_1582),
.B(n_1542),
.Y(n_1617)
);

INVx3_ASAP7_75t_L g1618 ( 
.A(n_1571),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1578),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1582),
.Y(n_1620)
);

INVx1_ASAP7_75t_SL g1621 ( 
.A(n_1576),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1605),
.B(n_1563),
.Y(n_1622)
);

AOI21xp5_ASAP7_75t_L g1623 ( 
.A1(n_1599),
.A2(n_1595),
.B(n_1594),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1601),
.Y(n_1624)
);

AOI221xp5_ASAP7_75t_L g1625 ( 
.A1(n_1610),
.A2(n_1545),
.B1(n_1566),
.B2(n_1569),
.C(n_1579),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1603),
.Y(n_1626)
);

OAI21xp5_ASAP7_75t_L g1627 ( 
.A1(n_1617),
.A2(n_1616),
.B(n_1607),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1603),
.Y(n_1628)
);

OAI31xp33_ASAP7_75t_L g1629 ( 
.A1(n_1606),
.A2(n_1566),
.A3(n_1569),
.B(n_1531),
.Y(n_1629)
);

INVx2_ASAP7_75t_SL g1630 ( 
.A(n_1597),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1612),
.Y(n_1631)
);

AND2x4_ASAP7_75t_L g1632 ( 
.A(n_1601),
.B(n_1576),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1600),
.B(n_1608),
.Y(n_1633)
);

OAI22xp5_ASAP7_75t_L g1634 ( 
.A1(n_1613),
.A2(n_1546),
.B1(n_1483),
.B2(n_1513),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1612),
.Y(n_1635)
);

OAI21xp33_ASAP7_75t_SL g1636 ( 
.A1(n_1601),
.A2(n_1593),
.B(n_1525),
.Y(n_1636)
);

OAI32xp33_ASAP7_75t_L g1637 ( 
.A1(n_1621),
.A2(n_1593),
.A3(n_1544),
.B1(n_1596),
.B2(n_1517),
.Y(n_1637)
);

HB1xp67_ASAP7_75t_L g1638 ( 
.A(n_1618),
.Y(n_1638)
);

NOR3xp33_ASAP7_75t_L g1639 ( 
.A(n_1620),
.B(n_1584),
.C(n_1581),
.Y(n_1639)
);

OAI21xp33_ASAP7_75t_L g1640 ( 
.A1(n_1597),
.A2(n_1551),
.B(n_1570),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1630),
.B(n_1624),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1632),
.B(n_1597),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1638),
.Y(n_1643)
);

NOR2xp33_ASAP7_75t_L g1644 ( 
.A(n_1622),
.B(n_1633),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_SL g1645 ( 
.A(n_1627),
.B(n_1618),
.Y(n_1645)
);

INVx3_ASAP7_75t_L g1646 ( 
.A(n_1632),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1626),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1628),
.Y(n_1648)
);

AOI22xp33_ASAP7_75t_L g1649 ( 
.A1(n_1625),
.A2(n_1611),
.B1(n_1620),
.B2(n_1513),
.Y(n_1649)
);

OR2x2_ASAP7_75t_L g1650 ( 
.A(n_1629),
.B(n_1614),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1631),
.Y(n_1651)
);

INVxp67_ASAP7_75t_L g1652 ( 
.A(n_1627),
.Y(n_1652)
);

A2O1A1Ixp33_ASAP7_75t_L g1653 ( 
.A1(n_1652),
.A2(n_1623),
.B(n_1644),
.C(n_1649),
.Y(n_1653)
);

A2O1A1Ixp33_ASAP7_75t_L g1654 ( 
.A1(n_1644),
.A2(n_1640),
.B(n_1634),
.C(n_1637),
.Y(n_1654)
);

A2O1A1Ixp33_ASAP7_75t_L g1655 ( 
.A1(n_1645),
.A2(n_1634),
.B(n_1639),
.C(n_1636),
.Y(n_1655)
);

NAND4xp25_ASAP7_75t_L g1656 ( 
.A(n_1641),
.B(n_1635),
.C(n_1614),
.D(n_1602),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_SL g1657 ( 
.A(n_1646),
.B(n_1611),
.Y(n_1657)
);

OAI211xp5_ASAP7_75t_L g1658 ( 
.A1(n_1645),
.A2(n_1619),
.B(n_1615),
.C(n_1618),
.Y(n_1658)
);

OAI221xp5_ASAP7_75t_L g1659 ( 
.A1(n_1650),
.A2(n_1619),
.B1(n_1615),
.B2(n_1609),
.C(n_1604),
.Y(n_1659)
);

NOR4xp25_ASAP7_75t_L g1660 ( 
.A(n_1646),
.B(n_1609),
.C(n_1604),
.D(n_1598),
.Y(n_1660)
);

AOI311xp33_ASAP7_75t_L g1661 ( 
.A1(n_1647),
.A2(n_1648),
.A3(n_1590),
.B(n_1592),
.C(n_1586),
.Y(n_1661)
);

AOI21xp5_ASAP7_75t_L g1662 ( 
.A1(n_1646),
.A2(n_1598),
.B(n_1588),
.Y(n_1662)
);

AOI22xp33_ASAP7_75t_L g1663 ( 
.A1(n_1659),
.A2(n_1642),
.B1(n_1643),
.B2(n_1651),
.Y(n_1663)
);

AOI211xp5_ASAP7_75t_L g1664 ( 
.A1(n_1655),
.A2(n_1653),
.B(n_1660),
.C(n_1654),
.Y(n_1664)
);

INVx3_ASAP7_75t_L g1665 ( 
.A(n_1658),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1657),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1662),
.Y(n_1667)
);

BUFx2_ASAP7_75t_L g1668 ( 
.A(n_1666),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1667),
.Y(n_1669)
);

NOR2xp33_ASAP7_75t_L g1670 ( 
.A(n_1665),
.B(n_1656),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1663),
.B(n_1643),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1663),
.B(n_1661),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1665),
.Y(n_1673)
);

A2O1A1Ixp33_ASAP7_75t_L g1674 ( 
.A1(n_1670),
.A2(n_1664),
.B(n_1651),
.C(n_1585),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1668),
.B(n_1529),
.Y(n_1675)
);

AOI31xp33_ASAP7_75t_L g1676 ( 
.A1(n_1671),
.A2(n_1369),
.A3(n_1596),
.B(n_1589),
.Y(n_1676)
);

OAI322xp33_ASAP7_75t_L g1677 ( 
.A1(n_1670),
.A2(n_1591),
.A3(n_1583),
.B1(n_1570),
.B2(n_1548),
.C1(n_1539),
.C2(n_1556),
.Y(n_1677)
);

OAI211xp5_ASAP7_75t_SL g1678 ( 
.A1(n_1673),
.A2(n_1583),
.B(n_1544),
.C(n_1539),
.Y(n_1678)
);

AND4x1_ASAP7_75t_L g1679 ( 
.A(n_1674),
.B(n_1669),
.C(n_1672),
.D(n_1369),
.Y(n_1679)
);

NOR4xp75_ASAP7_75t_SL g1680 ( 
.A(n_1676),
.B(n_1478),
.C(n_1544),
.D(n_1558),
.Y(n_1680)
);

NOR2xp67_ASAP7_75t_SL g1681 ( 
.A(n_1675),
.B(n_1398),
.Y(n_1681)
);

NAND2x1p5_ASAP7_75t_L g1682 ( 
.A(n_1679),
.B(n_1402),
.Y(n_1682)
);

OAI322xp33_ASAP7_75t_L g1683 ( 
.A1(n_1682),
.A2(n_1680),
.A3(n_1681),
.B1(n_1678),
.B2(n_1677),
.C1(n_1539),
.C2(n_1548),
.Y(n_1683)
);

XOR2xp5_ASAP7_75t_L g1684 ( 
.A(n_1683),
.B(n_1404),
.Y(n_1684)
);

HB1xp67_ASAP7_75t_L g1685 ( 
.A(n_1683),
.Y(n_1685)
);

OAI21xp5_ASAP7_75t_L g1686 ( 
.A1(n_1684),
.A2(n_1544),
.B(n_1548),
.Y(n_1686)
);

OAI22xp5_ASAP7_75t_L g1687 ( 
.A1(n_1685),
.A2(n_1549),
.B1(n_1556),
.B2(n_1517),
.Y(n_1687)
);

OAI22xp5_ASAP7_75t_L g1688 ( 
.A1(n_1687),
.A2(n_1686),
.B1(n_1549),
.B2(n_1556),
.Y(n_1688)
);

AND2x4_ASAP7_75t_L g1689 ( 
.A(n_1686),
.B(n_1558),
.Y(n_1689)
);

AOI21xp5_ASAP7_75t_L g1690 ( 
.A1(n_1688),
.A2(n_1559),
.B(n_1558),
.Y(n_1690)
);

NAND4xp25_ASAP7_75t_SL g1691 ( 
.A(n_1690),
.B(n_1689),
.C(n_1559),
.D(n_1535),
.Y(n_1691)
);

AOI21xp5_ASAP7_75t_L g1692 ( 
.A1(n_1691),
.A2(n_1559),
.B(n_1535),
.Y(n_1692)
);

AO21x2_ASAP7_75t_L g1693 ( 
.A1(n_1692),
.A2(n_1550),
.B(n_1555),
.Y(n_1693)
);

AOI31xp33_ASAP7_75t_L g1694 ( 
.A1(n_1693),
.A2(n_1404),
.A3(n_1535),
.B(n_1375),
.Y(n_1694)
);

AOI211xp5_ASAP7_75t_L g1695 ( 
.A1(n_1694),
.A2(n_1509),
.B(n_1503),
.C(n_1510),
.Y(n_1695)
);


endmodule