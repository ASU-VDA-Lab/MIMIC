module real_jpeg_6844_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_215;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_373;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g81 ( 
.A(n_0),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_1),
.A2(n_124),
.B1(n_128),
.B2(n_129),
.Y(n_123)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_1),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_1),
.A2(n_169),
.B1(n_170),
.B2(n_171),
.Y(n_168)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_1),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_1),
.A2(n_177),
.B1(n_179),
.B2(n_180),
.Y(n_176)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_1),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_1),
.A2(n_171),
.B1(n_184),
.B2(n_263),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_2),
.A2(n_79),
.B1(n_82),
.B2(n_83),
.Y(n_78)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_2),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_2),
.A2(n_82),
.B1(n_183),
.B2(n_184),
.Y(n_182)
);

OAI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_2),
.A2(n_82),
.B1(n_201),
.B2(n_204),
.Y(n_200)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_3),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_3),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_3),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_4),
.Y(n_373)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_5),
.Y(n_138)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_6),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_6),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_6),
.Y(n_190)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_6),
.Y(n_232)
);

BUFx5_ASAP7_75t_L g265 ( 
.A(n_6),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_6),
.B(n_10),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_7),
.A2(n_55),
.B1(n_59),
.B2(n_60),
.Y(n_54)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_7),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_7),
.A2(n_59),
.B1(n_80),
.B2(n_120),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_10),
.A2(n_49),
.B1(n_50),
.B2(n_51),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_10),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_10),
.A2(n_50),
.B1(n_100),
.B2(n_104),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_10),
.A2(n_50),
.B1(n_156),
.B2(n_157),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_10),
.A2(n_50),
.B1(n_55),
.B2(n_235),
.Y(n_234)
);

O2A1O1Ixp33_ASAP7_75t_L g253 ( 
.A1(n_10),
.A2(n_254),
.B(n_255),
.C(n_259),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_10),
.B(n_88),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_10),
.B(n_289),
.C(n_290),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_10),
.B(n_166),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_10),
.B(n_149),
.C(n_311),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_10),
.B(n_25),
.Y(n_326)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_11),
.Y(n_170)
);

INVx3_ASAP7_75t_L g369 ( 
.A(n_12),
.Y(n_369)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_13),
.Y(n_92)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_13),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_13),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_367),
.B(n_370),
.Y(n_14)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_215),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_213),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_191),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_18),
.B(n_191),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_115),
.C(n_161),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_19),
.A2(n_20),
.B1(n_115),
.B2(n_116),
.Y(n_240)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_76),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_53),
.B2(n_75),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_23),
.A2(n_53),
.B(n_76),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_47),
.B(n_48),
.Y(n_23)
);

OA22x2_ASAP7_75t_L g167 ( 
.A1(n_24),
.A2(n_47),
.B1(n_48),
.B2(n_168),
.Y(n_167)
);

OA22x2_ASAP7_75t_L g195 ( 
.A1(n_24),
.A2(n_47),
.B1(n_48),
.B2(n_168),
.Y(n_195)
);

OR2x2_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_37),
.Y(n_24)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_28),
.B1(n_31),
.B2(n_34),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_27),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_27),
.Y(n_129)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_27),
.Y(n_152)
);

BUFx5_ASAP7_75t_L g159 ( 
.A(n_27),
.Y(n_159)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_27),
.Y(n_203)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_28),
.Y(n_254)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx4_ASAP7_75t_L g256 ( 
.A(n_30),
.Y(n_256)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_33),
.Y(n_148)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_38),
.A2(n_40),
.B1(n_42),
.B2(n_44),
.Y(n_37)
);

INVx2_ASAP7_75t_SL g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI21xp33_ASAP7_75t_L g255 ( 
.A1(n_50),
.A2(n_256),
.B(n_257),
.Y(n_255)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_51),
.Y(n_169)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_53),
.B(n_77),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_53),
.A2(n_75),
.B1(n_77),
.B2(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_64),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_54),
.Y(n_186)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_55),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_58),
.Y(n_95)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx8_ASAP7_75t_L g183 ( 
.A(n_62),
.Y(n_183)
);

BUFx8_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g264 ( 
.A(n_63),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g292 ( 
.A(n_63),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_64),
.B(n_234),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_65),
.B(n_73),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_65),
.A2(n_182),
.B1(n_186),
.B2(n_187),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_66),
.B(n_234),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_66),
.A2(n_234),
.B1(n_262),
.B2(n_265),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_66),
.A2(n_234),
.B1(n_262),
.B2(n_278),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_70),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_69),
.Y(n_185)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_72),
.Y(n_278)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_77),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_86),
.B(n_98),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_78),
.A2(n_86),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_81),
.Y(n_85)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_81),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g287 ( 
.A(n_81),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_83),
.A2(n_107),
.B1(n_111),
.B2(n_113),
.Y(n_106)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_85),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_85),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_85),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_85),
.Y(n_179)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_87),
.A2(n_99),
.B1(n_105),
.B2(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_87),
.B(n_105),
.Y(n_208)
);

OA22x2_ASAP7_75t_L g228 ( 
.A1(n_87),
.A2(n_99),
.B1(n_105),
.B2(n_176),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_87),
.A2(n_99),
.B(n_105),
.Y(n_338)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_106),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_90),
.B1(n_93),
.B2(n_96),
.Y(n_88)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_92),
.Y(n_97)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_105),
.Y(n_98)
);

INVx5_ASAP7_75t_SL g100 ( 
.A(n_101),
.Y(n_100)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_103),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_105),
.Y(n_118)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_108),
.Y(n_178)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_110),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_112),
.Y(n_114)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_121),
.B(n_160),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_117),
.B(n_121),
.Y(n_160)
);

AND2x2_ASAP7_75t_SL g207 ( 
.A(n_119),
.B(n_208),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_121),
.B(n_167),
.C(n_252),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_121),
.A2(n_323),
.B1(n_324),
.B2(n_327),
.Y(n_322)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_121),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_121),
.A2(n_167),
.B1(n_222),
.B2(n_327),
.Y(n_352)
);

OA22x2_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_130),
.B1(n_131),
.B2(n_154),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

AO22x2_ASAP7_75t_L g164 ( 
.A1(n_123),
.A2(n_155),
.B1(n_165),
.B2(n_166),
.Y(n_164)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_127),
.Y(n_204)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_127),
.Y(n_258)
);

INVx6_ASAP7_75t_SL g156 ( 
.A(n_129),
.Y(n_156)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_130),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_130),
.B(n_131),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_131),
.B(n_146),
.Y(n_130)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_131),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_131),
.A2(n_199),
.B(n_205),
.Y(n_198)
);

AOI22x1_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_134),
.B1(n_139),
.B2(n_142),
.Y(n_131)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_138),
.Y(n_145)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_138),
.Y(n_149)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_147),
.A2(n_149),
.B1(n_150),
.B2(n_153),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

BUFx12f_ASAP7_75t_L g309 ( 
.A(n_148),
.Y(n_309)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_149),
.Y(n_153)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_155),
.B(n_165),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_155),
.B(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_160),
.A2(n_193),
.B1(n_194),
.B2(n_211),
.Y(n_192)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_160),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_161),
.A2(n_162),
.B1(n_239),
.B2(n_240),
.Y(n_238)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_167),
.C(n_172),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_163),
.A2(n_164),
.B1(n_167),
.B2(n_222),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_163),
.A2(n_164),
.B1(n_227),
.B2(n_228),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_163),
.A2(n_164),
.B1(n_337),
.B2(n_338),
.Y(n_336)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_164),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_164),
.B(n_227),
.C(n_306),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_164),
.B(n_210),
.C(n_338),
.Y(n_356)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_167),
.Y(n_222)
);

INVx8_ASAP7_75t_L g259 ( 
.A(n_170),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_172),
.B(n_221),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_173),
.B(n_181),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_173),
.A2(n_181),
.B1(n_249),
.B2(n_250),
.Y(n_248)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_173),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_173),
.A2(n_250),
.B1(n_319),
.B2(n_320),
.Y(n_318)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_174),
.A2(n_175),
.B1(n_299),
.B2(n_300),
.Y(n_298)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_181),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_182),
.A2(n_230),
.B(n_233),
.Y(n_229)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_212),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_196),
.B1(n_197),
.B2(n_210),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_195),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_195),
.B(n_226),
.C(n_236),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_195),
.A2(n_210),
.B1(n_236),
.B2(n_247),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_195),
.A2(n_210),
.B1(n_335),
.B2(n_336),
.Y(n_334)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_198),
.A2(n_206),
.B1(n_207),
.B2(n_209),
.Y(n_197)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_198),
.Y(n_209)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx6_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_207),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

OAI211xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_266),
.B(n_362),
.C(n_366),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_241),
.Y(n_217)
);

A2O1A1Ixp33_ASAP7_75t_L g362 ( 
.A1(n_218),
.A2(n_241),
.B(n_363),
.C(n_365),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_238),
.Y(n_218)
);

OR2x2_ASAP7_75t_L g366 ( 
.A(n_219),
.B(n_238),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_223),
.C(n_225),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_220),
.B(n_223),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_225),
.B(n_243),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_226),
.B(n_246),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_227),
.B(n_229),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_227),
.A2(n_228),
.B1(n_285),
.B2(n_293),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_227),
.B(n_293),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_227),
.A2(n_228),
.B1(n_229),
.B2(n_354),
.Y(n_353)
);

INVx2_ASAP7_75t_SL g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_229),
.Y(n_354)
);

INVx5_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_236),
.Y(n_247)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_242),
.B(n_244),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_242),
.B(n_244),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_248),
.C(n_251),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_245),
.B(n_248),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_250),
.B(n_261),
.C(n_299),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_250),
.B(n_319),
.C(n_321),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_251),
.B(n_348),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_252),
.B(n_352),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_260),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_253),
.A2(n_260),
.B1(n_261),
.B2(n_344),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_253),
.Y(n_344)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_260),
.A2(n_261),
.B1(n_297),
.B2(n_298),
.Y(n_296)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_261),
.B(n_280),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_261),
.B(n_280),
.Y(n_281)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

BUFx2_ASAP7_75t_L g275 ( 
.A(n_264),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_267),
.B(n_346),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_268),
.A2(n_331),
.B(n_345),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_316),
.B(n_330),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_270),
.A2(n_303),
.B(n_315),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_295),
.B(n_302),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_282),
.B(n_294),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_279),
.B(n_281),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_277),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_277),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_277),
.A2(n_283),
.B1(n_325),
.B2(n_326),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_283),
.B(n_284),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_283),
.B(n_325),
.C(n_327),
.Y(n_341)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_285),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_288),
.Y(n_285)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_287),
.Y(n_311)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx5_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_296),
.B(n_301),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_296),
.B(n_301),
.Y(n_302)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_299),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_304),
.B(n_305),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_314),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_307),
.A2(n_308),
.B1(n_312),
.B2(n_313),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_307),
.B(n_313),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_308),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_312),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_317),
.B(n_329),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_317),
.B(n_329),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_318),
.A2(n_321),
.B1(n_322),
.B2(n_328),
.Y(n_317)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_318),
.Y(n_328)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_319),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

CKINVDCx14_ASAP7_75t_R g325 ( 
.A(n_326),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_333),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_332),
.B(n_333),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_339),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_334),
.B(n_341),
.C(n_342),
.Y(n_358)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_340),
.A2(n_341),
.B1(n_342),
.B2(n_343),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_SL g346 ( 
.A1(n_347),
.A2(n_349),
.B(n_357),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_347),
.B(n_349),
.C(n_364),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_353),
.C(n_355),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_351),
.B(n_360),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_353),
.A2(n_355),
.B1(n_356),
.B2(n_361),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_353),
.Y(n_361)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_359),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_358),
.B(n_359),
.Y(n_364)
);

BUFx4f_ASAP7_75t_SL g367 ( 
.A(n_368),
.Y(n_367)
);

INVx13_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx5_ASAP7_75t_L g372 ( 
.A(n_369),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_373),
.Y(n_370)
);

BUFx12f_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);


endmodule