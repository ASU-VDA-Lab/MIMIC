module fake_jpeg_31472_n_46 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_46);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_46;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_2),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_4),
.Y(n_8)
);

INVx3_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_SL g10 ( 
.A(n_5),
.B(n_3),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

BUFx3_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

AOI22xp5_ASAP7_75t_SL g14 ( 
.A1(n_7),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_14)
);

OR2x2_ASAP7_75t_L g25 ( 
.A(n_14),
.B(n_16),
.Y(n_25)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_10),
.B(n_0),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_10),
.B(n_5),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_17),
.B(n_6),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_13),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_18),
.A2(n_19),
.B1(n_7),
.B2(n_8),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g19 ( 
.A1(n_9),
.A2(n_1),
.B1(n_6),
.B2(n_12),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_20),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_23),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_24),
.B(n_18),
.C(n_14),
.Y(n_28)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

INVxp67_ASAP7_75t_SL g33 ( 
.A(n_27),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_28),
.A2(n_25),
.B1(n_24),
.B2(n_16),
.Y(n_34)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_29),
.A2(n_31),
.B1(n_23),
.B2(n_27),
.Y(n_32)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

OAI322xp33_ASAP7_75t_L g36 ( 
.A1(n_32),
.A2(n_30),
.A3(n_8),
.B1(n_7),
.B2(n_25),
.C1(n_34),
.C2(n_33),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_35),
.C(n_32),
.Y(n_38)
);

XOR2xp5_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_25),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_38),
.Y(n_40)
);

XNOR2x2_ASAP7_75t_SL g37 ( 
.A(n_35),
.B(n_22),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_37),
.B(n_8),
.Y(n_39)
);

AOI322xp5_ASAP7_75t_L g42 ( 
.A1(n_39),
.A2(n_11),
.A3(n_9),
.B1(n_13),
.B2(n_20),
.C1(n_21),
.C2(n_12),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_38),
.B(n_11),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_41),
.B(n_9),
.Y(n_43)
);

OAI21x1_ASAP7_75t_L g44 ( 
.A1(n_42),
.A2(n_43),
.B(n_40),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_44),
.B(n_12),
.C(n_13),
.Y(n_45)
);

NAND2x1_ASAP7_75t_L g46 ( 
.A(n_45),
.B(n_20),
.Y(n_46)
);


endmodule