module fake_jpeg_13655_n_349 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_349);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_349;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx8_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_16),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_6),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_10),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_5),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_21),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_44),
.B(n_21),
.Y(n_74)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_46),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_18),
.B(n_9),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_47),
.B(n_72),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_49),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_17),
.Y(n_50)
);

AOI21xp33_ASAP7_75t_L g91 ( 
.A1(n_50),
.A2(n_51),
.B(n_57),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_18),
.B(n_16),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_52),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_53),
.Y(n_94)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_55),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_26),
.A2(n_9),
.B1(n_1),
.B2(n_2),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_56),
.A2(n_43),
.B1(n_38),
.B2(n_35),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_19),
.B(n_11),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_59),
.Y(n_112)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_61),
.Y(n_111)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_62),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_64),
.Y(n_107)
);

HAxp5_ASAP7_75t_SL g65 ( 
.A(n_42),
.B(n_0),
.CON(n_65),
.SN(n_65)
);

CKINVDCx5p33_ASAP7_75t_R g95 ( 
.A(n_65),
.Y(n_95)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_37),
.Y(n_66)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_66),
.Y(n_118)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_17),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_67),
.Y(n_88)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_68),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_19),
.B(n_16),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_3),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_25),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_70),
.Y(n_110)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_71),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_22),
.B(n_10),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_42),
.B(n_0),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_73),
.B(n_33),
.C(n_40),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_74),
.B(n_83),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_50),
.A2(n_24),
.B1(n_36),
.B2(n_33),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_75),
.A2(n_84),
.B1(n_86),
.B2(n_6),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_77),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_78),
.B(n_117),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_81),
.B(n_98),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_50),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_73),
.A2(n_24),
.B1(n_36),
.B2(n_45),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_73),
.A2(n_24),
.B1(n_36),
.B2(n_38),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_SL g87 ( 
.A(n_53),
.Y(n_87)
);

INVx2_ASAP7_75t_SL g123 ( 
.A(n_87),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_89),
.A2(n_29),
.B1(n_55),
.B2(n_52),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_53),
.A2(n_27),
.B1(n_41),
.B2(n_40),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_90),
.A2(n_96),
.B1(n_99),
.B2(n_3),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_65),
.A2(n_41),
.B1(n_39),
.B2(n_34),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_54),
.Y(n_97)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_97),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_60),
.B(n_22),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_46),
.A2(n_20),
.B1(n_39),
.B2(n_34),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_61),
.A2(n_43),
.B1(n_35),
.B2(n_31),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_100),
.A2(n_103),
.B1(n_15),
.B2(n_88),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_62),
.A2(n_29),
.B1(n_27),
.B2(n_20),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_64),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_104),
.B(n_105),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_70),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_68),
.B(n_31),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_108),
.B(n_114),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_71),
.B(n_30),
.Y(n_114)
);

INVx6_ASAP7_75t_SL g116 ( 
.A(n_66),
.Y(n_116)
);

INVx6_ASAP7_75t_SL g127 ( 
.A(n_116),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_48),
.B(n_30),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_63),
.B(n_28),
.Y(n_119)
);

NAND3xp33_ASAP7_75t_SL g140 ( 
.A(n_119),
.B(n_121),
.C(n_8),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_49),
.B(n_28),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_116),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_124),
.B(n_144),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_125),
.A2(n_136),
.B1(n_132),
.B2(n_123),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_95),
.A2(n_59),
.B1(n_17),
.B2(n_7),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_126),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_128),
.Y(n_196)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_85),
.Y(n_129)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_129),
.Y(n_199)
);

OR2x2_ASAP7_75t_L g170 ( 
.A(n_132),
.B(n_140),
.Y(n_170)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_106),
.Y(n_133)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_133),
.Y(n_166)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_80),
.Y(n_135)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_135),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_89),
.A2(n_8),
.B1(n_12),
.B2(n_13),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_113),
.Y(n_137)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_137),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g138 ( 
.A(n_118),
.Y(n_138)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_138),
.Y(n_188)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_85),
.Y(n_139)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_139),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_118),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_141),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_95),
.A2(n_8),
.B1(n_12),
.B2(n_13),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_143),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_103),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_78),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_145),
.A2(n_147),
.B1(n_143),
.B2(n_126),
.Y(n_197)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_111),
.Y(n_146)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_146),
.Y(n_171)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_113),
.Y(n_148)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_148),
.Y(n_172)
);

NAND2x1_ASAP7_75t_SL g149 ( 
.A(n_110),
.B(n_111),
.Y(n_149)
);

AND2x2_ASAP7_75t_SL g183 ( 
.A(n_149),
.B(n_76),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_88),
.A2(n_110),
.B1(n_101),
.B2(n_77),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_150),
.A2(n_160),
.B1(n_97),
.B2(n_123),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_93),
.A2(n_115),
.B1(n_92),
.B2(n_120),
.Y(n_151)
);

OAI22xp33_ASAP7_75t_L g180 ( 
.A1(n_151),
.A2(n_156),
.B1(n_94),
.B2(n_76),
.Y(n_180)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_93),
.Y(n_153)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_153),
.Y(n_179)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_102),
.B(n_81),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_154),
.B(n_159),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_79),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_155),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_115),
.A2(n_92),
.B1(n_120),
.B2(n_79),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_80),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_157),
.B(n_107),
.Y(n_165)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_107),
.Y(n_158)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_158),
.Y(n_184)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_109),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_101),
.A2(n_94),
.B1(n_97),
.B2(n_76),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_109),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_161),
.B(n_149),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_165),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_122),
.B(n_91),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_167),
.B(n_177),
.Y(n_216)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_168),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_142),
.B(n_112),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_173),
.B(n_175),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_142),
.B(n_162),
.C(n_131),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_174),
.B(n_189),
.C(n_198),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_142),
.B(n_112),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_134),
.B(n_82),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g220 ( 
.A1(n_180),
.A2(n_176),
.B1(n_183),
.B2(n_187),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_144),
.B(n_82),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_181),
.B(n_182),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_136),
.B(n_82),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_183),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_185),
.A2(n_199),
.B(n_186),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_137),
.B(n_148),
.C(n_154),
.Y(n_189)
);

OAI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_190),
.A2(n_170),
.B1(n_196),
.B2(n_198),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_147),
.A2(n_133),
.B1(n_124),
.B2(n_153),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_192),
.A2(n_123),
.B1(n_157),
.B2(n_161),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_127),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_193),
.B(n_127),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_149),
.B(n_129),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_194),
.B(n_135),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_197),
.A2(n_152),
.B1(n_155),
.B2(n_196),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_145),
.B(n_146),
.C(n_139),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_201),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_178),
.B(n_174),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_202),
.B(n_209),
.Y(n_258)
);

BUFx12f_ASAP7_75t_L g203 ( 
.A(n_193),
.Y(n_203)
);

INVx13_ASAP7_75t_L g236 ( 
.A(n_203),
.Y(n_236)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_204),
.Y(n_239)
);

OR2x2_ASAP7_75t_L g205 ( 
.A(n_168),
.B(n_152),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_205),
.B(n_215),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_190),
.A2(n_155),
.B1(n_159),
.B2(n_158),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_208),
.B(n_218),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_189),
.B(n_130),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_211),
.B(n_222),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_212),
.A2(n_223),
.B(n_230),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_164),
.A2(n_182),
.B1(n_181),
.B2(n_195),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_214),
.A2(n_220),
.B1(n_225),
.B2(n_213),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_163),
.B(n_188),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_166),
.B(n_167),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_217),
.B(n_224),
.Y(n_240)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_166),
.Y(n_219)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_219),
.Y(n_242)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_186),
.Y(n_221)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_221),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_173),
.B(n_175),
.C(n_183),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_222),
.B(n_200),
.C(n_211),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_194),
.A2(n_170),
.B(n_169),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_184),
.B(n_169),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_180),
.A2(n_172),
.B1(n_176),
.B2(n_184),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_172),
.B(n_191),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_226),
.B(n_227),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_179),
.B(n_171),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_179),
.B(n_171),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_228),
.B(n_207),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_199),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_229),
.Y(n_234)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_186),
.Y(n_232)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_232),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_235),
.A2(n_208),
.B1(n_223),
.B2(n_206),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_215),
.B(n_217),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_237),
.B(n_216),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_238),
.B(n_254),
.C(n_209),
.Y(n_265)
);

INVx13_ASAP7_75t_L g243 ( 
.A(n_203),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_243),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_201),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_244),
.B(n_250),
.Y(n_271)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_219),
.Y(n_247)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_247),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_249),
.B(n_255),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_227),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_251),
.B(n_240),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_SL g254 ( 
.A(n_216),
.B(n_200),
.C(n_202),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_231),
.B(n_210),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_224),
.Y(n_256)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_256),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_231),
.B(n_210),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_257),
.B(n_250),
.Y(n_267)
);

INVx13_ASAP7_75t_L g259 ( 
.A(n_203),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_259),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_261),
.A2(n_262),
.B1(n_273),
.B2(n_274),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_246),
.A2(n_204),
.B1(n_206),
.B2(n_212),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_264),
.B(n_266),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_265),
.B(n_268),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_234),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_267),
.B(n_280),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_238),
.B(n_205),
.C(n_214),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_241),
.A2(n_205),
.B(n_230),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_270),
.B(n_278),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_246),
.A2(n_229),
.B1(n_232),
.B2(n_221),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_239),
.A2(n_203),
.B1(n_226),
.B2(n_228),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_239),
.A2(n_237),
.B1(n_255),
.B2(n_257),
.Y(n_275)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_275),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_235),
.A2(n_244),
.B1(n_256),
.B2(n_248),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_276),
.A2(n_252),
.B1(n_249),
.B2(n_247),
.Y(n_285)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_242),
.Y(n_279)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_279),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_233),
.A2(n_241),
.B(n_240),
.Y(n_280)
);

AO22x1_ASAP7_75t_L g281 ( 
.A1(n_234),
.A2(n_233),
.B1(n_248),
.B2(n_242),
.Y(n_281)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_281),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_285),
.A2(n_279),
.B1(n_269),
.B2(n_262),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_271),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_286),
.B(n_298),
.Y(n_300)
);

OAI21xp33_ASAP7_75t_L g290 ( 
.A1(n_267),
.A2(n_252),
.B(n_254),
.Y(n_290)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_290),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_280),
.A2(n_251),
.B1(n_258),
.B2(n_245),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_291),
.A2(n_294),
.B1(n_268),
.B2(n_281),
.Y(n_303)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_277),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_292),
.B(n_293),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_260),
.B(n_245),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_277),
.A2(n_258),
.B1(n_253),
.B2(n_243),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_263),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_296),
.B(n_272),
.Y(n_306)
);

INVxp33_ASAP7_75t_SL g298 ( 
.A(n_276),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_291),
.B(n_278),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_301),
.B(n_310),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_295),
.B(n_260),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_302),
.B(n_307),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_303),
.B(n_304),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_297),
.B(n_265),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_282),
.B(n_261),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_305),
.B(n_285),
.Y(n_320)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_306),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_283),
.B(n_274),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_283),
.B(n_269),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_309),
.B(n_311),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_282),
.B(n_281),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_284),
.B(n_270),
.C(n_273),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_312),
.B(n_284),
.C(n_288),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_315),
.B(n_319),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_299),
.B(n_292),
.Y(n_316)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_316),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_300),
.B(n_294),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_320),
.B(n_317),
.C(n_318),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_308),
.B(n_296),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_322),
.B(n_289),
.Y(n_328)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_312),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g330 ( 
.A(n_323),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_321),
.B(n_303),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_324),
.B(n_325),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_315),
.B(n_310),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_327),
.B(n_331),
.Y(n_338)
);

OR2x2_ASAP7_75t_L g333 ( 
.A(n_328),
.B(n_329),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_314),
.A2(n_289),
.B1(n_316),
.B2(n_293),
.Y(n_329)
);

OAI21x1_ASAP7_75t_L g331 ( 
.A1(n_317),
.A2(n_305),
.B(n_301),
.Y(n_331)
);

INVx11_ASAP7_75t_L g335 ( 
.A(n_330),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_335),
.B(n_336),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_325),
.B(n_318),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_326),
.B(n_320),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_337),
.B(n_332),
.C(n_304),
.Y(n_341)
);

AOI221xp5_ASAP7_75t_L g339 ( 
.A1(n_335),
.A2(n_332),
.B1(n_329),
.B2(n_313),
.C(n_287),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_339),
.A2(n_342),
.B(n_333),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_341),
.B(n_334),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_337),
.A2(n_236),
.B(n_243),
.Y(n_342)
);

AOI21x1_ASAP7_75t_L g345 ( 
.A1(n_343),
.A2(n_344),
.B(n_340),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_345),
.A2(n_338),
.B(n_333),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_346),
.B(n_287),
.C(n_259),
.Y(n_347)
);

O2A1O1Ixp33_ASAP7_75t_SL g348 ( 
.A1(n_347),
.A2(n_236),
.B(n_259),
.C(n_253),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_348),
.B(n_236),
.Y(n_349)
);


endmodule