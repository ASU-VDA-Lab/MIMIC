module real_jpeg_4265_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_393;
wire n_221;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_120;
wire n_155;
wire n_405;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_546;
wire n_285;
wire n_531;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_534;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_545;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp33_ASAP7_75t_L g274 ( 
.A1(n_0),
.A2(n_275),
.B1(n_278),
.B2(n_279),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_0),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g372 ( 
.A1(n_0),
.A2(n_278),
.B1(n_373),
.B2(n_375),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_0),
.A2(n_76),
.B1(n_278),
.B2(n_407),
.Y(n_406)
);

OAI22xp33_ASAP7_75t_L g468 ( 
.A1(n_0),
.A2(n_278),
.B1(n_343),
.B2(n_469),
.Y(n_468)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_1),
.A2(n_89),
.B1(n_93),
.B2(n_96),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_1),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_1),
.A2(n_96),
.B1(n_144),
.B2(n_145),
.Y(n_143)
);

OAI22xp33_ASAP7_75t_SL g384 ( 
.A1(n_1),
.A2(n_96),
.B1(n_184),
.B2(n_385),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_1),
.A2(n_96),
.B1(n_421),
.B2(n_423),
.Y(n_420)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_2),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_2),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_2),
.Y(n_236)
);

INVx8_ASAP7_75t_L g246 ( 
.A(n_2),
.Y(n_246)
);

BUFx5_ASAP7_75t_L g280 ( 
.A(n_2),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_2),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_2),
.Y(n_428)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_3),
.A2(n_99),
.B1(n_102),
.B2(n_106),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_3),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_3),
.A2(n_106),
.B1(n_135),
.B2(n_138),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_3),
.A2(n_106),
.B1(n_146),
.B2(n_153),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_3),
.A2(n_106),
.B1(n_314),
.B2(n_353),
.Y(n_391)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_4),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_4),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_4),
.Y(n_153)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_4),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_4),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_4),
.Y(n_442)
);

INVx6_ASAP7_75t_L g471 ( 
.A(n_4),
.Y(n_471)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_5),
.A2(n_165),
.B1(n_166),
.B2(n_167),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_5),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_5),
.B(n_131),
.C(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_5),
.B(n_77),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_5),
.B(n_200),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_5),
.B(n_133),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_5),
.B(n_101),
.Y(n_266)
);

OAI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_6),
.A2(n_184),
.B1(n_185),
.B2(n_186),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_6),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_6),
.A2(n_185),
.B1(n_258),
.B2(n_260),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_L g368 ( 
.A1(n_6),
.A2(n_185),
.B1(n_304),
.B2(n_369),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_6),
.A2(n_185),
.B1(n_343),
.B2(n_416),
.Y(n_415)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g335 ( 
.A(n_7),
.Y(n_335)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_9),
.A2(n_170),
.B1(n_172),
.B2(n_173),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_9),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_9),
.A2(n_172),
.B1(n_202),
.B2(n_205),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_9),
.A2(n_172),
.B1(n_269),
.B2(n_270),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_9),
.A2(n_153),
.B1(n_172),
.B2(n_364),
.Y(n_363)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_10),
.Y(n_117)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_10),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_10),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_10),
.Y(n_131)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_11),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_12),
.Y(n_126)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_12),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_12),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_13),
.A2(n_58),
.B1(n_60),
.B2(n_61),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_13),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g351 ( 
.A1(n_13),
.A2(n_61),
.B1(n_313),
.B2(n_352),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_13),
.A2(n_61),
.B1(n_398),
.B2(n_400),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_13),
.A2(n_61),
.B1(n_454),
.B2(n_456),
.Y(n_453)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_14),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_15),
.A2(n_20),
.B1(n_23),
.B2(n_24),
.Y(n_19)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_16),
.A2(n_36),
.B1(n_52),
.B2(n_54),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_16),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g312 ( 
.A1(n_16),
.A2(n_54),
.B1(n_313),
.B2(n_315),
.Y(n_312)
);

OAI22xp33_ASAP7_75t_SL g393 ( 
.A1(n_16),
.A2(n_54),
.B1(n_210),
.B2(n_394),
.Y(n_393)
);

AOI22xp33_ASAP7_75t_SL g411 ( 
.A1(n_16),
.A2(n_54),
.B1(n_269),
.B2(n_412),
.Y(n_411)
);

AOI22xp33_ASAP7_75t_L g209 ( 
.A1(n_17),
.A2(n_210),
.B1(n_211),
.B2(n_212),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_17),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_17),
.A2(n_211),
.B1(n_229),
.B2(n_232),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g300 ( 
.A1(n_17),
.A2(n_211),
.B1(n_301),
.B2(n_304),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_17),
.A2(n_52),
.B1(n_211),
.B2(n_441),
.Y(n_440)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_22),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_546),
.B(n_549),
.Y(n_24)
);

AO21x1_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_154),
.B(n_545),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_151),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_27),
.B(n_151),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_142),
.C(n_148),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g540 ( 
.A1(n_28),
.A2(n_29),
.B1(n_541),
.B2(n_542),
.Y(n_540)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_62),
.C(n_107),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_SL g532 ( 
.A(n_30),
.B(n_533),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_31),
.A2(n_51),
.B1(n_55),
.B2(n_57),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_31),
.A2(n_55),
.B1(n_57),
.B2(n_143),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_31),
.A2(n_55),
.B1(n_143),
.B2(n_152),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g414 ( 
.A1(n_31),
.A2(n_362),
.B(n_415),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_L g439 ( 
.A1(n_31),
.A2(n_55),
.B1(n_415),
.B2(n_440),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g517 ( 
.A1(n_31),
.A2(n_51),
.B1(n_55),
.B2(n_518),
.Y(n_517)
);

INVx2_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

AOI21xp5_ASAP7_75t_L g359 ( 
.A1(n_32),
.A2(n_360),
.B(n_361),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_32),
.B(n_363),
.Y(n_472)
);

OAI21xp5_ASAP7_75t_L g547 ( 
.A1(n_32),
.A2(n_56),
.B(n_548),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_42),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_36),
.B1(n_38),
.B2(n_39),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_38),
.Y(n_144)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_40),
.A2(n_43),
.B1(n_46),
.B2(n_49),
.Y(n_42)
);

INVx6_ASAP7_75t_L g337 ( 
.A(n_40),
.Y(n_337)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_45),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_45),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_45),
.Y(n_105)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx4_ASAP7_75t_L g269 ( 
.A(n_48),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_48),
.Y(n_270)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OAI21xp33_ASAP7_75t_SL g360 ( 
.A1(n_52),
.A2(n_167),
.B(n_340),
.Y(n_360)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_55),
.B(n_167),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g482 ( 
.A1(n_55),
.A2(n_440),
.B(n_472),
.Y(n_482)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_56),
.B(n_363),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_56),
.B(n_468),
.Y(n_467)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_58),
.Y(n_60)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_62),
.A2(n_107),
.B1(n_108),
.B2(n_534),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_62),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_88),
.B1(n_97),
.B2(n_98),
.Y(n_62)
);

INVx3_ASAP7_75t_SL g149 ( 
.A(n_63),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_63),
.A2(n_97),
.B1(n_300),
.B2(n_368),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_63),
.A2(n_97),
.B1(n_406),
.B2(n_411),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g521 ( 
.A1(n_63),
.A2(n_88),
.B1(n_97),
.B2(n_522),
.Y(n_521)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_77),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_69),
.B1(n_73),
.B2(n_75),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_71),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_72),
.Y(n_95)
);

BUFx5_ASAP7_75t_L g282 ( 
.A(n_72),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_72),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_72),
.Y(n_410)
);

NAND2xp33_ASAP7_75t_SL g289 ( 
.A(n_73),
.B(n_137),
.Y(n_289)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_77),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_77),
.A2(n_149),
.B(n_150),
.Y(n_148)
);

AOI22x1_ASAP7_75t_L g443 ( 
.A1(n_77),
.A2(n_149),
.B1(n_308),
.B2(n_444),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_77),
.A2(n_149),
.B1(n_452),
.B2(n_453),
.Y(n_451)
);

AO22x2_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_79),
.B1(n_82),
.B2(n_85),
.Y(n_77)
);

INVx4_ASAP7_75t_SL g212 ( 
.A(n_79),
.Y(n_212)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_81),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_81),
.Y(n_114)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_81),
.Y(n_137)
);

INVx11_ASAP7_75t_L g141 ( 
.A(n_81),
.Y(n_141)
);

BUFx5_ASAP7_75t_L g177 ( 
.A(n_81),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_81),
.Y(n_399)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_83),
.Y(n_120)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_83),
.Y(n_374)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx4_ASAP7_75t_L g288 ( 
.A(n_87),
.Y(n_288)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx5_ASAP7_75t_L g306 ( 
.A(n_92),
.Y(n_306)
);

BUFx3_ASAP7_75t_L g413 ( 
.A(n_92),
.Y(n_413)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_97),
.B(n_268),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_97),
.A2(n_300),
.B(n_307),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_98),
.Y(n_150)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_100),
.Y(n_99)
);

INVx6_ASAP7_75t_SL g100 ( 
.A(n_101),
.Y(n_100)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_105),
.Y(n_264)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_105),
.Y(n_329)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_105),
.Y(n_339)
);

INVx3_ASAP7_75t_L g370 ( 
.A(n_105),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_107),
.A2(n_108),
.B1(n_520),
.B2(n_521),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_107),
.B(n_517),
.C(n_520),
.Y(n_528)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_109),
.A2(n_132),
.B(n_134),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_109),
.A2(n_164),
.B(n_168),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_109),
.A2(n_132),
.B1(n_209),
.B2(n_257),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_109),
.A2(n_168),
.B(n_257),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_109),
.A2(n_132),
.B1(n_372),
.B2(n_433),
.Y(n_432)
);

INVx2_ASAP7_75t_SL g109 ( 
.A(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_110),
.B(n_169),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_110),
.A2(n_133),
.B1(n_393),
.B2(n_397),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_110),
.A2(n_133),
.B1(n_397),
.B2(n_420),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_110),
.A2(n_133),
.B1(n_420),
.B2(n_459),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_121),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_115),
.B1(n_118),
.B2(n_120),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx3_ASAP7_75t_L g396 ( 
.A(n_114),
.Y(n_396)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx5_ASAP7_75t_SL g210 ( 
.A(n_120),
.Y(n_210)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_121),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_121),
.A2(n_209),
.B(n_213),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_124),
.B1(n_127),
.B2(n_130),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_124),
.Y(n_205)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g184 ( 
.A(n_126),
.Y(n_184)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_126),
.Y(n_204)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx8_ASAP7_75t_L g233 ( 
.A(n_128),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_129),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_129),
.Y(n_190)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_132),
.A2(n_213),
.B(n_372),
.Y(n_371)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_133),
.B(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_134),
.Y(n_459)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx4_ASAP7_75t_L g422 ( 
.A(n_137),
.Y(n_422)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_138),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_140),
.Y(n_285)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_141),
.Y(n_166)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_141),
.Y(n_171)
);

INVx6_ASAP7_75t_L g403 ( 
.A(n_141),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g542 ( 
.A(n_142),
.B(n_148),
.Y(n_542)
);

INVx8_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx8_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_149),
.A2(n_263),
.B(n_267),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_149),
.B(n_308),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g484 ( 
.A1(n_149),
.A2(n_267),
.B(n_485),
.Y(n_484)
);

OR2x2_ASAP7_75t_L g546 ( 
.A(n_151),
.B(n_547),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_151),
.B(n_547),
.Y(n_550)
);

CKINVDCx20_ASAP7_75t_R g548 ( 
.A(n_152),
.Y(n_548)
);

BUFx3_ASAP7_75t_L g365 ( 
.A(n_153),
.Y(n_365)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_153),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_539),
.B(n_544),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_156),
.A2(n_511),
.B(n_536),
.Y(n_155)
);

OAI311xp33_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_378),
.A3(n_487),
.B1(n_505),
.C1(n_510),
.Y(n_156)
);

AOI21x1_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_320),
.B(n_377),
.Y(n_157)
);

AO21x1_ASAP7_75t_SL g158 ( 
.A1(n_159),
.A2(n_291),
.B(n_319),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_160),
.A2(n_251),
.B(n_290),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_216),
.B(n_250),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_181),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_162),
.B(n_181),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_163),
.B(n_174),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_163),
.A2(n_174),
.B1(n_175),
.B2(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_163),
.Y(n_248)
);

INVx11_ASAP7_75t_L g173 ( 
.A(n_166),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_167),
.A2(n_191),
.B(n_198),
.Y(n_225)
);

OAI21xp33_ASAP7_75t_SL g263 ( 
.A1(n_167),
.A2(n_264),
.B(n_265),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_167),
.B(n_341),
.Y(n_340)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx5_ASAP7_75t_L g259 ( 
.A(n_171),
.Y(n_259)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_173),
.Y(n_375)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_178),
.Y(n_175)
);

INVx3_ASAP7_75t_SL g176 ( 
.A(n_177),
.Y(n_176)
);

INVx5_ASAP7_75t_L g424 ( 
.A(n_177),
.Y(n_424)
);

BUFx3_ASAP7_75t_L g315 ( 
.A(n_179),
.Y(n_315)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_180),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_206),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_182),
.B(n_207),
.C(n_215),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_191),
.B(n_198),
.Y(n_182)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_183),
.Y(n_243)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx4_ASAP7_75t_SL g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_188),
.Y(n_279)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx5_ASAP7_75t_L g197 ( 
.A(n_190),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_190),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_191),
.A2(n_346),
.B1(n_347),
.B2(n_350),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_191),
.A2(n_384),
.B1(n_388),
.B2(n_391),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_SL g425 ( 
.A1(n_191),
.A2(n_391),
.B(n_426),
.Y(n_425)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_192),
.B(n_201),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_192),
.A2(n_242),
.B1(n_243),
.B2(n_244),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_192),
.A2(n_274),
.B1(n_312),
.B2(n_316),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_192),
.A2(n_351),
.B1(n_435),
.B2(n_436),
.Y(n_434)
);

OR2x2_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_195),
.Y(n_192)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_201),
.Y(n_198)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_204),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_207),
.A2(n_208),
.B1(n_214),
.B2(n_215),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_210),
.Y(n_260)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_240),
.B(n_249),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_226),
.B(n_239),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_225),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_224),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_221),
.Y(n_220)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

BUFx5_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

BUFx8_ASAP7_75t_L g277 ( 
.A(n_223),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_227),
.B(n_238),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_227),
.B(n_238),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_234),
.B(n_237),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_228),
.Y(n_242)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx3_ASAP7_75t_SL g234 ( 
.A(n_235),
.Y(n_234)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_236),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_237),
.A2(n_273),
.B(n_280),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_247),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_241),
.B(n_247),
.Y(n_249)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_246),
.Y(n_349)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_246),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_252),
.B(n_253),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_271),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_255),
.A2(n_256),
.B1(n_261),
.B2(n_262),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_256),
.B(n_261),
.C(n_271),
.Y(n_292)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVxp33_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

AOI32xp33_ASAP7_75t_L g281 ( 
.A1(n_266),
.A2(n_282),
.A3(n_283),
.B1(n_286),
.B2(n_289),
.Y(n_281)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_268),
.Y(n_308)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_270),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_281),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_272),
.B(n_281),
.Y(n_297)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

BUFx2_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx8_ASAP7_75t_L g353 ( 
.A(n_277),
.Y(n_353)
);

BUFx2_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx4_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx8_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_292),
.B(n_293),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_294),
.A2(n_295),
.B1(n_298),
.B2(n_318),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_SL g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_296),
.B(n_297),
.C(n_318),
.Y(n_321)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_298),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_SL g298 ( 
.A(n_299),
.B(n_309),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_299),
.B(n_310),
.C(n_311),
.Y(n_354)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

BUFx12f_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_303),
.Y(n_455)
);

INVx4_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_312),
.Y(n_346)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_322),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g377 ( 
.A(n_321),
.B(n_322),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_357),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_324),
.A2(n_354),
.B1(n_355),
.B2(n_356),
.Y(n_323)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_324),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_325),
.A2(n_326),
.B1(n_344),
.B2(n_345),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_326),
.B(n_344),
.Y(n_483)
);

OAI32xp33_ASAP7_75t_L g326 ( 
.A1(n_327),
.A2(n_330),
.A3(n_333),
.B1(n_336),
.B2(n_340),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_338),
.Y(n_336)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx3_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx8_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx4_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_354),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_354),
.B(n_355),
.C(n_357),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_358),
.A2(n_359),
.B1(n_366),
.B2(n_376),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_358),
.B(n_367),
.C(n_371),
.Y(n_496)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_366),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_SL g366 ( 
.A(n_367),
.B(n_371),
.Y(n_366)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_368),
.Y(n_485)
);

INVx4_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

NAND2xp33_ASAP7_75t_SL g378 ( 
.A(n_379),
.B(n_473),
.Y(n_378)
);

A2O1A1Ixp33_ASAP7_75t_SL g505 ( 
.A1(n_379),
.A2(n_473),
.B(n_506),
.C(n_509),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_445),
.Y(n_379)
);

OR2x2_ASAP7_75t_L g510 ( 
.A(n_380),
.B(n_445),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_417),
.C(n_430),
.Y(n_380)
);

FAx1_ASAP7_75t_SL g486 ( 
.A(n_381),
.B(n_417),
.CI(n_430),
.CON(n_486),
.SN(n_486)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_404),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_382),
.B(n_405),
.C(n_414),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_392),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_383),
.B(n_392),
.Y(n_479)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_384),
.Y(n_435)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx6_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx3_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_393),
.Y(n_433)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx5_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

BUFx2_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVx8_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_414),
.Y(n_404)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_406),
.Y(n_444)
);

INVx1_ASAP7_75t_SL g407 ( 
.A(n_408),
.Y(n_407)
);

INVx5_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx3_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g452 ( 
.A(n_411),
.Y(n_452)
);

INVx4_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_418),
.A2(n_419),
.B1(n_425),
.B2(n_429),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_419),
.B(n_425),
.Y(n_463)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_425),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_425),
.A2(n_429),
.B1(n_465),
.B2(n_466),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_L g514 ( 
.A1(n_425),
.A2(n_463),
.B(n_466),
.Y(n_514)
);

INVx4_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

INVx4_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_438),
.C(n_443),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_431),
.B(n_477),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_432),
.B(n_434),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_432),
.B(n_434),
.Y(n_495)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_438),
.A2(n_439),
.B1(n_443),
.B2(n_478),
.Y(n_477)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx4_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_443),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_447),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_446),
.B(n_449),
.C(n_461),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_448),
.A2(n_449),
.B1(n_461),
.B2(n_462),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

AOI21xp5_ASAP7_75t_L g449 ( 
.A1(n_450),
.A2(n_457),
.B(n_460),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_451),
.B(n_458),
.Y(n_460)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_453),
.Y(n_522)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

INVxp67_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

FAx1_ASAP7_75t_SL g513 ( 
.A(n_460),
.B(n_514),
.CI(n_515),
.CON(n_513),
.SN(n_513)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_460),
.B(n_514),
.C(n_515),
.Y(n_535)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_463),
.B(n_464),
.Y(n_462)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_472),
.Y(n_466)
);

INVxp67_ASAP7_75t_L g518 ( 
.A(n_468),
.Y(n_518)
);

INVx1_ASAP7_75t_SL g469 ( 
.A(n_470),
.Y(n_469)
);

INVx8_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_474),
.B(n_486),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_474),
.B(n_486),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_475),
.B(n_479),
.C(n_480),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_475),
.A2(n_476),
.B1(n_479),
.B2(n_499),
.Y(n_498)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_479),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_480),
.B(n_498),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_481),
.B(n_483),
.C(n_484),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g492 ( 
.A1(n_481),
.A2(n_482),
.B1(n_484),
.B2(n_493),
.Y(n_492)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_483),
.B(n_492),
.Y(n_491)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_484),
.Y(n_493)
);

BUFx24_ASAP7_75t_SL g551 ( 
.A(n_486),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_488),
.B(n_500),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_L g506 ( 
.A1(n_489),
.A2(n_507),
.B(n_508),
.Y(n_506)
);

NOR2x1_ASAP7_75t_L g489 ( 
.A(n_490),
.B(n_497),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_490),
.B(n_497),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_491),
.B(n_494),
.C(n_496),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_491),
.B(n_503),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_494),
.A2(n_495),
.B1(n_496),
.B2(n_504),
.Y(n_503)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_496),
.Y(n_504)
);

OR2x2_ASAP7_75t_L g500 ( 
.A(n_501),
.B(n_502),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_501),
.B(n_502),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_512),
.B(n_525),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_SL g512 ( 
.A(n_513),
.B(n_524),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_513),
.B(n_524),
.Y(n_537)
);

BUFx24_ASAP7_75t_SL g553 ( 
.A(n_513),
.Y(n_553)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_516),
.A2(n_517),
.B1(n_519),
.B2(n_523),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_516),
.A2(n_517),
.B1(n_531),
.B2(n_532),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_516),
.B(n_527),
.C(n_531),
.Y(n_543)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_519),
.Y(n_523)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_L g536 ( 
.A1(n_525),
.A2(n_537),
.B(n_538),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_SL g525 ( 
.A(n_526),
.B(n_535),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_526),
.B(n_535),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_L g526 ( 
.A1(n_527),
.A2(n_528),
.B1(n_529),
.B2(n_530),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_528),
.Y(n_527)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_530),
.Y(n_529)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_532),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_540),
.B(n_543),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_540),
.B(n_543),
.Y(n_544)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_542),
.Y(n_541)
);

CKINVDCx14_ASAP7_75t_R g549 ( 
.A(n_550),
.Y(n_549)
);


endmodule