module fake_aes_6575_n_662 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_662);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_662;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVxp33_ASAP7_75t_SL g78 ( .A(n_75), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_2), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_76), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_57), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_26), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_8), .Y(n_83) );
INVx2_ASAP7_75t_L g84 ( .A(n_15), .Y(n_84) );
INVxp33_ASAP7_75t_SL g85 ( .A(n_33), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_29), .Y(n_86) );
INVxp33_ASAP7_75t_SL g87 ( .A(n_20), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_28), .Y(n_88) );
INVx2_ASAP7_75t_SL g89 ( .A(n_44), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_30), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_45), .Y(n_91) );
BUFx6f_ASAP7_75t_L g92 ( .A(n_72), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_47), .Y(n_93) );
CKINVDCx14_ASAP7_75t_R g94 ( .A(n_68), .Y(n_94) );
INVxp33_ASAP7_75t_SL g95 ( .A(n_9), .Y(n_95) );
BUFx3_ASAP7_75t_L g96 ( .A(n_55), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_19), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_71), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_0), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_23), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_43), .Y(n_101) );
INVxp33_ASAP7_75t_L g102 ( .A(n_62), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_42), .Y(n_103) );
CKINVDCx14_ASAP7_75t_R g104 ( .A(n_65), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_49), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_14), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_69), .Y(n_107) );
INVxp67_ASAP7_75t_SL g108 ( .A(n_53), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_59), .Y(n_109) );
BUFx6f_ASAP7_75t_L g110 ( .A(n_34), .Y(n_110) );
INVxp33_ASAP7_75t_SL g111 ( .A(n_31), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_48), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_21), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_60), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_1), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_50), .Y(n_116) );
INVxp67_ASAP7_75t_SL g117 ( .A(n_46), .Y(n_117) );
INVx2_ASAP7_75t_L g118 ( .A(n_40), .Y(n_118) );
INVxp67_ASAP7_75t_L g119 ( .A(n_22), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_11), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_14), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_67), .Y(n_122) );
CKINVDCx16_ASAP7_75t_R g123 ( .A(n_70), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_39), .Y(n_124) );
BUFx2_ASAP7_75t_SL g125 ( .A(n_4), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_77), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_109), .Y(n_127) );
OAI22xp5_ASAP7_75t_SL g128 ( .A1(n_106), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_89), .B(n_3), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_123), .Y(n_130) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_92), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_94), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_84), .Y(n_133) );
HB1xp67_ASAP7_75t_L g134 ( .A(n_79), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_84), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_104), .Y(n_136) );
INVx3_ASAP7_75t_L g137 ( .A(n_79), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_83), .Y(n_138) );
AND2x4_ASAP7_75t_L g139 ( .A(n_83), .B(n_3), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_97), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_97), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_99), .Y(n_142) );
NAND2xp5_ASAP7_75t_SL g143 ( .A(n_89), .B(n_4), .Y(n_143) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_92), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_120), .B(n_5), .Y(n_145) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_92), .Y(n_146) );
INVxp67_ASAP7_75t_L g147 ( .A(n_125), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_109), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_99), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g150 ( .A(n_78), .Y(n_150) );
CKINVDCx16_ASAP7_75t_R g151 ( .A(n_96), .Y(n_151) );
CKINVDCx20_ASAP7_75t_R g152 ( .A(n_125), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_113), .Y(n_153) );
NOR2xp33_ASAP7_75t_L g154 ( .A(n_87), .B(n_5), .Y(n_154) );
CKINVDCx5p33_ASAP7_75t_R g155 ( .A(n_85), .Y(n_155) );
CKINVDCx5p33_ASAP7_75t_R g156 ( .A(n_111), .Y(n_156) );
BUFx2_ASAP7_75t_L g157 ( .A(n_113), .Y(n_157) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_92), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_115), .Y(n_159) );
CKINVDCx5p33_ASAP7_75t_R g160 ( .A(n_90), .Y(n_160) );
NAND2xp33_ASAP7_75t_R g161 ( .A(n_95), .B(n_27), .Y(n_161) );
INVxp67_ASAP7_75t_L g162 ( .A(n_115), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_121), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_121), .Y(n_164) );
CKINVDCx20_ASAP7_75t_R g165 ( .A(n_91), .Y(n_165) );
BUFx2_ASAP7_75t_L g166 ( .A(n_96), .Y(n_166) );
AOI22xp5_ASAP7_75t_L g167 ( .A1(n_102), .A2(n_6), .B1(n_7), .B2(n_8), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_80), .Y(n_168) );
CKINVDCx5p33_ASAP7_75t_R g169 ( .A(n_105), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_137), .Y(n_170) );
BUFx3_ASAP7_75t_L g171 ( .A(n_166), .Y(n_171) );
AND2x4_ASAP7_75t_L g172 ( .A(n_139), .B(n_126), .Y(n_172) );
AND2x6_ASAP7_75t_L g173 ( .A(n_139), .B(n_126), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_137), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_137), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_146), .Y(n_176) );
OAI221xp5_ASAP7_75t_L g177 ( .A1(n_162), .A2(n_119), .B1(n_108), .B2(n_117), .C(n_103), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_127), .Y(n_178) );
AND2x6_ASAP7_75t_L g179 ( .A(n_139), .B(n_124), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_127), .Y(n_180) );
BUFx3_ASAP7_75t_L g181 ( .A(n_160), .Y(n_181) );
OR2x2_ASAP7_75t_L g182 ( .A(n_157), .B(n_124), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_151), .B(n_116), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_146), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_148), .Y(n_185) );
AND2x4_ASAP7_75t_L g186 ( .A(n_134), .B(n_122), .Y(n_186) );
BUFx6f_ASAP7_75t_L g187 ( .A(n_131), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_168), .B(n_118), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_146), .Y(n_189) );
AOI22xp33_ASAP7_75t_L g190 ( .A1(n_138), .A2(n_122), .B1(n_80), .B2(n_114), .Y(n_190) );
INVx3_ASAP7_75t_L g191 ( .A(n_148), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_140), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_141), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_150), .B(n_101), .Y(n_194) );
BUFx2_ASAP7_75t_L g195 ( .A(n_132), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_146), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_142), .Y(n_197) );
OAI22xp33_ASAP7_75t_L g198 ( .A1(n_167), .A2(n_98), .B1(n_114), .B2(n_112), .Y(n_198) );
INVx4_ASAP7_75t_L g199 ( .A(n_131), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_131), .Y(n_200) );
AND2x2_ASAP7_75t_L g201 ( .A(n_149), .B(n_98), .Y(n_201) );
INVx4_ASAP7_75t_L g202 ( .A(n_131), .Y(n_202) );
INVx3_ASAP7_75t_L g203 ( .A(n_153), .Y(n_203) );
AOI22x1_ASAP7_75t_L g204 ( .A1(n_159), .A2(n_93), .B1(n_112), .B2(n_82), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_132), .B(n_93), .Y(n_205) );
BUFx6f_ASAP7_75t_L g206 ( .A(n_131), .Y(n_206) );
OAI22xp5_ASAP7_75t_L g207 ( .A1(n_152), .A2(n_81), .B1(n_82), .B2(n_107), .Y(n_207) );
AND2x2_ASAP7_75t_L g208 ( .A(n_163), .B(n_100), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_164), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_133), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_135), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_144), .Y(n_212) );
INVx4_ASAP7_75t_L g213 ( .A(n_144), .Y(n_213) );
BUFx6f_ASAP7_75t_L g214 ( .A(n_144), .Y(n_214) );
BUFx2_ASAP7_75t_L g215 ( .A(n_136), .Y(n_215) );
AO22x2_ASAP7_75t_L g216 ( .A1(n_129), .A2(n_107), .B1(n_103), .B2(n_100), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g217 ( .A(n_150), .B(n_118), .Y(n_217) );
BUFx10_ASAP7_75t_L g218 ( .A(n_136), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_144), .Y(n_219) );
INVx3_ASAP7_75t_L g220 ( .A(n_144), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_158), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_158), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_158), .Y(n_223) );
AND2x2_ASAP7_75t_L g224 ( .A(n_147), .B(n_88), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_160), .B(n_88), .Y(n_225) );
AND2x2_ASAP7_75t_L g226 ( .A(n_169), .B(n_86), .Y(n_226) );
INVxp33_ASAP7_75t_L g227 ( .A(n_154), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_158), .Y(n_228) );
NAND3x1_ASAP7_75t_L g229 ( .A(n_145), .B(n_81), .C(n_86), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_158), .Y(n_230) );
BUFx6f_ASAP7_75t_L g231 ( .A(n_143), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_169), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_128), .Y(n_233) );
NAND2x1p5_ASAP7_75t_L g234 ( .A(n_181), .B(n_92), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_170), .Y(n_235) );
AND2x4_ASAP7_75t_SL g236 ( .A(n_218), .B(n_165), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_170), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_174), .Y(n_238) );
OR2x2_ASAP7_75t_L g239 ( .A(n_171), .B(n_130), .Y(n_239) );
NAND2xp33_ASAP7_75t_R g240 ( .A(n_195), .B(n_215), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_186), .B(n_155), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_186), .B(n_155), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_186), .B(n_156), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_174), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_175), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_227), .B(n_156), .Y(n_246) );
BUFx2_ASAP7_75t_L g247 ( .A(n_171), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_186), .B(n_130), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_175), .Y(n_249) );
INVx3_ASAP7_75t_L g250 ( .A(n_191), .Y(n_250) );
NOR3xp33_ASAP7_75t_SL g251 ( .A(n_198), .B(n_161), .C(n_152), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_203), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g253 ( .A(n_217), .B(n_110), .Y(n_253) );
NAND2x1p5_ASAP7_75t_L g254 ( .A(n_181), .B(n_110), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_203), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_191), .Y(n_256) );
AND3x1_ASAP7_75t_SL g257 ( .A(n_233), .B(n_9), .C(n_10), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_191), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_224), .B(n_110), .Y(n_259) );
HB1xp67_ASAP7_75t_L g260 ( .A(n_195), .Y(n_260) );
INVx5_ASAP7_75t_L g261 ( .A(n_173), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g262 ( .A(n_194), .B(n_110), .Y(n_262) );
INVx3_ASAP7_75t_L g263 ( .A(n_191), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_203), .Y(n_264) );
INVx3_ASAP7_75t_L g265 ( .A(n_173), .Y(n_265) );
BUFx8_ASAP7_75t_SL g266 ( .A(n_215), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_224), .B(n_110), .Y(n_267) );
INVx5_ASAP7_75t_L g268 ( .A(n_173), .Y(n_268) );
HB1xp67_ASAP7_75t_L g269 ( .A(n_182), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_210), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_210), .Y(n_271) );
NAND2xp5_ASAP7_75t_SL g272 ( .A(n_231), .B(n_36), .Y(n_272) );
HB1xp67_ASAP7_75t_L g273 ( .A(n_182), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_211), .Y(n_274) );
OR2x2_ASAP7_75t_L g275 ( .A(n_207), .B(n_10), .Y(n_275) );
NOR2xp33_ASAP7_75t_R g276 ( .A(n_218), .B(n_11), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_211), .Y(n_277) );
AND2x2_ASAP7_75t_SL g278 ( .A(n_172), .B(n_12), .Y(n_278) );
NAND2xp33_ASAP7_75t_SL g279 ( .A(n_231), .B(n_12), .Y(n_279) );
HB1xp67_ASAP7_75t_L g280 ( .A(n_183), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_178), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_178), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_180), .Y(n_283) );
BUFx3_ASAP7_75t_L g284 ( .A(n_173), .Y(n_284) );
BUFx3_ASAP7_75t_L g285 ( .A(n_173), .Y(n_285) );
BUFx3_ASAP7_75t_L g286 ( .A(n_173), .Y(n_286) );
NOR2xp33_ASAP7_75t_SL g287 ( .A(n_218), .B(n_13), .Y(n_287) );
XOR2xp5_ASAP7_75t_L g288 ( .A(n_232), .B(n_13), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_180), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_185), .Y(n_290) );
A2O1A1Ixp33_ASAP7_75t_L g291 ( .A1(n_192), .A2(n_15), .B(n_16), .C(n_17), .Y(n_291) );
BUFx6f_ASAP7_75t_L g292 ( .A(n_173), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_192), .B(n_16), .Y(n_293) );
NOR2xp33_ASAP7_75t_L g294 ( .A(n_205), .B(n_41), .Y(n_294) );
OR2x6_ASAP7_75t_L g295 ( .A(n_216), .B(n_17), .Y(n_295) );
INVx1_ASAP7_75t_SL g296 ( .A(n_226), .Y(n_296) );
INVx6_ASAP7_75t_L g297 ( .A(n_231), .Y(n_297) );
NOR2xp33_ASAP7_75t_R g298 ( .A(n_218), .B(n_18), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_193), .B(n_18), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_185), .Y(n_300) );
AND2x2_ASAP7_75t_L g301 ( .A(n_201), .B(n_19), .Y(n_301) );
INVx1_ASAP7_75t_SL g302 ( .A(n_247), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_237), .Y(n_303) );
INVxp67_ASAP7_75t_SL g304 ( .A(n_292), .Y(n_304) );
AOI21xp5_ASAP7_75t_L g305 ( .A1(n_252), .A2(n_172), .B(n_225), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_237), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_245), .Y(n_307) );
AOI22xp5_ASAP7_75t_L g308 ( .A1(n_278), .A2(n_179), .B1(n_226), .B2(n_232), .Y(n_308) );
AOI22xp5_ASAP7_75t_L g309 ( .A1(n_278), .A2(n_179), .B1(n_233), .B2(n_216), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_245), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_270), .Y(n_311) );
BUFx3_ASAP7_75t_L g312 ( .A(n_292), .Y(n_312) );
NOR2xp33_ASAP7_75t_L g313 ( .A(n_241), .B(n_177), .Y(n_313) );
AND2x4_ASAP7_75t_L g314 ( .A(n_284), .B(n_201), .Y(n_314) );
BUFx8_ASAP7_75t_L g315 ( .A(n_239), .Y(n_315) );
INVx1_ASAP7_75t_SL g316 ( .A(n_260), .Y(n_316) );
BUFx6f_ASAP7_75t_L g317 ( .A(n_292), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_271), .Y(n_318) );
AND2x4_ASAP7_75t_L g319 ( .A(n_284), .B(n_208), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_274), .Y(n_320) );
BUFx6f_ASAP7_75t_L g321 ( .A(n_292), .Y(n_321) );
INVx2_ASAP7_75t_SL g322 ( .A(n_285), .Y(n_322) );
AOI22xp33_ASAP7_75t_L g323 ( .A1(n_295), .A2(n_179), .B1(n_216), .B2(n_172), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_281), .Y(n_324) );
NOR2x1_ASAP7_75t_SL g325 ( .A(n_295), .B(n_209), .Y(n_325) );
INVx3_ASAP7_75t_L g326 ( .A(n_285), .Y(n_326) );
AOI22xp5_ASAP7_75t_L g327 ( .A1(n_296), .A2(n_179), .B1(n_216), .B2(n_172), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_277), .Y(n_328) );
AOI22xp5_ASAP7_75t_L g329 ( .A1(n_246), .A2(n_179), .B1(n_229), .B2(n_231), .Y(n_329) );
INVx3_ASAP7_75t_L g330 ( .A(n_286), .Y(n_330) );
AND2x4_ASAP7_75t_L g331 ( .A(n_286), .B(n_208), .Y(n_331) );
BUFx6f_ASAP7_75t_L g332 ( .A(n_261), .Y(n_332) );
BUFx4f_ASAP7_75t_SL g333 ( .A(n_239), .Y(n_333) );
O2A1O1Ixp33_ASAP7_75t_L g334 ( .A1(n_269), .A2(n_209), .B(n_193), .C(n_197), .Y(n_334) );
NAND2xp5_ASAP7_75t_SL g335 ( .A(n_261), .B(n_231), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_301), .Y(n_336) );
CKINVDCx11_ASAP7_75t_R g337 ( .A(n_295), .Y(n_337) );
BUFx3_ASAP7_75t_L g338 ( .A(n_261), .Y(n_338) );
CKINVDCx20_ASAP7_75t_R g339 ( .A(n_266), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_301), .Y(n_340) );
O2A1O1Ixp5_ASAP7_75t_L g341 ( .A1(n_272), .A2(n_188), .B(n_197), .C(n_202), .Y(n_341) );
BUFx2_ASAP7_75t_L g342 ( .A(n_295), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_281), .Y(n_343) );
BUFx2_ASAP7_75t_L g344 ( .A(n_276), .Y(n_344) );
NOR2xp33_ASAP7_75t_L g345 ( .A(n_242), .B(n_179), .Y(n_345) );
INVx5_ASAP7_75t_L g346 ( .A(n_261), .Y(n_346) );
AOI21xp5_ASAP7_75t_L g347 ( .A1(n_255), .A2(n_204), .B(n_190), .Y(n_347) );
OAI22xp33_ASAP7_75t_L g348 ( .A1(n_275), .A2(n_240), .B1(n_273), .B2(n_287), .Y(n_348) );
OR2x2_ASAP7_75t_L g349 ( .A(n_236), .B(n_20), .Y(n_349) );
INVx4_ASAP7_75t_L g350 ( .A(n_261), .Y(n_350) );
BUFx6f_ASAP7_75t_L g351 ( .A(n_268), .Y(n_351) );
NOR2x1_ASAP7_75t_SL g352 ( .A(n_268), .B(n_179), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_235), .Y(n_353) );
BUFx6f_ASAP7_75t_L g354 ( .A(n_268), .Y(n_354) );
AOI22xp33_ASAP7_75t_L g355 ( .A1(n_337), .A2(n_275), .B1(n_243), .B2(n_248), .Y(n_355) );
AND2x4_ASAP7_75t_L g356 ( .A(n_314), .B(n_268), .Y(n_356) );
NOR2x1_ASAP7_75t_SL g357 ( .A(n_346), .B(n_268), .Y(n_357) );
INVx2_ASAP7_75t_SL g358 ( .A(n_315), .Y(n_358) );
BUFx2_ASAP7_75t_L g359 ( .A(n_315), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_353), .Y(n_360) );
INVxp67_ASAP7_75t_SL g361 ( .A(n_323), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_353), .Y(n_362) );
OR2x6_ASAP7_75t_L g363 ( .A(n_342), .B(n_234), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_303), .Y(n_364) );
OR2x6_ASAP7_75t_SL g365 ( .A(n_337), .B(n_266), .Y(n_365) );
OAI221xp5_ASAP7_75t_L g366 ( .A1(n_309), .A2(n_251), .B1(n_240), .B2(n_291), .C(n_299), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_324), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g368 ( .A(n_333), .B(n_280), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_303), .Y(n_369) );
OR2x2_ASAP7_75t_L g370 ( .A(n_316), .B(n_236), .Y(n_370) );
NAND2xp33_ASAP7_75t_SL g371 ( .A(n_342), .B(n_276), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_306), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_306), .Y(n_373) );
AOI21x1_ASAP7_75t_L g374 ( .A1(n_347), .A2(n_272), .B(n_267), .Y(n_374) );
AOI22xp33_ASAP7_75t_L g375 ( .A1(n_348), .A2(n_298), .B1(n_264), .B2(n_279), .Y(n_375) );
BUFx2_ASAP7_75t_L g376 ( .A(n_315), .Y(n_376) );
A2O1A1Ixp33_ASAP7_75t_L g377 ( .A1(n_305), .A2(n_293), .B(n_294), .C(n_262), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_336), .B(n_300), .Y(n_378) );
OR2x2_ASAP7_75t_L g379 ( .A(n_302), .B(n_288), .Y(n_379) );
OAI22xp5_ASAP7_75t_L g380 ( .A1(n_327), .A2(n_234), .B1(n_254), .B2(n_283), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_324), .Y(n_381) );
NOR2x1_ASAP7_75t_SL g382 ( .A(n_346), .B(n_290), .Y(n_382) );
INVxp67_ASAP7_75t_SL g383 ( .A(n_325), .Y(n_383) );
NAND3x1_ASAP7_75t_L g384 ( .A(n_308), .B(n_257), .C(n_298), .Y(n_384) );
CKINVDCx5p33_ASAP7_75t_R g385 ( .A(n_339), .Y(n_385) );
BUFx2_ASAP7_75t_SL g386 ( .A(n_346), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_307), .Y(n_387) );
AOI221xp5_ASAP7_75t_L g388 ( .A1(n_355), .A2(n_313), .B1(n_334), .B2(n_340), .C(n_318), .Y(n_388) );
AOI22xp33_ASAP7_75t_SL g389 ( .A1(n_359), .A2(n_344), .B1(n_349), .B2(n_339), .Y(n_389) );
AOI22xp33_ASAP7_75t_L g390 ( .A1(n_361), .A2(n_349), .B1(n_345), .B2(n_344), .Y(n_390) );
AOI22xp5_ASAP7_75t_L g391 ( .A1(n_361), .A2(n_329), .B1(n_279), .B2(n_229), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_378), .B(n_311), .Y(n_392) );
CKINVDCx5p33_ASAP7_75t_R g393 ( .A(n_365), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_360), .Y(n_394) );
BUFx2_ASAP7_75t_L g395 ( .A(n_363), .Y(n_395) );
OAI221xp5_ASAP7_75t_L g396 ( .A1(n_366), .A2(n_291), .B1(n_320), .B2(n_328), .C(n_259), .Y(n_396) );
NOR2xp33_ASAP7_75t_L g397 ( .A(n_379), .B(n_314), .Y(n_397) );
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_366), .A2(n_319), .B1(n_314), .B2(n_331), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_364), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_378), .B(n_343), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_360), .B(n_343), .Y(n_401) );
OAI22xp33_ASAP7_75t_L g402 ( .A1(n_365), .A2(n_310), .B1(n_307), .B2(n_254), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_362), .B(n_310), .Y(n_403) );
OAI22xp5_ASAP7_75t_L g404 ( .A1(n_380), .A2(n_289), .B1(n_282), .B2(n_331), .Y(n_404) );
AOI22xp33_ASAP7_75t_L g405 ( .A1(n_376), .A2(n_319), .B1(n_263), .B2(n_250), .Y(n_405) );
OAI22xp33_ASAP7_75t_L g406 ( .A1(n_370), .A2(n_204), .B1(n_322), .B2(n_265), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_364), .Y(n_407) );
AOI21xp5_ASAP7_75t_L g408 ( .A1(n_377), .A2(n_341), .B(n_253), .Y(n_408) );
OAI211xp5_ASAP7_75t_L g409 ( .A1(n_375), .A2(n_250), .B(n_263), .C(n_335), .Y(n_409) );
OAI22xp5_ASAP7_75t_L g410 ( .A1(n_362), .A2(n_322), .B1(n_312), .B2(n_321), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_364), .Y(n_411) );
OA21x2_ASAP7_75t_L g412 ( .A1(n_374), .A2(n_244), .B(n_238), .Y(n_412) );
OR2x2_ASAP7_75t_L g413 ( .A(n_367), .B(n_250), .Y(n_413) );
INVx3_ASAP7_75t_L g414 ( .A(n_399), .Y(n_414) );
OAI21xp5_ASAP7_75t_L g415 ( .A1(n_391), .A2(n_384), .B(n_371), .Y(n_415) );
OAI22xp33_ASAP7_75t_L g416 ( .A1(n_404), .A2(n_358), .B1(n_363), .B2(n_383), .Y(n_416) );
OAI211xp5_ASAP7_75t_L g417 ( .A1(n_389), .A2(n_368), .B(n_385), .C(n_335), .Y(n_417) );
AND2x6_ASAP7_75t_SL g418 ( .A(n_393), .B(n_363), .Y(n_418) );
OR2x6_ASAP7_75t_L g419 ( .A(n_395), .B(n_386), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_399), .Y(n_420) );
BUFx3_ASAP7_75t_L g421 ( .A(n_395), .Y(n_421) );
INVxp67_ASAP7_75t_L g422 ( .A(n_397), .Y(n_422) );
NAND2x1_ASAP7_75t_L g423 ( .A(n_399), .B(n_369), .Y(n_423) );
CKINVDCx16_ASAP7_75t_R g424 ( .A(n_401), .Y(n_424) );
CKINVDCx5p33_ASAP7_75t_R g425 ( .A(n_392), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_407), .Y(n_426) );
OR2x2_ASAP7_75t_L g427 ( .A(n_394), .B(n_367), .Y(n_427) );
OAI22xp5_ASAP7_75t_L g428 ( .A1(n_398), .A2(n_384), .B1(n_381), .B2(n_372), .Y(n_428) );
OAI22xp5_ASAP7_75t_L g429 ( .A1(n_390), .A2(n_384), .B1(n_381), .B2(n_372), .Y(n_429) );
CKINVDCx20_ASAP7_75t_R g430 ( .A(n_400), .Y(n_430) );
OAI33xp33_ASAP7_75t_L g431 ( .A1(n_402), .A2(n_230), .A3(n_212), .B1(n_219), .B2(n_228), .B3(n_249), .Y(n_431) );
AO21x2_ASAP7_75t_L g432 ( .A1(n_408), .A2(n_374), .B(n_387), .Y(n_432) );
OAI22xp33_ASAP7_75t_L g433 ( .A1(n_391), .A2(n_387), .B1(n_369), .B2(n_373), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_407), .Y(n_434) );
AOI22xp33_ASAP7_75t_L g435 ( .A1(n_388), .A2(n_356), .B1(n_386), .B2(n_373), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_401), .B(n_372), .Y(n_436) );
BUFx3_ASAP7_75t_L g437 ( .A(n_407), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_403), .B(n_369), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_411), .Y(n_439) );
OR2x2_ASAP7_75t_L g440 ( .A(n_394), .B(n_356), .Y(n_440) );
OAI22xp5_ASAP7_75t_L g441 ( .A1(n_400), .A2(n_356), .B1(n_312), .B2(n_321), .Y(n_441) );
AO21x2_ASAP7_75t_L g442 ( .A1(n_408), .A2(n_382), .B(n_352), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_411), .Y(n_443) );
CKINVDCx5p33_ASAP7_75t_R g444 ( .A(n_392), .Y(n_444) );
AOI222xp33_ASAP7_75t_L g445 ( .A1(n_396), .A2(n_382), .B1(n_357), .B2(n_258), .C1(n_256), .C2(n_304), .Y(n_445) );
AND2x2_ASAP7_75t_SL g446 ( .A(n_424), .B(n_411), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_424), .B(n_403), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_420), .Y(n_448) );
OAI22xp5_ASAP7_75t_L g449 ( .A1(n_430), .A2(n_396), .B1(n_409), .B2(n_413), .Y(n_449) );
HB1xp67_ASAP7_75t_L g450 ( .A(n_425), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_420), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_436), .B(n_412), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_426), .Y(n_453) );
OAI33xp33_ASAP7_75t_L g454 ( .A1(n_444), .A2(n_406), .A3(n_413), .B1(n_410), .B2(n_230), .B3(n_228), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_426), .Y(n_455) );
AOI221xp5_ASAP7_75t_L g456 ( .A1(n_422), .A2(n_405), .B1(n_409), .B2(n_410), .C(n_213), .Y(n_456) );
HB1xp67_ASAP7_75t_L g457 ( .A(n_438), .Y(n_457) );
INVx1_ASAP7_75t_SL g458 ( .A(n_437), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_438), .B(n_412), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_434), .B(n_412), .Y(n_460) );
HB1xp67_ASAP7_75t_L g461 ( .A(n_437), .Y(n_461) );
HB1xp67_ASAP7_75t_L g462 ( .A(n_437), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_434), .B(n_412), .Y(n_463) );
OAI31xp33_ASAP7_75t_L g464 ( .A1(n_416), .A2(n_428), .A3(n_429), .B(n_417), .Y(n_464) );
NAND2xp5_ASAP7_75t_SL g465 ( .A(n_415), .B(n_346), .Y(n_465) );
NAND4xp25_ASAP7_75t_L g466 ( .A(n_435), .B(n_21), .C(n_199), .D(n_213), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_434), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_439), .B(n_24), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_439), .B(n_25), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_439), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_443), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_443), .Y(n_472) );
NAND3xp33_ASAP7_75t_L g473 ( .A(n_445), .B(n_214), .C(n_206), .Y(n_473) );
BUFx2_ASAP7_75t_L g474 ( .A(n_419), .Y(n_474) );
OR2x2_ASAP7_75t_SL g475 ( .A(n_427), .B(n_351), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_443), .B(n_32), .Y(n_476) );
OAI31xp33_ASAP7_75t_L g477 ( .A1(n_433), .A2(n_265), .A3(n_338), .B(n_330), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_427), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_414), .Y(n_479) );
OAI33xp33_ASAP7_75t_L g480 ( .A1(n_440), .A2(n_212), .A3(n_219), .B1(n_196), .B2(n_189), .B3(n_184), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_414), .B(n_297), .Y(n_481) );
INVx2_ASAP7_75t_SL g482 ( .A(n_419), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_414), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_414), .B(n_35), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_432), .Y(n_485) );
HB1xp67_ASAP7_75t_L g486 ( .A(n_440), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_423), .Y(n_487) );
INVx2_ASAP7_75t_SL g488 ( .A(n_419), .Y(n_488) );
BUFx3_ASAP7_75t_L g489 ( .A(n_419), .Y(n_489) );
INVx2_ASAP7_75t_SL g490 ( .A(n_419), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_432), .Y(n_491) );
NAND3xp33_ASAP7_75t_L g492 ( .A(n_445), .B(n_214), .C(n_206), .Y(n_492) );
AOI33xp33_ASAP7_75t_L g493 ( .A1(n_418), .A2(n_196), .A3(n_184), .B1(n_189), .B2(n_176), .B3(n_223), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_421), .B(n_37), .Y(n_494) );
NAND2xp33_ASAP7_75t_SL g495 ( .A(n_474), .B(n_423), .Y(n_495) );
CKINVDCx16_ASAP7_75t_R g496 ( .A(n_450), .Y(n_496) );
AOI221xp5_ASAP7_75t_L g497 ( .A1(n_449), .A2(n_431), .B1(n_421), .B2(n_441), .C(n_432), .Y(n_497) );
AO21x2_ASAP7_75t_L g498 ( .A1(n_473), .A2(n_442), .B(n_200), .Y(n_498) );
BUFx2_ASAP7_75t_L g499 ( .A(n_475), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_478), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_460), .B(n_421), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_457), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_486), .Y(n_503) );
INVx2_ASAP7_75t_SL g504 ( .A(n_461), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_460), .B(n_442), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_463), .B(n_442), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_447), .B(n_418), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_475), .Y(n_508) );
HB1xp67_ASAP7_75t_L g509 ( .A(n_447), .Y(n_509) );
OR2x2_ASAP7_75t_L g510 ( .A(n_452), .B(n_38), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_448), .Y(n_511) );
NAND4xp25_ASAP7_75t_L g512 ( .A(n_464), .B(n_199), .C(n_202), .D(n_213), .Y(n_512) );
OR2x2_ASAP7_75t_L g513 ( .A(n_452), .B(n_51), .Y(n_513) );
CKINVDCx16_ASAP7_75t_R g514 ( .A(n_489), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_467), .Y(n_515) );
INVxp67_ASAP7_75t_SL g516 ( .A(n_462), .Y(n_516) );
INVxp67_ASAP7_75t_L g517 ( .A(n_446), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_451), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_467), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_451), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_466), .B(n_52), .Y(n_521) );
OAI211xp5_ASAP7_75t_SL g522 ( .A1(n_464), .A2(n_176), .B(n_223), .C(n_222), .Y(n_522) );
NOR2x1_ASAP7_75t_L g523 ( .A(n_473), .B(n_350), .Y(n_523) );
HB1xp67_ASAP7_75t_L g524 ( .A(n_446), .Y(n_524) );
CKINVDCx5p33_ASAP7_75t_R g525 ( .A(n_446), .Y(n_525) );
NAND5xp2_ASAP7_75t_L g526 ( .A(n_456), .B(n_357), .C(n_56), .D(n_58), .E(n_61), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_453), .Y(n_527) );
OAI31xp33_ASAP7_75t_L g528 ( .A1(n_492), .A2(n_265), .A3(n_338), .B(n_330), .Y(n_528) );
INVx2_ASAP7_75t_SL g529 ( .A(n_489), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_463), .B(n_54), .Y(n_530) );
INVx2_ASAP7_75t_L g531 ( .A(n_467), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_471), .B(n_63), .Y(n_532) );
AND2x4_ASAP7_75t_L g533 ( .A(n_489), .B(n_64), .Y(n_533) );
NAND2xp33_ASAP7_75t_R g534 ( .A(n_474), .B(n_66), .Y(n_534) );
BUFx2_ASAP7_75t_L g535 ( .A(n_494), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_455), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_455), .B(n_297), .Y(n_537) );
HB1xp67_ASAP7_75t_L g538 ( .A(n_470), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_470), .B(n_73), .Y(n_539) );
BUFx2_ASAP7_75t_L g540 ( .A(n_494), .Y(n_540) );
OR2x6_ASAP7_75t_L g541 ( .A(n_482), .B(n_488), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_471), .B(n_74), .Y(n_542) );
OAI21xp5_ASAP7_75t_SL g543 ( .A1(n_499), .A2(n_492), .B(n_490), .Y(n_543) );
NOR2xp67_ASAP7_75t_L g544 ( .A(n_504), .B(n_482), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_502), .B(n_472), .Y(n_545) );
AOI211xp5_ASAP7_75t_L g546 ( .A1(n_499), .A2(n_465), .B(n_490), .C(n_488), .Y(n_546) );
OAI21xp33_ASAP7_75t_L g547 ( .A1(n_508), .A2(n_493), .B(n_487), .Y(n_547) );
A2O1A1O1Ixp25_ASAP7_75t_L g548 ( .A1(n_507), .A2(n_487), .B(n_479), .C(n_483), .D(n_454), .Y(n_548) );
NOR3xp33_ASAP7_75t_L g549 ( .A(n_521), .B(n_480), .C(n_481), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_509), .B(n_458), .Y(n_550) );
OAI22xp5_ASAP7_75t_L g551 ( .A1(n_535), .A2(n_458), .B1(n_459), .B2(n_471), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_503), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_500), .B(n_483), .Y(n_553) );
NAND3xp33_ASAP7_75t_SL g554 ( .A(n_528), .B(n_477), .C(n_484), .Y(n_554) );
NOR3xp33_ASAP7_75t_L g555 ( .A(n_521), .B(n_481), .C(n_484), .Y(n_555) );
HB1xp67_ASAP7_75t_L g556 ( .A(n_538), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_540), .B(n_491), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_504), .B(n_491), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_501), .B(n_485), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_501), .B(n_485), .Y(n_560) );
OR2x2_ASAP7_75t_L g561 ( .A(n_516), .B(n_476), .Y(n_561) );
INVx2_ASAP7_75t_SL g562 ( .A(n_541), .Y(n_562) );
AOI21xp33_ASAP7_75t_L g563 ( .A1(n_534), .A2(n_476), .B(n_469), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_511), .Y(n_564) );
NOR2xp33_ASAP7_75t_L g565 ( .A(n_496), .B(n_517), .Y(n_565) );
CKINVDCx14_ASAP7_75t_R g566 ( .A(n_525), .Y(n_566) );
INVxp33_ASAP7_75t_L g567 ( .A(n_523), .Y(n_567) );
AOI322xp5_ASAP7_75t_L g568 ( .A1(n_495), .A2(n_469), .A3(n_468), .B1(n_222), .B2(n_221), .C1(n_326), .C2(n_220), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_514), .B(n_468), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_518), .B(n_199), .Y(n_570) );
OAI31xp33_ASAP7_75t_SL g571 ( .A1(n_526), .A2(n_346), .A3(n_221), .B(n_350), .Y(n_571) );
AOI21xp33_ASAP7_75t_L g572 ( .A1(n_534), .A2(n_187), .B(n_206), .Y(n_572) );
NAND2x1p5_ASAP7_75t_L g573 ( .A(n_533), .B(n_317), .Y(n_573) );
OR2x2_ASAP7_75t_L g574 ( .A(n_505), .B(n_199), .Y(n_574) );
AOI222xp33_ASAP7_75t_L g575 ( .A1(n_497), .A2(n_202), .B1(n_187), .B2(n_206), .C1(n_214), .C2(n_326), .Y(n_575) );
OAI21xp33_ASAP7_75t_L g576 ( .A1(n_506), .A2(n_187), .B(n_206), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_520), .B(n_202), .Y(n_577) );
AOI32xp33_ASAP7_75t_L g578 ( .A1(n_495), .A2(n_350), .A3(n_220), .B1(n_317), .B2(n_321), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_527), .Y(n_579) );
NOR2x1_ASAP7_75t_SL g580 ( .A(n_541), .B(n_354), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_506), .B(n_187), .Y(n_581) );
OAI22xp5_ASAP7_75t_SL g582 ( .A1(n_525), .A2(n_321), .B1(n_317), .B2(n_354), .Y(n_582) );
AOI22xp5_ASAP7_75t_L g583 ( .A1(n_524), .A2(n_317), .B1(n_351), .B2(n_332), .Y(n_583) );
AO21x1_ASAP7_75t_L g584 ( .A1(n_533), .A2(n_187), .B(n_214), .Y(n_584) );
INVx1_ASAP7_75t_SL g585 ( .A(n_530), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_536), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_559), .B(n_541), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_556), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_556), .Y(n_589) );
NOR3xp33_ASAP7_75t_L g590 ( .A(n_547), .B(n_522), .C(n_512), .Y(n_590) );
INVx1_ASAP7_75t_SL g591 ( .A(n_550), .Y(n_591) );
INVxp67_ASAP7_75t_SL g592 ( .A(n_558), .Y(n_592) );
INVx1_ASAP7_75t_SL g593 ( .A(n_585), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_560), .B(n_541), .Y(n_594) );
NAND2xp5_ASAP7_75t_SL g595 ( .A(n_578), .B(n_533), .Y(n_595) );
NOR3xp33_ASAP7_75t_SL g596 ( .A(n_543), .B(n_539), .C(n_537), .Y(n_596) );
XOR2xp5_ASAP7_75t_L g597 ( .A(n_566), .B(n_513), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_552), .Y(n_598) );
OAI21xp33_ASAP7_75t_L g599 ( .A1(n_567), .A2(n_529), .B(n_513), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_564), .Y(n_600) );
NAND2xp67_ASAP7_75t_L g601 ( .A(n_548), .B(n_542), .Y(n_601) );
INVx3_ASAP7_75t_L g602 ( .A(n_562), .Y(n_602) );
INVx2_ASAP7_75t_SL g603 ( .A(n_562), .Y(n_603) );
NOR2xp33_ASAP7_75t_L g604 ( .A(n_565), .B(n_510), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_579), .Y(n_605) );
INVx1_ASAP7_75t_SL g606 ( .A(n_569), .Y(n_606) );
NOR2xp33_ASAP7_75t_L g607 ( .A(n_565), .B(n_510), .Y(n_607) );
BUFx2_ASAP7_75t_L g608 ( .A(n_566), .Y(n_608) );
NOR3xp33_ASAP7_75t_SL g609 ( .A(n_554), .B(n_498), .C(n_542), .Y(n_609) );
INVxp67_ASAP7_75t_SL g610 ( .A(n_544), .Y(n_610) );
NAND3xp33_ASAP7_75t_L g611 ( .A(n_575), .B(n_532), .C(n_531), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_586), .B(n_519), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_545), .Y(n_613) );
INVxp67_ASAP7_75t_L g614 ( .A(n_580), .Y(n_614) );
NOR3x1_ASAP7_75t_L g615 ( .A(n_554), .B(n_498), .C(n_532), .Y(n_615) );
INVx1_ASAP7_75t_SL g616 ( .A(n_608), .Y(n_616) );
AOI22xp5_ASAP7_75t_L g617 ( .A1(n_604), .A2(n_555), .B1(n_549), .B2(n_551), .Y(n_617) );
INVxp67_ASAP7_75t_L g618 ( .A(n_588), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_589), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_592), .B(n_557), .Y(n_620) );
AND2x2_ASAP7_75t_L g621 ( .A(n_591), .B(n_567), .Y(n_621) );
OAI22xp5_ASAP7_75t_L g622 ( .A1(n_597), .A2(n_546), .B1(n_563), .B2(n_573), .Y(n_622) );
XOR2xp5_ASAP7_75t_L g623 ( .A(n_606), .B(n_574), .Y(n_623) );
NAND3xp33_ASAP7_75t_L g624 ( .A(n_609), .B(n_571), .C(n_568), .Y(n_624) );
AOI222xp33_ASAP7_75t_L g625 ( .A1(n_607), .A2(n_553), .B1(n_581), .B2(n_570), .C1(n_577), .C2(n_582), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_600), .Y(n_626) );
CKINVDCx20_ASAP7_75t_R g627 ( .A(n_593), .Y(n_627) );
AOI221xp5_ASAP7_75t_L g628 ( .A1(n_613), .A2(n_572), .B1(n_561), .B2(n_576), .C(n_515), .Y(n_628) );
AOI22xp33_ASAP7_75t_L g629 ( .A1(n_590), .A2(n_498), .B1(n_584), .B2(n_515), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_605), .Y(n_630) );
XNOR2xp5_ASAP7_75t_L g631 ( .A(n_601), .B(n_573), .Y(n_631) );
NAND2xp5_ASAP7_75t_SL g632 ( .A(n_614), .B(n_583), .Y(n_632) );
AND2x2_ASAP7_75t_L g633 ( .A(n_587), .B(n_214), .Y(n_633) );
A2O1A1Ixp33_ASAP7_75t_L g634 ( .A1(n_595), .A2(n_332), .B(n_354), .C(n_351), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_617), .B(n_601), .Y(n_635) );
NOR2xp33_ASAP7_75t_R g636 ( .A(n_627), .B(n_607), .Y(n_636) );
NOR2xp33_ASAP7_75t_L g637 ( .A(n_616), .B(n_598), .Y(n_637) );
NOR2xp33_ASAP7_75t_R g638 ( .A(n_631), .B(n_602), .Y(n_638) );
HB1xp67_ASAP7_75t_L g639 ( .A(n_618), .Y(n_639) );
A2O1A1Ixp33_ASAP7_75t_L g640 ( .A1(n_634), .A2(n_610), .B(n_595), .C(n_596), .Y(n_640) );
AND2x4_ASAP7_75t_L g641 ( .A(n_621), .B(n_602), .Y(n_641) );
NAND2xp33_ASAP7_75t_SL g642 ( .A(n_622), .B(n_603), .Y(n_642) );
OAI21xp5_ASAP7_75t_SL g643 ( .A1(n_634), .A2(n_599), .B(n_611), .Y(n_643) );
AOI21xp33_ASAP7_75t_SL g644 ( .A1(n_624), .A2(n_615), .B(n_587), .Y(n_644) );
NOR3xp33_ASAP7_75t_L g645 ( .A(n_632), .B(n_612), .C(n_594), .Y(n_645) );
AOI21xp33_ASAP7_75t_SL g646 ( .A1(n_625), .A2(n_354), .B(n_623), .Y(n_646) );
OAI211xp5_ASAP7_75t_L g647 ( .A1(n_629), .A2(n_628), .B(n_633), .C(n_620), .Y(n_647) );
NAND4xp25_ASAP7_75t_L g648 ( .A(n_629), .B(n_619), .C(n_630), .D(n_626), .Y(n_648) );
O2A1O1Ixp33_ASAP7_75t_L g649 ( .A1(n_634), .A2(n_616), .B(n_622), .C(n_450), .Y(n_649) );
NAND3xp33_ASAP7_75t_SL g650 ( .A(n_634), .B(n_627), .C(n_617), .Y(n_650) );
CKINVDCx5p33_ASAP7_75t_R g651 ( .A(n_636), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_639), .Y(n_652) );
XNOR2x1_ASAP7_75t_L g653 ( .A(n_635), .B(n_650), .Y(n_653) );
CKINVDCx5p33_ASAP7_75t_R g654 ( .A(n_638), .Y(n_654) );
NOR3xp33_ASAP7_75t_L g655 ( .A(n_652), .B(n_642), .C(n_649), .Y(n_655) );
NAND3xp33_ASAP7_75t_L g656 ( .A(n_653), .B(n_654), .C(n_651), .Y(n_656) );
NAND3x1_ASAP7_75t_L g657 ( .A(n_653), .B(n_645), .C(n_637), .Y(n_657) );
AOI21xp5_ASAP7_75t_L g658 ( .A1(n_656), .A2(n_640), .B(n_646), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_655), .Y(n_659) );
OAI22xp5_ASAP7_75t_SL g660 ( .A1(n_659), .A2(n_657), .B1(n_641), .B2(n_644), .Y(n_660) );
AOI22xp33_ASAP7_75t_L g661 ( .A1(n_660), .A2(n_658), .B1(n_648), .B2(n_645), .Y(n_661) );
AOI21xp5_ASAP7_75t_L g662 ( .A1(n_661), .A2(n_643), .B(n_647), .Y(n_662) );
endmodule