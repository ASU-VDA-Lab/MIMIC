module fake_jpeg_4072_n_344 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_344);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_344;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx2_ASAP7_75t_SL g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_37),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_39),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_27),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_17),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_28),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_17),
.B(n_15),
.Y(n_42)
);

AO22x1_ASAP7_75t_L g51 ( 
.A1(n_42),
.A2(n_48),
.B1(n_26),
.B2(n_35),
.Y(n_51)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

BUFx10_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx3_ASAP7_75t_SL g48 ( 
.A(n_26),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_49),
.B(n_54),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_51),
.B(n_53),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_32),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_41),
.A2(n_24),
.B1(n_23),
.B2(n_29),
.Y(n_56)
);

A2O1A1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_56),
.A2(n_30),
.B(n_29),
.C(n_39),
.Y(n_95)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_43),
.A2(n_23),
.B1(n_24),
.B2(n_26),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_58),
.A2(n_19),
.B1(n_22),
.B2(n_21),
.Y(n_77)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_59),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_63),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_43),
.A2(n_23),
.B1(n_32),
.B2(n_30),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_64),
.A2(n_71),
.B1(n_19),
.B2(n_21),
.Y(n_90)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx4_ASAP7_75t_SL g83 ( 
.A(n_68),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_42),
.B(n_19),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_69),
.B(n_26),
.Y(n_76)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

AO22x2_ASAP7_75t_L g71 ( 
.A1(n_42),
.A2(n_34),
.B1(n_31),
.B2(n_35),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_72),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_74),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_76),
.B(n_92),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_77),
.A2(n_86),
.B1(n_54),
.B2(n_65),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_61),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_79),
.B(n_80),
.Y(n_106)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_85),
.B(n_86),
.Y(n_110)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_36),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_87),
.B(n_22),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_90),
.A2(n_95),
.B1(n_21),
.B2(n_33),
.Y(n_125)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_73),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_91),
.B(n_94),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_71),
.Y(n_92)
);

BUFx10_ASAP7_75t_L g94 ( 
.A(n_59),
.Y(n_94)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_44),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_60),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_98),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_50),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_99),
.Y(n_109)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_101),
.B(n_111),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_76),
.B(n_53),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_102),
.B(n_104),
.Y(n_130)
);

OA21x2_ASAP7_75t_L g103 ( 
.A1(n_87),
.A2(n_71),
.B(n_56),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_103),
.A2(n_93),
.B(n_38),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_93),
.B(n_64),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_71),
.C(n_44),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_107),
.B(n_120),
.C(n_88),
.Y(n_133)
);

BUFx24_ASAP7_75t_SL g108 ( 
.A(n_81),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_108),
.Y(n_142)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_99),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_112),
.Y(n_137)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_84),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_113),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_114),
.Y(n_155)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_83),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_116),
.B(n_121),
.Y(n_140)
);

AO22x1_ASAP7_75t_SL g117 ( 
.A1(n_92),
.A2(n_49),
.B1(n_47),
.B2(n_65),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_117),
.A2(n_119),
.B1(n_80),
.B2(n_75),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_22),
.Y(n_118)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_118),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_83),
.B(n_44),
.C(n_68),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_122),
.B(n_125),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_99),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_123),
.Y(n_156)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_75),
.Y(n_124)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_124),
.Y(n_152)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_85),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_127),
.Y(n_143)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_94),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_128),
.B(n_129),
.Y(n_134)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_94),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_131),
.A2(n_141),
.B(n_150),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_133),
.B(n_114),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_122),
.B(n_93),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_135),
.B(n_136),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_115),
.B(n_100),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_103),
.A2(n_66),
.B1(n_52),
.B2(n_97),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_138),
.B(n_153),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_107),
.A2(n_52),
.B1(n_70),
.B2(n_88),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_139),
.A2(n_149),
.B1(n_157),
.B2(n_116),
.Y(n_166)
);

AND2x2_ASAP7_75t_SL g141 ( 
.A(n_115),
.B(n_47),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_115),
.B(n_100),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_144),
.B(n_145),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_102),
.B(n_78),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_120),
.B(n_104),
.C(n_125),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_147),
.B(n_126),
.C(n_129),
.Y(n_177)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_110),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_148),
.B(n_113),
.Y(n_175)
);

AO22x2_ASAP7_75t_L g149 ( 
.A1(n_117),
.A2(n_103),
.B1(n_118),
.B2(n_62),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_117),
.A2(n_33),
.B(n_28),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_103),
.A2(n_97),
.B1(n_96),
.B2(n_91),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_149),
.A2(n_117),
.B1(n_111),
.B2(n_124),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_158),
.A2(n_166),
.B1(n_176),
.B2(n_155),
.Y(n_194)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_134),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_159),
.B(n_162),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_160),
.B(n_173),
.Y(n_192)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_134),
.Y(n_162)
);

BUFx5_ASAP7_75t_L g163 ( 
.A(n_141),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_163),
.Y(n_206)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_151),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_164),
.B(n_170),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_130),
.B(n_105),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_169),
.B(n_172),
.Y(n_189)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_145),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_149),
.A2(n_105),
.B1(n_101),
.B2(n_128),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_171),
.A2(n_31),
.B(n_34),
.Y(n_207)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_151),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_135),
.B(n_106),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_140),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_174),
.B(n_178),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_175),
.Y(n_204)
);

AO21x2_ASAP7_75t_L g176 ( 
.A1(n_149),
.A2(n_31),
.B(n_34),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_177),
.B(n_185),
.Y(n_198)
);

OAI32xp33_ASAP7_75t_L g178 ( 
.A1(n_149),
.A2(n_78),
.A3(n_82),
.B1(n_31),
.B2(n_34),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_146),
.B(n_113),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_179),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_140),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_180),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_139),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_181),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_131),
.A2(n_123),
.B(n_112),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_182),
.A2(n_155),
.B(n_132),
.Y(n_195)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_143),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_183),
.Y(n_212)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_130),
.Y(n_184)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_184),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_133),
.B(n_109),
.C(n_127),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_136),
.B(n_109),
.Y(n_186)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_186),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_176),
.A2(n_149),
.B1(n_157),
.B2(n_141),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_187),
.A2(n_191),
.B1(n_201),
.B2(n_205),
.Y(n_224)
);

XNOR2x2_ASAP7_75t_SL g188 ( 
.A(n_163),
.B(n_141),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_188),
.A2(n_18),
.B(n_35),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_176),
.A2(n_138),
.B1(n_153),
.B2(n_147),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_190),
.A2(n_194),
.B1(n_199),
.B2(n_170),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_176),
.A2(n_150),
.B1(n_132),
.B2(n_144),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_195),
.A2(n_209),
.B(n_167),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_176),
.A2(n_154),
.B1(n_148),
.B2(n_137),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_161),
.A2(n_154),
.B1(n_156),
.B2(n_137),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_169),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_202),
.B(n_211),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_165),
.B(n_156),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_203),
.B(n_173),
.C(n_168),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_161),
.A2(n_146),
.B1(n_67),
.B2(n_152),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_207),
.A2(n_165),
.B(n_174),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_182),
.A2(n_152),
.B(n_18),
.Y(n_209)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_186),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_215),
.A2(n_225),
.B1(n_196),
.B2(n_202),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_217),
.A2(n_228),
.B(n_239),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_212),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_218),
.B(n_219),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_213),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_205),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_220),
.B(n_240),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_189),
.B(n_184),
.Y(n_221)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_221),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_222),
.A2(n_227),
.B(n_18),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_192),
.B(n_160),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_223),
.B(n_230),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_199),
.A2(n_185),
.B1(n_167),
.B2(n_159),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_189),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_226),
.B(n_229),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_195),
.A2(n_168),
.B(n_171),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_210),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_214),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_192),
.B(n_177),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_203),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_231),
.B(n_235),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_214),
.B(n_172),
.Y(n_232)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_232),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_233),
.B(n_237),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_198),
.B(n_166),
.C(n_178),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_234),
.B(n_187),
.C(n_209),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_197),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_204),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_236),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_198),
.B(n_201),
.Y(n_237)
);

OAI21xp33_ASAP7_75t_L g238 ( 
.A1(n_188),
.A2(n_11),
.B(n_15),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_238),
.B(n_191),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_204),
.B(n_142),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_200),
.Y(n_240)
);

AO21x1_ASAP7_75t_L g265 ( 
.A1(n_241),
.A2(n_25),
.B(n_1),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_242),
.B(n_217),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_224),
.A2(n_208),
.B1(n_190),
.B2(n_200),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_244),
.A2(n_248),
.B1(n_257),
.B2(n_220),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_245),
.B(n_251),
.C(n_255),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_223),
.B(n_206),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_246),
.B(n_264),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_224),
.A2(n_207),
.B1(n_211),
.B2(n_196),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_250),
.A2(n_216),
.B1(n_25),
.B2(n_2),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_230),
.B(n_193),
.C(n_143),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_237),
.B(n_193),
.C(n_143),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_233),
.B(n_152),
.C(n_67),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_258),
.B(n_260),
.C(n_234),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_222),
.A2(n_8),
.B(n_14),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_10),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_225),
.B(n_25),
.C(n_20),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_227),
.B(n_35),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_265),
.B(n_228),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_266),
.A2(n_284),
.B1(n_260),
.B2(n_265),
.Y(n_285)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_249),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_267),
.B(n_271),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_243),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_268),
.A2(n_245),
.B(n_258),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_SL g269 ( 
.A(n_250),
.B(n_215),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_269),
.B(n_283),
.Y(n_293)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_270),
.Y(n_290)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_261),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_263),
.B(n_226),
.Y(n_272)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_272),
.Y(n_291)
);

BUFx24_ASAP7_75t_SL g273 ( 
.A(n_262),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_273),
.B(n_276),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_274),
.B(n_246),
.Y(n_289)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_248),
.Y(n_276)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_277),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_252),
.B(n_221),
.Y(n_279)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_279),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_280),
.B(n_281),
.C(n_247),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_251),
.B(n_247),
.C(n_255),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_257),
.A2(n_231),
.B1(n_236),
.B2(n_241),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_282),
.B(n_8),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_256),
.A2(n_25),
.B1(n_1),
.B2(n_2),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_285),
.A2(n_292),
.B1(n_0),
.B2(n_1),
.Y(n_306)
);

AOI21x1_ASAP7_75t_SL g286 ( 
.A1(n_269),
.A2(n_244),
.B(n_253),
.Y(n_286)
);

OR2x2_ASAP7_75t_L g308 ( 
.A(n_286),
.B(n_6),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_287),
.A2(n_299),
.B(n_280),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_288),
.B(n_0),
.C(n_3),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_289),
.B(n_298),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_268),
.A2(n_264),
.B1(n_242),
.B2(n_254),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_278),
.B(n_254),
.Y(n_298)
);

AOI21xp33_ASAP7_75t_L g299 ( 
.A1(n_275),
.A2(n_7),
.B(n_12),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_300),
.B(n_10),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_301),
.B(n_311),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_291),
.B(n_290),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_302),
.A2(n_303),
.B(n_304),
.Y(n_324)
);

NOR2xp67_ASAP7_75t_SL g303 ( 
.A(n_286),
.B(n_275),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_287),
.A2(n_281),
.B(n_278),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_305),
.B(n_310),
.C(n_312),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_SL g321 ( 
.A(n_306),
.B(n_308),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_288),
.B(n_8),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_307),
.B(n_9),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_296),
.B(n_6),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_309),
.A2(n_313),
.B(n_9),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_285),
.A2(n_292),
.B1(n_297),
.B2(n_294),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_298),
.B(n_0),
.C(n_3),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_289),
.B(n_3),
.C(n_4),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_308),
.B(n_295),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_317),
.A2(n_321),
.B(n_316),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_307),
.B(n_293),
.Y(n_318)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_318),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_310),
.B(n_293),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_319),
.B(n_322),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_320),
.B(n_6),
.C(n_11),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_313),
.B(n_3),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_323),
.A2(n_312),
.B(n_5),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_315),
.B(n_314),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_326),
.B(n_328),
.Y(n_337)
);

OR2x2_ASAP7_75t_L g327 ( 
.A(n_324),
.B(n_314),
.Y(n_327)
);

NOR2xp67_ASAP7_75t_L g333 ( 
.A(n_327),
.B(n_317),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_330),
.B(n_331),
.Y(n_334)
);

OAI21x1_ASAP7_75t_SL g332 ( 
.A1(n_321),
.A2(n_12),
.B(n_14),
.Y(n_332)
);

OAI21xp33_ASAP7_75t_L g336 ( 
.A1(n_332),
.A2(n_12),
.B(n_14),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_333),
.B(n_335),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_330),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_336),
.Y(n_339)
);

AOI21x1_ASAP7_75t_L g340 ( 
.A1(n_338),
.A2(n_337),
.B(n_334),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_325),
.C(n_329),
.Y(n_341)
);

BUFx24_ASAP7_75t_SL g342 ( 
.A(n_341),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_342),
.A2(n_339),
.B(n_4),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_343),
.B(n_4),
.Y(n_344)
);


endmodule