module fake_netlist_6_1191_n_3364 (n_52, n_591, n_435, n_1, n_91, n_793, n_326, n_801, n_256, n_853, n_440, n_587, n_695, n_507, n_909, n_580, n_762, n_881, n_875, n_209, n_367, n_465, n_680, n_741, n_760, n_590, n_625, n_63, n_661, n_223, n_278, n_341, n_362, n_148, n_226, n_828, n_161, n_22, n_208, n_462, n_68, n_607, n_671, n_726, n_316, n_419, n_28, n_304, n_212, n_700, n_50, n_694, n_7, n_740, n_578, n_703, n_144, n_365, n_125, n_168, n_384, n_297, n_595, n_627, n_524, n_342, n_77, n_820, n_783, n_106, n_725, n_358, n_160, n_751, n_449, n_131, n_749, n_798, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_575, n_677, n_805, n_396, n_495, n_815, n_350, n_78, n_84, n_585, n_732, n_568, n_392, n_840, n_442, n_480, n_142, n_874, n_724, n_143, n_382, n_673, n_180, n_62, n_628, n_883, n_557, n_823, n_349, n_643, n_233, n_617, n_698, n_898, n_845, n_255, n_807, n_739, n_284, n_400, n_140, n_337, n_865, n_893, n_214, n_485, n_67, n_15, n_443, n_246, n_892, n_768, n_38, n_471, n_289, n_421, n_781, n_424, n_789, n_615, n_59, n_181, n_182, n_238, n_573, n_769, n_202, n_320, n_108, n_639, n_676, n_327, n_794, n_727, n_894, n_369, n_597, n_685, n_280, n_287, n_832, n_353, n_610, n_555, n_389, n_814, n_415, n_830, n_65, n_230, n_605, n_461, n_873, n_141, n_383, n_826, n_669, n_200, n_447, n_176, n_872, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_718, n_747, n_852, n_667, n_71, n_74, n_229, n_542, n_847, n_644, n_682, n_851, n_621, n_305, n_72, n_721, n_750, n_532, n_742, n_173, n_535, n_691, n_250, n_372, n_468, n_544, n_901, n_111, n_504, n_314, n_378, n_413, n_377, n_791, n_35, n_183, n_510, n_837, n_836, n_79, n_863, n_375, n_601, n_338, n_522, n_466, n_704, n_748, n_506, n_56, n_763, n_360, n_603, n_119, n_235, n_536, n_895, n_866, n_622, n_147, n_191, n_340, n_710, n_387, n_452, n_616, n_658, n_744, n_39, n_344, n_73, n_581, n_428, n_761, n_785, n_746, n_609, n_765, n_432, n_641, n_822, n_693, n_101, n_167, n_631, n_174, n_127, n_516, n_153, n_720, n_525, n_758, n_842, n_611, n_156, n_491, n_878, n_145, n_42, n_133, n_656, n_772, n_96, n_8, n_843, n_797, n_666, n_371, n_795, n_770, n_567, n_899, n_189, n_738, n_405, n_213, n_538, n_294, n_302, n_499, n_380, n_838, n_129, n_705, n_647, n_197, n_11, n_137, n_17, n_343, n_844, n_448, n_886, n_20, n_494, n_539, n_493, n_397, n_155, n_109, n_614, n_529, n_445, n_425, n_684, n_122, n_888, n_45, n_454, n_34, n_218, n_638, n_70, n_234, n_910, n_37, n_486, n_381, n_82, n_27, n_236, n_653, n_887, n_752, n_908, n_112, n_172, n_713, n_648, n_657, n_576, n_472, n_270, n_239, n_126, n_414, n_97, n_563, n_58, n_782, n_490, n_803, n_290, n_220, n_809, n_118, n_224, n_48, n_25, n_93, n_839, n_80, n_734, n_708, n_196, n_402, n_352, n_668, n_478, n_626, n_574, n_779, n_9, n_800, n_460, n_107, n_907, n_854, n_6, n_417, n_14, n_446, n_498, n_662, n_89, n_374, n_659, n_709, n_870, n_366, n_904, n_777, n_407, n_450, n_103, n_808, n_867, n_272, n_526, n_185, n_712, n_348, n_711, n_579, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_559, n_53, n_370, n_44, n_458, n_232, n_650, n_16, n_163, n_717, n_46, n_330, n_771, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_551, n_154, n_699, n_456, n_564, n_98, n_260, n_265, n_313, n_451, n_624, n_824, n_279, n_686, n_796, n_252, n_757, n_228, n_565, n_594, n_719, n_356, n_577, n_166, n_184, n_552, n_619, n_885, n_216, n_455, n_896, n_83, n_521, n_363, n_572, n_395, n_813, n_592, n_745, n_654, n_323, n_829, n_606, n_393, n_818, n_411, n_503, n_716, n_152, n_623, n_92, n_884, n_599, n_513, n_855, n_776, n_321, n_645, n_331, n_105, n_227, n_132, n_868, n_570, n_731, n_859, n_406, n_483, n_735, n_102, n_204, n_482, n_755, n_474, n_527, n_261, n_608, n_620, n_420, n_683, n_630, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_792, n_880, n_476, n_714, n_2, n_291, n_219, n_543, n_889, n_357, n_150, n_264, n_263, n_589, n_860, n_481, n_788, n_819, n_821, n_325, n_767, n_804, n_329, n_464, n_600, n_831, n_802, n_561, n_33, n_477, n_549, n_533, n_408, n_806, n_864, n_879, n_61, n_237, n_584, n_244, n_399, n_76, n_243, n_124, n_548, n_905, n_94, n_282, n_436, n_833, n_116, n_211, n_523, n_117, n_175, n_322, n_707, n_345, n_409, n_231, n_354, n_689, n_40, n_799, n_505, n_240, n_756, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_558, n_810, n_635, n_95, n_787, n_311, n_10, n_403, n_723, n_253, n_634, n_583, n_596, n_123, n_136, n_546, n_562, n_249, n_201, n_386, n_764, n_556, n_159, n_157, n_162, n_692, n_733, n_754, n_115, n_487, n_550, n_128, n_241, n_30, n_275, n_553, n_43, n_652, n_849, n_560, n_753, n_642, n_276, n_569, n_441, n_221, n_811, n_882, n_444, n_586, n_423, n_146, n_737, n_318, n_303, n_511, n_715, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_418, n_113, n_618, n_790, n_582, n_4, n_199, n_138, n_266, n_296, n_861, n_674, n_857, n_871, n_775, n_571, n_268, n_271, n_404, n_651, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_679, n_5, n_453, n_612, n_633, n_665, n_902, n_333, n_588, n_215, n_178, n_247, n_225, n_308, n_309, n_759, n_355, n_426, n_317, n_149, n_632, n_702, n_431, n_90, n_347, n_812, n_24, n_459, n_54, n_502, n_328, n_672, n_534, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_780, n_773, n_675, n_903, n_85, n_99, n_257, n_730, n_655, n_13, n_706, n_786, n_670, n_203, n_286, n_254, n_207, n_834, n_242, n_835, n_19, n_47, n_690, n_29, n_850, n_75, n_401, n_324, n_743, n_766, n_816, n_335, n_430, n_463, n_545, n_489, n_877, n_205, n_604, n_848, n_120, n_251, n_301, n_274, n_636, n_825, n_728, n_681, n_729, n_110, n_151, n_876, n_774, n_412, n_640, n_81, n_660, n_36, n_26, n_55, n_267, n_438, n_339, n_784, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_598, n_422, n_696, n_906, n_688, n_722, n_862, n_135, n_165, n_351, n_869, n_437, n_259, n_177, n_540, n_593, n_514, n_646, n_528, n_391, n_457, n_687, n_697, n_364, n_890, n_637, n_295, n_385, n_701, n_817, n_629, n_388, n_190, n_858, n_262, n_484, n_613, n_736, n_187, n_897, n_900, n_846, n_501, n_841, n_531, n_827, n_60, n_361, n_508, n_663, n_856, n_379, n_170, n_778, n_332, n_891, n_336, n_12, n_398, n_410, n_566, n_554, n_602, n_194, n_664, n_171, n_678, n_192, n_57, n_169, n_51, n_649, n_283, n_3364);

input n_52;
input n_591;
input n_435;
input n_1;
input n_91;
input n_793;
input n_326;
input n_801;
input n_256;
input n_853;
input n_440;
input n_587;
input n_695;
input n_507;
input n_909;
input n_580;
input n_762;
input n_881;
input n_875;
input n_209;
input n_367;
input n_465;
input n_680;
input n_741;
input n_760;
input n_590;
input n_625;
input n_63;
input n_661;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_828;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_607;
input n_671;
input n_726;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_700;
input n_50;
input n_694;
input n_7;
input n_740;
input n_578;
input n_703;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_595;
input n_627;
input n_524;
input n_342;
input n_77;
input n_820;
input n_783;
input n_106;
input n_725;
input n_358;
input n_160;
input n_751;
input n_449;
input n_131;
input n_749;
input n_798;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_575;
input n_677;
input n_805;
input n_396;
input n_495;
input n_815;
input n_350;
input n_78;
input n_84;
input n_585;
input n_732;
input n_568;
input n_392;
input n_840;
input n_442;
input n_480;
input n_142;
input n_874;
input n_724;
input n_143;
input n_382;
input n_673;
input n_180;
input n_62;
input n_628;
input n_883;
input n_557;
input n_823;
input n_349;
input n_643;
input n_233;
input n_617;
input n_698;
input n_898;
input n_845;
input n_255;
input n_807;
input n_739;
input n_284;
input n_400;
input n_140;
input n_337;
input n_865;
input n_893;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_892;
input n_768;
input n_38;
input n_471;
input n_289;
input n_421;
input n_781;
input n_424;
input n_789;
input n_615;
input n_59;
input n_181;
input n_182;
input n_238;
input n_573;
input n_769;
input n_202;
input n_320;
input n_108;
input n_639;
input n_676;
input n_327;
input n_794;
input n_727;
input n_894;
input n_369;
input n_597;
input n_685;
input n_280;
input n_287;
input n_832;
input n_353;
input n_610;
input n_555;
input n_389;
input n_814;
input n_415;
input n_830;
input n_65;
input n_230;
input n_605;
input n_461;
input n_873;
input n_141;
input n_383;
input n_826;
input n_669;
input n_200;
input n_447;
input n_176;
input n_872;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_718;
input n_747;
input n_852;
input n_667;
input n_71;
input n_74;
input n_229;
input n_542;
input n_847;
input n_644;
input n_682;
input n_851;
input n_621;
input n_305;
input n_72;
input n_721;
input n_750;
input n_532;
input n_742;
input n_173;
input n_535;
input n_691;
input n_250;
input n_372;
input n_468;
input n_544;
input n_901;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_791;
input n_35;
input n_183;
input n_510;
input n_837;
input n_836;
input n_79;
input n_863;
input n_375;
input n_601;
input n_338;
input n_522;
input n_466;
input n_704;
input n_748;
input n_506;
input n_56;
input n_763;
input n_360;
input n_603;
input n_119;
input n_235;
input n_536;
input n_895;
input n_866;
input n_622;
input n_147;
input n_191;
input n_340;
input n_710;
input n_387;
input n_452;
input n_616;
input n_658;
input n_744;
input n_39;
input n_344;
input n_73;
input n_581;
input n_428;
input n_761;
input n_785;
input n_746;
input n_609;
input n_765;
input n_432;
input n_641;
input n_822;
input n_693;
input n_101;
input n_167;
input n_631;
input n_174;
input n_127;
input n_516;
input n_153;
input n_720;
input n_525;
input n_758;
input n_842;
input n_611;
input n_156;
input n_491;
input n_878;
input n_145;
input n_42;
input n_133;
input n_656;
input n_772;
input n_96;
input n_8;
input n_843;
input n_797;
input n_666;
input n_371;
input n_795;
input n_770;
input n_567;
input n_899;
input n_189;
input n_738;
input n_405;
input n_213;
input n_538;
input n_294;
input n_302;
input n_499;
input n_380;
input n_838;
input n_129;
input n_705;
input n_647;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_844;
input n_448;
input n_886;
input n_20;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_109;
input n_614;
input n_529;
input n_445;
input n_425;
input n_684;
input n_122;
input n_888;
input n_45;
input n_454;
input n_34;
input n_218;
input n_638;
input n_70;
input n_234;
input n_910;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_653;
input n_887;
input n_752;
input n_908;
input n_112;
input n_172;
input n_713;
input n_648;
input n_657;
input n_576;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_563;
input n_58;
input n_782;
input n_490;
input n_803;
input n_290;
input n_220;
input n_809;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_839;
input n_80;
input n_734;
input n_708;
input n_196;
input n_402;
input n_352;
input n_668;
input n_478;
input n_626;
input n_574;
input n_779;
input n_9;
input n_800;
input n_460;
input n_107;
input n_907;
input n_854;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_662;
input n_89;
input n_374;
input n_659;
input n_709;
input n_870;
input n_366;
input n_904;
input n_777;
input n_407;
input n_450;
input n_103;
input n_808;
input n_867;
input n_272;
input n_526;
input n_185;
input n_712;
input n_348;
input n_711;
input n_579;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_559;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_650;
input n_16;
input n_163;
input n_717;
input n_46;
input n_330;
input n_771;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_551;
input n_154;
input n_699;
input n_456;
input n_564;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_624;
input n_824;
input n_279;
input n_686;
input n_796;
input n_252;
input n_757;
input n_228;
input n_565;
input n_594;
input n_719;
input n_356;
input n_577;
input n_166;
input n_184;
input n_552;
input n_619;
input n_885;
input n_216;
input n_455;
input n_896;
input n_83;
input n_521;
input n_363;
input n_572;
input n_395;
input n_813;
input n_592;
input n_745;
input n_654;
input n_323;
input n_829;
input n_606;
input n_393;
input n_818;
input n_411;
input n_503;
input n_716;
input n_152;
input n_623;
input n_92;
input n_884;
input n_599;
input n_513;
input n_855;
input n_776;
input n_321;
input n_645;
input n_331;
input n_105;
input n_227;
input n_132;
input n_868;
input n_570;
input n_731;
input n_859;
input n_406;
input n_483;
input n_735;
input n_102;
input n_204;
input n_482;
input n_755;
input n_474;
input n_527;
input n_261;
input n_608;
input n_620;
input n_420;
input n_683;
input n_630;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_792;
input n_880;
input n_476;
input n_714;
input n_2;
input n_291;
input n_219;
input n_543;
input n_889;
input n_357;
input n_150;
input n_264;
input n_263;
input n_589;
input n_860;
input n_481;
input n_788;
input n_819;
input n_821;
input n_325;
input n_767;
input n_804;
input n_329;
input n_464;
input n_600;
input n_831;
input n_802;
input n_561;
input n_33;
input n_477;
input n_549;
input n_533;
input n_408;
input n_806;
input n_864;
input n_879;
input n_61;
input n_237;
input n_584;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_548;
input n_905;
input n_94;
input n_282;
input n_436;
input n_833;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_707;
input n_345;
input n_409;
input n_231;
input n_354;
input n_689;
input n_40;
input n_799;
input n_505;
input n_240;
input n_756;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_558;
input n_810;
input n_635;
input n_95;
input n_787;
input n_311;
input n_10;
input n_403;
input n_723;
input n_253;
input n_634;
input n_583;
input n_596;
input n_123;
input n_136;
input n_546;
input n_562;
input n_249;
input n_201;
input n_386;
input n_764;
input n_556;
input n_159;
input n_157;
input n_162;
input n_692;
input n_733;
input n_754;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_30;
input n_275;
input n_553;
input n_43;
input n_652;
input n_849;
input n_560;
input n_753;
input n_642;
input n_276;
input n_569;
input n_441;
input n_221;
input n_811;
input n_882;
input n_444;
input n_586;
input n_423;
input n_146;
input n_737;
input n_318;
input n_303;
input n_511;
input n_715;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_418;
input n_113;
input n_618;
input n_790;
input n_582;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_861;
input n_674;
input n_857;
input n_871;
input n_775;
input n_571;
input n_268;
input n_271;
input n_404;
input n_651;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_679;
input n_5;
input n_453;
input n_612;
input n_633;
input n_665;
input n_902;
input n_333;
input n_588;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_759;
input n_355;
input n_426;
input n_317;
input n_149;
input n_632;
input n_702;
input n_431;
input n_90;
input n_347;
input n_812;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_672;
input n_534;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_780;
input n_773;
input n_675;
input n_903;
input n_85;
input n_99;
input n_257;
input n_730;
input n_655;
input n_13;
input n_706;
input n_786;
input n_670;
input n_203;
input n_286;
input n_254;
input n_207;
input n_834;
input n_242;
input n_835;
input n_19;
input n_47;
input n_690;
input n_29;
input n_850;
input n_75;
input n_401;
input n_324;
input n_743;
input n_766;
input n_816;
input n_335;
input n_430;
input n_463;
input n_545;
input n_489;
input n_877;
input n_205;
input n_604;
input n_848;
input n_120;
input n_251;
input n_301;
input n_274;
input n_636;
input n_825;
input n_728;
input n_681;
input n_729;
input n_110;
input n_151;
input n_876;
input n_774;
input n_412;
input n_640;
input n_81;
input n_660;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_784;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_598;
input n_422;
input n_696;
input n_906;
input n_688;
input n_722;
input n_862;
input n_135;
input n_165;
input n_351;
input n_869;
input n_437;
input n_259;
input n_177;
input n_540;
input n_593;
input n_514;
input n_646;
input n_528;
input n_391;
input n_457;
input n_687;
input n_697;
input n_364;
input n_890;
input n_637;
input n_295;
input n_385;
input n_701;
input n_817;
input n_629;
input n_388;
input n_190;
input n_858;
input n_262;
input n_484;
input n_613;
input n_736;
input n_187;
input n_897;
input n_900;
input n_846;
input n_501;
input n_841;
input n_531;
input n_827;
input n_60;
input n_361;
input n_508;
input n_663;
input n_856;
input n_379;
input n_170;
input n_778;
input n_332;
input n_891;
input n_336;
input n_12;
input n_398;
input n_410;
input n_566;
input n_554;
input n_602;
input n_194;
input n_664;
input n_171;
input n_678;
input n_192;
input n_57;
input n_169;
input n_51;
input n_649;
input n_283;

output n_3364;

wire n_992;
wire n_2542;
wire n_1671;
wire n_2817;
wire n_1613;
wire n_1458;
wire n_1234;
wire n_2576;
wire n_3254;
wire n_1199;
wire n_1674;
wire n_1027;
wire n_1351;
wire n_3266;
wire n_1189;
wire n_3152;
wire n_1212;
wire n_2157;
wire n_3335;
wire n_2332;
wire n_1307;
wire n_3178;
wire n_2003;
wire n_1038;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_2534;
wire n_3089;
wire n_3301;
wire n_1357;
wire n_1853;
wire n_2451;
wire n_1738;
wire n_2243;
wire n_1575;
wire n_1854;
wire n_2324;
wire n_3088;
wire n_1923;
wire n_3257;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_3222;
wire n_1708;
wire n_1151;
wire n_2977;
wire n_1739;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_2847;
wire n_1402;
wire n_2557;
wire n_1691;
wire n_1688;
wire n_3332;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_2405;
wire n_1160;
wire n_2647;
wire n_1238;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_2997;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_2521;
wire n_3046;
wire n_2956;
wire n_1553;
wire n_1099;
wire n_2491;
wire n_1264;
wire n_1192;
wire n_1844;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_2382;
wire n_2672;
wire n_3030;
wire n_2291;
wire n_2299;
wire n_3340;
wire n_1371;
wire n_1285;
wire n_2886;
wire n_2974;
wire n_1985;
wire n_2989;
wire n_2838;
wire n_2184;
wire n_2982;
wire n_1803;
wire n_1172;
wire n_2509;
wire n_2513;
wire n_3282;
wire n_1590;
wire n_2645;
wire n_1532;
wire n_2313;
wire n_2628;
wire n_3071;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_2926;
wire n_1704;
wire n_1078;
wire n_1711;
wire n_2247;
wire n_3106;
wire n_1140;
wire n_2630;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_3275;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_3031;
wire n_3345;
wire n_2074;
wire n_2447;
wire n_2919;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_3080;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_1874;
wire n_3165;
wire n_1119;
wire n_2865;
wire n_2825;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_2510;
wire n_1541;
wire n_1300;
wire n_2480;
wire n_2739;
wire n_3023;
wire n_3232;
wire n_1313;
wire n_2791;
wire n_3251;
wire n_1056;
wire n_3316;
wire n_2212;
wire n_3048;
wire n_1455;
wire n_2418;
wire n_2864;
wire n_1163;
wire n_2729;
wire n_3063;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_943;
wire n_1798;
wire n_1550;
wire n_2703;
wire n_2786;
wire n_1591;
wire n_3122;
wire n_2806;
wire n_1344;
wire n_3261;
wire n_2730;
wire n_2495;
wire n_940;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_2603;
wire n_2660;
wire n_3028;
wire n_2981;
wire n_3076;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_1471;
wire n_953;
wire n_1094;
wire n_3077;
wire n_1345;
wire n_1820;
wire n_2873;
wire n_3107;
wire n_2880;
wire n_3225;
wire n_2394;
wire n_2108;
wire n_1421;
wire n_2836;
wire n_1936;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_2378;
wire n_1660;
wire n_1961;
wire n_3047;
wire n_1280;
wire n_2655;
wire n_1400;
wire n_2625;
wire n_3296;
wire n_2843;
wire n_1467;
wire n_3297;
wire n_976;
wire n_3067;
wire n_2155;
wire n_2686;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1526;
wire n_1560;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_2996;
wire n_2599;
wire n_2985;
wire n_1978;
wire n_2085;
wire n_917;
wire n_3347;
wire n_2370;
wire n_2612;
wire n_1446;
wire n_2591;
wire n_1815;
wire n_2214;
wire n_3351;
wire n_913;
wire n_1658;
wire n_2593;
wire n_3269;
wire n_1230;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_2613;
wire n_1333;
wire n_2496;
wire n_2708;
wire n_3313;
wire n_1648;
wire n_3189;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2725;
wire n_2277;
wire n_3164;
wire n_1558;
wire n_1732;
wire n_2300;
wire n_1986;
wire n_2397;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_2907;
wire n_2735;
wire n_1843;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_2778;
wire n_2850;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_1441;
wire n_1309;
wire n_1123;
wire n_2104;
wire n_1381;
wire n_2961;
wire n_1699;
wire n_916;
wire n_2093;
wire n_2633;
wire n_2207;
wire n_1970;
wire n_2770;
wire n_2101;
wire n_2696;
wire n_2059;
wire n_2198;
wire n_3319;
wire n_2669;
wire n_2925;
wire n_2073;
wire n_2273;
wire n_2546;
wire n_3272;
wire n_3193;
wire n_2522;
wire n_2792;
wire n_1328;
wire n_1957;
wire n_2917;
wire n_2616;
wire n_3118;
wire n_3315;
wire n_1907;
wire n_2529;
wire n_1162;
wire n_1530;
wire n_939;
wire n_1543;
wire n_2811;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_982;
wire n_2674;
wire n_2832;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_932;
wire n_2831;
wire n_2998;
wire n_3317;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_1873;
wire n_1866;
wire n_1680;
wire n_993;
wire n_2692;
wire n_3248;
wire n_2031;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_2941;
wire n_1278;
wire n_2455;
wire n_2876;
wire n_2654;
wire n_3036;
wire n_2469;
wire n_1064;
wire n_3099;
wire n_1396;
wire n_2355;
wire n_966;
wire n_2908;
wire n_3168;
wire n_2751;
wire n_2764;
wire n_3357;
wire n_1663;
wire n_2895;
wire n_2009;
wire n_1793;
wire n_2922;
wire n_1233;
wire n_1289;
wire n_2714;
wire n_2245;
wire n_3055;
wire n_3092;
wire n_2068;
wire n_1107;
wire n_2866;
wire n_2457;
wire n_3294;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_2821;
wire n_1875;
wire n_1865;
wire n_2459;
wire n_1701;
wire n_1111;
wire n_1713;
wire n_2971;
wire n_2678;
wire n_1251;
wire n_1265;
wire n_2711;
wire n_1726;
wire n_1950;
wire n_1563;
wire n_1912;
wire n_2434;
wire n_1982;
wire n_2878;
wire n_3012;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_2818;
wire n_2428;
wire n_3247;
wire n_3069;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_2664;
wire n_1664;
wire n_1722;
wire n_2641;
wire n_3022;
wire n_3052;
wire n_1165;
wire n_2749;
wire n_2008;
wire n_3298;
wire n_2192;
wire n_3281;
wire n_2254;
wire n_2345;
wire n_3346;
wire n_1926;
wire n_1175;
wire n_3273;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_2965;
wire n_1747;
wire n_3058;
wire n_1012;
wire n_2624;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2350;
wire n_2804;
wire n_2453;
wire n_2193;
wire n_2676;
wire n_1655;
wire n_928;
wire n_1214;
wire n_1801;
wire n_2347;
wire n_1886;
wire n_2092;
wire n_1654;
wire n_1157;
wire n_1750;
wire n_2994;
wire n_1462;
wire n_3153;
wire n_1188;
wire n_1752;
wire n_1813;
wire n_2514;
wire n_2206;
wire n_2810;
wire n_2967;
wire n_2319;
wire n_2519;
wire n_2916;
wire n_1063;
wire n_1588;
wire n_2963;
wire n_2947;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_3145;
wire n_1624;
wire n_1124;
wire n_2096;
wire n_2980;
wire n_1965;
wire n_2476;
wire n_3280;
wire n_1515;
wire n_961;
wire n_1317;
wire n_1082;
wire n_3227;
wire n_2733;
wire n_2824;
wire n_3289;
wire n_2377;
wire n_3271;
wire n_2178;
wire n_950;
wire n_2812;
wire n_2644;
wire n_2036;
wire n_3326;
wire n_2976;
wire n_2152;
wire n_1709;
wire n_3009;
wire n_2652;
wire n_2411;
wire n_2525;
wire n_1825;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_2657;
wire n_1792;
wire n_2067;
wire n_2136;
wire n_2921;
wire n_2409;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_2687;
wire n_3237;
wire n_949;
wire n_1630;
wire n_2887;
wire n_2075;
wire n_2194;
wire n_2972;
wire n_2619;
wire n_3139;
wire n_2763;
wire n_2762;
wire n_1987;
wire n_968;
wire n_1369;
wire n_2271;
wire n_1008;
wire n_3192;
wire n_1546;
wire n_2583;
wire n_2606;
wire n_2279;
wire n_1033;
wire n_1052;
wire n_2794;
wire n_1296;
wire n_2663;
wire n_1990;
wire n_3352;
wire n_2391;
wire n_2431;
wire n_3073;
wire n_2987;
wire n_2938;
wire n_2150;
wire n_1294;
wire n_2943;
wire n_1420;
wire n_2078;
wire n_1634;
wire n_3252;
wire n_2932;
wire n_1767;
wire n_1779;
wire n_1465;
wire n_3253;
wire n_3337;
wire n_3209;
wire n_2622;
wire n_1858;
wire n_1044;
wire n_2658;
wire n_2665;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_3021;
wire n_1391;
wire n_1523;
wire n_2558;
wire n_2893;
wire n_2775;
wire n_1208;
wire n_2750;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2954;
wire n_2728;
wire n_2349;
wire n_3128;
wire n_2684;
wire n_2712;
wire n_1072;
wire n_3146;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_1100;
wire n_1487;
wire n_2691;
wire n_2913;
wire n_1756;
wire n_3183;
wire n_1128;
wire n_2493;
wire n_2230;
wire n_2705;
wire n_1969;
wire n_2690;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_1952;
wire n_2573;
wire n_2646;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_2535;
wire n_2631;
wire n_1364;
wire n_3078;
wire n_2436;
wire n_2870;
wire n_1249;
wire n_2706;
wire n_1293;
wire n_2693;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_3159;
wire n_1451;
wire n_963;
wire n_2767;
wire n_1839;
wire n_2341;
wire n_1765;
wire n_2707;
wire n_3240;
wire n_1514;
wire n_1863;
wire n_3037;
wire n_1646;
wire n_3293;
wire n_1714;
wire n_1139;
wire n_3179;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_2537;
wire n_2897;
wire n_2554;
wire n_996;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_2747;
wire n_3171;
wire n_1913;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_2853;
wire n_1808;
wire n_3053;
wire n_948;
wire n_3358;
wire n_2517;
wire n_2713;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_2765;
wire n_2861;
wire n_3158;
wire n_1788;
wire n_1999;
wire n_2731;
wire n_2643;
wire n_2590;
wire n_3150;
wire n_3018;
wire n_3353;
wire n_1469;
wire n_2060;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_3133;
wire n_2002;
wire n_2650;
wire n_2138;
wire n_1492;
wire n_987;
wire n_2414;
wire n_1340;
wire n_3014;
wire n_3166;
wire n_1771;
wire n_2316;
wire n_3104;
wire n_3148;
wire n_2262;
wire n_3229;
wire n_3348;
wire n_1707;
wire n_2239;
wire n_3082;
wire n_1432;
wire n_2208;
wire n_989;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_2689;
wire n_2933;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_2717;
wire n_1246;
wire n_1878;
wire n_2574;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_2842;
wire n_2675;
wire n_1426;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_2473;
wire n_1022;
wire n_2069;
wire n_2307;
wire n_2362;
wire n_2667;
wire n_2539;
wire n_2698;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_3312;
wire n_1571;
wire n_1809;
wire n_3119;
wire n_2948;
wire n_1577;
wire n_2958;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_947;
wire n_2936;
wire n_3224;
wire n_1117;
wire n_2489;
wire n_1087;
wire n_1448;
wire n_3173;
wire n_1992;
wire n_1049;
wire n_3223;
wire n_2771;
wire n_2445;
wire n_3020;
wire n_2057;
wire n_2103;
wire n_3140;
wire n_3185;
wire n_2605;
wire n_1666;
wire n_2772;
wire n_1505;
wire n_1717;
wire n_926;
wire n_1817;
wire n_2449;
wire n_927;
wire n_2610;
wire n_3129;
wire n_1849;
wire n_2848;
wire n_919;
wire n_2868;
wire n_1698;
wire n_2231;
wire n_929;
wire n_2520;
wire n_1228;
wire n_2857;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_1299;
wire n_2896;
wire n_2718;
wire n_3019;
wire n_2639;
wire n_1183;
wire n_1436;
wire n_2898;
wire n_2251;
wire n_1384;
wire n_2494;
wire n_2959;
wire n_2501;
wire n_3203;
wire n_3325;
wire n_2238;
wire n_2368;
wire n_1070;
wire n_2403;
wire n_3342;
wire n_2837;
wire n_998;
wire n_3200;
wire n_1665;
wire n_3259;
wire n_2524;
wire n_3167;
wire n_1383;
wire n_2460;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_2338;
wire n_3324;
wire n_3341;
wire n_1073;
wire n_1000;
wire n_1195;
wire n_3025;
wire n_2137;
wire n_1626;
wire n_3191;
wire n_1507;
wire n_2482;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_3006;
wire n_2481;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_3056;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_2424;
wire n_3201;
wire n_1142;
wire n_2849;
wire n_1475;
wire n_1774;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_2354;
wire n_2682;
wire n_3032;
wire n_3103;
wire n_2589;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_2661;
wire n_2877;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_931;
wire n_1021;
wire n_1207;
wire n_2442;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_1250;
wire n_958;
wire n_3331;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_3087;
wire n_3072;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_2773;
wire n_2545;
wire n_2432;
wire n_2710;
wire n_1478;
wire n_1310;
wire n_3142;
wire n_2966;
wire n_2294;
wire n_1363;
wire n_2581;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_1314;
wire n_964;
wire n_1837;
wire n_2218;
wire n_2788;
wire n_3196;
wire n_2435;
wire n_954;
wire n_2504;
wire n_2797;
wire n_2623;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2892;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_2748;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2860;
wire n_3327;
wire n_2330;
wire n_1457;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_2701;
wire n_2475;
wire n_2511;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_2416;
wire n_2745;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_1877;
wire n_3144;
wire n_3211;
wire n_3244;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_2784;
wire n_2209;
wire n_2301;
wire n_3287;
wire n_2387;
wire n_3322;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_3270;
wire n_2618;
wire n_2025;
wire n_2357;
wire n_2846;
wire n_2464;
wire n_3265;
wire n_1125;
wire n_970;
wire n_3306;
wire n_2488;
wire n_2224;
wire n_1980;
wire n_1159;
wire n_995;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_3026;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_3090;
wire n_3033;
wire n_1252;
wire n_1784;
wire n_3311;
wire n_1223;
wire n_2990;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_2115;
wire n_2410;
wire n_2552;
wire n_1053;
wire n_3302;
wire n_2374;
wire n_1681;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2929;
wire n_2780;
wire n_3226;
wire n_3323;
wire n_2596;
wire n_2274;
wire n_3163;
wire n_1153;
wire n_1618;
wire n_1531;
wire n_2828;
wire n_1185;
wire n_2384;
wire n_1745;
wire n_914;
wire n_3127;
wire n_2724;
wire n_1831;
wire n_2585;
wire n_2621;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2601;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_2502;
wire n_2801;
wire n_2920;
wire n_1901;
wire n_920;
wire n_1374;
wire n_2556;
wire n_2648;
wire n_3212;
wire n_1315;
wire n_1647;
wire n_2575;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_3188;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_2889;
wire n_3243;
wire n_1617;
wire n_3260;
wire n_1470;
wire n_2550;
wire n_3093;
wire n_3175;
wire n_3214;
wire n_1243;
wire n_2732;
wire n_2928;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_2822;
wire n_1425;
wire n_3169;
wire n_3205;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_3284;
wire n_983;
wire n_3109;
wire n_2023;
wire n_3354;
wire n_2572;
wire n_2204;
wire n_1520;
wire n_2720;
wire n_3126;
wire n_2159;
wire n_1390;
wire n_2289;
wire n_1077;
wire n_1733;
wire n_2315;
wire n_1419;
wire n_2863;
wire n_3299;
wire n_2955;
wire n_2995;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_3051;
wire n_1437;
wire n_3360;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2859;
wire n_2202;
wire n_2049;
wire n_1331;
wire n_2627;
wire n_956;
wire n_960;
wire n_2276;
wire n_3234;
wire n_2803;
wire n_2100;
wire n_3314;
wire n_2993;
wire n_1668;
wire n_2777;
wire n_1134;
wire n_3016;
wire n_3004;
wire n_3202;
wire n_2830;
wire n_2781;
wire n_3220;
wire n_1129;
wire n_2829;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_1869;
wire n_2911;
wire n_1764;
wire n_1429;
wire n_2826;
wire n_1610;
wire n_3084;
wire n_1889;
wire n_2379;
wire n_2016;
wire n_1905;
wire n_2343;
wire n_1593;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_2942;
wire n_1079;
wire n_2515;
wire n_1744;
wire n_2139;
wire n_2142;
wire n_1551;
wire n_2448;
wire n_1103;
wire n_2875;
wire n_2555;
wire n_3338;
wire n_2219;
wire n_1203;
wire n_2851;
wire n_2327;
wire n_951;
wire n_2201;
wire n_952;
wire n_999;
wire n_1254;
wire n_2841;
wire n_3349;
wire n_2420;
wire n_2984;
wire n_994;
wire n_2263;
wire n_3291;
wire n_2304;
wire n_1508;
wire n_2487;
wire n_974;
wire n_2983;
wire n_2240;
wire n_2656;
wire n_2278;
wire n_2538;
wire n_3276;
wire n_2597;
wire n_2375;
wire n_3113;
wire n_3194;
wire n_3250;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_2756;
wire n_1871;
wire n_2924;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_2884;
wire n_1549;
wire n_1510;
wire n_3120;
wire n_1468;
wire n_2855;
wire n_1859;
wire n_2102;
wire n_2563;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_1270;
wire n_2549;
wire n_1187;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2544;
wire n_2381;
wire n_2052;
wire n_1847;
wire n_2302;
wire n_1667;
wire n_1206;
wire n_3230;
wire n_1037;
wire n_1397;
wire n_3236;
wire n_1279;
wire n_1115;
wire n_1499;
wire n_2755;
wire n_3141;
wire n_923;
wire n_1409;
wire n_1841;
wire n_2637;
wire n_2823;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_3112;
wire n_2819;
wire n_3195;
wire n_2526;
wire n_3041;
wire n_2423;
wire n_1057;
wire n_3277;
wire n_3108;
wire n_2548;
wire n_991;
wire n_2785;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_2636;
wire n_3131;
wire n_2439;
wire n_1818;
wire n_1108;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_2088;
wire n_1611;
wire n_2740;
wire n_1601;
wire n_3011;
wire n_1960;
wire n_2694;
wire n_2061;
wire n_1686;
wire n_2757;
wire n_2337;
wire n_2401;
wire n_1356;
wire n_1589;
wire n_3042;
wire n_3213;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_2607;
wire n_1740;
wire n_2737;
wire n_1497;
wire n_2890;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_3228;
wire n_1320;
wire n_2716;
wire n_3249;
wire n_3081;
wire n_2452;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_3010;
wire n_2499;
wire n_3043;
wire n_1622;
wire n_1586;
wire n_2543;
wire n_2264;
wire n_1694;
wire n_1535;
wire n_3137;
wire n_2486;
wire n_3132;
wire n_2571;
wire n_3138;
wire n_1596;
wire n_3177;
wire n_1190;
wire n_1734;
wire n_3172;
wire n_2902;
wire n_3217;
wire n_1983;
wire n_1938;
wire n_2498;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_2472;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_3238;
wire n_2235;
wire n_2988;
wire n_3136;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_2894;
wire n_2790;
wire n_2037;
wire n_2808;
wire n_2298;
wire n_2326;
wire n_1539;
wire n_1043;
wire n_3040;
wire n_1797;
wire n_3279;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_1870;
wire n_2964;
wire n_1692;
wire n_1084;
wire n_1171;
wire n_2169;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_3262;
wire n_2904;
wire n_2244;
wire n_3013;
wire n_3356;
wire n_2586;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_1642;
wire n_1352;
wire n_2789;
wire n_3105;
wire n_3210;
wire n_2872;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2699;
wire n_2200;
wire n_3029;
wire n_1046;
wire n_2560;
wire n_1940;
wire n_1979;
wire n_2760;
wire n_2704;
wire n_3329;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_2738;
wire n_1405;
wire n_972;
wire n_2376;
wire n_1406;
wire n_2766;
wire n_1332;
wire n_2670;
wire n_2700;
wire n_962;
wire n_1041;
wire n_2346;
wire n_3134;
wire n_1569;
wire n_936;
wire n_3045;
wire n_3115;
wire n_1883;
wire n_1288;
wire n_3318;
wire n_1186;
wire n_1062;
wire n_3278;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2970;
wire n_2882;
wire n_3320;
wire n_2541;
wire n_2940;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_1823;
wire n_2479;
wire n_3050;
wire n_3350;
wire n_2782;
wire n_1974;
wire n_2673;
wire n_2456;
wire n_1720;
wire n_2527;
wire n_934;
wire n_1637;
wire n_2635;
wire n_3307;
wire n_1407;
wire n_1795;
wire n_2768;
wire n_2871;
wire n_2688;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_3003;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2753;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_3292;
wire n_1545;
wire n_2007;
wire n_3121;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_3184;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_1846;
wire n_3245;
wire n_3075;
wire n_2406;
wire n_2390;
wire n_959;
wire n_2310;
wire n_2506;
wire n_2141;
wire n_2562;
wire n_2642;
wire n_1343;
wire n_1522;
wire n_2734;
wire n_1782;
wire n_2383;
wire n_2626;
wire n_1676;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_1319;
wire n_2986;
wire n_1900;
wire n_3246;
wire n_1548;
wire n_3044;
wire n_2973;
wire n_1155;
wire n_2536;
wire n_2196;
wire n_2629;
wire n_1633;
wire n_2195;
wire n_3208;
wire n_2809;
wire n_3007;
wire n_2172;
wire n_2835;
wire n_1416;
wire n_1528;
wire n_2820;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_3355;
wire n_2454;
wire n_2114;
wire n_3074;
wire n_3174;
wire n_1086;
wire n_1066;
wire n_3102;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_2561;
wire n_3321;
wire n_2567;
wire n_2322;
wire n_2962;
wire n_2727;
wire n_2154;
wire n_2939;
wire n_1906;
wire n_1484;
wire n_2992;
wire n_3305;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_2533;
wire n_3157;
wire n_1758;
wire n_3221;
wire n_3267;
wire n_2283;
wire n_2869;
wire n_2422;
wire n_1925;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_2759;
wire n_2945;
wire n_3061;
wire n_2361;
wire n_1373;
wire n_1292;
wire n_2266;
wire n_2960;
wire n_3005;
wire n_2427;
wire n_3151;
wire n_1029;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_2611;
wire n_2901;
wire n_3258;
wire n_1706;
wire n_1498;
wire n_3143;
wire n_2653;
wire n_2417;
wire n_3000;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_2189;
wire n_2680;
wire n_2246;
wire n_1047;
wire n_3149;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_3156;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_2834;
wire n_3207;
wire n_2668;
wire n_2441;
wire n_1257;
wire n_3008;
wire n_1751;
wire n_2840;
wire n_3197;
wire n_3242;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_1045;
wire n_1650;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_1872;
wire n_3091;
wire n_2695;
wire n_3124;
wire n_1746;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1949;
wire n_2888;
wire n_2761;
wire n_2885;
wire n_2793;
wire n_2715;
wire n_2923;
wire n_1804;
wire n_2671;
wire n_1727;
wire n_2508;
wire n_1019;
wire n_2054;
wire n_2845;
wire n_1337;
wire n_3097;
wire n_2062;
wire n_2041;
wire n_2975;
wire n_1477;
wire n_1360;
wire n_2839;
wire n_1860;
wire n_2856;
wire n_1904;
wire n_2874;
wire n_1200;
wire n_2070;
wire n_2588;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2944;
wire n_2614;
wire n_2126;
wire n_1154;
wire n_3308;
wire n_1600;
wire n_1113;
wire n_2833;
wire n_2253;
wire n_2758;
wire n_2366;
wire n_1098;
wire n_2937;
wire n_1329;
wire n_2045;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_3300;
wire n_2978;
wire n_2066;
wire n_1476;
wire n_2516;
wire n_1001;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_2903;
wire n_2827;
wire n_1177;
wire n_3216;
wire n_1150;
wire n_3190;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_1023;
wire n_1882;
wire n_2951;
wire n_1076;
wire n_1118;
wire n_2949;
wire n_1807;
wire n_1007;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_1592;
wire n_1759;
wire n_2719;
wire n_1814;
wire n_1631;
wire n_1377;
wire n_1879;
wire n_1542;
wire n_2587;
wire n_3199;
wire n_2931;
wire n_3339;
wire n_1678;
wire n_2569;
wire n_2400;
wire n_1716;
wire n_1256;
wire n_1953;
wire n_933;
wire n_3343;
wire n_3303;
wire n_978;
wire n_2752;
wire n_3135;
wire n_1976;
wire n_2905;
wire n_1291;
wire n_1217;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_3160;
wire n_1065;
wire n_2796;
wire n_3255;
wire n_2507;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_2815;
wire n_1204;
wire n_3034;
wire n_1132;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_955;
wire n_1379;
wire n_2528;
wire n_2814;
wire n_2787;
wire n_1338;
wire n_1097;
wire n_2969;
wire n_2395;
wire n_935;
wire n_3027;
wire n_1554;
wire n_3231;
wire n_1130;
wire n_3083;
wire n_2979;
wire n_1810;
wire n_2953;
wire n_2380;
wire n_1120;
wire n_1583;
wire n_3049;
wire n_1730;
wire n_2295;
wire n_2746;
wire n_2946;
wire n_1643;
wire n_2020;
wire n_2500;
wire n_2269;
wire n_1729;
wire n_2290;
wire n_2048;
wire n_2005;
wire n_2565;
wire n_1389;
wire n_1105;
wire n_3117;
wire n_1461;
wire n_2076;
wire n_2736;
wire n_2883;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_2935;
wire n_3015;
wire n_2175;
wire n_2182;
wire n_2910;
wire n_1283;
wire n_2385;
wire n_918;
wire n_1848;
wire n_1114;
wire n_1785;
wire n_1147;
wire n_3268;
wire n_1754;
wire n_2149;
wire n_3057;
wire n_3154;
wire n_2396;
wire n_1506;
wire n_2584;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_1227;
wire n_2450;
wire n_2485;
wire n_2284;
wire n_2566;
wire n_2287;
wire n_971;
wire n_2702;
wire n_3241;
wire n_946;
wire n_2906;
wire n_1303;
wire n_2769;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_2438;
wire n_2914;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_2463;
wire n_3363;
wire n_2881;
wire n_1677;
wire n_1116;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_3064;
wire n_1780;
wire n_3100;
wire n_1689;
wire n_2180;
wire n_2858;
wire n_3062;
wire n_2679;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_1501;
wire n_1221;
wire n_3334;
wire n_1245;
wire n_3215;
wire n_3336;
wire n_2952;
wire n_1017;
wire n_3068;
wire n_2117;
wire n_2234;
wire n_2779;
wire n_2685;
wire n_1083;
wire n_1561;
wire n_2741;
wire n_3114;
wire n_930;
wire n_2275;
wire n_1112;
wire n_2465;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_1737;
wire n_2430;
wire n_1414;
wire n_2649;
wire n_2721;
wire n_944;
wire n_2034;
wire n_1028;
wire n_2106;
wire n_2862;
wire n_2265;
wire n_2615;
wire n_2683;
wire n_1922;
wire n_2032;
wire n_2744;
wire n_1011;
wire n_2474;
wire n_1566;
wire n_1215;
wire n_2444;
wire n_2437;
wire n_2743;
wire n_1973;
wire n_3181;
wire n_2267;
wire n_3035;
wire n_990;
wire n_1500;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_3204;
wire n_1104;
wire n_1058;
wire n_2312;
wire n_1122;
wire n_1253;
wire n_1266;
wire n_2242;
wire n_3362;
wire n_1509;
wire n_3328;
wire n_1693;
wire n_2934;
wire n_3290;
wire n_1109;
wire n_2222;
wire n_3256;
wire n_1276;
wire n_3176;
wire n_3309;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_2466;
wire n_2915;
wire n_2530;
wire n_1148;
wire n_2188;
wire n_2505;
wire n_1989;
wire n_1161;
wire n_2609;
wire n_1085;
wire n_2802;
wire n_2999;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_1584;
wire n_2425;
wire n_924;
wire n_1582;
wire n_2318;
wire n_3286;
wire n_2408;
wire n_1149;
wire n_3170;
wire n_1184;
wire n_2483;
wire n_2950;
wire n_1972;
wire n_3060;
wire n_3304;
wire n_2592;
wire n_1525;
wire n_3098;
wire n_2594;
wire n_2666;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_2564;
wire n_1816;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_1362;
wire n_1156;
wire n_3123;
wire n_984;
wire n_2600;
wire n_1829;
wire n_2035;
wire n_3024;
wire n_1450;
wire n_1638;
wire n_3038;
wire n_3086;
wire n_2033;
wire n_1789;
wire n_2531;
wire n_1770;
wire n_3285;
wire n_2523;
wire n_1218;
wire n_2413;
wire n_1482;
wire n_3361;
wire n_981;
wire n_1349;
wire n_1144;
wire n_2071;
wire n_3219;
wire n_2429;
wire n_3130;
wire n_985;
wire n_2233;
wire n_2440;
wire n_2723;
wire n_3233;
wire n_997;
wire n_1710;
wire n_2800;
wire n_2161;
wire n_1301;
wire n_2805;
wire n_3310;
wire n_980;
wire n_2681;
wire n_1306;
wire n_3264;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_3096;
wire n_2360;
wire n_2047;
wire n_2651;
wire n_2095;
wire n_3239;
wire n_1609;
wire n_2174;
wire n_3161;
wire n_2799;
wire n_3344;
wire n_2334;
wire n_3295;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_3066;
wire n_1574;
wire n_2426;
wire n_2490;
wire n_2844;
wire n_3101;
wire n_2478;
wire n_2303;
wire n_1619;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_1133;
wire n_1194;
wire n_2742;
wire n_2640;
wire n_1051;
wire n_1552;
wire n_2918;
wire n_3288;
wire n_1996;
wire n_2367;
wire n_2867;
wire n_3198;
wire n_1039;
wire n_1442;
wire n_2726;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_3125;
wire n_1158;
wire n_2909;
wire n_2248;
wire n_941;
wire n_975;
wire n_3206;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_2662;
wire n_3116;
wire n_3147;
wire n_1753;
wire n_3095;
wire n_3180;
wire n_3359;
wire n_2795;
wire n_2471;
wire n_3187;
wire n_2540;
wire n_973;
wire n_2807;
wire n_1921;
wire n_3218;
wire n_3330;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2217;
wire n_2197;
wire n_2065;
wire n_2879;
wire n_967;
wire n_2215;
wire n_2461;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_2968;
wire n_1629;
wire n_1170;
wire n_2221;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_2553;
wire n_1040;
wire n_915;
wire n_3059;
wire n_1166;
wire n_2038;
wire n_2891;
wire n_1131;
wire n_2634;
wire n_1761;
wire n_2709;
wire n_3155;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_3110;
wire n_1632;
wire n_1890;
wire n_3017;
wire n_1805;
wire n_2477;
wire n_1888;
wire n_1557;
wire n_2280;
wire n_1833;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2697;
wire n_3235;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_3001;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_2512;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_2927;
wire n_1836;
wire n_2774;
wire n_3039;
wire n_1226;
wire n_3162;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_3094;
wire n_2899;
wire n_3274;
wire n_3333;
wire n_3186;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_1059;
wire n_1197;
wire n_3065;
wire n_2632;
wire n_2579;
wire n_2105;
wire n_3079;
wire n_2098;
wire n_3085;
wire n_1423;
wire n_2813;
wire n_1935;
wire n_2027;
wire n_3070;
wire n_2223;
wire n_2091;
wire n_3263;
wire n_2991;
wire n_1915;
wire n_1621;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_1449;
wire n_2912;
wire n_2659;
wire n_2930;
wire n_1025;
wire n_2419;
wire n_3111;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_2677;
wire n_1013;
wire n_3182;
wire n_1259;
wire n_3054;
wire n_3283;
wire n_2183;
wire n_3002;
wire n_1538;
wire n_1742;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_296),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_837),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_509),
.Y(n_913)
);

BUFx3_ASAP7_75t_L g914 ( 
.A(n_276),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_727),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_561),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_501),
.Y(n_917)
);

BUFx5_ASAP7_75t_L g918 ( 
.A(n_66),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_783),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_111),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_1),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_651),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_91),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_885),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_440),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_821),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_592),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_774),
.Y(n_928)
);

CKINVDCx20_ASAP7_75t_R g929 ( 
.A(n_777),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_881),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_845),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_848),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_753),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_745),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_886),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_672),
.Y(n_936)
);

INVx1_ASAP7_75t_SL g937 ( 
.A(n_796),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_225),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_229),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_533),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_781),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_295),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_309),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_542),
.Y(n_944)
);

CKINVDCx20_ASAP7_75t_R g945 ( 
.A(n_849),
.Y(n_945)
);

CKINVDCx20_ASAP7_75t_R g946 ( 
.A(n_760),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_296),
.Y(n_947)
);

CKINVDCx20_ASAP7_75t_R g948 ( 
.A(n_571),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_235),
.Y(n_949)
);

BUFx2_ASAP7_75t_L g950 ( 
.A(n_518),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_109),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_673),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_830),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_812),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_56),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_688),
.Y(n_956)
);

CKINVDCx20_ASAP7_75t_R g957 ( 
.A(n_200),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_522),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_453),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_879),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_160),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_290),
.Y(n_962)
);

BUFx2_ASAP7_75t_L g963 ( 
.A(n_459),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_201),
.Y(n_964)
);

CKINVDCx16_ASAP7_75t_R g965 ( 
.A(n_836),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_481),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_482),
.Y(n_967)
);

BUFx10_ASAP7_75t_L g968 ( 
.A(n_221),
.Y(n_968)
);

CKINVDCx20_ASAP7_75t_R g969 ( 
.A(n_880),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_530),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_444),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_785),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_811),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_632),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_64),
.Y(n_975)
);

CKINVDCx16_ASAP7_75t_R g976 ( 
.A(n_697),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_445),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_717),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_536),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_658),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_852),
.Y(n_981)
);

BUFx10_ASAP7_75t_L g982 ( 
.A(n_788),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_778),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_858),
.Y(n_984)
);

BUFx6f_ASAP7_75t_L g985 ( 
.A(n_121),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_383),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_477),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_546),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_701),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_270),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_99),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_424),
.Y(n_992)
);

INVx1_ASAP7_75t_SL g993 ( 
.A(n_68),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_823),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_251),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_868),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_360),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_817),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_589),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_298),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_457),
.Y(n_1001)
);

CKINVDCx14_ASAP7_75t_R g1002 ( 
.A(n_141),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_414),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_548),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_875),
.Y(n_1005)
);

CKINVDCx20_ASAP7_75t_R g1006 ( 
.A(n_767),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_841),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_862),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_310),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_606),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_138),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_69),
.Y(n_1012)
);

CKINVDCx20_ASAP7_75t_R g1013 ( 
.A(n_253),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_376),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_865),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_204),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_358),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_605),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_857),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_496),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_720),
.Y(n_1021)
);

CKINVDCx20_ASAP7_75t_R g1022 ( 
.A(n_504),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_854),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_310),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_631),
.Y(n_1025)
);

CKINVDCx16_ASAP7_75t_R g1026 ( 
.A(n_295),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_151),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_738),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_356),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_338),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_152),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_408),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_855),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_838),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_765),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_866),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_800),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_792),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_178),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_721),
.Y(n_1040)
);

BUFx3_ASAP7_75t_L g1041 ( 
.A(n_901),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_863),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_29),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_264),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_409),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_789),
.Y(n_1046)
);

CKINVDCx14_ASAP7_75t_R g1047 ( 
.A(n_703),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_103),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_56),
.Y(n_1049)
);

CKINVDCx20_ASAP7_75t_R g1050 ( 
.A(n_769),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_103),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_527),
.Y(n_1052)
);

BUFx2_ASAP7_75t_SL g1053 ( 
.A(n_452),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_877),
.Y(n_1054)
);

CKINVDCx20_ASAP7_75t_R g1055 ( 
.A(n_864),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_822),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_813),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_742),
.Y(n_1058)
);

BUFx3_ASAP7_75t_L g1059 ( 
.A(n_876),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_495),
.Y(n_1060)
);

CKINVDCx20_ASAP7_75t_R g1061 ( 
.A(n_24),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_331),
.Y(n_1062)
);

INVxp67_ASAP7_75t_L g1063 ( 
.A(n_775),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_867),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_195),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_768),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_790),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_366),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_488),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_544),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_805),
.Y(n_1071)
);

BUFx6f_ASAP7_75t_L g1072 ( 
.A(n_41),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_335),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_748),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_276),
.Y(n_1075)
);

BUFx10_ASAP7_75t_L g1076 ( 
.A(n_814),
.Y(n_1076)
);

BUFx6f_ASAP7_75t_L g1077 ( 
.A(n_588),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_871),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_60),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_893),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_861),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_583),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_595),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_844),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_516),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_464),
.Y(n_1086)
);

BUFx10_ASAP7_75t_L g1087 ( 
.A(n_184),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_828),
.Y(n_1088)
);

INVxp67_ASAP7_75t_L g1089 ( 
.A(n_773),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_640),
.Y(n_1090)
);

CKINVDCx20_ASAP7_75t_R g1091 ( 
.A(n_190),
.Y(n_1091)
);

BUFx2_ASAP7_75t_L g1092 ( 
.A(n_840),
.Y(n_1092)
);

CKINVDCx20_ASAP7_75t_R g1093 ( 
.A(n_856),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_456),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_98),
.Y(n_1095)
);

CKINVDCx20_ASAP7_75t_R g1096 ( 
.A(n_809),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_11),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_455),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_873),
.Y(n_1099)
);

CKINVDCx20_ASAP7_75t_R g1100 ( 
.A(n_806),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_882),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_299),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_349),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_794),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_33),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_490),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_535),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_354),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_897),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_468),
.Y(n_1110)
);

INVx1_ASAP7_75t_SL g1111 ( 
.A(n_870),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_782),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_416),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_793),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_776),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_802),
.Y(n_1116)
);

CKINVDCx16_ASAP7_75t_R g1117 ( 
.A(n_134),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_869),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_556),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_393),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_647),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_750),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_630),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_302),
.Y(n_1124)
);

CKINVDCx20_ASAP7_75t_R g1125 ( 
.A(n_612),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_59),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_287),
.Y(n_1127)
);

INVx1_ASAP7_75t_SL g1128 ( 
.A(n_514),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_396),
.Y(n_1129)
);

BUFx6f_ASAP7_75t_L g1130 ( 
.A(n_121),
.Y(n_1130)
);

INVx2_ASAP7_75t_SL g1131 ( 
.A(n_826),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_135),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_804),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_851),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_839),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_693),
.Y(n_1136)
);

BUFx3_ASAP7_75t_L g1137 ( 
.A(n_404),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_582),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_39),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_115),
.Y(n_1140)
);

CKINVDCx20_ASAP7_75t_R g1141 ( 
.A(n_172),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_480),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_872),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_307),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_76),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_158),
.Y(n_1146)
);

CKINVDCx14_ASAP7_75t_R g1147 ( 
.A(n_705),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_699),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_18),
.Y(n_1149)
);

BUFx6f_ASAP7_75t_L g1150 ( 
.A(n_379),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_14),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_334),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_832),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_569),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_874),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_61),
.Y(n_1156)
);

CKINVDCx20_ASAP7_75t_R g1157 ( 
.A(n_324),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_853),
.Y(n_1158)
);

CKINVDCx20_ASAP7_75t_R g1159 ( 
.A(n_364),
.Y(n_1159)
);

BUFx6f_ASAP7_75t_L g1160 ( 
.A(n_427),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_859),
.Y(n_1161)
);

BUFx3_ASAP7_75t_L g1162 ( 
.A(n_803),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_764),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_402),
.Y(n_1164)
);

CKINVDCx20_ASAP7_75t_R g1165 ( 
.A(n_824),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_559),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_75),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_512),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_674),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_169),
.Y(n_1170)
);

CKINVDCx14_ASAP7_75t_R g1171 ( 
.A(n_33),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_348),
.Y(n_1172)
);

CKINVDCx20_ASAP7_75t_R g1173 ( 
.A(n_317),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_277),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_338),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_529),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_390),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_377),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_829),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_160),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_831),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_644),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_391),
.Y(n_1183)
);

BUFx5_ASAP7_75t_L g1184 ( 
.A(n_786),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_67),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_787),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_791),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_807),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_463),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_810),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_691),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_611),
.Y(n_1192)
);

CKINVDCx16_ASAP7_75t_R g1193 ( 
.A(n_220),
.Y(n_1193)
);

CKINVDCx20_ASAP7_75t_R g1194 ( 
.A(n_114),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_454),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_352),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_423),
.Y(n_1197)
);

HB1xp67_ASAP7_75t_L g1198 ( 
.A(n_827),
.Y(n_1198)
);

BUFx6f_ASAP7_75t_L g1199 ( 
.A(n_835),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_32),
.Y(n_1200)
);

INVxp67_ASAP7_75t_L g1201 ( 
.A(n_446),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_119),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_627),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_225),
.Y(n_1204)
);

CKINVDCx20_ASAP7_75t_R g1205 ( 
.A(n_883),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_415),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_551),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_833),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_493),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_834),
.Y(n_1210)
);

INVx1_ASAP7_75t_SL g1211 ( 
.A(n_797),
.Y(n_1211)
);

CKINVDCx20_ASAP7_75t_R g1212 ( 
.A(n_256),
.Y(n_1212)
);

CKINVDCx20_ASAP7_75t_R g1213 ( 
.A(n_600),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_168),
.Y(n_1214)
);

CKINVDCx20_ASAP7_75t_R g1215 ( 
.A(n_405),
.Y(n_1215)
);

BUFx2_ASAP7_75t_L g1216 ( 
.A(n_431),
.Y(n_1216)
);

CKINVDCx20_ASAP7_75t_R g1217 ( 
.A(n_798),
.Y(n_1217)
);

INVx1_ASAP7_75t_SL g1218 ( 
.A(n_425),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_795),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_843),
.Y(n_1220)
);

CKINVDCx20_ASAP7_75t_R g1221 ( 
.A(n_780),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_825),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_200),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_648),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_348),
.Y(n_1225)
);

CKINVDCx20_ASAP7_75t_R g1226 ( 
.A(n_389),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_232),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_676),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_784),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_850),
.Y(n_1230)
);

BUFx5_ASAP7_75t_L g1231 ( 
.A(n_454),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_808),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_740),
.Y(n_1233)
);

CKINVDCx20_ASAP7_75t_R g1234 ( 
.A(n_92),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_10),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_178),
.Y(n_1236)
);

CKINVDCx20_ASAP7_75t_R g1237 ( 
.A(n_695),
.Y(n_1237)
);

CKINVDCx20_ASAP7_75t_R g1238 ( 
.A(n_446),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_120),
.Y(n_1239)
);

CKINVDCx20_ASAP7_75t_R g1240 ( 
.A(n_10),
.Y(n_1240)
);

INVx1_ASAP7_75t_SL g1241 ( 
.A(n_884),
.Y(n_1241)
);

CKINVDCx5p33_ASAP7_75t_R g1242 ( 
.A(n_842),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_510),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_878),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_903),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_219),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_448),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_173),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_97),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_646),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_78),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_847),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_152),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_801),
.Y(n_1254)
);

CKINVDCx20_ASAP7_75t_R g1255 ( 
.A(n_365),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_165),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_860),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_815),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_706),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_472),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_355),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_779),
.Y(n_1262)
);

INVxp67_ASAP7_75t_L g1263 ( 
.A(n_322),
.Y(n_1263)
);

CKINVDCx20_ASAP7_75t_R g1264 ( 
.A(n_237),
.Y(n_1264)
);

BUFx6f_ASAP7_75t_L g1265 ( 
.A(n_521),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_322),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_846),
.Y(n_1267)
);

INVx1_ASAP7_75t_SL g1268 ( 
.A(n_47),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_13),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_528),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_412),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_188),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_289),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_799),
.Y(n_1274)
);

INVx1_ASAP7_75t_SL g1275 ( 
.A(n_737),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_663),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_887),
.Y(n_1277)
);

CKINVDCx20_ASAP7_75t_R g1278 ( 
.A(n_694),
.Y(n_1278)
);

CKINVDCx5p33_ASAP7_75t_R g1279 ( 
.A(n_820),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_711),
.Y(n_1280)
);

HB1xp67_ASAP7_75t_L g1281 ( 
.A(n_378),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_315),
.Y(n_1282)
);

INVxp67_ASAP7_75t_SL g1283 ( 
.A(n_816),
.Y(n_1283)
);

CKINVDCx20_ASAP7_75t_R g1284 ( 
.A(n_818),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_623),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_44),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_29),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_819),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_918),
.Y(n_1289)
);

BUFx3_ASAP7_75t_L g1290 ( 
.A(n_982),
.Y(n_1290)
);

INVxp67_ASAP7_75t_SL g1291 ( 
.A(n_1198),
.Y(n_1291)
);

CKINVDCx20_ASAP7_75t_R g1292 ( 
.A(n_929),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_918),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_918),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_918),
.Y(n_1295)
);

CKINVDCx16_ASAP7_75t_R g1296 ( 
.A(n_1026),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_918),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1231),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1231),
.Y(n_1299)
);

BUFx6f_ASAP7_75t_L g1300 ( 
.A(n_985),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_912),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_913),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1231),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1231),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1231),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_985),
.Y(n_1306)
);

HB1xp67_ASAP7_75t_L g1307 ( 
.A(n_1117),
.Y(n_1307)
);

HB1xp67_ASAP7_75t_L g1308 ( 
.A(n_1193),
.Y(n_1308)
);

INVxp67_ASAP7_75t_L g1309 ( 
.A(n_1216),
.Y(n_1309)
);

BUFx3_ASAP7_75t_L g1310 ( 
.A(n_982),
.Y(n_1310)
);

INVxp67_ASAP7_75t_L g1311 ( 
.A(n_1281),
.Y(n_1311)
);

CKINVDCx20_ASAP7_75t_R g1312 ( 
.A(n_945),
.Y(n_1312)
);

NOR2xp67_ASAP7_75t_L g1313 ( 
.A(n_1201),
.B(n_0),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_985),
.Y(n_1314)
);

BUFx3_ASAP7_75t_L g1315 ( 
.A(n_1076),
.Y(n_1315)
);

BUFx3_ASAP7_75t_L g1316 ( 
.A(n_1076),
.Y(n_1316)
);

BUFx6f_ASAP7_75t_L g1317 ( 
.A(n_1072),
.Y(n_1317)
);

CKINVDCx16_ASAP7_75t_R g1318 ( 
.A(n_965),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1072),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1072),
.Y(n_1320)
);

INVxp67_ASAP7_75t_L g1321 ( 
.A(n_968),
.Y(n_1321)
);

INVxp33_ASAP7_75t_SL g1322 ( 
.A(n_911),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_916),
.Y(n_1323)
);

CKINVDCx20_ASAP7_75t_R g1324 ( 
.A(n_946),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1130),
.Y(n_1325)
);

INVxp67_ASAP7_75t_L g1326 ( 
.A(n_968),
.Y(n_1326)
);

INVxp33_ASAP7_75t_SL g1327 ( 
.A(n_920),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1130),
.Y(n_1328)
);

NOR2xp33_ASAP7_75t_L g1329 ( 
.A(n_950),
.B(n_963),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_922),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1130),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1150),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_924),
.Y(n_1333)
);

BUFx6f_ASAP7_75t_L g1334 ( 
.A(n_1150),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1150),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1160),
.Y(n_1336)
);

INVxp67_ASAP7_75t_L g1337 ( 
.A(n_1087),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1160),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1160),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_914),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1137),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_921),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_942),
.Y(n_1343)
);

HB1xp67_ASAP7_75t_L g1344 ( 
.A(n_923),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1184),
.Y(n_1345)
);

HB1xp67_ASAP7_75t_L g1346 ( 
.A(n_938),
.Y(n_1346)
);

INVxp33_ASAP7_75t_SL g1347 ( 
.A(n_939),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_947),
.Y(n_1348)
);

CKINVDCx16_ASAP7_75t_R g1349 ( 
.A(n_976),
.Y(n_1349)
);

INVxp67_ASAP7_75t_SL g1350 ( 
.A(n_1092),
.Y(n_1350)
);

CKINVDCx20_ASAP7_75t_R g1351 ( 
.A(n_948),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_949),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_959),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_964),
.Y(n_1354)
);

BUFx3_ASAP7_75t_L g1355 ( 
.A(n_1041),
.Y(n_1355)
);

CKINVDCx16_ASAP7_75t_R g1356 ( 
.A(n_1002),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_971),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_977),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1000),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1300),
.Y(n_1360)
);

OAI22xp5_ASAP7_75t_L g1361 ( 
.A1(n_1329),
.A2(n_1350),
.B1(n_1309),
.B2(n_1291),
.Y(n_1361)
);

NOR2xp33_ASAP7_75t_SL g1362 ( 
.A(n_1356),
.B(n_969),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1344),
.B(n_1047),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_1300),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1317),
.Y(n_1365)
);

INVx3_ASAP7_75t_L g1366 ( 
.A(n_1317),
.Y(n_1366)
);

HB1xp67_ASAP7_75t_L g1367 ( 
.A(n_1307),
.Y(n_1367)
);

BUFx6f_ASAP7_75t_L g1368 ( 
.A(n_1334),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1334),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1306),
.Y(n_1370)
);

INVx6_ASAP7_75t_L g1371 ( 
.A(n_1290),
.Y(n_1371)
);

OAI22xp5_ASAP7_75t_L g1372 ( 
.A1(n_1308),
.A2(n_1171),
.B1(n_1147),
.B2(n_1263),
.Y(n_1372)
);

INVx3_ASAP7_75t_L g1373 ( 
.A(n_1355),
.Y(n_1373)
);

AND2x4_ASAP7_75t_L g1374 ( 
.A(n_1310),
.B(n_1059),
.Y(n_1374)
);

OAI21x1_ASAP7_75t_L g1375 ( 
.A1(n_1345),
.A2(n_932),
.B(n_917),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1314),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1319),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1320),
.Y(n_1378)
);

BUFx6f_ASAP7_75t_L g1379 ( 
.A(n_1325),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1301),
.B(n_1131),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1302),
.B(n_1323),
.Y(n_1381)
);

OAI22x1_ASAP7_75t_L g1382 ( 
.A1(n_1321),
.A2(n_1218),
.B1(n_1268),
.B2(n_993),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1330),
.B(n_1333),
.Y(n_1383)
);

CKINVDCx16_ASAP7_75t_R g1384 ( 
.A(n_1296),
.Y(n_1384)
);

HB1xp67_ASAP7_75t_L g1385 ( 
.A(n_1315),
.Y(n_1385)
);

AOI22xp5_ASAP7_75t_L g1386 ( 
.A1(n_1318),
.A2(n_1349),
.B1(n_1311),
.B2(n_1327),
.Y(n_1386)
);

BUFx6f_ASAP7_75t_L g1387 ( 
.A(n_1328),
.Y(n_1387)
);

BUFx6f_ASAP7_75t_L g1388 ( 
.A(n_1331),
.Y(n_1388)
);

INVx2_ASAP7_75t_SL g1389 ( 
.A(n_1316),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1332),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1335),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1336),
.Y(n_1392)
);

BUFx2_ASAP7_75t_L g1393 ( 
.A(n_1326),
.Y(n_1393)
);

AOI22xp5_ASAP7_75t_L g1394 ( 
.A1(n_1322),
.A2(n_1347),
.B1(n_1337),
.B2(n_1346),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1338),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1340),
.B(n_1162),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1339),
.Y(n_1397)
);

NOR2xp33_ASAP7_75t_L g1398 ( 
.A(n_1341),
.B(n_937),
.Y(n_1398)
);

INVx2_ASAP7_75t_SL g1399 ( 
.A(n_1342),
.Y(n_1399)
);

HB1xp67_ASAP7_75t_L g1400 ( 
.A(n_1343),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1289),
.B(n_940),
.Y(n_1401)
);

INVx4_ASAP7_75t_L g1402 ( 
.A(n_1293),
.Y(n_1402)
);

BUFx3_ASAP7_75t_L g1403 ( 
.A(n_1294),
.Y(n_1403)
);

INVx6_ASAP7_75t_L g1404 ( 
.A(n_1348),
.Y(n_1404)
);

BUFx6f_ASAP7_75t_L g1405 ( 
.A(n_1352),
.Y(n_1405)
);

BUFx6f_ASAP7_75t_L g1406 ( 
.A(n_1353),
.Y(n_1406)
);

AND2x4_ASAP7_75t_L g1407 ( 
.A(n_1354),
.B(n_1063),
.Y(n_1407)
);

INVx6_ASAP7_75t_L g1408 ( 
.A(n_1357),
.Y(n_1408)
);

BUFx6f_ASAP7_75t_L g1409 ( 
.A(n_1358),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1295),
.B(n_1297),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1298),
.Y(n_1411)
);

BUFx6f_ASAP7_75t_L g1412 ( 
.A(n_1359),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1299),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1409),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1412),
.Y(n_1415)
);

NAND2xp33_ASAP7_75t_R g1416 ( 
.A(n_1393),
.B(n_1374),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1402),
.B(n_1403),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1376),
.Y(n_1418)
);

NOR2xp33_ASAP7_75t_SL g1419 ( 
.A(n_1384),
.B(n_1362),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1411),
.Y(n_1420)
);

BUFx6f_ASAP7_75t_L g1421 ( 
.A(n_1368),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1377),
.Y(n_1422)
);

INVx3_ASAP7_75t_L g1423 ( 
.A(n_1366),
.Y(n_1423)
);

OAI22xp5_ASAP7_75t_L g1424 ( 
.A1(n_1381),
.A2(n_1313),
.B1(n_1022),
.B2(n_1050),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1413),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1405),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1395),
.Y(n_1427)
);

AND2x4_ASAP7_75t_L g1428 ( 
.A(n_1373),
.B(n_1006),
.Y(n_1428)
);

INVx1_ASAP7_75t_SL g1429 ( 
.A(n_1371),
.Y(n_1429)
);

BUFx6f_ASAP7_75t_L g1430 ( 
.A(n_1405),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1406),
.Y(n_1431)
);

HB1xp67_ASAP7_75t_L g1432 ( 
.A(n_1367),
.Y(n_1432)
);

AOI22xp5_ASAP7_75t_L g1433 ( 
.A1(n_1361),
.A2(n_1093),
.B1(n_1096),
.B2(n_1055),
.Y(n_1433)
);

NAND2x1_ASAP7_75t_L g1434 ( 
.A(n_1410),
.B(n_1077),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1406),
.Y(n_1435)
);

INVx1_ASAP7_75t_SL g1436 ( 
.A(n_1385),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1380),
.B(n_1363),
.Y(n_1437)
);

INVxp67_ASAP7_75t_L g1438 ( 
.A(n_1398),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1404),
.Y(n_1439)
);

OA21x2_ASAP7_75t_L g1440 ( 
.A1(n_1375),
.A2(n_1304),
.B(n_1303),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1408),
.Y(n_1441)
);

BUFx6f_ASAP7_75t_L g1442 ( 
.A(n_1379),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1383),
.B(n_1305),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1397),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_1360),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1400),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1399),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1370),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1389),
.B(n_1087),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1378),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1390),
.Y(n_1451)
);

BUFx6f_ASAP7_75t_L g1452 ( 
.A(n_1387),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1391),
.Y(n_1453)
);

BUFx6f_ASAP7_75t_L g1454 ( 
.A(n_1388),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1394),
.B(n_1292),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1392),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1364),
.Y(n_1457)
);

AOI22xp5_ASAP7_75t_L g1458 ( 
.A1(n_1372),
.A2(n_1125),
.B1(n_1165),
.B2(n_1100),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1401),
.B(n_1111),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1369),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1407),
.B(n_1312),
.Y(n_1461)
);

OAI22xp5_ASAP7_75t_SL g1462 ( 
.A1(n_1386),
.A2(n_1013),
.B1(n_1061),
.B2(n_957),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1396),
.B(n_1324),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1365),
.Y(n_1464)
);

BUFx6f_ASAP7_75t_L g1465 ( 
.A(n_1382),
.Y(n_1465)
);

NOR2xp33_ASAP7_75t_SL g1466 ( 
.A(n_1384),
.B(n_1205),
.Y(n_1466)
);

INVx3_ASAP7_75t_L g1467 ( 
.A(n_1368),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_SL g1468 ( 
.A(n_1363),
.B(n_1213),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1376),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1376),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1409),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1402),
.B(n_1128),
.Y(n_1472)
);

BUFx6f_ASAP7_75t_L g1473 ( 
.A(n_1368),
.Y(n_1473)
);

AOI22xp5_ASAP7_75t_L g1474 ( 
.A1(n_1361),
.A2(n_1217),
.B1(n_1237),
.B2(n_1221),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1376),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1376),
.Y(n_1476)
);

INVx1_ASAP7_75t_SL g1477 ( 
.A(n_1393),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1409),
.Y(n_1478)
);

INVxp67_ASAP7_75t_L g1479 ( 
.A(n_1393),
.Y(n_1479)
);

HB1xp67_ASAP7_75t_L g1480 ( 
.A(n_1373),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1376),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1409),
.Y(n_1482)
);

XOR2xp5_ASAP7_75t_L g1483 ( 
.A(n_1384),
.B(n_1351),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1409),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1376),
.Y(n_1485)
);

INVxp67_ASAP7_75t_L g1486 ( 
.A(n_1393),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1409),
.Y(n_1487)
);

INVx3_ASAP7_75t_L g1488 ( 
.A(n_1368),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1448),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1418),
.Y(n_1490)
);

INVxp67_ASAP7_75t_SL g1491 ( 
.A(n_1430),
.Y(n_1491)
);

BUFx3_ASAP7_75t_L g1492 ( 
.A(n_1430),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1438),
.B(n_1091),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1450),
.Y(n_1494)
);

AOI22xp5_ASAP7_75t_L g1495 ( 
.A1(n_1437),
.A2(n_1284),
.B1(n_1278),
.B2(n_1283),
.Y(n_1495)
);

NOR2xp33_ASAP7_75t_L g1496 ( 
.A(n_1443),
.B(n_1211),
.Y(n_1496)
);

NOR2xp33_ASAP7_75t_L g1497 ( 
.A(n_1479),
.B(n_1241),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_SL g1498 ( 
.A(n_1424),
.B(n_1275),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1449),
.B(n_1141),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_SL g1500 ( 
.A(n_1459),
.B(n_1274),
.Y(n_1500)
);

INVx3_ASAP7_75t_L g1501 ( 
.A(n_1421),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1422),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_SL g1503 ( 
.A(n_1472),
.B(n_1276),
.Y(n_1503)
);

BUFx4f_ASAP7_75t_L g1504 ( 
.A(n_1465),
.Y(n_1504)
);

INVx2_ASAP7_75t_SL g1505 ( 
.A(n_1428),
.Y(n_1505)
);

INVx4_ASAP7_75t_L g1506 ( 
.A(n_1442),
.Y(n_1506)
);

INVx3_ASAP7_75t_L g1507 ( 
.A(n_1421),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1427),
.Y(n_1508)
);

BUFx6f_ASAP7_75t_L g1509 ( 
.A(n_1473),
.Y(n_1509)
);

NOR2xp33_ASAP7_75t_L g1510 ( 
.A(n_1486),
.B(n_1089),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_SL g1511 ( 
.A(n_1463),
.B(n_1279),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1420),
.B(n_915),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1444),
.Y(n_1513)
);

AOI22xp33_ASAP7_75t_L g1514 ( 
.A1(n_1425),
.A2(n_1280),
.B1(n_1071),
.B2(n_1133),
.Y(n_1514)
);

BUFx2_ASAP7_75t_L g1515 ( 
.A(n_1432),
.Y(n_1515)
);

OAI22xp5_ASAP7_75t_L g1516 ( 
.A1(n_1433),
.A2(n_1153),
.B1(n_1176),
.B2(n_1037),
.Y(n_1516)
);

AOI22xp33_ASAP7_75t_L g1517 ( 
.A1(n_1440),
.A2(n_1250),
.B1(n_1258),
.B2(n_1053),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1469),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1470),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1475),
.Y(n_1520)
);

BUFx10_ASAP7_75t_L g1521 ( 
.A(n_1439),
.Y(n_1521)
);

BUFx8_ASAP7_75t_SL g1522 ( 
.A(n_1455),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_SL g1523 ( 
.A(n_1447),
.B(n_1285),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1476),
.Y(n_1524)
);

BUFx3_ASAP7_75t_L g1525 ( 
.A(n_1473),
.Y(n_1525)
);

NAND3xp33_ASAP7_75t_L g1526 ( 
.A(n_1446),
.B(n_951),
.C(n_943),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1481),
.Y(n_1527)
);

BUFx6f_ASAP7_75t_L g1528 ( 
.A(n_1442),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1451),
.Y(n_1529)
);

HB1xp67_ASAP7_75t_L g1530 ( 
.A(n_1477),
.Y(n_1530)
);

BUFx2_ASAP7_75t_L g1531 ( 
.A(n_1461),
.Y(n_1531)
);

NOR2xp33_ASAP7_75t_L g1532 ( 
.A(n_1436),
.B(n_1474),
.Y(n_1532)
);

AOI22xp33_ASAP7_75t_L g1533 ( 
.A1(n_1453),
.A2(n_1456),
.B1(n_1465),
.B2(n_1485),
.Y(n_1533)
);

NOR2xp33_ASAP7_75t_L g1534 ( 
.A(n_1468),
.B(n_955),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_SL g1535 ( 
.A(n_1419),
.B(n_1288),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1480),
.B(n_1157),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1445),
.Y(n_1537)
);

AND2x4_ASAP7_75t_L g1538 ( 
.A(n_1429),
.B(n_1029),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1457),
.Y(n_1539)
);

BUFx4f_ASAP7_75t_L g1540 ( 
.A(n_1452),
.Y(n_1540)
);

AOI22xp5_ASAP7_75t_L g1541 ( 
.A1(n_1416),
.A2(n_926),
.B1(n_928),
.B2(n_927),
.Y(n_1541)
);

OR2x6_ASAP7_75t_L g1542 ( 
.A(n_1462),
.B(n_1031),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1417),
.B(n_919),
.Y(n_1543)
);

BUFx2_ASAP7_75t_L g1544 ( 
.A(n_1483),
.Y(n_1544)
);

AND2x6_ASAP7_75t_L g1545 ( 
.A(n_1460),
.B(n_936),
.Y(n_1545)
);

AO21x2_ASAP7_75t_L g1546 ( 
.A1(n_1426),
.A2(n_952),
.B(n_944),
.Y(n_1546)
);

INVx1_ASAP7_75t_SL g1547 ( 
.A(n_1441),
.Y(n_1547)
);

NOR2xp33_ASAP7_75t_L g1548 ( 
.A(n_1458),
.B(n_961),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1464),
.Y(n_1549)
);

AOI22xp5_ASAP7_75t_L g1550 ( 
.A1(n_1466),
.A2(n_930),
.B1(n_933),
.B2(n_931),
.Y(n_1550)
);

INVxp67_ASAP7_75t_SL g1551 ( 
.A(n_1431),
.Y(n_1551)
);

NOR2x1p5_ASAP7_75t_L g1552 ( 
.A(n_1467),
.B(n_1269),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1435),
.B(n_958),
.Y(n_1553)
);

AOI22xp33_ASAP7_75t_L g1554 ( 
.A1(n_1434),
.A2(n_967),
.B1(n_983),
.B2(n_981),
.Y(n_1554)
);

NAND2x1p5_ASAP7_75t_L g1555 ( 
.A(n_1452),
.B(n_984),
.Y(n_1555)
);

INVx2_ASAP7_75t_L g1556 ( 
.A(n_1423),
.Y(n_1556)
);

AND2x6_ASAP7_75t_L g1557 ( 
.A(n_1414),
.B(n_994),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1415),
.Y(n_1558)
);

BUFx4f_ASAP7_75t_L g1559 ( 
.A(n_1454),
.Y(n_1559)
);

OR2x6_ASAP7_75t_L g1560 ( 
.A(n_1454),
.B(n_1073),
.Y(n_1560)
);

AO21x2_ASAP7_75t_L g1561 ( 
.A1(n_1471),
.A2(n_999),
.B(n_998),
.Y(n_1561)
);

INVxp67_ASAP7_75t_SL g1562 ( 
.A(n_1488),
.Y(n_1562)
);

HB1xp67_ASAP7_75t_L g1563 ( 
.A(n_1478),
.Y(n_1563)
);

BUFx6f_ASAP7_75t_L g1564 ( 
.A(n_1482),
.Y(n_1564)
);

OR2x6_ASAP7_75t_L g1565 ( 
.A(n_1484),
.B(n_1075),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1487),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_SL g1567 ( 
.A(n_1438),
.B(n_934),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1443),
.B(n_1007),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_SL g1569 ( 
.A(n_1438),
.B(n_1262),
.Y(n_1569)
);

BUFx6f_ASAP7_75t_L g1570 ( 
.A(n_1421),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_SL g1571 ( 
.A(n_1438),
.B(n_935),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_SL g1572 ( 
.A(n_1438),
.B(n_941),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1418),
.Y(n_1573)
);

BUFx6f_ASAP7_75t_L g1574 ( 
.A(n_1421),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1418),
.Y(n_1575)
);

INVx3_ASAP7_75t_L g1576 ( 
.A(n_1421),
.Y(n_1576)
);

OR2x6_ASAP7_75t_L g1577 ( 
.A(n_1428),
.B(n_1079),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1418),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1418),
.Y(n_1579)
);

AOI22xp33_ASAP7_75t_L g1580 ( 
.A1(n_1443),
.A2(n_1008),
.B1(n_1020),
.B2(n_1019),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1418),
.Y(n_1581)
);

NAND2xp33_ASAP7_75t_L g1582 ( 
.A(n_1437),
.B(n_953),
.Y(n_1582)
);

BUFx2_ASAP7_75t_L g1583 ( 
.A(n_1432),
.Y(n_1583)
);

AOI22xp33_ASAP7_75t_L g1584 ( 
.A1(n_1443),
.A2(n_1023),
.B1(n_1033),
.B2(n_1025),
.Y(n_1584)
);

BUFx6f_ASAP7_75t_L g1585 ( 
.A(n_1421),
.Y(n_1585)
);

AND2x6_ASAP7_75t_L g1586 ( 
.A(n_1437),
.B(n_1035),
.Y(n_1586)
);

INVxp67_ASAP7_75t_SL g1587 ( 
.A(n_1430),
.Y(n_1587)
);

CKINVDCx5p33_ASAP7_75t_R g1588 ( 
.A(n_1429),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1443),
.B(n_1042),
.Y(n_1589)
);

NOR3xp33_ASAP7_75t_L g1590 ( 
.A(n_1424),
.B(n_975),
.C(n_962),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1448),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_SL g1592 ( 
.A(n_1438),
.B(n_1259),
.Y(n_1592)
);

OAI22xp33_ASAP7_75t_L g1593 ( 
.A1(n_1438),
.A2(n_1083),
.B1(n_1115),
.B2(n_1069),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1418),
.Y(n_1594)
);

AOI22xp5_ASAP7_75t_SL g1595 ( 
.A1(n_1455),
.A2(n_1173),
.B1(n_1194),
.B2(n_1159),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_SL g1596 ( 
.A(n_1438),
.B(n_954),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1448),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_SL g1598 ( 
.A(n_1438),
.B(n_956),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1448),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1448),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1418),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1443),
.B(n_1064),
.Y(n_1602)
);

NOR2xp33_ASAP7_75t_L g1603 ( 
.A(n_1438),
.B(n_986),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1448),
.Y(n_1604)
);

INVx8_ASAP7_75t_L g1605 ( 
.A(n_1509),
.Y(n_1605)
);

NAND2xp33_ASAP7_75t_L g1606 ( 
.A(n_1586),
.B(n_1517),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1496),
.B(n_1067),
.Y(n_1607)
);

AOI221xp5_ASAP7_75t_L g1608 ( 
.A1(n_1548),
.A2(n_1095),
.B1(n_1144),
.B2(n_1145),
.C(n_1140),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1489),
.Y(n_1609)
);

INVx1_ASAP7_75t_SL g1610 ( 
.A(n_1530),
.Y(n_1610)
);

INVx1_ASAP7_75t_SL g1611 ( 
.A(n_1515),
.Y(n_1611)
);

AND2x4_ASAP7_75t_L g1612 ( 
.A(n_1506),
.B(n_1146),
.Y(n_1612)
);

NOR2xp33_ASAP7_75t_L g1613 ( 
.A(n_1532),
.B(n_1212),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1568),
.B(n_1081),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1494),
.Y(n_1615)
);

INVx2_ASAP7_75t_SL g1616 ( 
.A(n_1528),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_SL g1617 ( 
.A(n_1497),
.B(n_960),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1589),
.B(n_1099),
.Y(n_1618)
);

AOI22xp33_ASAP7_75t_L g1619 ( 
.A1(n_1590),
.A2(n_1104),
.B1(n_1112),
.B2(n_1109),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1602),
.B(n_1121),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_SL g1621 ( 
.A(n_1495),
.B(n_966),
.Y(n_1621)
);

AOI22xp5_ASAP7_75t_L g1622 ( 
.A1(n_1586),
.A2(n_1135),
.B1(n_1148),
.B2(n_1123),
.Y(n_1622)
);

NAND2xp33_ASAP7_75t_L g1623 ( 
.A(n_1586),
.B(n_1184),
.Y(n_1623)
);

HB1xp67_ASAP7_75t_L g1624 ( 
.A(n_1583),
.Y(n_1624)
);

BUFx3_ASAP7_75t_L g1625 ( 
.A(n_1528),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1603),
.B(n_1155),
.Y(n_1626)
);

NAND2x1_ASAP7_75t_L g1627 ( 
.A(n_1490),
.B(n_1077),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1529),
.Y(n_1628)
);

INVxp67_ASAP7_75t_L g1629 ( 
.A(n_1536),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1591),
.Y(n_1630)
);

NOR2xp67_ASAP7_75t_L g1631 ( 
.A(n_1588),
.B(n_970),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_SL g1632 ( 
.A(n_1499),
.B(n_972),
.Y(n_1632)
);

NOR2xp33_ASAP7_75t_SL g1633 ( 
.A(n_1531),
.B(n_1215),
.Y(n_1633)
);

OR2x2_ASAP7_75t_L g1634 ( 
.A(n_1493),
.B(n_1271),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_SL g1635 ( 
.A(n_1534),
.B(n_973),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1597),
.B(n_1158),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1599),
.B(n_1186),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1600),
.B(n_1187),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_SL g1639 ( 
.A(n_1604),
.B(n_1533),
.Y(n_1639)
);

XOR2xp5_ASAP7_75t_L g1640 ( 
.A(n_1595),
.B(n_1226),
.Y(n_1640)
);

INVx1_ASAP7_75t_SL g1641 ( 
.A(n_1492),
.Y(n_1641)
);

NOR2xp33_ASAP7_75t_L g1642 ( 
.A(n_1567),
.B(n_1234),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1543),
.B(n_1188),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1502),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1508),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_SL g1646 ( 
.A(n_1510),
.B(n_974),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1513),
.B(n_1189),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1518),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1519),
.B(n_1190),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1520),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1524),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1527),
.B(n_1191),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1573),
.B(n_1192),
.Y(n_1653)
);

BUFx4f_ASAP7_75t_L g1654 ( 
.A(n_1509),
.Y(n_1654)
);

NOR2xp33_ASAP7_75t_L g1655 ( 
.A(n_1569),
.B(n_1238),
.Y(n_1655)
);

INVx5_ASAP7_75t_L g1656 ( 
.A(n_1570),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1538),
.B(n_990),
.Y(n_1657)
);

BUFx6f_ASAP7_75t_L g1658 ( 
.A(n_1570),
.Y(n_1658)
);

BUFx3_ASAP7_75t_L g1659 ( 
.A(n_1540),
.Y(n_1659)
);

AND2x6_ASAP7_75t_L g1660 ( 
.A(n_1558),
.B(n_1220),
.Y(n_1660)
);

NOR2xp33_ASAP7_75t_L g1661 ( 
.A(n_1571),
.B(n_1240),
.Y(n_1661)
);

NOR2xp33_ASAP7_75t_L g1662 ( 
.A(n_1572),
.B(n_1255),
.Y(n_1662)
);

BUFx3_ASAP7_75t_L g1663 ( 
.A(n_1559),
.Y(n_1663)
);

INVxp33_ASAP7_75t_L g1664 ( 
.A(n_1574),
.Y(n_1664)
);

INVx2_ASAP7_75t_SL g1665 ( 
.A(n_1574),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1575),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1578),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1579),
.Y(n_1668)
);

INVx2_ASAP7_75t_SL g1669 ( 
.A(n_1585),
.Y(n_1669)
);

AOI22xp5_ASAP7_75t_L g1670 ( 
.A1(n_1582),
.A2(n_1229),
.B1(n_1232),
.B2(n_1222),
.Y(n_1670)
);

NAND3xp33_ASAP7_75t_L g1671 ( 
.A(n_1498),
.B(n_992),
.C(n_991),
.Y(n_1671)
);

NOR2xp33_ASAP7_75t_L g1672 ( 
.A(n_1592),
.B(n_1264),
.Y(n_1672)
);

OR2x2_ASAP7_75t_L g1673 ( 
.A(n_1544),
.B(n_1282),
.Y(n_1673)
);

NOR2xp33_ASAP7_75t_L g1674 ( 
.A(n_1596),
.B(n_995),
.Y(n_1674)
);

NOR2xp33_ASAP7_75t_L g1675 ( 
.A(n_1598),
.B(n_997),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_1581),
.Y(n_1676)
);

AOI22xp33_ASAP7_75t_L g1677 ( 
.A1(n_1516),
.A2(n_1267),
.B1(n_1270),
.B2(n_1252),
.Y(n_1677)
);

INVxp67_ASAP7_75t_L g1678 ( 
.A(n_1563),
.Y(n_1678)
);

INVx2_ASAP7_75t_SL g1679 ( 
.A(n_1585),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1594),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1601),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1539),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1580),
.B(n_1584),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1500),
.B(n_1277),
.Y(n_1684)
);

AND2x4_ASAP7_75t_L g1685 ( 
.A(n_1525),
.B(n_1149),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1503),
.B(n_978),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1537),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1549),
.Y(n_1688)
);

AOI22xp5_ASAP7_75t_L g1689 ( 
.A1(n_1511),
.A2(n_979),
.B1(n_987),
.B2(n_980),
.Y(n_1689)
);

INVx3_ASAP7_75t_L g1690 ( 
.A(n_1501),
.Y(n_1690)
);

INVx1_ASAP7_75t_SL g1691 ( 
.A(n_1547),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1505),
.B(n_1003),
.Y(n_1692)
);

NOR2xp33_ASAP7_75t_L g1693 ( 
.A(n_1535),
.B(n_1009),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1551),
.B(n_988),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1512),
.B(n_989),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1553),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1566),
.Y(n_1697)
);

INVx8_ASAP7_75t_L g1698 ( 
.A(n_1557),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1556),
.Y(n_1699)
);

AOI22xp5_ASAP7_75t_L g1700 ( 
.A1(n_1523),
.A2(n_996),
.B1(n_1004),
.B2(n_1001),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_SL g1701 ( 
.A(n_1550),
.B(n_1005),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1564),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1491),
.Y(n_1703)
);

BUFx4_ASAP7_75t_L g1704 ( 
.A(n_1504),
.Y(n_1704)
);

AOI22xp5_ASAP7_75t_L g1705 ( 
.A1(n_1526),
.A2(n_1010),
.B1(n_1018),
.B2(n_1015),
.Y(n_1705)
);

NOR2xp33_ASAP7_75t_L g1706 ( 
.A(n_1541),
.B(n_1011),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1587),
.B(n_1021),
.Y(n_1707)
);

AND2x4_ASAP7_75t_SL g1708 ( 
.A(n_1521),
.B(n_1077),
.Y(n_1708)
);

OAI22xp5_ASAP7_75t_L g1709 ( 
.A1(n_1514),
.A2(n_1034),
.B1(n_1036),
.B2(n_1028),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1577),
.B(n_1012),
.Y(n_1710)
);

INVxp67_ASAP7_75t_L g1711 ( 
.A(n_1577),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1564),
.Y(n_1712)
);

AOI22xp33_ASAP7_75t_L g1713 ( 
.A1(n_1542),
.A2(n_1184),
.B1(n_1265),
.B2(n_1199),
.Y(n_1713)
);

NOR2xp33_ASAP7_75t_L g1714 ( 
.A(n_1542),
.B(n_1014),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1546),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1562),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1561),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1545),
.B(n_1593),
.Y(n_1718)
);

NOR2xp33_ASAP7_75t_SL g1719 ( 
.A(n_1522),
.B(n_1038),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1545),
.B(n_1040),
.Y(n_1720)
);

INVx8_ASAP7_75t_L g1721 ( 
.A(n_1557),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_SL g1722 ( 
.A(n_1507),
.B(n_1576),
.Y(n_1722)
);

INVx2_ASAP7_75t_SL g1723 ( 
.A(n_1552),
.Y(n_1723)
);

CKINVDCx20_ASAP7_75t_R g1724 ( 
.A(n_1560),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1545),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1557),
.B(n_1046),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1554),
.B(n_1052),
.Y(n_1727)
);

NAND2xp33_ASAP7_75t_L g1728 ( 
.A(n_1555),
.B(n_1184),
.Y(n_1728)
);

NOR2xp33_ASAP7_75t_L g1729 ( 
.A(n_1565),
.B(n_1560),
.Y(n_1729)
);

OAI22xp5_ASAP7_75t_L g1730 ( 
.A1(n_1565),
.A2(n_1056),
.B1(n_1057),
.B2(n_1054),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1496),
.B(n_1058),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_SL g1732 ( 
.A(n_1496),
.B(n_1060),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1489),
.Y(n_1733)
);

NOR2xp33_ASAP7_75t_L g1734 ( 
.A(n_1532),
.B(n_1016),
.Y(n_1734)
);

AND2x6_ASAP7_75t_SL g1735 ( 
.A(n_1542),
.B(n_1256),
.Y(n_1735)
);

INVx2_ASAP7_75t_SL g1736 ( 
.A(n_1530),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1493),
.B(n_1017),
.Y(n_1737)
);

OAI22xp5_ASAP7_75t_L g1738 ( 
.A1(n_1496),
.A2(n_1070),
.B1(n_1074),
.B2(n_1066),
.Y(n_1738)
);

AO221x1_ASAP7_75t_L g1739 ( 
.A1(n_1593),
.A2(n_1177),
.B1(n_1183),
.B2(n_1180),
.C(n_1175),
.Y(n_1739)
);

NOR2xp33_ASAP7_75t_L g1740 ( 
.A(n_1532),
.B(n_1024),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1496),
.B(n_1078),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1490),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1489),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1489),
.Y(n_1744)
);

AO22x2_ASAP7_75t_L g1745 ( 
.A1(n_1516),
.A2(n_1206),
.B1(n_1214),
.B2(n_1185),
.Y(n_1745)
);

INVx2_ASAP7_75t_SL g1746 ( 
.A(n_1530),
.Y(n_1746)
);

NOR2xp33_ASAP7_75t_L g1747 ( 
.A(n_1532),
.B(n_1027),
.Y(n_1747)
);

AOI22xp33_ASAP7_75t_L g1748 ( 
.A1(n_1548),
.A2(n_1184),
.B1(n_1265),
.B2(n_1199),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1490),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1496),
.B(n_1080),
.Y(n_1750)
);

NOR2xp33_ASAP7_75t_L g1751 ( 
.A(n_1532),
.B(n_1032),
.Y(n_1751)
);

NOR2xp33_ASAP7_75t_SL g1752 ( 
.A(n_1530),
.B(n_1082),
.Y(n_1752)
);

OAI22xp5_ASAP7_75t_L g1753 ( 
.A1(n_1496),
.A2(n_1085),
.B1(n_1086),
.B2(n_1084),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1496),
.B(n_1088),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1490),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1489),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1496),
.B(n_1090),
.Y(n_1757)
);

INVx8_ASAP7_75t_L g1758 ( 
.A(n_1509),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1496),
.B(n_1101),
.Y(n_1759)
);

NOR2xp33_ASAP7_75t_R g1760 ( 
.A(n_1588),
.B(n_1106),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1496),
.B(n_1107),
.Y(n_1761)
);

NOR2xp33_ASAP7_75t_L g1762 ( 
.A(n_1532),
.B(n_1039),
.Y(n_1762)
);

INVx3_ASAP7_75t_L g1763 ( 
.A(n_1528),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1496),
.B(n_1110),
.Y(n_1764)
);

NAND2xp33_ASAP7_75t_L g1765 ( 
.A(n_1586),
.B(n_1114),
.Y(n_1765)
);

INVxp67_ASAP7_75t_L g1766 ( 
.A(n_1530),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1496),
.B(n_1116),
.Y(n_1767)
);

NAND3xp33_ASAP7_75t_L g1768 ( 
.A(n_1496),
.B(n_1044),
.C(n_1043),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1609),
.Y(n_1769)
);

OAI21x1_ASAP7_75t_L g1770 ( 
.A1(n_1715),
.A2(n_1235),
.B(n_1223),
.Y(n_1770)
);

OAI22xp5_ASAP7_75t_SL g1771 ( 
.A1(n_1640),
.A2(n_1132),
.B1(n_1152),
.B2(n_1094),
.Y(n_1771)
);

AOI22xp33_ASAP7_75t_SL g1772 ( 
.A1(n_1613),
.A2(n_1287),
.B1(n_1286),
.B2(n_1048),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_SL g1773 ( 
.A(n_1691),
.B(n_1736),
.Y(n_1773)
);

AOI22xp5_ASAP7_75t_L g1774 ( 
.A1(n_1734),
.A2(n_1119),
.B1(n_1122),
.B2(n_1118),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1740),
.B(n_1134),
.Y(n_1775)
);

AND2x2_ASAP7_75t_SL g1776 ( 
.A(n_1747),
.B(n_925),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1751),
.B(n_1136),
.Y(n_1777)
);

AOI21xp5_ASAP7_75t_L g1778 ( 
.A1(n_1606),
.A2(n_1265),
.B(n_1199),
.Y(n_1778)
);

BUFx6f_ASAP7_75t_L g1779 ( 
.A(n_1658),
.Y(n_1779)
);

NOR2xp33_ASAP7_75t_L g1780 ( 
.A(n_1762),
.B(n_1045),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_SL g1781 ( 
.A(n_1746),
.B(n_1138),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1644),
.Y(n_1782)
);

BUFx6f_ASAP7_75t_L g1783 ( 
.A(n_1658),
.Y(n_1783)
);

AND3x2_ASAP7_75t_SL g1784 ( 
.A(n_1702),
.B(n_1049),
.C(n_1030),
.Y(n_1784)
);

INVx4_ASAP7_75t_L g1785 ( 
.A(n_1605),
.Y(n_1785)
);

INVx4_ASAP7_75t_L g1786 ( 
.A(n_1605),
.Y(n_1786)
);

INVx3_ASAP7_75t_L g1787 ( 
.A(n_1758),
.Y(n_1787)
);

NOR2xp33_ASAP7_75t_L g1788 ( 
.A(n_1642),
.B(n_1062),
.Y(n_1788)
);

AND2x6_ASAP7_75t_SL g1789 ( 
.A(n_1714),
.B(n_1239),
.Y(n_1789)
);

AOI22xp5_ASAP7_75t_L g1790 ( 
.A1(n_1706),
.A2(n_1260),
.B1(n_1257),
.B2(n_1143),
.Y(n_1790)
);

INVxp67_ASAP7_75t_L g1791 ( 
.A(n_1624),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_SL g1792 ( 
.A(n_1610),
.B(n_1142),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1696),
.B(n_1154),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_1645),
.Y(n_1794)
);

BUFx6f_ASAP7_75t_L g1795 ( 
.A(n_1758),
.Y(n_1795)
);

BUFx2_ASAP7_75t_L g1796 ( 
.A(n_1611),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1737),
.B(n_1065),
.Y(n_1797)
);

BUFx2_ASAP7_75t_L g1798 ( 
.A(n_1766),
.Y(n_1798)
);

NAND2x1p5_ASAP7_75t_L g1799 ( 
.A(n_1656),
.B(n_1654),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1615),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1628),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_1676),
.Y(n_1802)
);

AOI221xp5_ASAP7_75t_SL g1803 ( 
.A1(n_1608),
.A2(n_1261),
.B1(n_1266),
.B2(n_1248),
.C(n_1247),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1607),
.B(n_1161),
.Y(n_1804)
);

INVx2_ASAP7_75t_L g1805 ( 
.A(n_1742),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1630),
.Y(n_1806)
);

INVx1_ASAP7_75t_SL g1807 ( 
.A(n_1704),
.Y(n_1807)
);

INVx2_ASAP7_75t_SL g1808 ( 
.A(n_1656),
.Y(n_1808)
);

BUFx6f_ASAP7_75t_L g1809 ( 
.A(n_1656),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1731),
.B(n_1163),
.Y(n_1810)
);

INVx2_ASAP7_75t_L g1811 ( 
.A(n_1749),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1655),
.B(n_1068),
.Y(n_1812)
);

NOR3xp33_ASAP7_75t_SL g1813 ( 
.A(n_1661),
.B(n_1098),
.C(n_1097),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1733),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1741),
.B(n_1166),
.Y(n_1815)
);

INVx4_ASAP7_75t_L g1816 ( 
.A(n_1659),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1662),
.B(n_1102),
.Y(n_1817)
);

BUFx6f_ASAP7_75t_L g1818 ( 
.A(n_1663),
.Y(n_1818)
);

AOI22xp5_ASAP7_75t_L g1819 ( 
.A1(n_1672),
.A2(n_1254),
.B1(n_1169),
.B2(n_1179),
.Y(n_1819)
);

INVx2_ASAP7_75t_L g1820 ( 
.A(n_1755),
.Y(n_1820)
);

NOR2x2_ASAP7_75t_L g1821 ( 
.A(n_1688),
.B(n_1712),
.Y(n_1821)
);

AOI22xp33_ASAP7_75t_L g1822 ( 
.A1(n_1626),
.A2(n_1181),
.B1(n_1182),
.B2(n_1168),
.Y(n_1822)
);

INVx3_ASAP7_75t_L g1823 ( 
.A(n_1625),
.Y(n_1823)
);

OR2x2_ASAP7_75t_L g1824 ( 
.A(n_1673),
.B(n_1105),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_SL g1825 ( 
.A(n_1633),
.B(n_1203),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1743),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1744),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_SL g1828 ( 
.A(n_1752),
.B(n_1207),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_SL g1829 ( 
.A(n_1718),
.B(n_1208),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1756),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_SL g1831 ( 
.A(n_1629),
.B(n_1209),
.Y(n_1831)
);

NAND2xp33_ASAP7_75t_L g1832 ( 
.A(n_1698),
.B(n_1210),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1682),
.Y(n_1833)
);

NOR2xp33_ASAP7_75t_L g1834 ( 
.A(n_1678),
.B(n_1108),
.Y(n_1834)
);

OR2x6_ASAP7_75t_L g1835 ( 
.A(n_1698),
.B(n_1272),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1750),
.B(n_1219),
.Y(n_1836)
);

AND2x6_ASAP7_75t_L g1837 ( 
.A(n_1725),
.B(n_1273),
.Y(n_1837)
);

AND2x4_ASAP7_75t_L g1838 ( 
.A(n_1641),
.B(n_1051),
.Y(n_1838)
);

INVx2_ASAP7_75t_SL g1839 ( 
.A(n_1763),
.Y(n_1839)
);

INVx2_ASAP7_75t_L g1840 ( 
.A(n_1687),
.Y(n_1840)
);

INVx5_ASAP7_75t_L g1841 ( 
.A(n_1735),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1697),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_SL g1843 ( 
.A(n_1768),
.B(n_1224),
.Y(n_1843)
);

CKINVDCx5p33_ASAP7_75t_R g1844 ( 
.A(n_1760),
.Y(n_1844)
);

INVx2_ASAP7_75t_L g1845 ( 
.A(n_1648),
.Y(n_1845)
);

AOI21xp5_ASAP7_75t_L g1846 ( 
.A1(n_1639),
.A2(n_1230),
.B(n_1228),
.Y(n_1846)
);

AOI22xp33_ASAP7_75t_L g1847 ( 
.A1(n_1683),
.A2(n_1242),
.B1(n_1243),
.B2(n_1233),
.Y(n_1847)
);

INVx5_ASAP7_75t_L g1848 ( 
.A(n_1616),
.Y(n_1848)
);

INVx3_ASAP7_75t_L g1849 ( 
.A(n_1690),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1754),
.B(n_1244),
.Y(n_1850)
);

AOI22xp5_ASAP7_75t_L g1851 ( 
.A1(n_1674),
.A2(n_1245),
.B1(n_1113),
.B2(n_1126),
.Y(n_1851)
);

BUFx6f_ASAP7_75t_L g1852 ( 
.A(n_1665),
.Y(n_1852)
);

NOR2xp33_ASAP7_75t_L g1853 ( 
.A(n_1757),
.B(n_1124),
.Y(n_1853)
);

BUFx2_ASAP7_75t_L g1854 ( 
.A(n_1724),
.Y(n_1854)
);

A2O1A1Ixp33_ASAP7_75t_L g1855 ( 
.A1(n_1675),
.A2(n_1120),
.B(n_1174),
.C(n_1103),
.Y(n_1855)
);

AOI21x1_ASAP7_75t_L g1856 ( 
.A1(n_1717),
.A2(n_1618),
.B(n_1614),
.Y(n_1856)
);

INVx3_ASAP7_75t_L g1857 ( 
.A(n_1669),
.Y(n_1857)
);

INVx2_ASAP7_75t_L g1858 ( 
.A(n_1650),
.Y(n_1858)
);

OR2x6_ASAP7_75t_L g1859 ( 
.A(n_1721),
.B(n_1679),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1651),
.Y(n_1860)
);

NOR2x1_ASAP7_75t_L g1861 ( 
.A(n_1671),
.B(n_1196),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1759),
.B(n_1127),
.Y(n_1862)
);

AOI22xp33_ASAP7_75t_L g1863 ( 
.A1(n_1619),
.A2(n_1139),
.B1(n_1151),
.B2(n_1129),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1657),
.B(n_1156),
.Y(n_1864)
);

INVx3_ASAP7_75t_L g1865 ( 
.A(n_1685),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1634),
.B(n_1164),
.Y(n_1866)
);

AND2x4_ASAP7_75t_L g1867 ( 
.A(n_1723),
.B(n_1711),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1761),
.B(n_1167),
.Y(n_1868)
);

NOR2x1_ASAP7_75t_L g1869 ( 
.A(n_1631),
.B(n_1170),
.Y(n_1869)
);

AND2x4_ASAP7_75t_L g1870 ( 
.A(n_1699),
.B(n_458),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1666),
.Y(n_1871)
);

INVx2_ASAP7_75t_SL g1872 ( 
.A(n_1612),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1764),
.B(n_1172),
.Y(n_1873)
);

OAI22xp33_ASAP7_75t_L g1874 ( 
.A1(n_1767),
.A2(n_1195),
.B1(n_1197),
.B2(n_1178),
.Y(n_1874)
);

INVx5_ASAP7_75t_L g1875 ( 
.A(n_1660),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1667),
.Y(n_1876)
);

AOI22xp33_ASAP7_75t_L g1877 ( 
.A1(n_1693),
.A2(n_1202),
.B1(n_1200),
.B2(n_1204),
.Y(n_1877)
);

HB1xp67_ASAP7_75t_L g1878 ( 
.A(n_1664),
.Y(n_1878)
);

CKINVDCx5p33_ASAP7_75t_R g1879 ( 
.A(n_1729),
.Y(n_1879)
);

AOI22xp33_ASAP7_75t_L g1880 ( 
.A1(n_1748),
.A2(n_1227),
.B1(n_1225),
.B2(n_1236),
.Y(n_1880)
);

INVx2_ASAP7_75t_L g1881 ( 
.A(n_1668),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_SL g1882 ( 
.A(n_1716),
.B(n_1246),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1680),
.Y(n_1883)
);

AOI22xp33_ASAP7_75t_L g1884 ( 
.A1(n_1621),
.A2(n_1251),
.B1(n_1249),
.B2(n_1253),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1732),
.B(n_0),
.Y(n_1885)
);

INVx2_ASAP7_75t_SL g1886 ( 
.A(n_1692),
.Y(n_1886)
);

AND2x2_ASAP7_75t_L g1887 ( 
.A(n_1776),
.B(n_1710),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1769),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1800),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_SL g1890 ( 
.A(n_1780),
.B(n_1719),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_SL g1891 ( 
.A(n_1886),
.B(n_1703),
.Y(n_1891)
);

HB1xp67_ASAP7_75t_L g1892 ( 
.A(n_1796),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1853),
.B(n_1617),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_L g1894 ( 
.A(n_1788),
.B(n_1646),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_SL g1895 ( 
.A(n_1879),
.B(n_1694),
.Y(n_1895)
);

OAI22xp5_ASAP7_75t_L g1896 ( 
.A1(n_1775),
.A2(n_1635),
.B1(n_1686),
.B2(n_1681),
.Y(n_1896)
);

AND2x4_ASAP7_75t_L g1897 ( 
.A(n_1785),
.B(n_1722),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1801),
.Y(n_1898)
);

INVx2_ASAP7_75t_L g1899 ( 
.A(n_1840),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1812),
.B(n_1636),
.Y(n_1900)
);

NOR2xp33_ASAP7_75t_R g1901 ( 
.A(n_1844),
.B(n_1721),
.Y(n_1901)
);

NOR2x1p5_ASAP7_75t_SL g1902 ( 
.A(n_1856),
.B(n_1623),
.Y(n_1902)
);

OR2x2_ASAP7_75t_L g1903 ( 
.A(n_1798),
.B(n_1637),
.Y(n_1903)
);

INVx3_ASAP7_75t_L g1904 ( 
.A(n_1816),
.Y(n_1904)
);

AND2x4_ASAP7_75t_L g1905 ( 
.A(n_1786),
.B(n_1708),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1817),
.B(n_1638),
.Y(n_1906)
);

INVx2_ASAP7_75t_L g1907 ( 
.A(n_1806),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1814),
.Y(n_1908)
);

OR2x6_ASAP7_75t_L g1909 ( 
.A(n_1818),
.B(n_1745),
.Y(n_1909)
);

INVx4_ASAP7_75t_L g1910 ( 
.A(n_1818),
.Y(n_1910)
);

AND2x4_ASAP7_75t_L g1911 ( 
.A(n_1787),
.B(n_1632),
.Y(n_1911)
);

NAND2x1p5_ASAP7_75t_L g1912 ( 
.A(n_1795),
.B(n_1627),
.Y(n_1912)
);

INVx5_ASAP7_75t_L g1913 ( 
.A(n_1809),
.Y(n_1913)
);

NOR2xp33_ASAP7_75t_L g1914 ( 
.A(n_1791),
.B(n_1738),
.Y(n_1914)
);

HB1xp67_ASAP7_75t_L g1915 ( 
.A(n_1878),
.Y(n_1915)
);

INVx2_ASAP7_75t_L g1916 ( 
.A(n_1826),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_1777),
.B(n_1862),
.Y(n_1917)
);

OR2x6_ASAP7_75t_L g1918 ( 
.A(n_1799),
.B(n_1745),
.Y(n_1918)
);

INVx2_ASAP7_75t_L g1919 ( 
.A(n_1827),
.Y(n_1919)
);

INVx2_ASAP7_75t_L g1920 ( 
.A(n_1830),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_L g1921 ( 
.A(n_1868),
.B(n_1620),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1873),
.B(n_1660),
.Y(n_1922)
);

BUFx4f_ASAP7_75t_L g1923 ( 
.A(n_1795),
.Y(n_1923)
);

OAI21xp5_ASAP7_75t_L g1924 ( 
.A1(n_1829),
.A2(n_1778),
.B(n_1793),
.Y(n_1924)
);

INVx3_ASAP7_75t_L g1925 ( 
.A(n_1809),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1833),
.B(n_1660),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1842),
.B(n_1695),
.Y(n_1927)
);

BUFx3_ASAP7_75t_L g1928 ( 
.A(n_1779),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1797),
.B(n_1643),
.Y(n_1929)
);

INVx2_ASAP7_75t_L g1930 ( 
.A(n_1860),
.Y(n_1930)
);

NOR2xp33_ASAP7_75t_L g1931 ( 
.A(n_1773),
.B(n_1753),
.Y(n_1931)
);

AOI22xp33_ASAP7_75t_L g1932 ( 
.A1(n_1772),
.A2(n_1701),
.B1(n_1739),
.B2(n_1765),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_L g1933 ( 
.A(n_1804),
.B(n_1707),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1810),
.B(n_1684),
.Y(n_1934)
);

BUFx3_ASAP7_75t_L g1935 ( 
.A(n_1779),
.Y(n_1935)
);

INVx2_ASAP7_75t_L g1936 ( 
.A(n_1871),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1815),
.B(n_1689),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1836),
.B(n_1726),
.Y(n_1938)
);

AND2x4_ASAP7_75t_L g1939 ( 
.A(n_1867),
.B(n_1720),
.Y(n_1939)
);

INVx2_ASAP7_75t_L g1940 ( 
.A(n_1876),
.Y(n_1940)
);

OR2x6_ASAP7_75t_L g1941 ( 
.A(n_1859),
.B(n_1647),
.Y(n_1941)
);

AND2x4_ASAP7_75t_L g1942 ( 
.A(n_1872),
.B(n_1653),
.Y(n_1942)
);

CKINVDCx5p33_ASAP7_75t_R g1943 ( 
.A(n_1807),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1883),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1845),
.Y(n_1945)
);

AOI22xp5_ASAP7_75t_L g1946 ( 
.A1(n_1771),
.A2(n_1705),
.B1(n_1700),
.B2(n_1730),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_L g1947 ( 
.A(n_1850),
.B(n_1713),
.Y(n_1947)
);

INVx2_ASAP7_75t_SL g1948 ( 
.A(n_1848),
.Y(n_1948)
);

AND2x4_ASAP7_75t_L g1949 ( 
.A(n_1865),
.B(n_1649),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1858),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_L g1951 ( 
.A(n_1866),
.B(n_1652),
.Y(n_1951)
);

INVx2_ASAP7_75t_SL g1952 ( 
.A(n_1848),
.Y(n_1952)
);

NOR2xp33_ASAP7_75t_L g1953 ( 
.A(n_1834),
.B(n_1709),
.Y(n_1953)
);

BUFx2_ASAP7_75t_SL g1954 ( 
.A(n_1823),
.Y(n_1954)
);

INVx2_ASAP7_75t_L g1955 ( 
.A(n_1881),
.Y(n_1955)
);

BUFx6f_ASAP7_75t_L g1956 ( 
.A(n_1783),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1864),
.B(n_1670),
.Y(n_1957)
);

INVx2_ASAP7_75t_L g1958 ( 
.A(n_1782),
.Y(n_1958)
);

INVx3_ASAP7_75t_L g1959 ( 
.A(n_1783),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1794),
.B(n_1677),
.Y(n_1960)
);

INVx5_ASAP7_75t_L g1961 ( 
.A(n_1852),
.Y(n_1961)
);

INVx2_ASAP7_75t_L g1962 ( 
.A(n_1802),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_L g1963 ( 
.A(n_1805),
.B(n_1811),
.Y(n_1963)
);

INVx2_ASAP7_75t_L g1964 ( 
.A(n_1820),
.Y(n_1964)
);

NOR2xp33_ASAP7_75t_SL g1965 ( 
.A(n_1841),
.B(n_1727),
.Y(n_1965)
);

BUFx3_ASAP7_75t_L g1966 ( 
.A(n_1852),
.Y(n_1966)
);

INVx2_ASAP7_75t_L g1967 ( 
.A(n_1770),
.Y(n_1967)
);

INVx2_ASAP7_75t_L g1968 ( 
.A(n_1849),
.Y(n_1968)
);

INVx5_ASAP7_75t_L g1969 ( 
.A(n_1835),
.Y(n_1969)
);

HB1xp67_ASAP7_75t_L g1970 ( 
.A(n_1857),
.Y(n_1970)
);

AND2x4_ASAP7_75t_L g1971 ( 
.A(n_1839),
.B(n_1622),
.Y(n_1971)
);

INVx2_ASAP7_75t_L g1972 ( 
.A(n_1821),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1870),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_L g1974 ( 
.A(n_1874),
.B(n_1728),
.Y(n_1974)
);

AOI221xp5_ASAP7_75t_L g1975 ( 
.A1(n_1877),
.A2(n_3),
.B1(n_1),
.B2(n_2),
.C(n_4),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1885),
.Y(n_1976)
);

AOI22xp5_ASAP7_75t_L g1977 ( 
.A1(n_1790),
.A2(n_4),
.B1(n_2),
.B2(n_3),
.Y(n_1977)
);

HB1xp67_ASAP7_75t_L g1978 ( 
.A(n_1838),
.Y(n_1978)
);

INVx3_ASAP7_75t_L g1979 ( 
.A(n_1808),
.Y(n_1979)
);

BUFx12f_ASAP7_75t_L g1980 ( 
.A(n_1854),
.Y(n_1980)
);

BUFx2_ASAP7_75t_L g1981 ( 
.A(n_1837),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1803),
.B(n_5),
.Y(n_1982)
);

BUFx2_ASAP7_75t_L g1983 ( 
.A(n_1837),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1882),
.B(n_5),
.Y(n_1984)
);

BUFx2_ASAP7_75t_L g1985 ( 
.A(n_1837),
.Y(n_1985)
);

NOR2xp33_ASAP7_75t_L g1986 ( 
.A(n_1824),
.B(n_6),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_L g1987 ( 
.A(n_1813),
.B(n_6),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_SL g1988 ( 
.A(n_1875),
.B(n_7),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1861),
.Y(n_1989)
);

OAI22xp5_ASAP7_75t_L g1990 ( 
.A1(n_1847),
.A2(n_9),
.B1(n_7),
.B2(n_8),
.Y(n_1990)
);

BUFx3_ASAP7_75t_L g1991 ( 
.A(n_1841),
.Y(n_1991)
);

INVx1_ASAP7_75t_SL g1992 ( 
.A(n_1792),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1855),
.Y(n_1993)
);

AOI22x1_ASAP7_75t_L g1994 ( 
.A1(n_1846),
.A2(n_461),
.B1(n_462),
.B2(n_460),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1831),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1869),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1875),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_L g1998 ( 
.A(n_1851),
.B(n_8),
.Y(n_1998)
);

INVx4_ASAP7_75t_L g1999 ( 
.A(n_1835),
.Y(n_1999)
);

NOR2xp33_ASAP7_75t_L g2000 ( 
.A(n_1825),
.B(n_9),
.Y(n_2000)
);

NOR2xp33_ASAP7_75t_L g2001 ( 
.A(n_1781),
.B(n_11),
.Y(n_2001)
);

CKINVDCx20_ASAP7_75t_R g2002 ( 
.A(n_1828),
.Y(n_2002)
);

CKINVDCx5p33_ASAP7_75t_R g2003 ( 
.A(n_1789),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1843),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1784),
.Y(n_2005)
);

AOI21xp5_ASAP7_75t_L g2006 ( 
.A1(n_1832),
.A2(n_466),
.B(n_465),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1774),
.Y(n_2007)
);

INVx2_ASAP7_75t_L g2008 ( 
.A(n_1819),
.Y(n_2008)
);

NOR2xp33_ASAP7_75t_L g2009 ( 
.A(n_1884),
.B(n_12),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_L g2010 ( 
.A(n_1822),
.B(n_1880),
.Y(n_2010)
);

HB1xp67_ASAP7_75t_L g2011 ( 
.A(n_1863),
.Y(n_2011)
);

NAND3xp33_ASAP7_75t_L g2012 ( 
.A(n_1780),
.B(n_12),
.C(n_13),
.Y(n_2012)
);

CKINVDCx5p33_ASAP7_75t_R g2013 ( 
.A(n_1844),
.Y(n_2013)
);

AO31x2_ASAP7_75t_L g2014 ( 
.A1(n_1967),
.A2(n_469),
.A3(n_470),
.B(n_467),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1907),
.Y(n_2015)
);

AOI21x1_ASAP7_75t_L g2016 ( 
.A1(n_1922),
.A2(n_473),
.B(n_471),
.Y(n_2016)
);

AOI21xp5_ASAP7_75t_L g2017 ( 
.A1(n_1924),
.A2(n_905),
.B(n_904),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_SL g2018 ( 
.A(n_1894),
.B(n_1953),
.Y(n_2018)
);

OAI21xp5_ASAP7_75t_L g2019 ( 
.A1(n_1900),
.A2(n_1906),
.B(n_1893),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_L g2020 ( 
.A(n_1917),
.B(n_14),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_L g2021 ( 
.A(n_1921),
.B(n_1934),
.Y(n_2021)
);

OAI21xp5_ASAP7_75t_L g2022 ( 
.A1(n_1929),
.A2(n_15),
.B(n_16),
.Y(n_2022)
);

OAI21xp5_ASAP7_75t_L g2023 ( 
.A1(n_1933),
.A2(n_1951),
.B(n_1947),
.Y(n_2023)
);

OAI22xp5_ASAP7_75t_L g2024 ( 
.A1(n_1946),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.Y(n_2024)
);

OAI21x1_ASAP7_75t_L g2025 ( 
.A1(n_1994),
.A2(n_475),
.B(n_474),
.Y(n_2025)
);

AOI21xp5_ASAP7_75t_SL g2026 ( 
.A1(n_1937),
.A2(n_478),
.B(n_476),
.Y(n_2026)
);

AOI21xp5_ASAP7_75t_L g2027 ( 
.A1(n_1938),
.A2(n_894),
.B(n_892),
.Y(n_2027)
);

OAI21x1_ASAP7_75t_L g2028 ( 
.A1(n_1993),
.A2(n_483),
.B(n_479),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1916),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_L g2030 ( 
.A(n_1976),
.B(n_17),
.Y(n_2030)
);

AO31x2_ASAP7_75t_L g2031 ( 
.A1(n_1896),
.A2(n_485),
.A3(n_486),
.B(n_484),
.Y(n_2031)
);

OAI22xp5_ASAP7_75t_L g2032 ( 
.A1(n_1957),
.A2(n_20),
.B1(n_18),
.B2(n_19),
.Y(n_2032)
);

A2O1A1Ixp33_ASAP7_75t_L g2033 ( 
.A1(n_1931),
.A2(n_21),
.B(n_19),
.C(n_20),
.Y(n_2033)
);

OAI21x1_ASAP7_75t_L g2034 ( 
.A1(n_2006),
.A2(n_489),
.B(n_487),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_L g2035 ( 
.A(n_1927),
.B(n_21),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_1919),
.Y(n_2036)
);

AO32x2_ASAP7_75t_L g2037 ( 
.A1(n_1990),
.A2(n_24),
.A3(n_22),
.B1(n_23),
.B2(n_25),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_L g2038 ( 
.A(n_2011),
.B(n_22),
.Y(n_2038)
);

NAND2xp5_ASAP7_75t_SL g2039 ( 
.A(n_1887),
.B(n_23),
.Y(n_2039)
);

AOI21xp5_ASAP7_75t_L g2040 ( 
.A1(n_1974),
.A2(n_895),
.B(n_891),
.Y(n_2040)
);

AOI221xp5_ASAP7_75t_SL g2041 ( 
.A1(n_2009),
.A2(n_27),
.B1(n_25),
.B2(n_26),
.C(n_28),
.Y(n_2041)
);

AOI21xp5_ASAP7_75t_L g2042 ( 
.A1(n_1890),
.A2(n_898),
.B(n_896),
.Y(n_2042)
);

AO21x2_ASAP7_75t_L g2043 ( 
.A1(n_1982),
.A2(n_492),
.B(n_491),
.Y(n_2043)
);

HB1xp67_ASAP7_75t_L g2044 ( 
.A(n_1892),
.Y(n_2044)
);

OAI21x1_ASAP7_75t_L g2045 ( 
.A1(n_1926),
.A2(n_497),
.B(n_494),
.Y(n_2045)
);

A2O1A1Ixp33_ASAP7_75t_L g2046 ( 
.A1(n_2007),
.A2(n_28),
.B(n_26),
.C(n_27),
.Y(n_2046)
);

NOR2xp33_ASAP7_75t_L g2047 ( 
.A(n_1895),
.B(n_498),
.Y(n_2047)
);

O2A1O1Ixp5_ASAP7_75t_L g2048 ( 
.A1(n_1998),
.A2(n_32),
.B(n_30),
.C(n_31),
.Y(n_2048)
);

NAND2xp5_ASAP7_75t_SL g2049 ( 
.A(n_1965),
.B(n_30),
.Y(n_2049)
);

OAI21xp33_ASAP7_75t_L g2050 ( 
.A1(n_1986),
.A2(n_31),
.B(n_34),
.Y(n_2050)
);

OAI21x1_ASAP7_75t_SL g2051 ( 
.A1(n_1932),
.A2(n_34),
.B(n_35),
.Y(n_2051)
);

NAND2xp5_ASAP7_75t_L g2052 ( 
.A(n_1903),
.B(n_2008),
.Y(n_2052)
);

AOI221x1_ASAP7_75t_L g2053 ( 
.A1(n_2012),
.A2(n_37),
.B1(n_35),
.B2(n_36),
.C(n_38),
.Y(n_2053)
);

OAI21x1_ASAP7_75t_L g2054 ( 
.A1(n_1989),
.A2(n_500),
.B(n_499),
.Y(n_2054)
);

OAI21x1_ASAP7_75t_L g2055 ( 
.A1(n_2004),
.A2(n_503),
.B(n_502),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1920),
.Y(n_2056)
);

INVxp67_ASAP7_75t_L g2057 ( 
.A(n_1915),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_L g2058 ( 
.A(n_1992),
.B(n_36),
.Y(n_2058)
);

NOR2xp33_ASAP7_75t_L g2059 ( 
.A(n_1914),
.B(n_505),
.Y(n_2059)
);

OAI21x1_ASAP7_75t_L g2060 ( 
.A1(n_1996),
.A2(n_507),
.B(n_506),
.Y(n_2060)
);

AOI21xp5_ASAP7_75t_L g2061 ( 
.A1(n_1960),
.A2(n_909),
.B(n_908),
.Y(n_2061)
);

A2O1A1Ixp33_ASAP7_75t_L g2062 ( 
.A1(n_2000),
.A2(n_2001),
.B(n_2010),
.C(n_1995),
.Y(n_2062)
);

AOI21xp5_ASAP7_75t_L g2063 ( 
.A1(n_1891),
.A2(n_910),
.B(n_511),
.Y(n_2063)
);

A2O1A1Ixp33_ASAP7_75t_L g2064 ( 
.A1(n_1977),
.A2(n_39),
.B(n_37),
.C(n_38),
.Y(n_2064)
);

INVx3_ASAP7_75t_L g2065 ( 
.A(n_1904),
.Y(n_2065)
);

OAI21x1_ASAP7_75t_SL g2066 ( 
.A1(n_1984),
.A2(n_40),
.B(n_41),
.Y(n_2066)
);

AND2x2_ASAP7_75t_L g2067 ( 
.A(n_1972),
.B(n_40),
.Y(n_2067)
);

BUFx3_ASAP7_75t_L g2068 ( 
.A(n_1961),
.Y(n_2068)
);

CKINVDCx5p33_ASAP7_75t_R g2069 ( 
.A(n_2013),
.Y(n_2069)
);

BUFx2_ASAP7_75t_L g2070 ( 
.A(n_1978),
.Y(n_2070)
);

AND2x2_ASAP7_75t_L g2071 ( 
.A(n_2005),
.B(n_42),
.Y(n_2071)
);

AOI21x1_ASAP7_75t_L g2072 ( 
.A1(n_1944),
.A2(n_1889),
.B(n_1888),
.Y(n_2072)
);

AND2x2_ASAP7_75t_L g2073 ( 
.A(n_1899),
.B(n_42),
.Y(n_2073)
);

NAND2xp33_ASAP7_75t_SL g2074 ( 
.A(n_1901),
.B(n_43),
.Y(n_2074)
);

NAND2xp5_ASAP7_75t_SL g2075 ( 
.A(n_1969),
.B(n_43),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_1898),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_SL g2077 ( 
.A(n_1969),
.B(n_44),
.Y(n_2077)
);

NAND2xp5_ASAP7_75t_SL g2078 ( 
.A(n_1949),
.B(n_45),
.Y(n_2078)
);

OAI21x1_ASAP7_75t_L g2079 ( 
.A1(n_1963),
.A2(n_513),
.B(n_508),
.Y(n_2079)
);

OAI21x1_ASAP7_75t_L g2080 ( 
.A1(n_1930),
.A2(n_517),
.B(n_515),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_L g2081 ( 
.A(n_1955),
.B(n_45),
.Y(n_2081)
);

NOR2x1_ASAP7_75t_L g2082 ( 
.A(n_1954),
.B(n_519),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_1908),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_1936),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_L g2085 ( 
.A(n_1940),
.B(n_46),
.Y(n_2085)
);

AND2x2_ASAP7_75t_L g2086 ( 
.A(n_1958),
.B(n_46),
.Y(n_2086)
);

INVx4_ASAP7_75t_L g2087 ( 
.A(n_1961),
.Y(n_2087)
);

AOI21xp5_ASAP7_75t_SL g2088 ( 
.A1(n_1973),
.A2(n_523),
.B(n_520),
.Y(n_2088)
);

AOI31xp67_ASAP7_75t_L g2089 ( 
.A1(n_1902),
.A2(n_525),
.A3(n_526),
.B(n_524),
.Y(n_2089)
);

OAI21x1_ASAP7_75t_L g2090 ( 
.A1(n_1945),
.A2(n_532),
.B(n_531),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_1950),
.Y(n_2091)
);

BUFx6f_ASAP7_75t_L g2092 ( 
.A(n_1923),
.Y(n_2092)
);

OAI21xp5_ASAP7_75t_L g2093 ( 
.A1(n_1975),
.A2(n_1987),
.B(n_1942),
.Y(n_2093)
);

NAND2xp5_ASAP7_75t_L g2094 ( 
.A(n_2021),
.B(n_1962),
.Y(n_2094)
);

OR2x6_ASAP7_75t_SL g2095 ( 
.A(n_2038),
.B(n_2003),
.Y(n_2095)
);

AO21x2_ASAP7_75t_L g2096 ( 
.A1(n_2017),
.A2(n_1988),
.B(n_1997),
.Y(n_2096)
);

CKINVDCx11_ASAP7_75t_R g2097 ( 
.A(n_2092),
.Y(n_2097)
);

INVx2_ASAP7_75t_L g2098 ( 
.A(n_2015),
.Y(n_2098)
);

HB1xp67_ASAP7_75t_L g2099 ( 
.A(n_2044),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_L g2100 ( 
.A(n_2018),
.B(n_2023),
.Y(n_2100)
);

INVx2_ASAP7_75t_L g2101 ( 
.A(n_2029),
.Y(n_2101)
);

HB1xp67_ASAP7_75t_L g2102 ( 
.A(n_2057),
.Y(n_2102)
);

NOR3xp33_ASAP7_75t_L g2103 ( 
.A(n_2050),
.B(n_1999),
.C(n_1983),
.Y(n_2103)
);

AND2x4_ASAP7_75t_L g2104 ( 
.A(n_2070),
.B(n_1966),
.Y(n_2104)
);

INVx1_ASAP7_75t_SL g2105 ( 
.A(n_2052),
.Y(n_2105)
);

AOI22xp5_ASAP7_75t_L g2106 ( 
.A1(n_2059),
.A2(n_2002),
.B1(n_1911),
.B2(n_1939),
.Y(n_2106)
);

AND2x2_ASAP7_75t_L g2107 ( 
.A(n_2019),
.B(n_1909),
.Y(n_2107)
);

NAND2xp5_ASAP7_75t_L g2108 ( 
.A(n_2062),
.B(n_1964),
.Y(n_2108)
);

BUFx6f_ASAP7_75t_SL g2109 ( 
.A(n_2092),
.Y(n_2109)
);

INVx3_ASAP7_75t_L g2110 ( 
.A(n_2087),
.Y(n_2110)
);

INVx3_ASAP7_75t_L g2111 ( 
.A(n_2068),
.Y(n_2111)
);

AND2x6_ASAP7_75t_L g2112 ( 
.A(n_2082),
.B(n_1971),
.Y(n_2112)
);

INVx5_ASAP7_75t_L g2113 ( 
.A(n_2065),
.Y(n_2113)
);

AOI21xp5_ASAP7_75t_L g2114 ( 
.A1(n_2026),
.A2(n_1941),
.B(n_1918),
.Y(n_2114)
);

AOI22xp5_ASAP7_75t_L g2115 ( 
.A1(n_2047),
.A2(n_1981),
.B1(n_1985),
.B2(n_1943),
.Y(n_2115)
);

INVx2_ASAP7_75t_L g2116 ( 
.A(n_2036),
.Y(n_2116)
);

BUFx2_ASAP7_75t_L g2117 ( 
.A(n_2056),
.Y(n_2117)
);

INVx1_ASAP7_75t_SL g2118 ( 
.A(n_2069),
.Y(n_2118)
);

NOR2xp67_ASAP7_75t_L g2119 ( 
.A(n_2020),
.B(n_1970),
.Y(n_2119)
);

INVx2_ASAP7_75t_L g2120 ( 
.A(n_2084),
.Y(n_2120)
);

BUFx2_ASAP7_75t_L g2121 ( 
.A(n_2076),
.Y(n_2121)
);

INVx2_ASAP7_75t_L g2122 ( 
.A(n_2072),
.Y(n_2122)
);

INVx2_ASAP7_75t_L g2123 ( 
.A(n_2091),
.Y(n_2123)
);

AND2x4_ASAP7_75t_L g2124 ( 
.A(n_2083),
.B(n_1910),
.Y(n_2124)
);

INVx2_ASAP7_75t_L g2125 ( 
.A(n_2086),
.Y(n_2125)
);

AND2x2_ASAP7_75t_L g2126 ( 
.A(n_2073),
.B(n_1909),
.Y(n_2126)
);

INVx3_ASAP7_75t_L g2127 ( 
.A(n_2016),
.Y(n_2127)
);

INVx2_ASAP7_75t_SL g2128 ( 
.A(n_2067),
.Y(n_2128)
);

NAND2xp33_ASAP7_75t_L g2129 ( 
.A(n_2064),
.B(n_1913),
.Y(n_2129)
);

AOI221xp5_ASAP7_75t_L g2130 ( 
.A1(n_2024),
.A2(n_1991),
.B1(n_1968),
.B2(n_1897),
.C(n_1979),
.Y(n_2130)
);

AOI21xp5_ASAP7_75t_L g2131 ( 
.A1(n_2040),
.A2(n_1941),
.B(n_1918),
.Y(n_2131)
);

AOI21xp5_ASAP7_75t_L g2132 ( 
.A1(n_2022),
.A2(n_1912),
.B(n_1905),
.Y(n_2132)
);

AND2x2_ASAP7_75t_L g2133 ( 
.A(n_2093),
.B(n_1980),
.Y(n_2133)
);

OR2x2_ASAP7_75t_L g2134 ( 
.A(n_2039),
.B(n_1959),
.Y(n_2134)
);

BUFx6f_ASAP7_75t_L g2135 ( 
.A(n_2081),
.Y(n_2135)
);

INVx2_ASAP7_75t_SL g2136 ( 
.A(n_2058),
.Y(n_2136)
);

INVx2_ASAP7_75t_L g2137 ( 
.A(n_2085),
.Y(n_2137)
);

BUFx2_ASAP7_75t_L g2138 ( 
.A(n_2030),
.Y(n_2138)
);

OAI22xp5_ASAP7_75t_L g2139 ( 
.A1(n_2035),
.A2(n_1948),
.B1(n_1952),
.B2(n_1913),
.Y(n_2139)
);

BUFx4_ASAP7_75t_SL g2140 ( 
.A(n_2074),
.Y(n_2140)
);

INVx2_ASAP7_75t_L g2141 ( 
.A(n_2043),
.Y(n_2141)
);

NAND2x1p5_ASAP7_75t_L g2142 ( 
.A(n_2105),
.B(n_2113),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_2121),
.Y(n_2143)
);

NAND2xp5_ASAP7_75t_L g2144 ( 
.A(n_2100),
.B(n_2041),
.Y(n_2144)
);

OR2x2_ASAP7_75t_L g2145 ( 
.A(n_2099),
.B(n_2031),
.Y(n_2145)
);

AOI21xp5_ASAP7_75t_SL g2146 ( 
.A1(n_2114),
.A2(n_2033),
.B(n_2046),
.Y(n_2146)
);

NAND2xp5_ASAP7_75t_L g2147 ( 
.A(n_2138),
.B(n_2071),
.Y(n_2147)
);

NAND2xp5_ASAP7_75t_L g2148 ( 
.A(n_2137),
.B(n_2053),
.Y(n_2148)
);

AOI21xp5_ASAP7_75t_L g2149 ( 
.A1(n_2132),
.A2(n_2108),
.B(n_2131),
.Y(n_2149)
);

CKINVDCx5p33_ASAP7_75t_R g2150 ( 
.A(n_2097),
.Y(n_2150)
);

NAND2xp5_ASAP7_75t_L g2151 ( 
.A(n_2117),
.B(n_2078),
.Y(n_2151)
);

AND2x2_ASAP7_75t_L g2152 ( 
.A(n_2107),
.B(n_2031),
.Y(n_2152)
);

A2O1A1Ixp33_ASAP7_75t_SL g2153 ( 
.A1(n_2141),
.A2(n_2127),
.B(n_2103),
.C(n_2032),
.Y(n_2153)
);

CKINVDCx5p33_ASAP7_75t_R g2154 ( 
.A(n_2109),
.Y(n_2154)
);

AND2x2_ASAP7_75t_L g2155 ( 
.A(n_2126),
.B(n_2045),
.Y(n_2155)
);

A2O1A1Ixp33_ASAP7_75t_L g2156 ( 
.A1(n_2129),
.A2(n_2048),
.B(n_2049),
.C(n_2042),
.Y(n_2156)
);

AND2x2_ASAP7_75t_L g2157 ( 
.A(n_2125),
.B(n_2075),
.Y(n_2157)
);

INVx2_ASAP7_75t_L g2158 ( 
.A(n_2098),
.Y(n_2158)
);

NOR2xp67_ASAP7_75t_L g2159 ( 
.A(n_2113),
.B(n_2027),
.Y(n_2159)
);

CKINVDCx5p33_ASAP7_75t_R g2160 ( 
.A(n_2118),
.Y(n_2160)
);

AND2x2_ASAP7_75t_L g2161 ( 
.A(n_2133),
.B(n_2077),
.Y(n_2161)
);

CKINVDCx5p33_ASAP7_75t_R g2162 ( 
.A(n_2104),
.Y(n_2162)
);

NOR2x1_ASAP7_75t_SL g2163 ( 
.A(n_2096),
.B(n_2089),
.Y(n_2163)
);

NAND2xp5_ASAP7_75t_L g2164 ( 
.A(n_2102),
.B(n_2066),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_2122),
.Y(n_2165)
);

O2A1O1Ixp5_ASAP7_75t_L g2166 ( 
.A1(n_2139),
.A2(n_2061),
.B(n_2063),
.C(n_2037),
.Y(n_2166)
);

NOR2xp33_ASAP7_75t_L g2167 ( 
.A(n_2115),
.B(n_1925),
.Y(n_2167)
);

NAND2xp5_ASAP7_75t_L g2168 ( 
.A(n_2123),
.B(n_2051),
.Y(n_2168)
);

NAND2xp5_ASAP7_75t_L g2169 ( 
.A(n_2101),
.B(n_2014),
.Y(n_2169)
);

CKINVDCx5p33_ASAP7_75t_R g2170 ( 
.A(n_2140),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_2116),
.Y(n_2171)
);

AOI21xp5_ASAP7_75t_L g2172 ( 
.A1(n_2094),
.A2(n_2034),
.B(n_2025),
.Y(n_2172)
);

AOI21xp5_ASAP7_75t_L g2173 ( 
.A1(n_2119),
.A2(n_2088),
.B(n_2028),
.Y(n_2173)
);

AOI21xp5_ASAP7_75t_L g2174 ( 
.A1(n_2106),
.A2(n_2055),
.B(n_2054),
.Y(n_2174)
);

HB1xp67_ASAP7_75t_L g2175 ( 
.A(n_2120),
.Y(n_2175)
);

HB1xp67_ASAP7_75t_L g2176 ( 
.A(n_2135),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_2135),
.Y(n_2177)
);

OR2x2_ASAP7_75t_L g2178 ( 
.A(n_2136),
.B(n_2014),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_2134),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_2124),
.Y(n_2180)
);

AND2x2_ASAP7_75t_L g2181 ( 
.A(n_2128),
.B(n_2037),
.Y(n_2181)
);

NOR2xp33_ASAP7_75t_L g2182 ( 
.A(n_2095),
.B(n_1956),
.Y(n_2182)
);

INVx2_ASAP7_75t_SL g2183 ( 
.A(n_2111),
.Y(n_2183)
);

AOI21xp5_ASAP7_75t_SL g2184 ( 
.A1(n_2130),
.A2(n_2112),
.B(n_1935),
.Y(n_2184)
);

OR2x2_ASAP7_75t_L g2185 ( 
.A(n_2110),
.B(n_2079),
.Y(n_2185)
);

INVx2_ASAP7_75t_L g2186 ( 
.A(n_2112),
.Y(n_2186)
);

OAI21xp33_ASAP7_75t_L g2187 ( 
.A1(n_2112),
.A2(n_2060),
.B(n_2090),
.Y(n_2187)
);

AND2x2_ASAP7_75t_L g2188 ( 
.A(n_2107),
.B(n_2080),
.Y(n_2188)
);

A2O1A1Ixp33_ASAP7_75t_L g2189 ( 
.A1(n_2131),
.A2(n_1928),
.B(n_1956),
.C(n_49),
.Y(n_2189)
);

OA21x2_ASAP7_75t_L g2190 ( 
.A1(n_2141),
.A2(n_47),
.B(n_48),
.Y(n_2190)
);

NAND2xp5_ASAP7_75t_L g2191 ( 
.A(n_2105),
.B(n_48),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_2121),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_2175),
.Y(n_2193)
);

AO21x2_ASAP7_75t_L g2194 ( 
.A1(n_2163),
.A2(n_2149),
.B(n_2148),
.Y(n_2194)
);

OAI21x1_ASAP7_75t_L g2195 ( 
.A1(n_2172),
.A2(n_2174),
.B(n_2173),
.Y(n_2195)
);

AOI22xp33_ASAP7_75t_L g2196 ( 
.A1(n_2155),
.A2(n_51),
.B1(n_49),
.B2(n_50),
.Y(n_2196)
);

AOI21x1_ASAP7_75t_L g2197 ( 
.A1(n_2159),
.A2(n_50),
.B(n_51),
.Y(n_2197)
);

AO21x2_ASAP7_75t_L g2198 ( 
.A1(n_2169),
.A2(n_52),
.B(n_53),
.Y(n_2198)
);

INVx2_ASAP7_75t_L g2199 ( 
.A(n_2158),
.Y(n_2199)
);

INVx2_ASAP7_75t_L g2200 ( 
.A(n_2171),
.Y(n_2200)
);

OAI222xp33_ASAP7_75t_L g2201 ( 
.A1(n_2144),
.A2(n_54),
.B1(n_57),
.B2(n_52),
.C1(n_53),
.C2(n_55),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_2165),
.Y(n_2202)
);

INVx2_ASAP7_75t_L g2203 ( 
.A(n_2143),
.Y(n_2203)
);

AND2x2_ASAP7_75t_L g2204 ( 
.A(n_2179),
.B(n_54),
.Y(n_2204)
);

NAND2xp5_ASAP7_75t_L g2205 ( 
.A(n_2192),
.B(n_55),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_2145),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_2178),
.Y(n_2207)
);

INVx2_ASAP7_75t_L g2208 ( 
.A(n_2177),
.Y(n_2208)
);

INVx2_ASAP7_75t_L g2209 ( 
.A(n_2142),
.Y(n_2209)
);

INVx2_ASAP7_75t_L g2210 ( 
.A(n_2176),
.Y(n_2210)
);

AO21x1_ASAP7_75t_SL g2211 ( 
.A1(n_2187),
.A2(n_57),
.B(n_58),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_2190),
.Y(n_2212)
);

INVx2_ASAP7_75t_L g2213 ( 
.A(n_2164),
.Y(n_2213)
);

AND2x2_ASAP7_75t_L g2214 ( 
.A(n_2152),
.B(n_58),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_2190),
.Y(n_2215)
);

INVx2_ASAP7_75t_L g2216 ( 
.A(n_2180),
.Y(n_2216)
);

OAI21x1_ASAP7_75t_L g2217 ( 
.A1(n_2166),
.A2(n_537),
.B(n_534),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_2181),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_2185),
.Y(n_2219)
);

BUFx3_ASAP7_75t_L g2220 ( 
.A(n_2162),
.Y(n_2220)
);

INVx3_ASAP7_75t_L g2221 ( 
.A(n_2183),
.Y(n_2221)
);

AND2x4_ASAP7_75t_SL g2222 ( 
.A(n_2186),
.B(n_538),
.Y(n_2222)
);

INVx2_ASAP7_75t_L g2223 ( 
.A(n_2188),
.Y(n_2223)
);

OR2x2_ASAP7_75t_L g2224 ( 
.A(n_2147),
.B(n_59),
.Y(n_2224)
);

INVx2_ASAP7_75t_L g2225 ( 
.A(n_2168),
.Y(n_2225)
);

NAND2xp5_ASAP7_75t_L g2226 ( 
.A(n_2151),
.B(n_60),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_2157),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_2191),
.Y(n_2228)
);

INVx2_ASAP7_75t_L g2229 ( 
.A(n_2161),
.Y(n_2229)
);

AND2x2_ASAP7_75t_L g2230 ( 
.A(n_2182),
.B(n_61),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_2167),
.Y(n_2231)
);

OA21x2_ASAP7_75t_L g2232 ( 
.A1(n_2189),
.A2(n_70),
.B(n_62),
.Y(n_2232)
);

AND2x2_ASAP7_75t_L g2233 ( 
.A(n_2160),
.B(n_62),
.Y(n_2233)
);

INVx2_ASAP7_75t_L g2234 ( 
.A(n_2184),
.Y(n_2234)
);

HB1xp67_ASAP7_75t_L g2235 ( 
.A(n_2156),
.Y(n_2235)
);

BUFx2_ASAP7_75t_L g2236 ( 
.A(n_2150),
.Y(n_2236)
);

INVx2_ASAP7_75t_L g2237 ( 
.A(n_2146),
.Y(n_2237)
);

OAI21xp33_ASAP7_75t_SL g2238 ( 
.A1(n_2153),
.A2(n_63),
.B(n_64),
.Y(n_2238)
);

BUFx3_ASAP7_75t_L g2239 ( 
.A(n_2154),
.Y(n_2239)
);

AND2x2_ASAP7_75t_L g2240 ( 
.A(n_2170),
.B(n_63),
.Y(n_2240)
);

BUFx6f_ASAP7_75t_L g2241 ( 
.A(n_2183),
.Y(n_2241)
);

BUFx3_ASAP7_75t_L g2242 ( 
.A(n_2162),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_2175),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_2175),
.Y(n_2244)
);

INVx2_ASAP7_75t_L g2245 ( 
.A(n_2158),
.Y(n_2245)
);

AND2x2_ASAP7_75t_L g2246 ( 
.A(n_2179),
.B(n_65),
.Y(n_2246)
);

INVx2_ASAP7_75t_L g2247 ( 
.A(n_2158),
.Y(n_2247)
);

INVx1_ASAP7_75t_L g2248 ( 
.A(n_2175),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_2175),
.Y(n_2249)
);

BUFx6f_ASAP7_75t_L g2250 ( 
.A(n_2183),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_2175),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_2175),
.Y(n_2252)
);

INVx3_ASAP7_75t_L g2253 ( 
.A(n_2183),
.Y(n_2253)
);

INVx2_ASAP7_75t_L g2254 ( 
.A(n_2158),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_2175),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_2175),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_2175),
.Y(n_2257)
);

INVx2_ASAP7_75t_L g2258 ( 
.A(n_2158),
.Y(n_2258)
);

AND2x2_ASAP7_75t_L g2259 ( 
.A(n_2179),
.B(n_65),
.Y(n_2259)
);

OA21x2_ASAP7_75t_L g2260 ( 
.A1(n_2149),
.A2(n_74),
.B(n_66),
.Y(n_2260)
);

OAI21xp5_ASAP7_75t_L g2261 ( 
.A1(n_2149),
.A2(n_67),
.B(n_68),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_2175),
.Y(n_2262)
);

INVx2_ASAP7_75t_SL g2263 ( 
.A(n_2183),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_2175),
.Y(n_2264)
);

INVx2_ASAP7_75t_L g2265 ( 
.A(n_2158),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_2175),
.Y(n_2266)
);

INVx2_ASAP7_75t_L g2267 ( 
.A(n_2158),
.Y(n_2267)
);

OAI21xp5_ASAP7_75t_SL g2268 ( 
.A1(n_2149),
.A2(n_71),
.B(n_70),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_2207),
.Y(n_2269)
);

BUFx2_ASAP7_75t_L g2270 ( 
.A(n_2209),
.Y(n_2270)
);

HB1xp67_ASAP7_75t_L g2271 ( 
.A(n_2206),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_2200),
.Y(n_2272)
);

INVx2_ASAP7_75t_SL g2273 ( 
.A(n_2241),
.Y(n_2273)
);

INVx2_ASAP7_75t_L g2274 ( 
.A(n_2225),
.Y(n_2274)
);

INVxp67_ASAP7_75t_SL g2275 ( 
.A(n_2213),
.Y(n_2275)
);

AND2x2_ASAP7_75t_L g2276 ( 
.A(n_2229),
.B(n_69),
.Y(n_2276)
);

HB1xp67_ASAP7_75t_L g2277 ( 
.A(n_2219),
.Y(n_2277)
);

INVx2_ASAP7_75t_L g2278 ( 
.A(n_2208),
.Y(n_2278)
);

INVx2_ASAP7_75t_L g2279 ( 
.A(n_2193),
.Y(n_2279)
);

OR2x2_ASAP7_75t_L g2280 ( 
.A(n_2243),
.B(n_71),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_2244),
.Y(n_2281)
);

OR2x2_ASAP7_75t_L g2282 ( 
.A(n_2248),
.B(n_72),
.Y(n_2282)
);

NAND2xp5_ASAP7_75t_L g2283 ( 
.A(n_2249),
.B(n_72),
.Y(n_2283)
);

INVx1_ASAP7_75t_L g2284 ( 
.A(n_2251),
.Y(n_2284)
);

AND2x2_ASAP7_75t_L g2285 ( 
.A(n_2210),
.B(n_73),
.Y(n_2285)
);

BUFx3_ASAP7_75t_L g2286 ( 
.A(n_2236),
.Y(n_2286)
);

BUFx2_ASAP7_75t_L g2287 ( 
.A(n_2223),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_2252),
.Y(n_2288)
);

INVx2_ASAP7_75t_L g2289 ( 
.A(n_2255),
.Y(n_2289)
);

NAND2xp5_ASAP7_75t_L g2290 ( 
.A(n_2256),
.B(n_73),
.Y(n_2290)
);

AND2x4_ASAP7_75t_L g2291 ( 
.A(n_2227),
.B(n_74),
.Y(n_2291)
);

HB1xp67_ASAP7_75t_L g2292 ( 
.A(n_2257),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_2262),
.Y(n_2293)
);

INVx2_ASAP7_75t_L g2294 ( 
.A(n_2264),
.Y(n_2294)
);

INVx2_ASAP7_75t_L g2295 ( 
.A(n_2266),
.Y(n_2295)
);

INVx1_ASAP7_75t_L g2296 ( 
.A(n_2202),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_2199),
.Y(n_2297)
);

NAND2xp5_ASAP7_75t_L g2298 ( 
.A(n_2203),
.B(n_2231),
.Y(n_2298)
);

HB1xp67_ASAP7_75t_L g2299 ( 
.A(n_2212),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_2245),
.Y(n_2300)
);

INVx2_ASAP7_75t_L g2301 ( 
.A(n_2247),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_2254),
.Y(n_2302)
);

INVxp67_ASAP7_75t_L g2303 ( 
.A(n_2235),
.Y(n_2303)
);

AND2x2_ASAP7_75t_L g2304 ( 
.A(n_2218),
.B(n_75),
.Y(n_2304)
);

BUFx2_ASAP7_75t_SL g2305 ( 
.A(n_2239),
.Y(n_2305)
);

INVx1_ASAP7_75t_L g2306 ( 
.A(n_2258),
.Y(n_2306)
);

HB1xp67_ASAP7_75t_L g2307 ( 
.A(n_2215),
.Y(n_2307)
);

OR2x2_ASAP7_75t_L g2308 ( 
.A(n_2216),
.B(n_76),
.Y(n_2308)
);

INVx2_ASAP7_75t_L g2309 ( 
.A(n_2265),
.Y(n_2309)
);

INVx2_ASAP7_75t_L g2310 ( 
.A(n_2267),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_2194),
.Y(n_2311)
);

INVx2_ASAP7_75t_L g2312 ( 
.A(n_2263),
.Y(n_2312)
);

NAND2xp5_ASAP7_75t_L g2313 ( 
.A(n_2228),
.B(n_77),
.Y(n_2313)
);

AND2x2_ASAP7_75t_L g2314 ( 
.A(n_2221),
.B(n_77),
.Y(n_2314)
);

AND2x2_ASAP7_75t_L g2315 ( 
.A(n_2253),
.B(n_78),
.Y(n_2315)
);

AND2x2_ASAP7_75t_L g2316 ( 
.A(n_2241),
.B(n_79),
.Y(n_2316)
);

INVx2_ASAP7_75t_L g2317 ( 
.A(n_2250),
.Y(n_2317)
);

AO31x2_ASAP7_75t_L g2318 ( 
.A1(n_2234),
.A2(n_81),
.A3(n_79),
.B(n_80),
.Y(n_2318)
);

AND2x2_ASAP7_75t_L g2319 ( 
.A(n_2250),
.B(n_80),
.Y(n_2319)
);

HB1xp67_ASAP7_75t_L g2320 ( 
.A(n_2198),
.Y(n_2320)
);

OR2x2_ASAP7_75t_L g2321 ( 
.A(n_2224),
.B(n_81),
.Y(n_2321)
);

INVx1_ASAP7_75t_L g2322 ( 
.A(n_2205),
.Y(n_2322)
);

INVx2_ASAP7_75t_L g2323 ( 
.A(n_2195),
.Y(n_2323)
);

HB1xp67_ASAP7_75t_L g2324 ( 
.A(n_2224),
.Y(n_2324)
);

INVx2_ASAP7_75t_L g2325 ( 
.A(n_2204),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_L g2326 ( 
.A(n_2214),
.B(n_82),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_2246),
.Y(n_2327)
);

INVx2_ASAP7_75t_L g2328 ( 
.A(n_2259),
.Y(n_2328)
);

AND2x2_ASAP7_75t_L g2329 ( 
.A(n_2236),
.B(n_82),
.Y(n_2329)
);

AND2x2_ASAP7_75t_L g2330 ( 
.A(n_2220),
.B(n_83),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_2260),
.Y(n_2331)
);

INVx2_ASAP7_75t_L g2332 ( 
.A(n_2237),
.Y(n_2332)
);

OAI22xp5_ASAP7_75t_L g2333 ( 
.A1(n_2268),
.A2(n_85),
.B1(n_83),
.B2(n_84),
.Y(n_2333)
);

AND2x4_ASAP7_75t_SL g2334 ( 
.A(n_2233),
.B(n_906),
.Y(n_2334)
);

INVx2_ASAP7_75t_L g2335 ( 
.A(n_2217),
.Y(n_2335)
);

OR2x2_ASAP7_75t_L g2336 ( 
.A(n_2226),
.B(n_84),
.Y(n_2336)
);

NOR2x1p5_ASAP7_75t_L g2337 ( 
.A(n_2242),
.B(n_85),
.Y(n_2337)
);

INVx2_ASAP7_75t_L g2338 ( 
.A(n_2197),
.Y(n_2338)
);

AND2x2_ASAP7_75t_L g2339 ( 
.A(n_2230),
.B(n_86),
.Y(n_2339)
);

INVx1_ASAP7_75t_L g2340 ( 
.A(n_2232),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_2261),
.Y(n_2341)
);

INVx2_ASAP7_75t_L g2342 ( 
.A(n_2240),
.Y(n_2342)
);

BUFx6f_ASAP7_75t_L g2343 ( 
.A(n_2211),
.Y(n_2343)
);

AO31x2_ASAP7_75t_L g2344 ( 
.A1(n_2238),
.A2(n_88),
.A3(n_86),
.B(n_87),
.Y(n_2344)
);

AND2x2_ASAP7_75t_L g2345 ( 
.A(n_2222),
.B(n_2196),
.Y(n_2345)
);

INVx2_ASAP7_75t_L g2346 ( 
.A(n_2201),
.Y(n_2346)
);

INVx2_ASAP7_75t_L g2347 ( 
.A(n_2200),
.Y(n_2347)
);

AND2x4_ASAP7_75t_L g2348 ( 
.A(n_2209),
.B(n_87),
.Y(n_2348)
);

INVx2_ASAP7_75t_L g2349 ( 
.A(n_2200),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_2207),
.Y(n_2350)
);

INVx1_ASAP7_75t_L g2351 ( 
.A(n_2207),
.Y(n_2351)
);

INVx2_ASAP7_75t_L g2352 ( 
.A(n_2200),
.Y(n_2352)
);

INVx2_ASAP7_75t_L g2353 ( 
.A(n_2200),
.Y(n_2353)
);

OAI21xp5_ASAP7_75t_SL g2354 ( 
.A1(n_2268),
.A2(n_88),
.B(n_89),
.Y(n_2354)
);

AND2x2_ASAP7_75t_L g2355 ( 
.A(n_2229),
.B(n_89),
.Y(n_2355)
);

AND2x2_ASAP7_75t_L g2356 ( 
.A(n_2229),
.B(n_90),
.Y(n_2356)
);

INVx3_ASAP7_75t_L g2357 ( 
.A(n_2241),
.Y(n_2357)
);

AND2x2_ASAP7_75t_L g2358 ( 
.A(n_2229),
.B(n_90),
.Y(n_2358)
);

OR2x2_ASAP7_75t_L g2359 ( 
.A(n_2219),
.B(n_91),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_2207),
.Y(n_2360)
);

INVx4_ASAP7_75t_L g2361 ( 
.A(n_2236),
.Y(n_2361)
);

INVx2_ASAP7_75t_L g2362 ( 
.A(n_2200),
.Y(n_2362)
);

NAND2xp5_ASAP7_75t_L g2363 ( 
.A(n_2213),
.B(n_92),
.Y(n_2363)
);

BUFx3_ASAP7_75t_L g2364 ( 
.A(n_2236),
.Y(n_2364)
);

AND2x4_ASAP7_75t_L g2365 ( 
.A(n_2209),
.B(n_93),
.Y(n_2365)
);

INVx3_ASAP7_75t_L g2366 ( 
.A(n_2241),
.Y(n_2366)
);

AND2x2_ASAP7_75t_L g2367 ( 
.A(n_2270),
.B(n_93),
.Y(n_2367)
);

INVx1_ASAP7_75t_L g2368 ( 
.A(n_2299),
.Y(n_2368)
);

CKINVDCx20_ASAP7_75t_R g2369 ( 
.A(n_2286),
.Y(n_2369)
);

HB1xp67_ASAP7_75t_L g2370 ( 
.A(n_2307),
.Y(n_2370)
);

HB1xp67_ASAP7_75t_L g2371 ( 
.A(n_2320),
.Y(n_2371)
);

AND2x2_ASAP7_75t_L g2372 ( 
.A(n_2324),
.B(n_94),
.Y(n_2372)
);

CKINVDCx5p33_ASAP7_75t_R g2373 ( 
.A(n_2305),
.Y(n_2373)
);

OR2x6_ASAP7_75t_L g2374 ( 
.A(n_2361),
.B(n_94),
.Y(n_2374)
);

BUFx2_ASAP7_75t_L g2375 ( 
.A(n_2364),
.Y(n_2375)
);

AND2x2_ASAP7_75t_L g2376 ( 
.A(n_2312),
.B(n_95),
.Y(n_2376)
);

INVx2_ASAP7_75t_L g2377 ( 
.A(n_2332),
.Y(n_2377)
);

BUFx2_ASAP7_75t_L g2378 ( 
.A(n_2303),
.Y(n_2378)
);

INVx2_ASAP7_75t_SL g2379 ( 
.A(n_2357),
.Y(n_2379)
);

AND2x2_ASAP7_75t_L g2380 ( 
.A(n_2275),
.B(n_95),
.Y(n_2380)
);

BUFx2_ASAP7_75t_L g2381 ( 
.A(n_2292),
.Y(n_2381)
);

HB1xp67_ASAP7_75t_L g2382 ( 
.A(n_2277),
.Y(n_2382)
);

AOI22xp33_ASAP7_75t_L g2383 ( 
.A1(n_2341),
.A2(n_98),
.B1(n_96),
.B2(n_97),
.Y(n_2383)
);

INVx2_ASAP7_75t_L g2384 ( 
.A(n_2278),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_2271),
.Y(n_2385)
);

INVx2_ASAP7_75t_L g2386 ( 
.A(n_2274),
.Y(n_2386)
);

INVx2_ASAP7_75t_L g2387 ( 
.A(n_2347),
.Y(n_2387)
);

INVx1_ASAP7_75t_L g2388 ( 
.A(n_2296),
.Y(n_2388)
);

INVx2_ASAP7_75t_L g2389 ( 
.A(n_2349),
.Y(n_2389)
);

OR2x2_ASAP7_75t_L g2390 ( 
.A(n_2298),
.B(n_96),
.Y(n_2390)
);

INVx2_ASAP7_75t_L g2391 ( 
.A(n_2352),
.Y(n_2391)
);

NAND2xp5_ASAP7_75t_L g2392 ( 
.A(n_2322),
.B(n_99),
.Y(n_2392)
);

INVx1_ASAP7_75t_SL g2393 ( 
.A(n_2329),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_2269),
.Y(n_2394)
);

INVx1_ASAP7_75t_L g2395 ( 
.A(n_2350),
.Y(n_2395)
);

AND2x4_ASAP7_75t_L g2396 ( 
.A(n_2317),
.B(n_2273),
.Y(n_2396)
);

NAND2xp5_ASAP7_75t_L g2397 ( 
.A(n_2281),
.B(n_100),
.Y(n_2397)
);

AND2x2_ASAP7_75t_L g2398 ( 
.A(n_2287),
.B(n_100),
.Y(n_2398)
);

INVxp67_ASAP7_75t_R g2399 ( 
.A(n_2330),
.Y(n_2399)
);

INVx1_ASAP7_75t_L g2400 ( 
.A(n_2351),
.Y(n_2400)
);

INVx2_ASAP7_75t_L g2401 ( 
.A(n_2353),
.Y(n_2401)
);

OR2x2_ASAP7_75t_L g2402 ( 
.A(n_2279),
.B(n_101),
.Y(n_2402)
);

BUFx3_ASAP7_75t_L g2403 ( 
.A(n_2366),
.Y(n_2403)
);

NAND2xp5_ASAP7_75t_L g2404 ( 
.A(n_2284),
.B(n_101),
.Y(n_2404)
);

AOI22xp33_ASAP7_75t_L g2405 ( 
.A1(n_2346),
.A2(n_2333),
.B1(n_2340),
.B2(n_2343),
.Y(n_2405)
);

BUFx3_ASAP7_75t_L g2406 ( 
.A(n_2316),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_2360),
.Y(n_2407)
);

INVx4_ASAP7_75t_L g2408 ( 
.A(n_2348),
.Y(n_2408)
);

INVx2_ASAP7_75t_L g2409 ( 
.A(n_2362),
.Y(n_2409)
);

INVxp67_ASAP7_75t_SL g2410 ( 
.A(n_2311),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2272),
.Y(n_2411)
);

INVx2_ASAP7_75t_L g2412 ( 
.A(n_2289),
.Y(n_2412)
);

NOR2xp33_ASAP7_75t_L g2413 ( 
.A(n_2336),
.B(n_2321),
.Y(n_2413)
);

INVx2_ASAP7_75t_L g2414 ( 
.A(n_2294),
.Y(n_2414)
);

INVx1_ASAP7_75t_L g2415 ( 
.A(n_2288),
.Y(n_2415)
);

HB1xp67_ASAP7_75t_L g2416 ( 
.A(n_2331),
.Y(n_2416)
);

NOR2x1p5_ASAP7_75t_L g2417 ( 
.A(n_2343),
.B(n_102),
.Y(n_2417)
);

OR2x2_ASAP7_75t_L g2418 ( 
.A(n_2295),
.B(n_2293),
.Y(n_2418)
);

AND2x2_ASAP7_75t_L g2419 ( 
.A(n_2325),
.B(n_102),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_2297),
.Y(n_2420)
);

AND2x2_ASAP7_75t_L g2421 ( 
.A(n_2328),
.B(n_104),
.Y(n_2421)
);

BUFx6f_ASAP7_75t_L g2422 ( 
.A(n_2365),
.Y(n_2422)
);

HB1xp67_ASAP7_75t_L g2423 ( 
.A(n_2300),
.Y(n_2423)
);

AND2x2_ASAP7_75t_L g2424 ( 
.A(n_2327),
.B(n_104),
.Y(n_2424)
);

OR2x2_ASAP7_75t_SL g2425 ( 
.A(n_2342),
.B(n_2280),
.Y(n_2425)
);

AND2x2_ASAP7_75t_L g2426 ( 
.A(n_2301),
.B(n_105),
.Y(n_2426)
);

INVx1_ASAP7_75t_L g2427 ( 
.A(n_2302),
.Y(n_2427)
);

AND2x4_ASAP7_75t_SL g2428 ( 
.A(n_2319),
.B(n_105),
.Y(n_2428)
);

AND2x4_ASAP7_75t_L g2429 ( 
.A(n_2306),
.B(n_2309),
.Y(n_2429)
);

BUFx2_ASAP7_75t_L g2430 ( 
.A(n_2310),
.Y(n_2430)
);

INVx2_ASAP7_75t_L g2431 ( 
.A(n_2308),
.Y(n_2431)
);

AND2x2_ASAP7_75t_L g2432 ( 
.A(n_2359),
.B(n_106),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_2338),
.Y(n_2433)
);

AOI22xp33_ASAP7_75t_L g2434 ( 
.A1(n_2337),
.A2(n_2345),
.B1(n_2335),
.B2(n_2339),
.Y(n_2434)
);

INVx3_ASAP7_75t_L g2435 ( 
.A(n_2291),
.Y(n_2435)
);

INVx2_ASAP7_75t_L g2436 ( 
.A(n_2323),
.Y(n_2436)
);

INVx2_ASAP7_75t_L g2437 ( 
.A(n_2282),
.Y(n_2437)
);

AND2x2_ASAP7_75t_L g2438 ( 
.A(n_2285),
.B(n_2304),
.Y(n_2438)
);

INVx1_ASAP7_75t_L g2439 ( 
.A(n_2283),
.Y(n_2439)
);

INVx1_ASAP7_75t_L g2440 ( 
.A(n_2290),
.Y(n_2440)
);

AND2x2_ASAP7_75t_L g2441 ( 
.A(n_2276),
.B(n_2355),
.Y(n_2441)
);

AND2x2_ASAP7_75t_L g2442 ( 
.A(n_2356),
.B(n_106),
.Y(n_2442)
);

AND2x2_ASAP7_75t_L g2443 ( 
.A(n_2358),
.B(n_107),
.Y(n_2443)
);

HB1xp67_ASAP7_75t_L g2444 ( 
.A(n_2363),
.Y(n_2444)
);

INVx2_ASAP7_75t_L g2445 ( 
.A(n_2314),
.Y(n_2445)
);

INVx1_ASAP7_75t_L g2446 ( 
.A(n_2313),
.Y(n_2446)
);

INVxp33_ASAP7_75t_SL g2447 ( 
.A(n_2315),
.Y(n_2447)
);

INVx2_ASAP7_75t_L g2448 ( 
.A(n_2318),
.Y(n_2448)
);

AND2x2_ASAP7_75t_L g2449 ( 
.A(n_2326),
.B(n_107),
.Y(n_2449)
);

INVx2_ASAP7_75t_L g2450 ( 
.A(n_2318),
.Y(n_2450)
);

INVx1_ASAP7_75t_L g2451 ( 
.A(n_2344),
.Y(n_2451)
);

INVx2_ASAP7_75t_L g2452 ( 
.A(n_2344),
.Y(n_2452)
);

INVx1_ASAP7_75t_L g2453 ( 
.A(n_2354),
.Y(n_2453)
);

AND2x2_ASAP7_75t_L g2454 ( 
.A(n_2334),
.B(n_108),
.Y(n_2454)
);

INVx2_ASAP7_75t_L g2455 ( 
.A(n_2332),
.Y(n_2455)
);

HB1xp67_ASAP7_75t_L g2456 ( 
.A(n_2299),
.Y(n_2456)
);

INVx1_ASAP7_75t_L g2457 ( 
.A(n_2299),
.Y(n_2457)
);

AND2x2_ASAP7_75t_L g2458 ( 
.A(n_2270),
.B(n_108),
.Y(n_2458)
);

INVx1_ASAP7_75t_L g2459 ( 
.A(n_2299),
.Y(n_2459)
);

NAND2xp5_ASAP7_75t_L g2460 ( 
.A(n_2303),
.B(n_109),
.Y(n_2460)
);

INVx1_ASAP7_75t_L g2461 ( 
.A(n_2299),
.Y(n_2461)
);

INVx1_ASAP7_75t_L g2462 ( 
.A(n_2299),
.Y(n_2462)
);

NAND2xp33_ASAP7_75t_L g2463 ( 
.A(n_2343),
.B(n_110),
.Y(n_2463)
);

NAND2xp5_ASAP7_75t_L g2464 ( 
.A(n_2303),
.B(n_110),
.Y(n_2464)
);

INVx1_ASAP7_75t_L g2465 ( 
.A(n_2299),
.Y(n_2465)
);

BUFx2_ASAP7_75t_L g2466 ( 
.A(n_2361),
.Y(n_2466)
);

OR2x2_ASAP7_75t_L g2467 ( 
.A(n_2324),
.B(n_111),
.Y(n_2467)
);

INVx1_ASAP7_75t_L g2468 ( 
.A(n_2299),
.Y(n_2468)
);

INVx1_ASAP7_75t_L g2469 ( 
.A(n_2299),
.Y(n_2469)
);

INVxp67_ASAP7_75t_SL g2470 ( 
.A(n_2303),
.Y(n_2470)
);

OR2x2_ASAP7_75t_L g2471 ( 
.A(n_2324),
.B(n_112),
.Y(n_2471)
);

INVx2_ASAP7_75t_L g2472 ( 
.A(n_2332),
.Y(n_2472)
);

NOR2xp33_ASAP7_75t_L g2473 ( 
.A(n_2361),
.B(n_112),
.Y(n_2473)
);

INVx2_ASAP7_75t_L g2474 ( 
.A(n_2332),
.Y(n_2474)
);

INVx1_ASAP7_75t_L g2475 ( 
.A(n_2299),
.Y(n_2475)
);

AND2x2_ASAP7_75t_L g2476 ( 
.A(n_2270),
.B(n_113),
.Y(n_2476)
);

NAND3xp33_ASAP7_75t_L g2477 ( 
.A(n_2341),
.B(n_113),
.C(n_114),
.Y(n_2477)
);

INVx2_ASAP7_75t_L g2478 ( 
.A(n_2332),
.Y(n_2478)
);

AND2x4_ASAP7_75t_L g2479 ( 
.A(n_2286),
.B(n_115),
.Y(n_2479)
);

INVx2_ASAP7_75t_L g2480 ( 
.A(n_2332),
.Y(n_2480)
);

INVx2_ASAP7_75t_L g2481 ( 
.A(n_2332),
.Y(n_2481)
);

AND2x4_ASAP7_75t_L g2482 ( 
.A(n_2286),
.B(n_116),
.Y(n_2482)
);

NAND2xp5_ASAP7_75t_L g2483 ( 
.A(n_2303),
.B(n_116),
.Y(n_2483)
);

INVx1_ASAP7_75t_L g2484 ( 
.A(n_2299),
.Y(n_2484)
);

OAI21xp33_ASAP7_75t_SL g2485 ( 
.A1(n_2361),
.A2(n_117),
.B(n_118),
.Y(n_2485)
);

AOI22xp5_ASAP7_75t_L g2486 ( 
.A1(n_2354),
.A2(n_119),
.B1(n_117),
.B2(n_118),
.Y(n_2486)
);

INVxp67_ASAP7_75t_L g2487 ( 
.A(n_2324),
.Y(n_2487)
);

AND2x2_ASAP7_75t_L g2488 ( 
.A(n_2270),
.B(n_120),
.Y(n_2488)
);

NAND3xp33_ASAP7_75t_L g2489 ( 
.A(n_2341),
.B(n_122),
.C(n_123),
.Y(n_2489)
);

AND2x4_ASAP7_75t_L g2490 ( 
.A(n_2286),
.B(n_122),
.Y(n_2490)
);

AND2x4_ASAP7_75t_L g2491 ( 
.A(n_2286),
.B(n_123),
.Y(n_2491)
);

AND2x4_ASAP7_75t_L g2492 ( 
.A(n_2375),
.B(n_124),
.Y(n_2492)
);

NOR2x1_ASAP7_75t_L g2493 ( 
.A(n_2378),
.B(n_124),
.Y(n_2493)
);

INVx2_ASAP7_75t_L g2494 ( 
.A(n_2466),
.Y(n_2494)
);

INVx2_ASAP7_75t_SL g2495 ( 
.A(n_2373),
.Y(n_2495)
);

INVx1_ASAP7_75t_L g2496 ( 
.A(n_2388),
.Y(n_2496)
);

INVx2_ASAP7_75t_L g2497 ( 
.A(n_2418),
.Y(n_2497)
);

INVx1_ASAP7_75t_L g2498 ( 
.A(n_2394),
.Y(n_2498)
);

INVx1_ASAP7_75t_L g2499 ( 
.A(n_2395),
.Y(n_2499)
);

HB1xp67_ASAP7_75t_L g2500 ( 
.A(n_2382),
.Y(n_2500)
);

INVx2_ASAP7_75t_L g2501 ( 
.A(n_2377),
.Y(n_2501)
);

OR2x2_ASAP7_75t_L g2502 ( 
.A(n_2425),
.B(n_125),
.Y(n_2502)
);

INVx1_ASAP7_75t_L g2503 ( 
.A(n_2400),
.Y(n_2503)
);

INVx2_ASAP7_75t_L g2504 ( 
.A(n_2455),
.Y(n_2504)
);

INVx2_ASAP7_75t_L g2505 ( 
.A(n_2472),
.Y(n_2505)
);

INVx1_ASAP7_75t_L g2506 ( 
.A(n_2407),
.Y(n_2506)
);

NAND2xp5_ASAP7_75t_L g2507 ( 
.A(n_2470),
.B(n_125),
.Y(n_2507)
);

AND2x2_ASAP7_75t_L g2508 ( 
.A(n_2431),
.B(n_126),
.Y(n_2508)
);

INVx1_ASAP7_75t_L g2509 ( 
.A(n_2415),
.Y(n_2509)
);

INVx2_ASAP7_75t_L g2510 ( 
.A(n_2474),
.Y(n_2510)
);

AND2x4_ASAP7_75t_L g2511 ( 
.A(n_2379),
.B(n_2403),
.Y(n_2511)
);

INVx2_ASAP7_75t_SL g2512 ( 
.A(n_2422),
.Y(n_2512)
);

OR2x2_ASAP7_75t_L g2513 ( 
.A(n_2451),
.B(n_126),
.Y(n_2513)
);

INVx1_ASAP7_75t_L g2514 ( 
.A(n_2411),
.Y(n_2514)
);

INVx1_ASAP7_75t_L g2515 ( 
.A(n_2420),
.Y(n_2515)
);

AND2x2_ASAP7_75t_L g2516 ( 
.A(n_2444),
.B(n_127),
.Y(n_2516)
);

INVx1_ASAP7_75t_L g2517 ( 
.A(n_2427),
.Y(n_2517)
);

INVx1_ASAP7_75t_L g2518 ( 
.A(n_2423),
.Y(n_2518)
);

INVx4_ASAP7_75t_L g2519 ( 
.A(n_2374),
.Y(n_2519)
);

INVx2_ASAP7_75t_L g2520 ( 
.A(n_2478),
.Y(n_2520)
);

INVx2_ASAP7_75t_L g2521 ( 
.A(n_2480),
.Y(n_2521)
);

INVx1_ASAP7_75t_L g2522 ( 
.A(n_2433),
.Y(n_2522)
);

NAND2xp5_ASAP7_75t_L g2523 ( 
.A(n_2446),
.B(n_127),
.Y(n_2523)
);

HB1xp67_ASAP7_75t_L g2524 ( 
.A(n_2416),
.Y(n_2524)
);

BUFx2_ASAP7_75t_L g2525 ( 
.A(n_2381),
.Y(n_2525)
);

INVx1_ASAP7_75t_L g2526 ( 
.A(n_2385),
.Y(n_2526)
);

OR2x2_ASAP7_75t_L g2527 ( 
.A(n_2487),
.B(n_128),
.Y(n_2527)
);

INVx2_ASAP7_75t_L g2528 ( 
.A(n_2481),
.Y(n_2528)
);

NAND2xp5_ASAP7_75t_L g2529 ( 
.A(n_2439),
.B(n_2440),
.Y(n_2529)
);

INVx2_ASAP7_75t_L g2530 ( 
.A(n_2430),
.Y(n_2530)
);

AND2x4_ASAP7_75t_L g2531 ( 
.A(n_2437),
.B(n_128),
.Y(n_2531)
);

INVx1_ASAP7_75t_L g2532 ( 
.A(n_2452),
.Y(n_2532)
);

INVx2_ASAP7_75t_L g2533 ( 
.A(n_2429),
.Y(n_2533)
);

INVx2_ASAP7_75t_L g2534 ( 
.A(n_2384),
.Y(n_2534)
);

CKINVDCx11_ASAP7_75t_R g2535 ( 
.A(n_2369),
.Y(n_2535)
);

NAND2xp5_ASAP7_75t_L g2536 ( 
.A(n_2413),
.B(n_129),
.Y(n_2536)
);

INVx1_ASAP7_75t_L g2537 ( 
.A(n_2370),
.Y(n_2537)
);

NAND2x1p5_ASAP7_75t_L g2538 ( 
.A(n_2408),
.B(n_129),
.Y(n_2538)
);

NAND2xp5_ASAP7_75t_L g2539 ( 
.A(n_2380),
.B(n_130),
.Y(n_2539)
);

INVx2_ASAP7_75t_L g2540 ( 
.A(n_2387),
.Y(n_2540)
);

INVx1_ASAP7_75t_L g2541 ( 
.A(n_2456),
.Y(n_2541)
);

AND2x2_ASAP7_75t_SL g2542 ( 
.A(n_2463),
.B(n_130),
.Y(n_2542)
);

INVx2_ASAP7_75t_L g2543 ( 
.A(n_2389),
.Y(n_2543)
);

INVx1_ASAP7_75t_L g2544 ( 
.A(n_2368),
.Y(n_2544)
);

NAND2xp5_ASAP7_75t_L g2545 ( 
.A(n_2390),
.B(n_131),
.Y(n_2545)
);

HB1xp67_ASAP7_75t_L g2546 ( 
.A(n_2371),
.Y(n_2546)
);

AND2x2_ASAP7_75t_L g2547 ( 
.A(n_2393),
.B(n_131),
.Y(n_2547)
);

BUFx2_ASAP7_75t_L g2548 ( 
.A(n_2448),
.Y(n_2548)
);

NOR2x1_ASAP7_75t_L g2549 ( 
.A(n_2374),
.B(n_132),
.Y(n_2549)
);

AND2x2_ASAP7_75t_L g2550 ( 
.A(n_2396),
.B(n_132),
.Y(n_2550)
);

INVxp67_ASAP7_75t_SL g2551 ( 
.A(n_2450),
.Y(n_2551)
);

AND2x2_ASAP7_75t_L g2552 ( 
.A(n_2445),
.B(n_133),
.Y(n_2552)
);

INVx1_ASAP7_75t_L g2553 ( 
.A(n_2457),
.Y(n_2553)
);

INVx1_ASAP7_75t_L g2554 ( 
.A(n_2459),
.Y(n_2554)
);

INVx2_ASAP7_75t_L g2555 ( 
.A(n_2391),
.Y(n_2555)
);

INVx2_ASAP7_75t_L g2556 ( 
.A(n_2401),
.Y(n_2556)
);

INVx1_ASAP7_75t_SL g2557 ( 
.A(n_2428),
.Y(n_2557)
);

HB1xp67_ASAP7_75t_L g2558 ( 
.A(n_2461),
.Y(n_2558)
);

INVx1_ASAP7_75t_SL g2559 ( 
.A(n_2367),
.Y(n_2559)
);

INVx2_ASAP7_75t_L g2560 ( 
.A(n_2409),
.Y(n_2560)
);

BUFx3_ASAP7_75t_L g2561 ( 
.A(n_2422),
.Y(n_2561)
);

HB1xp67_ASAP7_75t_L g2562 ( 
.A(n_2462),
.Y(n_2562)
);

NAND2xp5_ASAP7_75t_L g2563 ( 
.A(n_2426),
.B(n_133),
.Y(n_2563)
);

AND2x2_ASAP7_75t_L g2564 ( 
.A(n_2399),
.B(n_134),
.Y(n_2564)
);

OR2x2_ASAP7_75t_L g2565 ( 
.A(n_2465),
.B(n_135),
.Y(n_2565)
);

INVx1_ASAP7_75t_L g2566 ( 
.A(n_2468),
.Y(n_2566)
);

NAND2xp5_ASAP7_75t_L g2567 ( 
.A(n_2397),
.B(n_136),
.Y(n_2567)
);

AND2x2_ASAP7_75t_L g2568 ( 
.A(n_2435),
.B(n_136),
.Y(n_2568)
);

INVxp67_ASAP7_75t_L g2569 ( 
.A(n_2453),
.Y(n_2569)
);

INVx2_ASAP7_75t_SL g2570 ( 
.A(n_2406),
.Y(n_2570)
);

INVx2_ASAP7_75t_L g2571 ( 
.A(n_2386),
.Y(n_2571)
);

INVx2_ASAP7_75t_L g2572 ( 
.A(n_2412),
.Y(n_2572)
);

INVx2_ASAP7_75t_L g2573 ( 
.A(n_2414),
.Y(n_2573)
);

AND2x2_ASAP7_75t_L g2574 ( 
.A(n_2438),
.B(n_137),
.Y(n_2574)
);

AND2x2_ASAP7_75t_L g2575 ( 
.A(n_2441),
.B(n_137),
.Y(n_2575)
);

INVx2_ASAP7_75t_L g2576 ( 
.A(n_2436),
.Y(n_2576)
);

AND2x2_ASAP7_75t_L g2577 ( 
.A(n_2469),
.B(n_2475),
.Y(n_2577)
);

NAND2xp5_ASAP7_75t_L g2578 ( 
.A(n_2404),
.B(n_2392),
.Y(n_2578)
);

INVx1_ASAP7_75t_L g2579 ( 
.A(n_2484),
.Y(n_2579)
);

INVx2_ASAP7_75t_L g2580 ( 
.A(n_2402),
.Y(n_2580)
);

OR2x2_ASAP7_75t_L g2581 ( 
.A(n_2467),
.B(n_138),
.Y(n_2581)
);

INVx1_ASAP7_75t_L g2582 ( 
.A(n_2410),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_2471),
.Y(n_2583)
);

NAND2xp5_ASAP7_75t_L g2584 ( 
.A(n_2458),
.B(n_2488),
.Y(n_2584)
);

AND2x4_ASAP7_75t_L g2585 ( 
.A(n_2476),
.B(n_139),
.Y(n_2585)
);

INVx2_ASAP7_75t_L g2586 ( 
.A(n_2376),
.Y(n_2586)
);

AND2x2_ASAP7_75t_L g2587 ( 
.A(n_2434),
.B(n_139),
.Y(n_2587)
);

AND2x2_ASAP7_75t_L g2588 ( 
.A(n_2398),
.B(n_140),
.Y(n_2588)
);

INVx1_ASAP7_75t_L g2589 ( 
.A(n_2372),
.Y(n_2589)
);

AND2x2_ASAP7_75t_L g2590 ( 
.A(n_2424),
.B(n_140),
.Y(n_2590)
);

AND2x4_ASAP7_75t_L g2591 ( 
.A(n_2419),
.B(n_141),
.Y(n_2591)
);

AND2x4_ASAP7_75t_L g2592 ( 
.A(n_2421),
.B(n_142),
.Y(n_2592)
);

AOI22xp33_ASAP7_75t_L g2593 ( 
.A1(n_2405),
.A2(n_2486),
.B1(n_2489),
.B2(n_2477),
.Y(n_2593)
);

OR2x2_ASAP7_75t_L g2594 ( 
.A(n_2460),
.B(n_142),
.Y(n_2594)
);

AND2x2_ASAP7_75t_L g2595 ( 
.A(n_2432),
.B(n_143),
.Y(n_2595)
);

NAND2xp5_ASAP7_75t_L g2596 ( 
.A(n_2464),
.B(n_143),
.Y(n_2596)
);

NAND2xp5_ASAP7_75t_L g2597 ( 
.A(n_2483),
.B(n_144),
.Y(n_2597)
);

INVx2_ASAP7_75t_SL g2598 ( 
.A(n_2479),
.Y(n_2598)
);

HB1xp67_ASAP7_75t_L g2599 ( 
.A(n_2447),
.Y(n_2599)
);

AOI22xp33_ASAP7_75t_L g2600 ( 
.A1(n_2417),
.A2(n_2383),
.B1(n_2473),
.B2(n_2449),
.Y(n_2600)
);

AND2x4_ASAP7_75t_SL g2601 ( 
.A(n_2482),
.B(n_144),
.Y(n_2601)
);

INVx1_ASAP7_75t_L g2602 ( 
.A(n_2442),
.Y(n_2602)
);

OR2x2_ASAP7_75t_L g2603 ( 
.A(n_2443),
.B(n_145),
.Y(n_2603)
);

AND2x2_ASAP7_75t_L g2604 ( 
.A(n_2490),
.B(n_145),
.Y(n_2604)
);

AND2x2_ASAP7_75t_L g2605 ( 
.A(n_2491),
.B(n_146),
.Y(n_2605)
);

OR2x2_ASAP7_75t_L g2606 ( 
.A(n_2454),
.B(n_146),
.Y(n_2606)
);

AND2x2_ASAP7_75t_L g2607 ( 
.A(n_2485),
.B(n_147),
.Y(n_2607)
);

INVx1_ASAP7_75t_L g2608 ( 
.A(n_2388),
.Y(n_2608)
);

INVx1_ASAP7_75t_L g2609 ( 
.A(n_2388),
.Y(n_2609)
);

INVx1_ASAP7_75t_L g2610 ( 
.A(n_2388),
.Y(n_2610)
);

INVx2_ASAP7_75t_L g2611 ( 
.A(n_2466),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_2388),
.Y(n_2612)
);

AND2x4_ASAP7_75t_L g2613 ( 
.A(n_2375),
.B(n_147),
.Y(n_2613)
);

INVx1_ASAP7_75t_L g2614 ( 
.A(n_2388),
.Y(n_2614)
);

AND2x4_ASAP7_75t_L g2615 ( 
.A(n_2375),
.B(n_148),
.Y(n_2615)
);

NOR2x1_ASAP7_75t_L g2616 ( 
.A(n_2378),
.B(n_148),
.Y(n_2616)
);

AND2x2_ASAP7_75t_L g2617 ( 
.A(n_2378),
.B(n_149),
.Y(n_2617)
);

OR2x2_ASAP7_75t_L g2618 ( 
.A(n_2425),
.B(n_149),
.Y(n_2618)
);

AND2x2_ASAP7_75t_L g2619 ( 
.A(n_2378),
.B(n_150),
.Y(n_2619)
);

NOR2xp33_ASAP7_75t_L g2620 ( 
.A(n_2453),
.B(n_150),
.Y(n_2620)
);

INVx1_ASAP7_75t_L g2621 ( 
.A(n_2388),
.Y(n_2621)
);

NOR2x1_ASAP7_75t_L g2622 ( 
.A(n_2378),
.B(n_151),
.Y(n_2622)
);

AND2x2_ASAP7_75t_L g2623 ( 
.A(n_2378),
.B(n_153),
.Y(n_2623)
);

NAND2xp5_ASAP7_75t_L g2624 ( 
.A(n_2470),
.B(n_153),
.Y(n_2624)
);

NAND2xp5_ASAP7_75t_L g2625 ( 
.A(n_2470),
.B(n_154),
.Y(n_2625)
);

INVx1_ASAP7_75t_L g2626 ( 
.A(n_2388),
.Y(n_2626)
);

AND2x2_ASAP7_75t_L g2627 ( 
.A(n_2378),
.B(n_154),
.Y(n_2627)
);

AND2x2_ASAP7_75t_L g2628 ( 
.A(n_2378),
.B(n_155),
.Y(n_2628)
);

INVx2_ASAP7_75t_L g2629 ( 
.A(n_2466),
.Y(n_2629)
);

HB1xp67_ASAP7_75t_L g2630 ( 
.A(n_2382),
.Y(n_2630)
);

AND2x2_ASAP7_75t_L g2631 ( 
.A(n_2378),
.B(n_155),
.Y(n_2631)
);

AND2x4_ASAP7_75t_L g2632 ( 
.A(n_2375),
.B(n_156),
.Y(n_2632)
);

INVx2_ASAP7_75t_L g2633 ( 
.A(n_2466),
.Y(n_2633)
);

INVx1_ASAP7_75t_L g2634 ( 
.A(n_2388),
.Y(n_2634)
);

INVx2_ASAP7_75t_L g2635 ( 
.A(n_2466),
.Y(n_2635)
);

AOI22xp33_ASAP7_75t_L g2636 ( 
.A1(n_2453),
.A2(n_158),
.B1(n_156),
.B2(n_157),
.Y(n_2636)
);

NAND2xp5_ASAP7_75t_L g2637 ( 
.A(n_2470),
.B(n_157),
.Y(n_2637)
);

NOR2xp33_ASAP7_75t_L g2638 ( 
.A(n_2453),
.B(n_159),
.Y(n_2638)
);

NAND2xp5_ASAP7_75t_L g2639 ( 
.A(n_2470),
.B(n_159),
.Y(n_2639)
);

BUFx12f_ASAP7_75t_L g2640 ( 
.A(n_2417),
.Y(n_2640)
);

HB1xp67_ASAP7_75t_L g2641 ( 
.A(n_2382),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_2388),
.Y(n_2642)
);

HB1xp67_ASAP7_75t_L g2643 ( 
.A(n_2382),
.Y(n_2643)
);

INVx1_ASAP7_75t_L g2644 ( 
.A(n_2388),
.Y(n_2644)
);

AND2x2_ASAP7_75t_L g2645 ( 
.A(n_2378),
.B(n_161),
.Y(n_2645)
);

AND2x2_ASAP7_75t_L g2646 ( 
.A(n_2378),
.B(n_161),
.Y(n_2646)
);

INVx2_ASAP7_75t_L g2647 ( 
.A(n_2466),
.Y(n_2647)
);

INVxp67_ASAP7_75t_SL g2648 ( 
.A(n_2470),
.Y(n_2648)
);

INVx1_ASAP7_75t_L g2649 ( 
.A(n_2388),
.Y(n_2649)
);

INVx2_ASAP7_75t_L g2650 ( 
.A(n_2466),
.Y(n_2650)
);

OR2x2_ASAP7_75t_L g2651 ( 
.A(n_2425),
.B(n_162),
.Y(n_2651)
);

INVx2_ASAP7_75t_L g2652 ( 
.A(n_2466),
.Y(n_2652)
);

INVx1_ASAP7_75t_L g2653 ( 
.A(n_2388),
.Y(n_2653)
);

AOI22xp33_ASAP7_75t_L g2654 ( 
.A1(n_2453),
.A2(n_164),
.B1(n_162),
.B2(n_163),
.Y(n_2654)
);

OR2x2_ASAP7_75t_L g2655 ( 
.A(n_2425),
.B(n_163),
.Y(n_2655)
);

AND2x4_ASAP7_75t_SL g2656 ( 
.A(n_2369),
.B(n_164),
.Y(n_2656)
);

INVx1_ASAP7_75t_L g2657 ( 
.A(n_2388),
.Y(n_2657)
);

NAND2xp5_ASAP7_75t_L g2658 ( 
.A(n_2470),
.B(n_165),
.Y(n_2658)
);

NAND2xp5_ASAP7_75t_L g2659 ( 
.A(n_2470),
.B(n_166),
.Y(n_2659)
);

INVx2_ASAP7_75t_L g2660 ( 
.A(n_2466),
.Y(n_2660)
);

OR2x2_ASAP7_75t_L g2661 ( 
.A(n_2425),
.B(n_166),
.Y(n_2661)
);

INVx2_ASAP7_75t_L g2662 ( 
.A(n_2466),
.Y(n_2662)
);

INVx2_ASAP7_75t_L g2663 ( 
.A(n_2466),
.Y(n_2663)
);

AND2x2_ASAP7_75t_L g2664 ( 
.A(n_2378),
.B(n_167),
.Y(n_2664)
);

OAI221xp5_ASAP7_75t_L g2665 ( 
.A1(n_2593),
.A2(n_2648),
.B1(n_2569),
.B2(n_2599),
.C(n_2600),
.Y(n_2665)
);

OAI21x1_ASAP7_75t_L g2666 ( 
.A1(n_2494),
.A2(n_167),
.B(n_168),
.Y(n_2666)
);

INVx1_ASAP7_75t_SL g2667 ( 
.A(n_2535),
.Y(n_2667)
);

INVx1_ASAP7_75t_L g2668 ( 
.A(n_2496),
.Y(n_2668)
);

OAI22xp5_ASAP7_75t_L g2669 ( 
.A1(n_2519),
.A2(n_2493),
.B1(n_2622),
.B2(n_2616),
.Y(n_2669)
);

INVx1_ASAP7_75t_L g2670 ( 
.A(n_2498),
.Y(n_2670)
);

OR2x2_ASAP7_75t_L g2671 ( 
.A(n_2497),
.B(n_169),
.Y(n_2671)
);

HB1xp67_ASAP7_75t_L g2672 ( 
.A(n_2524),
.Y(n_2672)
);

INVx2_ASAP7_75t_L g2673 ( 
.A(n_2561),
.Y(n_2673)
);

INVx1_ASAP7_75t_L g2674 ( 
.A(n_2499),
.Y(n_2674)
);

AOI33xp33_ASAP7_75t_L g2675 ( 
.A1(n_2636),
.A2(n_172),
.A3(n_174),
.B1(n_170),
.B2(n_171),
.B3(n_173),
.Y(n_2675)
);

AOI221xp5_ASAP7_75t_L g2676 ( 
.A1(n_2620),
.A2(n_174),
.B1(n_170),
.B2(n_171),
.C(n_175),
.Y(n_2676)
);

HB1xp67_ASAP7_75t_L g2677 ( 
.A(n_2525),
.Y(n_2677)
);

AND2x2_ASAP7_75t_L g2678 ( 
.A(n_2611),
.B(n_2629),
.Y(n_2678)
);

INVx1_ASAP7_75t_L g2679 ( 
.A(n_2503),
.Y(n_2679)
);

OR2x2_ASAP7_75t_L g2680 ( 
.A(n_2537),
.B(n_175),
.Y(n_2680)
);

INVx1_ASAP7_75t_SL g2681 ( 
.A(n_2640),
.Y(n_2681)
);

NOR2xp33_ASAP7_75t_L g2682 ( 
.A(n_2495),
.B(n_2570),
.Y(n_2682)
);

O2A1O1Ixp5_ASAP7_75t_SL g2683 ( 
.A1(n_2532),
.A2(n_179),
.B(n_176),
.C(n_177),
.Y(n_2683)
);

INVx1_ASAP7_75t_SL g2684 ( 
.A(n_2557),
.Y(n_2684)
);

INVx1_ASAP7_75t_L g2685 ( 
.A(n_2506),
.Y(n_2685)
);

OAI22xp33_ASAP7_75t_L g2686 ( 
.A1(n_2502),
.A2(n_179),
.B1(n_176),
.B2(n_177),
.Y(n_2686)
);

HB1xp67_ASAP7_75t_L g2687 ( 
.A(n_2500),
.Y(n_2687)
);

BUFx3_ASAP7_75t_L g2688 ( 
.A(n_2656),
.Y(n_2688)
);

INVx2_ASAP7_75t_L g2689 ( 
.A(n_2511),
.Y(n_2689)
);

INVx1_ASAP7_75t_L g2690 ( 
.A(n_2509),
.Y(n_2690)
);

INVx1_ASAP7_75t_SL g2691 ( 
.A(n_2564),
.Y(n_2691)
);

INVx2_ASAP7_75t_L g2692 ( 
.A(n_2633),
.Y(n_2692)
);

INVx1_ASAP7_75t_L g2693 ( 
.A(n_2608),
.Y(n_2693)
);

INVx1_ASAP7_75t_SL g2694 ( 
.A(n_2617),
.Y(n_2694)
);

AND2x2_ASAP7_75t_L g2695 ( 
.A(n_2635),
.B(n_180),
.Y(n_2695)
);

AOI211xp5_ASAP7_75t_SL g2696 ( 
.A1(n_2638),
.A2(n_182),
.B(n_180),
.C(n_181),
.Y(n_2696)
);

OR2x2_ASAP7_75t_L g2697 ( 
.A(n_2541),
.B(n_181),
.Y(n_2697)
);

INVx1_ASAP7_75t_L g2698 ( 
.A(n_2609),
.Y(n_2698)
);

INVx2_ASAP7_75t_L g2699 ( 
.A(n_2647),
.Y(n_2699)
);

AOI221xp5_ASAP7_75t_L g2700 ( 
.A1(n_2587),
.A2(n_184),
.B1(n_182),
.B2(n_183),
.C(n_185),
.Y(n_2700)
);

AOI22xp33_ASAP7_75t_L g2701 ( 
.A1(n_2580),
.A2(n_186),
.B1(n_183),
.B2(n_185),
.Y(n_2701)
);

AND2x2_ASAP7_75t_L g2702 ( 
.A(n_2650),
.B(n_2652),
.Y(n_2702)
);

AND2x2_ASAP7_75t_L g2703 ( 
.A(n_2660),
.B(n_186),
.Y(n_2703)
);

INVx1_ASAP7_75t_L g2704 ( 
.A(n_2610),
.Y(n_2704)
);

INVx1_ASAP7_75t_L g2705 ( 
.A(n_2612),
.Y(n_2705)
);

OAI211xp5_ASAP7_75t_SL g2706 ( 
.A1(n_2578),
.A2(n_189),
.B(n_187),
.C(n_188),
.Y(n_2706)
);

INVx2_ASAP7_75t_L g2707 ( 
.A(n_2662),
.Y(n_2707)
);

AOI211xp5_ASAP7_75t_L g2708 ( 
.A1(n_2618),
.A2(n_190),
.B(n_187),
.C(n_189),
.Y(n_2708)
);

INVx2_ASAP7_75t_L g2709 ( 
.A(n_2663),
.Y(n_2709)
);

INVx2_ASAP7_75t_L g2710 ( 
.A(n_2512),
.Y(n_2710)
);

CKINVDCx20_ASAP7_75t_R g2711 ( 
.A(n_2601),
.Y(n_2711)
);

INVx1_ASAP7_75t_L g2712 ( 
.A(n_2614),
.Y(n_2712)
);

INVx1_ASAP7_75t_L g2713 ( 
.A(n_2621),
.Y(n_2713)
);

BUFx2_ASAP7_75t_L g2714 ( 
.A(n_2630),
.Y(n_2714)
);

INVxp67_ASAP7_75t_SL g2715 ( 
.A(n_2549),
.Y(n_2715)
);

NAND4xp25_ASAP7_75t_L g2716 ( 
.A(n_2654),
.B(n_193),
.C(n_194),
.D(n_192),
.Y(n_2716)
);

INVx1_ASAP7_75t_L g2717 ( 
.A(n_2626),
.Y(n_2717)
);

INVx1_ASAP7_75t_L g2718 ( 
.A(n_2634),
.Y(n_2718)
);

AOI21x1_ASAP7_75t_L g2719 ( 
.A1(n_2651),
.A2(n_191),
.B(n_192),
.Y(n_2719)
);

OAI22xp33_ASAP7_75t_L g2720 ( 
.A1(n_2655),
.A2(n_194),
.B1(n_191),
.B2(n_193),
.Y(n_2720)
);

OAI33xp33_ASAP7_75t_L g2721 ( 
.A1(n_2582),
.A2(n_197),
.A3(n_199),
.B1(n_195),
.B2(n_196),
.B3(n_198),
.Y(n_2721)
);

BUFx3_ASAP7_75t_L g2722 ( 
.A(n_2492),
.Y(n_2722)
);

OAI31xp33_ASAP7_75t_L g2723 ( 
.A1(n_2661),
.A2(n_198),
.A3(n_196),
.B(n_197),
.Y(n_2723)
);

HB1xp67_ASAP7_75t_L g2724 ( 
.A(n_2641),
.Y(n_2724)
);

INVx3_ASAP7_75t_L g2725 ( 
.A(n_2613),
.Y(n_2725)
);

NAND2xp5_ASAP7_75t_SL g2726 ( 
.A(n_2542),
.B(n_199),
.Y(n_2726)
);

AND2x4_ASAP7_75t_L g2727 ( 
.A(n_2598),
.B(n_201),
.Y(n_2727)
);

INVx1_ASAP7_75t_L g2728 ( 
.A(n_2642),
.Y(n_2728)
);

INVx2_ASAP7_75t_L g2729 ( 
.A(n_2548),
.Y(n_2729)
);

NAND4xp25_ASAP7_75t_SL g2730 ( 
.A(n_2507),
.B(n_204),
.C(n_202),
.D(n_203),
.Y(n_2730)
);

OAI211xp5_ASAP7_75t_L g2731 ( 
.A1(n_2624),
.A2(n_205),
.B(n_202),
.C(n_203),
.Y(n_2731)
);

AND2x2_ASAP7_75t_L g2732 ( 
.A(n_2533),
.B(n_205),
.Y(n_2732)
);

AND2x2_ASAP7_75t_L g2733 ( 
.A(n_2530),
.B(n_206),
.Y(n_2733)
);

INVx1_ASAP7_75t_L g2734 ( 
.A(n_2644),
.Y(n_2734)
);

A2O1A1Ixp33_ASAP7_75t_SL g2735 ( 
.A1(n_2523),
.A2(n_208),
.B(n_206),
.C(n_207),
.Y(n_2735)
);

AOI33xp33_ASAP7_75t_L g2736 ( 
.A1(n_2607),
.A2(n_209),
.A3(n_211),
.B1(n_207),
.B2(n_208),
.B3(n_210),
.Y(n_2736)
);

INVx1_ASAP7_75t_SL g2737 ( 
.A(n_2619),
.Y(n_2737)
);

INVx1_ASAP7_75t_L g2738 ( 
.A(n_2649),
.Y(n_2738)
);

NAND2xp5_ASAP7_75t_L g2739 ( 
.A(n_2583),
.B(n_209),
.Y(n_2739)
);

HB1xp67_ASAP7_75t_L g2740 ( 
.A(n_2643),
.Y(n_2740)
);

CKINVDCx5p33_ASAP7_75t_R g2741 ( 
.A(n_2615),
.Y(n_2741)
);

BUFx2_ASAP7_75t_L g2742 ( 
.A(n_2546),
.Y(n_2742)
);

HB1xp67_ASAP7_75t_L g2743 ( 
.A(n_2548),
.Y(n_2743)
);

HB1xp67_ASAP7_75t_L g2744 ( 
.A(n_2558),
.Y(n_2744)
);

INVx1_ASAP7_75t_L g2745 ( 
.A(n_2653),
.Y(n_2745)
);

INVx5_ASAP7_75t_L g2746 ( 
.A(n_2623),
.Y(n_2746)
);

HB1xp67_ASAP7_75t_L g2747 ( 
.A(n_2562),
.Y(n_2747)
);

INVx5_ASAP7_75t_SL g2748 ( 
.A(n_2632),
.Y(n_2748)
);

AND2x2_ASAP7_75t_L g2749 ( 
.A(n_2559),
.B(n_210),
.Y(n_2749)
);

INVx1_ASAP7_75t_L g2750 ( 
.A(n_2657),
.Y(n_2750)
);

BUFx2_ASAP7_75t_L g2751 ( 
.A(n_2538),
.Y(n_2751)
);

BUFx3_ASAP7_75t_L g2752 ( 
.A(n_2591),
.Y(n_2752)
);

INVx1_ASAP7_75t_L g2753 ( 
.A(n_2514),
.Y(n_2753)
);

INVxp67_ASAP7_75t_L g2754 ( 
.A(n_2513),
.Y(n_2754)
);

AOI322xp5_ASAP7_75t_L g2755 ( 
.A1(n_2536),
.A2(n_216),
.A3(n_215),
.B1(n_213),
.B2(n_211),
.C1(n_212),
.C2(n_214),
.Y(n_2755)
);

INVx1_ASAP7_75t_L g2756 ( 
.A(n_2515),
.Y(n_2756)
);

AND2x2_ASAP7_75t_L g2757 ( 
.A(n_2577),
.B(n_212),
.Y(n_2757)
);

INVx2_ASAP7_75t_L g2758 ( 
.A(n_2586),
.Y(n_2758)
);

OA21x2_ASAP7_75t_L g2759 ( 
.A1(n_2551),
.A2(n_213),
.B(n_214),
.Y(n_2759)
);

OAI21x1_ASAP7_75t_L g2760 ( 
.A1(n_2518),
.A2(n_215),
.B(n_216),
.Y(n_2760)
);

AND2x2_ASAP7_75t_L g2761 ( 
.A(n_2589),
.B(n_217),
.Y(n_2761)
);

AND2x2_ASAP7_75t_L g2762 ( 
.A(n_2602),
.B(n_217),
.Y(n_2762)
);

AND2x2_ASAP7_75t_L g2763 ( 
.A(n_2501),
.B(n_218),
.Y(n_2763)
);

NOR4xp25_ASAP7_75t_L g2764 ( 
.A(n_2625),
.B(n_220),
.C(n_218),
.D(n_219),
.Y(n_2764)
);

INVx2_ASAP7_75t_L g2765 ( 
.A(n_2504),
.Y(n_2765)
);

NAND4xp75_ASAP7_75t_L g2766 ( 
.A(n_2627),
.B(n_223),
.C(n_221),
.D(n_222),
.Y(n_2766)
);

INVx4_ASAP7_75t_L g2767 ( 
.A(n_2585),
.Y(n_2767)
);

AND2x2_ASAP7_75t_L g2768 ( 
.A(n_2505),
.B(n_222),
.Y(n_2768)
);

NAND2x1_ASAP7_75t_L g2769 ( 
.A(n_2576),
.B(n_223),
.Y(n_2769)
);

INVx1_ASAP7_75t_L g2770 ( 
.A(n_2517),
.Y(n_2770)
);

OAI211xp5_ASAP7_75t_SL g2771 ( 
.A1(n_2529),
.A2(n_227),
.B(n_224),
.C(n_226),
.Y(n_2771)
);

AO21x2_ASAP7_75t_L g2772 ( 
.A1(n_2637),
.A2(n_224),
.B(n_226),
.Y(n_2772)
);

OAI221xp5_ASAP7_75t_L g2773 ( 
.A1(n_2639),
.A2(n_229),
.B1(n_227),
.B2(n_228),
.C(n_230),
.Y(n_2773)
);

OR2x2_ASAP7_75t_L g2774 ( 
.A(n_2572),
.B(n_228),
.Y(n_2774)
);

OR2x2_ASAP7_75t_L g2775 ( 
.A(n_2573),
.B(n_230),
.Y(n_2775)
);

INVx1_ASAP7_75t_L g2776 ( 
.A(n_2522),
.Y(n_2776)
);

AO21x2_ASAP7_75t_L g2777 ( 
.A1(n_2658),
.A2(n_231),
.B(n_232),
.Y(n_2777)
);

NAND3xp33_ASAP7_75t_SL g2778 ( 
.A(n_2659),
.B(n_231),
.C(n_233),
.Y(n_2778)
);

AO21x2_ASAP7_75t_L g2779 ( 
.A1(n_2628),
.A2(n_233),
.B(n_234),
.Y(n_2779)
);

OAI21x1_ASAP7_75t_L g2780 ( 
.A1(n_2510),
.A2(n_234),
.B(n_235),
.Y(n_2780)
);

INVx2_ASAP7_75t_L g2781 ( 
.A(n_2520),
.Y(n_2781)
);

AND2x2_ASAP7_75t_L g2782 ( 
.A(n_2521),
.B(n_236),
.Y(n_2782)
);

HB1xp67_ASAP7_75t_L g2783 ( 
.A(n_2528),
.Y(n_2783)
);

INVx2_ASAP7_75t_L g2784 ( 
.A(n_2534),
.Y(n_2784)
);

INVx1_ASAP7_75t_L g2785 ( 
.A(n_2526),
.Y(n_2785)
);

AOI22xp33_ASAP7_75t_L g2786 ( 
.A1(n_2544),
.A2(n_2554),
.B1(n_2566),
.B2(n_2553),
.Y(n_2786)
);

HB1xp67_ASAP7_75t_L g2787 ( 
.A(n_2540),
.Y(n_2787)
);

NAND2x1_ASAP7_75t_L g2788 ( 
.A(n_2759),
.B(n_2631),
.Y(n_2788)
);

NAND2xp5_ASAP7_75t_L g2789 ( 
.A(n_2715),
.B(n_2516),
.Y(n_2789)
);

OR2x2_ASAP7_75t_L g2790 ( 
.A(n_2714),
.B(n_2579),
.Y(n_2790)
);

NAND2x1p5_ASAP7_75t_L g2791 ( 
.A(n_2746),
.B(n_2645),
.Y(n_2791)
);

NAND2xp5_ASAP7_75t_L g2792 ( 
.A(n_2684),
.B(n_2646),
.Y(n_2792)
);

INVx2_ASAP7_75t_L g2793 ( 
.A(n_2722),
.Y(n_2793)
);

OR2x2_ASAP7_75t_L g2794 ( 
.A(n_2742),
.B(n_2694),
.Y(n_2794)
);

BUFx3_ASAP7_75t_L g2795 ( 
.A(n_2688),
.Y(n_2795)
);

AND2x2_ASAP7_75t_L g2796 ( 
.A(n_2746),
.B(n_2543),
.Y(n_2796)
);

HB1xp67_ASAP7_75t_L g2797 ( 
.A(n_2677),
.Y(n_2797)
);

NAND2xp5_ASAP7_75t_L g2798 ( 
.A(n_2746),
.B(n_2664),
.Y(n_2798)
);

NAND2xp5_ASAP7_75t_L g2799 ( 
.A(n_2691),
.B(n_2737),
.Y(n_2799)
);

OR2x2_ASAP7_75t_L g2800 ( 
.A(n_2692),
.B(n_2555),
.Y(n_2800)
);

INVx1_ASAP7_75t_L g2801 ( 
.A(n_2744),
.Y(n_2801)
);

NAND2xp5_ASAP7_75t_L g2802 ( 
.A(n_2687),
.B(n_2531),
.Y(n_2802)
);

INVx1_ASAP7_75t_L g2803 ( 
.A(n_2747),
.Y(n_2803)
);

INVx1_ASAP7_75t_L g2804 ( 
.A(n_2724),
.Y(n_2804)
);

INVx1_ASAP7_75t_L g2805 ( 
.A(n_2740),
.Y(n_2805)
);

AND2x2_ASAP7_75t_L g2806 ( 
.A(n_2689),
.B(n_2556),
.Y(n_2806)
);

NAND2xp5_ASAP7_75t_L g2807 ( 
.A(n_2772),
.B(n_2777),
.Y(n_2807)
);

AND2x4_ASAP7_75t_L g2808 ( 
.A(n_2767),
.B(n_2568),
.Y(n_2808)
);

INVx1_ASAP7_75t_L g2809 ( 
.A(n_2672),
.Y(n_2809)
);

AND2x2_ASAP7_75t_L g2810 ( 
.A(n_2673),
.B(n_2560),
.Y(n_2810)
);

INVx1_ASAP7_75t_L g2811 ( 
.A(n_2743),
.Y(n_2811)
);

AND2x2_ASAP7_75t_L g2812 ( 
.A(n_2710),
.B(n_2571),
.Y(n_2812)
);

NAND2x1p5_ASAP7_75t_L g2813 ( 
.A(n_2769),
.B(n_2550),
.Y(n_2813)
);

HB1xp67_ASAP7_75t_L g2814 ( 
.A(n_2759),
.Y(n_2814)
);

INVx2_ASAP7_75t_L g2815 ( 
.A(n_2725),
.Y(n_2815)
);

AND2x2_ASAP7_75t_L g2816 ( 
.A(n_2678),
.B(n_2574),
.Y(n_2816)
);

INVx1_ASAP7_75t_L g2817 ( 
.A(n_2668),
.Y(n_2817)
);

OR2x2_ASAP7_75t_L g2818 ( 
.A(n_2699),
.B(n_2527),
.Y(n_2818)
);

INVxp67_ASAP7_75t_L g2819 ( 
.A(n_2751),
.Y(n_2819)
);

NAND2xp5_ASAP7_75t_L g2820 ( 
.A(n_2754),
.B(n_2547),
.Y(n_2820)
);

AND2x2_ASAP7_75t_L g2821 ( 
.A(n_2702),
.B(n_2575),
.Y(n_2821)
);

OR2x2_ASAP7_75t_L g2822 ( 
.A(n_2707),
.B(n_2584),
.Y(n_2822)
);

OR2x2_ASAP7_75t_L g2823 ( 
.A(n_2709),
.B(n_2565),
.Y(n_2823)
);

NAND2xp5_ASAP7_75t_L g2824 ( 
.A(n_2779),
.B(n_2508),
.Y(n_2824)
);

NAND2xp5_ASAP7_75t_SL g2825 ( 
.A(n_2669),
.B(n_2592),
.Y(n_2825)
);

NAND2x1p5_ASAP7_75t_L g2826 ( 
.A(n_2667),
.B(n_2552),
.Y(n_2826)
);

OR2x2_ASAP7_75t_L g2827 ( 
.A(n_2758),
.B(n_2665),
.Y(n_2827)
);

AND2x2_ASAP7_75t_L g2828 ( 
.A(n_2682),
.B(n_2595),
.Y(n_2828)
);

AND2x2_ASAP7_75t_L g2829 ( 
.A(n_2748),
.B(n_2588),
.Y(n_2829)
);

INVx2_ASAP7_75t_L g2830 ( 
.A(n_2752),
.Y(n_2830)
);

INVx1_ASAP7_75t_SL g2831 ( 
.A(n_2711),
.Y(n_2831)
);

AND2x2_ASAP7_75t_L g2832 ( 
.A(n_2748),
.B(n_2590),
.Y(n_2832)
);

INVx2_ASAP7_75t_L g2833 ( 
.A(n_2681),
.Y(n_2833)
);

AND2x2_ASAP7_75t_L g2834 ( 
.A(n_2762),
.B(n_2604),
.Y(n_2834)
);

AND2x4_ASAP7_75t_L g2835 ( 
.A(n_2733),
.B(n_2605),
.Y(n_2835)
);

NAND2x1p5_ASAP7_75t_L g2836 ( 
.A(n_2726),
.B(n_2581),
.Y(n_2836)
);

OR2x2_ASAP7_75t_L g2837 ( 
.A(n_2765),
.B(n_2545),
.Y(n_2837)
);

AND2x2_ASAP7_75t_L g2838 ( 
.A(n_2761),
.B(n_2606),
.Y(n_2838)
);

NOR2xp33_ASAP7_75t_L g2839 ( 
.A(n_2739),
.B(n_2741),
.Y(n_2839)
);

INVx1_ASAP7_75t_L g2840 ( 
.A(n_2670),
.Y(n_2840)
);

OR2x2_ASAP7_75t_L g2841 ( 
.A(n_2781),
.B(n_2594),
.Y(n_2841)
);

INVx2_ASAP7_75t_L g2842 ( 
.A(n_2729),
.Y(n_2842)
);

AND2x4_ASAP7_75t_L g2843 ( 
.A(n_2695),
.B(n_2603),
.Y(n_2843)
);

INVx1_ASAP7_75t_L g2844 ( 
.A(n_2674),
.Y(n_2844)
);

NAND2xp5_ASAP7_75t_L g2845 ( 
.A(n_2764),
.B(n_2567),
.Y(n_2845)
);

INVx2_ASAP7_75t_L g2846 ( 
.A(n_2774),
.Y(n_2846)
);

NOR2xp67_ASAP7_75t_L g2847 ( 
.A(n_2783),
.B(n_2539),
.Y(n_2847)
);

INVx2_ASAP7_75t_L g2848 ( 
.A(n_2795),
.Y(n_2848)
);

HB1xp67_ASAP7_75t_L g2849 ( 
.A(n_2797),
.Y(n_2849)
);

INVx1_ASAP7_75t_L g2850 ( 
.A(n_2804),
.Y(n_2850)
);

INVx1_ASAP7_75t_L g2851 ( 
.A(n_2805),
.Y(n_2851)
);

AND2x4_ASAP7_75t_L g2852 ( 
.A(n_2831),
.B(n_2833),
.Y(n_2852)
);

AND2x2_ASAP7_75t_L g2853 ( 
.A(n_2829),
.B(n_2784),
.Y(n_2853)
);

OAI31xp33_ASAP7_75t_L g2854 ( 
.A1(n_2807),
.A2(n_2696),
.A3(n_2731),
.B(n_2706),
.Y(n_2854)
);

AOI22xp5_ASAP7_75t_L g2855 ( 
.A1(n_2819),
.A2(n_2771),
.B1(n_2721),
.B2(n_2730),
.Y(n_2855)
);

INVx1_ASAP7_75t_L g2856 ( 
.A(n_2809),
.Y(n_2856)
);

AND2x2_ASAP7_75t_L g2857 ( 
.A(n_2832),
.B(n_2787),
.Y(n_2857)
);

INVx2_ASAP7_75t_L g2858 ( 
.A(n_2791),
.Y(n_2858)
);

OR2x2_ASAP7_75t_L g2859 ( 
.A(n_2794),
.B(n_2786),
.Y(n_2859)
);

NAND2xp5_ASAP7_75t_L g2860 ( 
.A(n_2843),
.B(n_2708),
.Y(n_2860)
);

INVx1_ASAP7_75t_L g2861 ( 
.A(n_2801),
.Y(n_2861)
);

INVx1_ASAP7_75t_L g2862 ( 
.A(n_2803),
.Y(n_2862)
);

NAND2xp5_ASAP7_75t_L g2863 ( 
.A(n_2838),
.B(n_2686),
.Y(n_2863)
);

AND2x2_ASAP7_75t_L g2864 ( 
.A(n_2826),
.B(n_2749),
.Y(n_2864)
);

INVx1_ASAP7_75t_SL g2865 ( 
.A(n_2828),
.Y(n_2865)
);

INVx2_ASAP7_75t_L g2866 ( 
.A(n_2808),
.Y(n_2866)
);

INVx2_ASAP7_75t_L g2867 ( 
.A(n_2793),
.Y(n_2867)
);

INVx3_ASAP7_75t_L g2868 ( 
.A(n_2835),
.Y(n_2868)
);

INVx1_ASAP7_75t_L g2869 ( 
.A(n_2814),
.Y(n_2869)
);

INVx1_ASAP7_75t_L g2870 ( 
.A(n_2811),
.Y(n_2870)
);

AND2x2_ASAP7_75t_L g2871 ( 
.A(n_2816),
.B(n_2757),
.Y(n_2871)
);

INVx1_ASAP7_75t_L g2872 ( 
.A(n_2799),
.Y(n_2872)
);

INVx2_ASAP7_75t_L g2873 ( 
.A(n_2813),
.Y(n_2873)
);

INVx2_ASAP7_75t_L g2874 ( 
.A(n_2830),
.Y(n_2874)
);

INVx1_ASAP7_75t_L g2875 ( 
.A(n_2790),
.Y(n_2875)
);

INVx1_ASAP7_75t_L g2876 ( 
.A(n_2846),
.Y(n_2876)
);

INVx1_ASAP7_75t_L g2877 ( 
.A(n_2837),
.Y(n_2877)
);

NAND2xp5_ASAP7_75t_L g2878 ( 
.A(n_2834),
.B(n_2720),
.Y(n_2878)
);

NAND2xp5_ASAP7_75t_L g2879 ( 
.A(n_2847),
.B(n_2703),
.Y(n_2879)
);

NOR2xp33_ASAP7_75t_R g2880 ( 
.A(n_2868),
.B(n_2778),
.Y(n_2880)
);

AOI221xp5_ASAP7_75t_SL g2881 ( 
.A1(n_2869),
.A2(n_2845),
.B1(n_2825),
.B2(n_2773),
.C(n_2827),
.Y(n_2881)
);

INVx1_ASAP7_75t_L g2882 ( 
.A(n_2849),
.Y(n_2882)
);

INVx1_ASAP7_75t_L g2883 ( 
.A(n_2875),
.Y(n_2883)
);

AND2x2_ASAP7_75t_L g2884 ( 
.A(n_2864),
.B(n_2821),
.Y(n_2884)
);

INVx1_ASAP7_75t_SL g2885 ( 
.A(n_2865),
.Y(n_2885)
);

INVx1_ASAP7_75t_L g2886 ( 
.A(n_2870),
.Y(n_2886)
);

AND2x2_ASAP7_75t_L g2887 ( 
.A(n_2848),
.B(n_2815),
.Y(n_2887)
);

OR2x2_ASAP7_75t_L g2888 ( 
.A(n_2863),
.B(n_2789),
.Y(n_2888)
);

AND2x2_ASAP7_75t_L g2889 ( 
.A(n_2852),
.B(n_2857),
.Y(n_2889)
);

INVx1_ASAP7_75t_SL g2890 ( 
.A(n_2879),
.Y(n_2890)
);

AND2x2_ASAP7_75t_L g2891 ( 
.A(n_2873),
.B(n_2810),
.Y(n_2891)
);

OR2x2_ASAP7_75t_L g2892 ( 
.A(n_2878),
.B(n_2788),
.Y(n_2892)
);

NAND4xp75_ASAP7_75t_L g2893 ( 
.A(n_2854),
.B(n_2676),
.C(n_2723),
.D(n_2700),
.Y(n_2893)
);

NAND2xp5_ASAP7_75t_L g2894 ( 
.A(n_2871),
.B(n_2792),
.Y(n_2894)
);

INVx1_ASAP7_75t_L g2895 ( 
.A(n_2850),
.Y(n_2895)
);

INVxp67_ASAP7_75t_L g2896 ( 
.A(n_2860),
.Y(n_2896)
);

OR2x2_ASAP7_75t_L g2897 ( 
.A(n_2859),
.B(n_2788),
.Y(n_2897)
);

AND2x4_ASAP7_75t_L g2898 ( 
.A(n_2866),
.B(n_2798),
.Y(n_2898)
);

AND2x2_ASAP7_75t_L g2899 ( 
.A(n_2853),
.B(n_2806),
.Y(n_2899)
);

AND2x2_ASAP7_75t_L g2900 ( 
.A(n_2889),
.B(n_2858),
.Y(n_2900)
);

INVx2_ASAP7_75t_L g2901 ( 
.A(n_2884),
.Y(n_2901)
);

INVx2_ASAP7_75t_SL g2902 ( 
.A(n_2899),
.Y(n_2902)
);

AND2x2_ASAP7_75t_L g2903 ( 
.A(n_2887),
.B(n_2891),
.Y(n_2903)
);

NOR3xp33_ASAP7_75t_L g2904 ( 
.A(n_2896),
.B(n_2872),
.C(n_2867),
.Y(n_2904)
);

INVx1_ASAP7_75t_L g2905 ( 
.A(n_2882),
.Y(n_2905)
);

INVx2_ASAP7_75t_L g2906 ( 
.A(n_2898),
.Y(n_2906)
);

NAND2xp5_ASAP7_75t_L g2907 ( 
.A(n_2885),
.B(n_2855),
.Y(n_2907)
);

AND2x4_ASAP7_75t_L g2908 ( 
.A(n_2883),
.B(n_2874),
.Y(n_2908)
);

INVx1_ASAP7_75t_L g2909 ( 
.A(n_2894),
.Y(n_2909)
);

AND2x2_ASAP7_75t_L g2910 ( 
.A(n_2900),
.B(n_2890),
.Y(n_2910)
);

OR2x2_ASAP7_75t_L g2911 ( 
.A(n_2902),
.B(n_2897),
.Y(n_2911)
);

OAI22xp5_ASAP7_75t_L g2912 ( 
.A1(n_2907),
.A2(n_2893),
.B1(n_2892),
.B2(n_2888),
.Y(n_2912)
);

HB1xp67_ASAP7_75t_L g2913 ( 
.A(n_2906),
.Y(n_2913)
);

INVx1_ASAP7_75t_L g2914 ( 
.A(n_2901),
.Y(n_2914)
);

AOI22xp5_ASAP7_75t_L g2915 ( 
.A1(n_2903),
.A2(n_2881),
.B1(n_2839),
.B2(n_2796),
.Y(n_2915)
);

AOI221xp5_ASAP7_75t_L g2916 ( 
.A1(n_2904),
.A2(n_2861),
.B1(n_2862),
.B2(n_2856),
.C(n_2851),
.Y(n_2916)
);

XOR2x2_ASAP7_75t_L g2917 ( 
.A(n_2909),
.B(n_2766),
.Y(n_2917)
);

NAND2xp5_ASAP7_75t_L g2918 ( 
.A(n_2908),
.B(n_2876),
.Y(n_2918)
);

AND2x2_ASAP7_75t_L g2919 ( 
.A(n_2910),
.B(n_2877),
.Y(n_2919)
);

INVx1_ASAP7_75t_L g2920 ( 
.A(n_2913),
.Y(n_2920)
);

INVx1_ASAP7_75t_L g2921 ( 
.A(n_2911),
.Y(n_2921)
);

INVx1_ASAP7_75t_L g2922 ( 
.A(n_2918),
.Y(n_2922)
);

INVx1_ASAP7_75t_L g2923 ( 
.A(n_2914),
.Y(n_2923)
);

INVx1_ASAP7_75t_L g2924 ( 
.A(n_2917),
.Y(n_2924)
);

NOR3xp33_ASAP7_75t_L g2925 ( 
.A(n_2912),
.B(n_2905),
.C(n_2895),
.Y(n_2925)
);

NAND2xp5_ASAP7_75t_L g2926 ( 
.A(n_2915),
.B(n_2880),
.Y(n_2926)
);

NAND2xp5_ASAP7_75t_L g2927 ( 
.A(n_2916),
.B(n_2820),
.Y(n_2927)
);

AND2x2_ASAP7_75t_L g2928 ( 
.A(n_2910),
.B(n_2812),
.Y(n_2928)
);

AND2x2_ASAP7_75t_L g2929 ( 
.A(n_2910),
.B(n_2842),
.Y(n_2929)
);

AND2x2_ASAP7_75t_L g2930 ( 
.A(n_2910),
.B(n_2886),
.Y(n_2930)
);

NAND2xp5_ASAP7_75t_L g2931 ( 
.A(n_2910),
.B(n_2802),
.Y(n_2931)
);

OR2x2_ASAP7_75t_L g2932 ( 
.A(n_2911),
.B(n_2822),
.Y(n_2932)
);

NAND2xp5_ASAP7_75t_L g2933 ( 
.A(n_2910),
.B(n_2824),
.Y(n_2933)
);

NAND2xp5_ASAP7_75t_L g2934 ( 
.A(n_2910),
.B(n_2836),
.Y(n_2934)
);

HB1xp67_ASAP7_75t_L g2935 ( 
.A(n_2911),
.Y(n_2935)
);

AND2x4_ASAP7_75t_L g2936 ( 
.A(n_2910),
.B(n_2841),
.Y(n_2936)
);

AND2x2_ASAP7_75t_L g2937 ( 
.A(n_2928),
.B(n_2818),
.Y(n_2937)
);

NOR2x1_ASAP7_75t_L g2938 ( 
.A(n_2921),
.B(n_2680),
.Y(n_2938)
);

AND2x2_ASAP7_75t_L g2939 ( 
.A(n_2929),
.B(n_2823),
.Y(n_2939)
);

OAI22xp5_ASAP7_75t_L g2940 ( 
.A1(n_2935),
.A2(n_2800),
.B1(n_2785),
.B2(n_2817),
.Y(n_2940)
);

OR2x2_ASAP7_75t_L g2941 ( 
.A(n_2932),
.B(n_2840),
.Y(n_2941)
);

OR2x2_ASAP7_75t_L g2942 ( 
.A(n_2933),
.B(n_2844),
.Y(n_2942)
);

INVx1_ASAP7_75t_L g2943 ( 
.A(n_2919),
.Y(n_2943)
);

NAND3xp33_ASAP7_75t_L g2944 ( 
.A(n_2925),
.B(n_2755),
.C(n_2701),
.Y(n_2944)
);

NAND2xp5_ASAP7_75t_L g2945 ( 
.A(n_2936),
.B(n_2679),
.Y(n_2945)
);

INVx1_ASAP7_75t_L g2946 ( 
.A(n_2931),
.Y(n_2946)
);

AOI22xp5_ASAP7_75t_L g2947 ( 
.A1(n_2924),
.A2(n_2716),
.B1(n_2776),
.B2(n_2690),
.Y(n_2947)
);

OR2x2_ASAP7_75t_L g2948 ( 
.A(n_2920),
.B(n_2697),
.Y(n_2948)
);

INVx2_ASAP7_75t_L g2949 ( 
.A(n_2930),
.Y(n_2949)
);

INVx1_ASAP7_75t_L g2950 ( 
.A(n_2934),
.Y(n_2950)
);

INVx1_ASAP7_75t_L g2951 ( 
.A(n_2923),
.Y(n_2951)
);

AND2x2_ASAP7_75t_L g2952 ( 
.A(n_2922),
.B(n_2685),
.Y(n_2952)
);

INVx2_ASAP7_75t_L g2953 ( 
.A(n_2926),
.Y(n_2953)
);

NOR4xp25_ASAP7_75t_SL g2954 ( 
.A(n_2927),
.B(n_2698),
.C(n_2704),
.D(n_2693),
.Y(n_2954)
);

INVxp67_ASAP7_75t_SL g2955 ( 
.A(n_2935),
.Y(n_2955)
);

NAND2xp5_ASAP7_75t_L g2956 ( 
.A(n_2935),
.B(n_2705),
.Y(n_2956)
);

NOR3xp33_ASAP7_75t_L g2957 ( 
.A(n_2955),
.B(n_2597),
.C(n_2596),
.Y(n_2957)
);

O2A1O1Ixp33_ASAP7_75t_L g2958 ( 
.A1(n_2943),
.A2(n_2735),
.B(n_2775),
.C(n_2671),
.Y(n_2958)
);

AND4x1_ASAP7_75t_L g2959 ( 
.A(n_2938),
.B(n_2736),
.C(n_2675),
.D(n_2732),
.Y(n_2959)
);

NAND2xp5_ASAP7_75t_L g2960 ( 
.A(n_2939),
.B(n_2770),
.Y(n_2960)
);

INVx1_ASAP7_75t_L g2961 ( 
.A(n_2937),
.Y(n_2961)
);

INVxp33_ASAP7_75t_L g2962 ( 
.A(n_2949),
.Y(n_2962)
);

NAND4xp25_ASAP7_75t_L g2963 ( 
.A(n_2950),
.B(n_2563),
.C(n_2768),
.D(n_2763),
.Y(n_2963)
);

INVx2_ASAP7_75t_L g2964 ( 
.A(n_2948),
.Y(n_2964)
);

NAND3xp33_ASAP7_75t_SL g2965 ( 
.A(n_2954),
.B(n_2782),
.C(n_2683),
.Y(n_2965)
);

NAND4xp25_ASAP7_75t_L g2966 ( 
.A(n_2953),
.B(n_2727),
.C(n_2734),
.D(n_2712),
.Y(n_2966)
);

NOR2xp33_ASAP7_75t_L g2967 ( 
.A(n_2944),
.B(n_2719),
.Y(n_2967)
);

NOR3xp33_ASAP7_75t_L g2968 ( 
.A(n_2946),
.B(n_2760),
.C(n_2666),
.Y(n_2968)
);

NAND3xp33_ASAP7_75t_L g2969 ( 
.A(n_2956),
.B(n_2717),
.C(n_2713),
.Y(n_2969)
);

AOI31xp33_ASAP7_75t_L g2970 ( 
.A1(n_2941),
.A2(n_2728),
.A3(n_2738),
.B(n_2718),
.Y(n_2970)
);

OAI21xp33_ASAP7_75t_SL g2971 ( 
.A1(n_2945),
.A2(n_2951),
.B(n_2952),
.Y(n_2971)
);

INVx1_ASAP7_75t_L g2972 ( 
.A(n_2940),
.Y(n_2972)
);

INVx1_ASAP7_75t_L g2973 ( 
.A(n_2942),
.Y(n_2973)
);

NAND2xp5_ASAP7_75t_L g2974 ( 
.A(n_2947),
.B(n_2745),
.Y(n_2974)
);

OAI21xp5_ASAP7_75t_SL g2975 ( 
.A1(n_2944),
.A2(n_2753),
.B(n_2750),
.Y(n_2975)
);

NAND2xp5_ASAP7_75t_L g2976 ( 
.A(n_2955),
.B(n_2756),
.Y(n_2976)
);

OR2x2_ASAP7_75t_L g2977 ( 
.A(n_2955),
.B(n_2780),
.Y(n_2977)
);

NAND2xp5_ASAP7_75t_L g2978 ( 
.A(n_2961),
.B(n_236),
.Y(n_2978)
);

NAND4xp25_ASAP7_75t_L g2979 ( 
.A(n_2967),
.B(n_239),
.C(n_237),
.D(n_238),
.Y(n_2979)
);

INVx1_ASAP7_75t_L g2980 ( 
.A(n_2977),
.Y(n_2980)
);

NAND3xp33_ASAP7_75t_L g2981 ( 
.A(n_2972),
.B(n_238),
.C(n_239),
.Y(n_2981)
);

NAND2xp5_ASAP7_75t_SL g2982 ( 
.A(n_2958),
.B(n_240),
.Y(n_2982)
);

AOI221xp5_ASAP7_75t_L g2983 ( 
.A1(n_2965),
.A2(n_242),
.B1(n_240),
.B2(n_241),
.C(n_243),
.Y(n_2983)
);

AOI22xp5_ASAP7_75t_L g2984 ( 
.A1(n_2957),
.A2(n_243),
.B1(n_241),
.B2(n_242),
.Y(n_2984)
);

NOR4xp25_ASAP7_75t_L g2985 ( 
.A(n_2971),
.B(n_246),
.C(n_244),
.D(n_245),
.Y(n_2985)
);

NAND2xp5_ASAP7_75t_L g2986 ( 
.A(n_2959),
.B(n_244),
.Y(n_2986)
);

NAND3xp33_ASAP7_75t_L g2987 ( 
.A(n_2976),
.B(n_2964),
.C(n_2973),
.Y(n_2987)
);

O2A1O1Ixp33_ASAP7_75t_L g2988 ( 
.A1(n_2962),
.A2(n_247),
.B(n_245),
.C(n_246),
.Y(n_2988)
);

AOI21x1_ASAP7_75t_L g2989 ( 
.A1(n_2974),
.A2(n_249),
.B(n_248),
.Y(n_2989)
);

OA22x2_ASAP7_75t_L g2990 ( 
.A1(n_2975),
.A2(n_249),
.B1(n_247),
.B2(n_248),
.Y(n_2990)
);

NOR2xp33_ASAP7_75t_L g2991 ( 
.A(n_2963),
.B(n_250),
.Y(n_2991)
);

NAND4xp25_ASAP7_75t_L g2992 ( 
.A(n_2960),
.B(n_252),
.C(n_250),
.D(n_251),
.Y(n_2992)
);

AND3x1_ASAP7_75t_L g2993 ( 
.A(n_2968),
.B(n_252),
.C(n_253),
.Y(n_2993)
);

NOR3xp33_ASAP7_75t_L g2994 ( 
.A(n_2966),
.B(n_256),
.C(n_255),
.Y(n_2994)
);

NAND2xp5_ASAP7_75t_SL g2995 ( 
.A(n_2970),
.B(n_254),
.Y(n_2995)
);

NOR3xp33_ASAP7_75t_L g2996 ( 
.A(n_2969),
.B(n_257),
.C(n_255),
.Y(n_2996)
);

BUFx2_ASAP7_75t_L g2997 ( 
.A(n_2961),
.Y(n_2997)
);

NAND2xp5_ASAP7_75t_L g2998 ( 
.A(n_2961),
.B(n_254),
.Y(n_2998)
);

NAND2xp5_ASAP7_75t_L g2999 ( 
.A(n_2961),
.B(n_257),
.Y(n_2999)
);

NAND3xp33_ASAP7_75t_L g3000 ( 
.A(n_2961),
.B(n_258),
.C(n_259),
.Y(n_3000)
);

OAI21xp5_ASAP7_75t_L g3001 ( 
.A1(n_2962),
.A2(n_260),
.B(n_259),
.Y(n_3001)
);

AND2x2_ASAP7_75t_L g3002 ( 
.A(n_2961),
.B(n_258),
.Y(n_3002)
);

NAND4xp75_ASAP7_75t_L g3003 ( 
.A(n_2971),
.B(n_262),
.C(n_260),
.D(n_261),
.Y(n_3003)
);

AOI21xp33_ASAP7_75t_L g3004 ( 
.A1(n_2962),
.A2(n_261),
.B(n_262),
.Y(n_3004)
);

AOI211xp5_ASAP7_75t_L g3005 ( 
.A1(n_2962),
.A2(n_265),
.B(n_263),
.C(n_264),
.Y(n_3005)
);

NAND3xp33_ASAP7_75t_SL g3006 ( 
.A(n_2961),
.B(n_263),
.C(n_265),
.Y(n_3006)
);

NAND4xp25_ASAP7_75t_SL g3007 ( 
.A(n_2961),
.B(n_268),
.C(n_266),
.D(n_267),
.Y(n_3007)
);

NAND4xp75_ASAP7_75t_L g3008 ( 
.A(n_2971),
.B(n_268),
.C(n_266),
.D(n_267),
.Y(n_3008)
);

AND2x2_ASAP7_75t_L g3009 ( 
.A(n_2961),
.B(n_269),
.Y(n_3009)
);

OAI22xp33_ASAP7_75t_L g3010 ( 
.A1(n_2962),
.A2(n_271),
.B1(n_269),
.B2(n_270),
.Y(n_3010)
);

OAI211xp5_ASAP7_75t_SL g3011 ( 
.A1(n_2961),
.A2(n_273),
.B(n_271),
.C(n_272),
.Y(n_3011)
);

NAND3xp33_ASAP7_75t_L g3012 ( 
.A(n_2961),
.B(n_272),
.C(n_273),
.Y(n_3012)
);

OAI211xp5_ASAP7_75t_L g3013 ( 
.A1(n_2971),
.A2(n_277),
.B(n_274),
.C(n_275),
.Y(n_3013)
);

INVxp67_ASAP7_75t_L g3014 ( 
.A(n_2961),
.Y(n_3014)
);

NAND4xp75_ASAP7_75t_L g3015 ( 
.A(n_2971),
.B(n_278),
.C(n_274),
.D(n_275),
.Y(n_3015)
);

INVx1_ASAP7_75t_L g3016 ( 
.A(n_2977),
.Y(n_3016)
);

NOR2xp33_ASAP7_75t_L g3017 ( 
.A(n_2962),
.B(n_278),
.Y(n_3017)
);

NOR3xp33_ASAP7_75t_L g3018 ( 
.A(n_2987),
.B(n_279),
.C(n_280),
.Y(n_3018)
);

INVx1_ASAP7_75t_L g3019 ( 
.A(n_2997),
.Y(n_3019)
);

INVx1_ASAP7_75t_L g3020 ( 
.A(n_3002),
.Y(n_3020)
);

OAI22xp5_ASAP7_75t_L g3021 ( 
.A1(n_3014),
.A2(n_281),
.B1(n_279),
.B2(n_280),
.Y(n_3021)
);

AOI21xp5_ASAP7_75t_L g3022 ( 
.A1(n_2982),
.A2(n_281),
.B(n_282),
.Y(n_3022)
);

INVxp67_ASAP7_75t_L g3023 ( 
.A(n_2993),
.Y(n_3023)
);

OAI221xp5_ASAP7_75t_L g3024 ( 
.A1(n_2983),
.A2(n_2985),
.B1(n_2994),
.B2(n_3013),
.C(n_2986),
.Y(n_3024)
);

OAI211xp5_ASAP7_75t_L g3025 ( 
.A1(n_2995),
.A2(n_284),
.B(n_282),
.C(n_283),
.Y(n_3025)
);

INVx1_ASAP7_75t_L g3026 ( 
.A(n_3009),
.Y(n_3026)
);

OAI221xp5_ASAP7_75t_L g3027 ( 
.A1(n_2996),
.A2(n_285),
.B1(n_283),
.B2(n_284),
.C(n_286),
.Y(n_3027)
);

OAI21xp5_ASAP7_75t_L g3028 ( 
.A1(n_3017),
.A2(n_285),
.B(n_286),
.Y(n_3028)
);

AOI22xp5_ASAP7_75t_L g3029 ( 
.A1(n_2991),
.A2(n_289),
.B1(n_287),
.B2(n_288),
.Y(n_3029)
);

AOI211xp5_ASAP7_75t_L g3030 ( 
.A1(n_2981),
.A2(n_291),
.B(n_288),
.C(n_290),
.Y(n_3030)
);

OR2x2_ASAP7_75t_L g3031 ( 
.A(n_2979),
.B(n_291),
.Y(n_3031)
);

OAI22xp5_ASAP7_75t_L g3032 ( 
.A1(n_2984),
.A2(n_294),
.B1(n_292),
.B2(n_293),
.Y(n_3032)
);

AOI211xp5_ASAP7_75t_L g3033 ( 
.A1(n_3006),
.A2(n_294),
.B(n_292),
.C(n_293),
.Y(n_3033)
);

NAND2xp5_ASAP7_75t_L g3034 ( 
.A(n_3010),
.B(n_297),
.Y(n_3034)
);

INVx1_ASAP7_75t_L g3035 ( 
.A(n_2990),
.Y(n_3035)
);

NOR2x1_ASAP7_75t_L g3036 ( 
.A(n_3003),
.B(n_297),
.Y(n_3036)
);

INVx1_ASAP7_75t_L g3037 ( 
.A(n_2989),
.Y(n_3037)
);

INVx1_ASAP7_75t_L g3038 ( 
.A(n_3008),
.Y(n_3038)
);

AOI221xp5_ASAP7_75t_L g3039 ( 
.A1(n_2980),
.A2(n_3016),
.B1(n_2998),
.B2(n_2999),
.C(n_2978),
.Y(n_3039)
);

HB1xp67_ASAP7_75t_L g3040 ( 
.A(n_3015),
.Y(n_3040)
);

NAND2xp33_ASAP7_75t_L g3041 ( 
.A(n_3000),
.B(n_298),
.Y(n_3041)
);

INVx2_ASAP7_75t_SL g3042 ( 
.A(n_3012),
.Y(n_3042)
);

INVx1_ASAP7_75t_L g3043 ( 
.A(n_2988),
.Y(n_3043)
);

AOI221xp5_ASAP7_75t_L g3044 ( 
.A1(n_3004),
.A2(n_301),
.B1(n_299),
.B2(n_300),
.C(n_302),
.Y(n_3044)
);

NOR2xp33_ASAP7_75t_L g3045 ( 
.A(n_2992),
.B(n_300),
.Y(n_3045)
);

AOI21xp5_ASAP7_75t_L g3046 ( 
.A1(n_3001),
.A2(n_301),
.B(n_303),
.Y(n_3046)
);

NAND4xp75_ASAP7_75t_L g3047 ( 
.A(n_3007),
.B(n_305),
.C(n_303),
.D(n_304),
.Y(n_3047)
);

AND2x4_ASAP7_75t_SL g3048 ( 
.A(n_3011),
.B(n_304),
.Y(n_3048)
);

NOR3xp33_ASAP7_75t_L g3049 ( 
.A(n_3005),
.B(n_305),
.C(n_306),
.Y(n_3049)
);

OAI22xp5_ASAP7_75t_L g3050 ( 
.A1(n_3014),
.A2(n_308),
.B1(n_306),
.B2(n_307),
.Y(n_3050)
);

INVx1_ASAP7_75t_L g3051 ( 
.A(n_2997),
.Y(n_3051)
);

INVx1_ASAP7_75t_L g3052 ( 
.A(n_2997),
.Y(n_3052)
);

NAND3x1_ASAP7_75t_SL g3053 ( 
.A(n_2983),
.B(n_308),
.C(n_309),
.Y(n_3053)
);

AOI22xp5_ASAP7_75t_L g3054 ( 
.A1(n_3014),
.A2(n_313),
.B1(n_311),
.B2(n_312),
.Y(n_3054)
);

OAI222xp33_ASAP7_75t_L g3055 ( 
.A1(n_3014),
.A2(n_313),
.B1(n_315),
.B2(n_311),
.C1(n_312),
.C2(n_314),
.Y(n_3055)
);

AND2x2_ASAP7_75t_L g3056 ( 
.A(n_2997),
.B(n_314),
.Y(n_3056)
);

NAND4xp75_ASAP7_75t_L g3057 ( 
.A(n_2983),
.B(n_318),
.C(n_316),
.D(n_317),
.Y(n_3057)
);

NAND4xp75_ASAP7_75t_L g3058 ( 
.A(n_2983),
.B(n_319),
.C(n_316),
.D(n_318),
.Y(n_3058)
);

NAND2xp5_ASAP7_75t_L g3059 ( 
.A(n_3002),
.B(n_319),
.Y(n_3059)
);

OAI21xp33_ASAP7_75t_L g3060 ( 
.A1(n_3014),
.A2(n_320),
.B(n_321),
.Y(n_3060)
);

NAND2xp5_ASAP7_75t_L g3061 ( 
.A(n_3002),
.B(n_320),
.Y(n_3061)
);

INVx1_ASAP7_75t_L g3062 ( 
.A(n_2997),
.Y(n_3062)
);

INVx1_ASAP7_75t_L g3063 ( 
.A(n_2997),
.Y(n_3063)
);

INVx1_ASAP7_75t_L g3064 ( 
.A(n_2997),
.Y(n_3064)
);

O2A1O1Ixp33_ASAP7_75t_L g3065 ( 
.A1(n_2995),
.A2(n_324),
.B(n_321),
.C(n_323),
.Y(n_3065)
);

XNOR2xp5_ASAP7_75t_L g3066 ( 
.A(n_2993),
.B(n_323),
.Y(n_3066)
);

NAND2xp5_ASAP7_75t_L g3067 ( 
.A(n_3002),
.B(n_325),
.Y(n_3067)
);

INVx1_ASAP7_75t_L g3068 ( 
.A(n_3056),
.Y(n_3068)
);

NOR4xp25_ASAP7_75t_L g3069 ( 
.A(n_3024),
.B(n_327),
.C(n_325),
.D(n_326),
.Y(n_3069)
);

AND3x4_ASAP7_75t_L g3070 ( 
.A(n_3036),
.B(n_326),
.C(n_327),
.Y(n_3070)
);

AND2x2_ASAP7_75t_L g3071 ( 
.A(n_3048),
.B(n_328),
.Y(n_3071)
);

AOI21xp5_ASAP7_75t_L g3072 ( 
.A1(n_3041),
.A2(n_328),
.B(n_329),
.Y(n_3072)
);

AND2x2_ASAP7_75t_L g3073 ( 
.A(n_3019),
.B(n_329),
.Y(n_3073)
);

INVx2_ASAP7_75t_L g3074 ( 
.A(n_3047),
.Y(n_3074)
);

AND2x2_ASAP7_75t_SL g3075 ( 
.A(n_3051),
.B(n_330),
.Y(n_3075)
);

AND2x2_ASAP7_75t_L g3076 ( 
.A(n_3052),
.B(n_3062),
.Y(n_3076)
);

INVx1_ASAP7_75t_L g3077 ( 
.A(n_3066),
.Y(n_3077)
);

NOR3x1_ASAP7_75t_L g3078 ( 
.A(n_3057),
.B(n_330),
.C(n_331),
.Y(n_3078)
);

NOR3xp33_ASAP7_75t_L g3079 ( 
.A(n_3039),
.B(n_341),
.C(n_332),
.Y(n_3079)
);

NOR2x1_ASAP7_75t_L g3080 ( 
.A(n_3037),
.B(n_332),
.Y(n_3080)
);

NAND3xp33_ASAP7_75t_L g3081 ( 
.A(n_3033),
.B(n_333),
.C(n_334),
.Y(n_3081)
);

NOR2xp67_ASAP7_75t_L g3082 ( 
.A(n_3023),
.B(n_335),
.Y(n_3082)
);

BUFx2_ASAP7_75t_L g3083 ( 
.A(n_3063),
.Y(n_3083)
);

NAND4xp75_ASAP7_75t_L g3084 ( 
.A(n_3064),
.B(n_337),
.C(n_333),
.D(n_336),
.Y(n_3084)
);

AND2x4_ASAP7_75t_L g3085 ( 
.A(n_3020),
.B(n_336),
.Y(n_3085)
);

INVx1_ASAP7_75t_L g3086 ( 
.A(n_3059),
.Y(n_3086)
);

NAND3x1_ASAP7_75t_L g3087 ( 
.A(n_3061),
.B(n_337),
.C(n_339),
.Y(n_3087)
);

NOR2xp33_ASAP7_75t_L g3088 ( 
.A(n_3060),
.B(n_339),
.Y(n_3088)
);

INVxp67_ASAP7_75t_SL g3089 ( 
.A(n_3065),
.Y(n_3089)
);

INVx1_ASAP7_75t_L g3090 ( 
.A(n_3067),
.Y(n_3090)
);

NOR2x1_ASAP7_75t_L g3091 ( 
.A(n_3055),
.B(n_340),
.Y(n_3091)
);

NOR2x1_ASAP7_75t_L g3092 ( 
.A(n_3038),
.B(n_340),
.Y(n_3092)
);

AND2x2_ASAP7_75t_L g3093 ( 
.A(n_3035),
.B(n_341),
.Y(n_3093)
);

NOR2xp67_ASAP7_75t_L g3094 ( 
.A(n_3025),
.B(n_3040),
.Y(n_3094)
);

NAND4xp75_ASAP7_75t_L g3095 ( 
.A(n_3022),
.B(n_344),
.C(n_342),
.D(n_343),
.Y(n_3095)
);

NOR2x1_ASAP7_75t_L g3096 ( 
.A(n_3028),
.B(n_342),
.Y(n_3096)
);

NAND3x1_ASAP7_75t_L g3097 ( 
.A(n_3018),
.B(n_343),
.C(n_344),
.Y(n_3097)
);

NOR2x1_ASAP7_75t_L g3098 ( 
.A(n_3031),
.B(n_345),
.Y(n_3098)
);

NAND3xp33_ASAP7_75t_L g3099 ( 
.A(n_3030),
.B(n_345),
.C(n_346),
.Y(n_3099)
);

NOR2x1_ASAP7_75t_L g3100 ( 
.A(n_3058),
.B(n_346),
.Y(n_3100)
);

AOI21xp5_ASAP7_75t_L g3101 ( 
.A1(n_3046),
.A2(n_347),
.B(n_349),
.Y(n_3101)
);

NOR3xp33_ASAP7_75t_L g3102 ( 
.A(n_3043),
.B(n_357),
.C(n_347),
.Y(n_3102)
);

OR2x2_ASAP7_75t_L g3103 ( 
.A(n_3034),
.B(n_350),
.Y(n_3103)
);

NOR3xp33_ASAP7_75t_L g3104 ( 
.A(n_3045),
.B(n_358),
.C(n_350),
.Y(n_3104)
);

NAND4xp75_ASAP7_75t_L g3105 ( 
.A(n_3042),
.B(n_353),
.C(n_351),
.D(n_352),
.Y(n_3105)
);

INVx2_ASAP7_75t_L g3106 ( 
.A(n_3026),
.Y(n_3106)
);

INVx2_ASAP7_75t_L g3107 ( 
.A(n_3054),
.Y(n_3107)
);

INVxp33_ASAP7_75t_SL g3108 ( 
.A(n_3029),
.Y(n_3108)
);

AND2x4_ASAP7_75t_L g3109 ( 
.A(n_3049),
.B(n_351),
.Y(n_3109)
);

NAND2xp5_ASAP7_75t_L g3110 ( 
.A(n_3044),
.B(n_353),
.Y(n_3110)
);

BUFx12f_ASAP7_75t_L g3111 ( 
.A(n_3053),
.Y(n_3111)
);

NAND2xp5_ASAP7_75t_SL g3112 ( 
.A(n_3032),
.B(n_354),
.Y(n_3112)
);

INVx1_ASAP7_75t_L g3113 ( 
.A(n_3027),
.Y(n_3113)
);

NAND4xp75_ASAP7_75t_L g3114 ( 
.A(n_3021),
.B(n_357),
.C(n_355),
.D(n_356),
.Y(n_3114)
);

NOR2xp33_ASAP7_75t_L g3115 ( 
.A(n_3050),
.B(n_359),
.Y(n_3115)
);

NAND4xp75_ASAP7_75t_L g3116 ( 
.A(n_3036),
.B(n_361),
.C(n_359),
.D(n_360),
.Y(n_3116)
);

NOR4xp75_ASAP7_75t_L g3117 ( 
.A(n_3024),
.B(n_363),
.C(n_361),
.D(n_362),
.Y(n_3117)
);

NOR3xp33_ASAP7_75t_L g3118 ( 
.A(n_3039),
.B(n_370),
.C(n_362),
.Y(n_3118)
);

NOR2xp33_ASAP7_75t_L g3119 ( 
.A(n_3023),
.B(n_363),
.Y(n_3119)
);

OAI211xp5_ASAP7_75t_L g3120 ( 
.A1(n_3025),
.A2(n_366),
.B(n_364),
.C(n_365),
.Y(n_3120)
);

OR2x2_ASAP7_75t_L g3121 ( 
.A(n_3019),
.B(n_367),
.Y(n_3121)
);

NOR3xp33_ASAP7_75t_SL g3122 ( 
.A(n_3024),
.B(n_367),
.C(n_368),
.Y(n_3122)
);

NOR3xp33_ASAP7_75t_L g3123 ( 
.A(n_3039),
.B(n_376),
.C(n_368),
.Y(n_3123)
);

OR2x2_ASAP7_75t_L g3124 ( 
.A(n_3019),
.B(n_369),
.Y(n_3124)
);

NAND2xp5_ASAP7_75t_L g3125 ( 
.A(n_3056),
.B(n_369),
.Y(n_3125)
);

NOR2x1_ASAP7_75t_L g3126 ( 
.A(n_3037),
.B(n_370),
.Y(n_3126)
);

NAND3x1_ASAP7_75t_SL g3127 ( 
.A(n_3036),
.B(n_371),
.C(n_372),
.Y(n_3127)
);

CKINVDCx12_ASAP7_75t_R g3128 ( 
.A(n_3056),
.Y(n_3128)
);

INVx2_ASAP7_75t_L g3129 ( 
.A(n_3056),
.Y(n_3129)
);

NAND2xp5_ASAP7_75t_L g3130 ( 
.A(n_3056),
.B(n_371),
.Y(n_3130)
);

NAND2xp5_ASAP7_75t_L g3131 ( 
.A(n_3075),
.B(n_373),
.Y(n_3131)
);

INVxp67_ASAP7_75t_L g3132 ( 
.A(n_3073),
.Y(n_3132)
);

NOR2x1_ASAP7_75t_L g3133 ( 
.A(n_3084),
.B(n_372),
.Y(n_3133)
);

NOR2xp33_ASAP7_75t_L g3134 ( 
.A(n_3083),
.B(n_373),
.Y(n_3134)
);

OAI221xp5_ASAP7_75t_L g3135 ( 
.A1(n_3069),
.A2(n_377),
.B1(n_374),
.B2(n_375),
.C(n_378),
.Y(n_3135)
);

NAND2xp5_ASAP7_75t_L g3136 ( 
.A(n_3082),
.B(n_375),
.Y(n_3136)
);

NAND4xp25_ASAP7_75t_L g3137 ( 
.A(n_3094),
.B(n_380),
.C(n_374),
.D(n_379),
.Y(n_3137)
);

XNOR2xp5_ASAP7_75t_SL g3138 ( 
.A(n_3068),
.B(n_381),
.Y(n_3138)
);

NOR4xp75_ASAP7_75t_L g3139 ( 
.A(n_3097),
.B(n_382),
.C(n_380),
.D(n_381),
.Y(n_3139)
);

NAND2xp33_ASAP7_75t_SL g3140 ( 
.A(n_3070),
.B(n_382),
.Y(n_3140)
);

NAND4xp25_ASAP7_75t_L g3141 ( 
.A(n_3078),
.B(n_385),
.C(n_383),
.D(n_384),
.Y(n_3141)
);

AOI211xp5_ASAP7_75t_L g3142 ( 
.A1(n_3120),
.A2(n_3119),
.B(n_3102),
.C(n_3118),
.Y(n_3142)
);

NOR3xp33_ASAP7_75t_SL g3143 ( 
.A(n_3112),
.B(n_384),
.C(n_385),
.Y(n_3143)
);

NOR2xp67_ASAP7_75t_L g3144 ( 
.A(n_3111),
.B(n_386),
.Y(n_3144)
);

OAI221xp5_ASAP7_75t_L g3145 ( 
.A1(n_3079),
.A2(n_388),
.B1(n_386),
.B2(n_387),
.C(n_389),
.Y(n_3145)
);

AOI22xp5_ASAP7_75t_L g3146 ( 
.A1(n_3076),
.A2(n_390),
.B1(n_387),
.B2(n_388),
.Y(n_3146)
);

AOI22xp5_ASAP7_75t_L g3147 ( 
.A1(n_3071),
.A2(n_393),
.B1(n_391),
.B2(n_392),
.Y(n_3147)
);

INVx1_ASAP7_75t_L g3148 ( 
.A(n_3121),
.Y(n_3148)
);

AOI22xp5_ASAP7_75t_L g3149 ( 
.A1(n_3093),
.A2(n_395),
.B1(n_392),
.B2(n_394),
.Y(n_3149)
);

OR2x2_ASAP7_75t_L g3150 ( 
.A(n_3125),
.B(n_394),
.Y(n_3150)
);

NOR2x1_ASAP7_75t_L g3151 ( 
.A(n_3116),
.B(n_395),
.Y(n_3151)
);

OR2x2_ASAP7_75t_L g3152 ( 
.A(n_3130),
.B(n_396),
.Y(n_3152)
);

INVx1_ASAP7_75t_L g3153 ( 
.A(n_3124),
.Y(n_3153)
);

INVx1_ASAP7_75t_L g3154 ( 
.A(n_3085),
.Y(n_3154)
);

INVx1_ASAP7_75t_L g3155 ( 
.A(n_3085),
.Y(n_3155)
);

INVxp67_ASAP7_75t_SL g3156 ( 
.A(n_3087),
.Y(n_3156)
);

NOR2x1_ASAP7_75t_L g3157 ( 
.A(n_3105),
.B(n_397),
.Y(n_3157)
);

OAI21xp33_ASAP7_75t_L g3158 ( 
.A1(n_3108),
.A2(n_3122),
.B(n_3077),
.Y(n_3158)
);

AND3x4_ASAP7_75t_L g3159 ( 
.A(n_3091),
.B(n_397),
.C(n_398),
.Y(n_3159)
);

NOR3xp33_ASAP7_75t_SL g3160 ( 
.A(n_3081),
.B(n_398),
.C(n_399),
.Y(n_3160)
);

NOR3xp33_ASAP7_75t_L g3161 ( 
.A(n_3127),
.B(n_401),
.C(n_400),
.Y(n_3161)
);

NAND2xp5_ASAP7_75t_L g3162 ( 
.A(n_3092),
.B(n_400),
.Y(n_3162)
);

AOI322xp5_ASAP7_75t_L g3163 ( 
.A1(n_3089),
.A2(n_405),
.A3(n_404),
.B1(n_402),
.B2(n_406),
.C1(n_401),
.C2(n_403),
.Y(n_3163)
);

NOR2x1_ASAP7_75t_L g3164 ( 
.A(n_3080),
.B(n_399),
.Y(n_3164)
);

HB1xp67_ASAP7_75t_L g3165 ( 
.A(n_3117),
.Y(n_3165)
);

AOI22xp5_ASAP7_75t_L g3166 ( 
.A1(n_3106),
.A2(n_407),
.B1(n_403),
.B2(n_406),
.Y(n_3166)
);

AND2x4_ASAP7_75t_L g3167 ( 
.A(n_3126),
.B(n_407),
.Y(n_3167)
);

AOI31xp33_ASAP7_75t_L g3168 ( 
.A1(n_3100),
.A2(n_410),
.A3(n_408),
.B(n_409),
.Y(n_3168)
);

NAND3xp33_ASAP7_75t_L g3169 ( 
.A(n_3123),
.B(n_410),
.C(n_411),
.Y(n_3169)
);

BUFx2_ASAP7_75t_L g3170 ( 
.A(n_3098),
.Y(n_3170)
);

NAND5xp2_ASAP7_75t_L g3171 ( 
.A(n_3113),
.B(n_413),
.C(n_415),
.D(n_412),
.E(n_414),
.Y(n_3171)
);

AOI221xp5_ASAP7_75t_L g3172 ( 
.A1(n_3115),
.A2(n_416),
.B1(n_411),
.B2(n_413),
.C(n_417),
.Y(n_3172)
);

NOR2xp67_ASAP7_75t_L g3173 ( 
.A(n_3099),
.B(n_417),
.Y(n_3173)
);

AND3x4_ASAP7_75t_L g3174 ( 
.A(n_3096),
.B(n_418),
.C(n_419),
.Y(n_3174)
);

AND2x2_ASAP7_75t_L g3175 ( 
.A(n_3129),
.B(n_418),
.Y(n_3175)
);

NAND4xp75_ASAP7_75t_L g3176 ( 
.A(n_3110),
.B(n_421),
.C(n_419),
.D(n_420),
.Y(n_3176)
);

NOR2xp33_ASAP7_75t_L g3177 ( 
.A(n_3095),
.B(n_420),
.Y(n_3177)
);

NAND4xp25_ASAP7_75t_L g3178 ( 
.A(n_3074),
.B(n_423),
.C(n_421),
.D(n_422),
.Y(n_3178)
);

NOR2x1_ASAP7_75t_SL g3179 ( 
.A(n_3114),
.B(n_424),
.Y(n_3179)
);

NOR3xp33_ASAP7_75t_SL g3180 ( 
.A(n_3072),
.B(n_422),
.C(n_425),
.Y(n_3180)
);

AOI31xp33_ASAP7_75t_L g3181 ( 
.A1(n_3103),
.A2(n_428),
.A3(n_426),
.B(n_427),
.Y(n_3181)
);

NAND2xp5_ASAP7_75t_L g3182 ( 
.A(n_3088),
.B(n_428),
.Y(n_3182)
);

NOR3xp33_ASAP7_75t_L g3183 ( 
.A(n_3104),
.B(n_430),
.C(n_429),
.Y(n_3183)
);

AOI221xp5_ASAP7_75t_L g3184 ( 
.A1(n_3101),
.A2(n_430),
.B1(n_426),
.B2(n_429),
.C(n_431),
.Y(n_3184)
);

NOR2xp33_ASAP7_75t_L g3185 ( 
.A(n_3128),
.B(n_432),
.Y(n_3185)
);

OR2x2_ASAP7_75t_L g3186 ( 
.A(n_3107),
.B(n_432),
.Y(n_3186)
);

NOR3xp33_ASAP7_75t_L g3187 ( 
.A(n_3086),
.B(n_435),
.C(n_434),
.Y(n_3187)
);

NAND3xp33_ASAP7_75t_L g3188 ( 
.A(n_3109),
.B(n_3090),
.C(n_433),
.Y(n_3188)
);

HB1xp67_ASAP7_75t_L g3189 ( 
.A(n_3109),
.Y(n_3189)
);

OR2x2_ASAP7_75t_L g3190 ( 
.A(n_3069),
.B(n_433),
.Y(n_3190)
);

INVx1_ASAP7_75t_L g3191 ( 
.A(n_3073),
.Y(n_3191)
);

XOR2xp5_ASAP7_75t_L g3192 ( 
.A(n_3116),
.B(n_434),
.Y(n_3192)
);

NAND2xp5_ASAP7_75t_L g3193 ( 
.A(n_3144),
.B(n_435),
.Y(n_3193)
);

INVxp67_ASAP7_75t_L g3194 ( 
.A(n_3171),
.Y(n_3194)
);

XNOR2x1_ASAP7_75t_L g3195 ( 
.A(n_3159),
.B(n_436),
.Y(n_3195)
);

OAI22x1_ASAP7_75t_L g3196 ( 
.A1(n_3174),
.A2(n_438),
.B1(n_439),
.B2(n_437),
.Y(n_3196)
);

INVx1_ASAP7_75t_SL g3197 ( 
.A(n_3139),
.Y(n_3197)
);

INVx1_ASAP7_75t_L g3198 ( 
.A(n_3138),
.Y(n_3198)
);

AOI22xp5_ASAP7_75t_L g3199 ( 
.A1(n_3140),
.A2(n_444),
.B1(n_453),
.B2(n_436),
.Y(n_3199)
);

OR2x2_ASAP7_75t_L g3200 ( 
.A(n_3137),
.B(n_437),
.Y(n_3200)
);

NAND2xp5_ASAP7_75t_L g3201 ( 
.A(n_3175),
.B(n_438),
.Y(n_3201)
);

XOR2x1_ASAP7_75t_L g3202 ( 
.A(n_3167),
.B(n_439),
.Y(n_3202)
);

AOI22xp5_ASAP7_75t_L g3203 ( 
.A1(n_3185),
.A2(n_450),
.B1(n_440),
.B2(n_442),
.Y(n_3203)
);

INVx1_ASAP7_75t_L g3204 ( 
.A(n_3167),
.Y(n_3204)
);

INVx2_ASAP7_75t_L g3205 ( 
.A(n_3186),
.Y(n_3205)
);

INVxp67_ASAP7_75t_SL g3206 ( 
.A(n_3164),
.Y(n_3206)
);

AO22x1_ASAP7_75t_L g3207 ( 
.A1(n_3151),
.A2(n_443),
.B1(n_441),
.B2(n_442),
.Y(n_3207)
);

AND2x4_ASAP7_75t_L g3208 ( 
.A(n_3154),
.B(n_441),
.Y(n_3208)
);

INVx1_ASAP7_75t_L g3209 ( 
.A(n_3192),
.Y(n_3209)
);

OAI22xp5_ASAP7_75t_L g3210 ( 
.A1(n_3190),
.A2(n_3135),
.B1(n_3169),
.B2(n_3156),
.Y(n_3210)
);

XNOR2xp5_ASAP7_75t_L g3211 ( 
.A(n_3165),
.B(n_3176),
.Y(n_3211)
);

INVx1_ASAP7_75t_SL g3212 ( 
.A(n_3170),
.Y(n_3212)
);

INVx2_ASAP7_75t_L g3213 ( 
.A(n_3150),
.Y(n_3213)
);

OAI22xp5_ASAP7_75t_SL g3214 ( 
.A1(n_3155),
.A2(n_447),
.B1(n_443),
.B2(n_445),
.Y(n_3214)
);

AND2x4_ASAP7_75t_L g3215 ( 
.A(n_3191),
.B(n_3132),
.Y(n_3215)
);

INVx1_ASAP7_75t_L g3216 ( 
.A(n_3136),
.Y(n_3216)
);

INVx1_ASAP7_75t_L g3217 ( 
.A(n_3131),
.Y(n_3217)
);

OAI22xp5_ASAP7_75t_L g3218 ( 
.A1(n_3145),
.A2(n_449),
.B1(n_447),
.B2(n_448),
.Y(n_3218)
);

XNOR2x1_ASAP7_75t_L g3219 ( 
.A(n_3133),
.B(n_449),
.Y(n_3219)
);

INVx1_ASAP7_75t_L g3220 ( 
.A(n_3134),
.Y(n_3220)
);

INVx1_ASAP7_75t_L g3221 ( 
.A(n_3168),
.Y(n_3221)
);

NAND4xp75_ASAP7_75t_L g3222 ( 
.A(n_3157),
.B(n_452),
.C(n_450),
.D(n_451),
.Y(n_3222)
);

INVx1_ASAP7_75t_L g3223 ( 
.A(n_3162),
.Y(n_3223)
);

INVx1_ASAP7_75t_L g3224 ( 
.A(n_3181),
.Y(n_3224)
);

INVx3_ASAP7_75t_L g3225 ( 
.A(n_3152),
.Y(n_3225)
);

NAND4xp75_ASAP7_75t_L g3226 ( 
.A(n_3173),
.B(n_456),
.C(n_451),
.D(n_455),
.Y(n_3226)
);

XNOR2xp5_ASAP7_75t_L g3227 ( 
.A(n_3141),
.B(n_539),
.Y(n_3227)
);

NOR2x1_ASAP7_75t_L g3228 ( 
.A(n_3178),
.B(n_540),
.Y(n_3228)
);

NAND2xp5_ASAP7_75t_L g3229 ( 
.A(n_3161),
.B(n_541),
.Y(n_3229)
);

OAI31xp67_ASAP7_75t_L g3230 ( 
.A1(n_3158),
.A2(n_547),
.A3(n_543),
.B(n_545),
.Y(n_3230)
);

INVx1_ASAP7_75t_L g3231 ( 
.A(n_3179),
.Y(n_3231)
);

INVxp67_ASAP7_75t_L g3232 ( 
.A(n_3177),
.Y(n_3232)
);

AND3x4_ASAP7_75t_L g3233 ( 
.A(n_3143),
.B(n_560),
.C(n_549),
.Y(n_3233)
);

NAND4xp75_ASAP7_75t_L g3234 ( 
.A(n_3182),
.B(n_900),
.C(n_902),
.D(n_899),
.Y(n_3234)
);

OR2x2_ASAP7_75t_L g3235 ( 
.A(n_3148),
.B(n_550),
.Y(n_3235)
);

NAND2xp5_ASAP7_75t_L g3236 ( 
.A(n_3147),
.B(n_552),
.Y(n_3236)
);

OR2x2_ASAP7_75t_L g3237 ( 
.A(n_3153),
.B(n_553),
.Y(n_3237)
);

OAI22xp5_ASAP7_75t_SL g3238 ( 
.A1(n_3188),
.A2(n_557),
.B1(n_554),
.B2(n_555),
.Y(n_3238)
);

INVx1_ASAP7_75t_L g3239 ( 
.A(n_3189),
.Y(n_3239)
);

AND2x2_ASAP7_75t_L g3240 ( 
.A(n_3160),
.B(n_558),
.Y(n_3240)
);

OAI22xp5_ASAP7_75t_L g3241 ( 
.A1(n_3142),
.A2(n_564),
.B1(n_562),
.B2(n_563),
.Y(n_3241)
);

INVx1_ASAP7_75t_L g3242 ( 
.A(n_3180),
.Y(n_3242)
);

AOI211xp5_ASAP7_75t_SL g3243 ( 
.A1(n_3210),
.A2(n_3239),
.B(n_3194),
.C(n_3231),
.Y(n_3243)
);

OAI21xp5_ASAP7_75t_L g3244 ( 
.A1(n_3195),
.A2(n_3183),
.B(n_3184),
.Y(n_3244)
);

INVx2_ASAP7_75t_L g3245 ( 
.A(n_3202),
.Y(n_3245)
);

OA22x2_ASAP7_75t_L g3246 ( 
.A1(n_3199),
.A2(n_3149),
.B1(n_3146),
.B2(n_3166),
.Y(n_3246)
);

AO22x2_ASAP7_75t_L g3247 ( 
.A1(n_3222),
.A2(n_3187),
.B1(n_3172),
.B2(n_3163),
.Y(n_3247)
);

OAI21xp33_ASAP7_75t_L g3248 ( 
.A1(n_3212),
.A2(n_3211),
.B(n_3197),
.Y(n_3248)
);

OAI22xp5_ASAP7_75t_L g3249 ( 
.A1(n_3200),
.A2(n_567),
.B1(n_565),
.B2(n_566),
.Y(n_3249)
);

INVx2_ASAP7_75t_L g3250 ( 
.A(n_3208),
.Y(n_3250)
);

BUFx6f_ASAP7_75t_L g3251 ( 
.A(n_3215),
.Y(n_3251)
);

OR2x6_ASAP7_75t_L g3252 ( 
.A(n_3204),
.B(n_568),
.Y(n_3252)
);

INVx1_ASAP7_75t_L g3253 ( 
.A(n_3193),
.Y(n_3253)
);

INVxp67_ASAP7_75t_SL g3254 ( 
.A(n_3196),
.Y(n_3254)
);

HB1xp67_ASAP7_75t_L g3255 ( 
.A(n_3226),
.Y(n_3255)
);

AOI22xp5_ASAP7_75t_L g3256 ( 
.A1(n_3233),
.A2(n_573),
.B1(n_570),
.B2(n_572),
.Y(n_3256)
);

AOI221xp5_ASAP7_75t_L g3257 ( 
.A1(n_3207),
.A2(n_576),
.B1(n_574),
.B2(n_575),
.C(n_577),
.Y(n_3257)
);

CKINVDCx20_ASAP7_75t_R g3258 ( 
.A(n_3209),
.Y(n_3258)
);

AND3x2_ASAP7_75t_L g3259 ( 
.A(n_3206),
.B(n_580),
.C(n_579),
.Y(n_3259)
);

INVx1_ASAP7_75t_SL g3260 ( 
.A(n_3219),
.Y(n_3260)
);

HB1xp67_ASAP7_75t_L g3261 ( 
.A(n_3214),
.Y(n_3261)
);

XNOR2xp5_ASAP7_75t_L g3262 ( 
.A(n_3227),
.B(n_3228),
.Y(n_3262)
);

AOI22xp5_ASAP7_75t_L g3263 ( 
.A1(n_3221),
.A2(n_584),
.B1(n_578),
.B2(n_581),
.Y(n_3263)
);

AOI221x1_ASAP7_75t_L g3264 ( 
.A1(n_3224),
.A2(n_587),
.B1(n_585),
.B2(n_586),
.C(n_590),
.Y(n_3264)
);

XNOR2xp5_ASAP7_75t_L g3265 ( 
.A(n_3242),
.B(n_591),
.Y(n_3265)
);

NAND2xp5_ASAP7_75t_L g3266 ( 
.A(n_3203),
.B(n_593),
.Y(n_3266)
);

OA21x2_ASAP7_75t_L g3267 ( 
.A1(n_3201),
.A2(n_594),
.B(n_596),
.Y(n_3267)
);

NAND2xp5_ASAP7_75t_L g3268 ( 
.A(n_3240),
.B(n_597),
.Y(n_3268)
);

HB1xp67_ASAP7_75t_L g3269 ( 
.A(n_3234),
.Y(n_3269)
);

OAI22xp5_ASAP7_75t_SL g3270 ( 
.A1(n_3198),
.A2(n_601),
.B1(n_598),
.B2(n_599),
.Y(n_3270)
);

INVx5_ASAP7_75t_L g3271 ( 
.A(n_3225),
.Y(n_3271)
);

AOI21xp5_ASAP7_75t_L g3272 ( 
.A1(n_3229),
.A2(n_602),
.B(n_603),
.Y(n_3272)
);

OAI211xp5_ASAP7_75t_L g3273 ( 
.A1(n_3232),
.A2(n_889),
.B(n_890),
.C(n_888),
.Y(n_3273)
);

INVx1_ASAP7_75t_SL g3274 ( 
.A(n_3235),
.Y(n_3274)
);

INVx2_ASAP7_75t_L g3275 ( 
.A(n_3237),
.Y(n_3275)
);

AND2x2_ASAP7_75t_L g3276 ( 
.A(n_3205),
.B(n_604),
.Y(n_3276)
);

NAND3xp33_ASAP7_75t_L g3277 ( 
.A(n_3218),
.B(n_607),
.C(n_608),
.Y(n_3277)
);

OAI22xp5_ASAP7_75t_L g3278 ( 
.A1(n_3220),
.A2(n_613),
.B1(n_609),
.B2(n_610),
.Y(n_3278)
);

INVx1_ASAP7_75t_L g3279 ( 
.A(n_3236),
.Y(n_3279)
);

OAI22x1_ASAP7_75t_L g3280 ( 
.A1(n_3213),
.A2(n_616),
.B1(n_614),
.B2(n_615),
.Y(n_3280)
);

AND3x2_ASAP7_75t_L g3281 ( 
.A(n_3223),
.B(n_619),
.C(n_618),
.Y(n_3281)
);

HB1xp67_ASAP7_75t_L g3282 ( 
.A(n_3238),
.Y(n_3282)
);

NAND2xp5_ASAP7_75t_L g3283 ( 
.A(n_3216),
.B(n_3217),
.Y(n_3283)
);

AND2x2_ASAP7_75t_L g3284 ( 
.A(n_3230),
.B(n_617),
.Y(n_3284)
);

INVx1_ASAP7_75t_L g3285 ( 
.A(n_3241),
.Y(n_3285)
);

INVx2_ASAP7_75t_L g3286 ( 
.A(n_3202),
.Y(n_3286)
);

AOI22xp5_ASAP7_75t_L g3287 ( 
.A1(n_3258),
.A2(n_622),
.B1(n_620),
.B2(n_621),
.Y(n_3287)
);

INVx1_ASAP7_75t_L g3288 ( 
.A(n_3251),
.Y(n_3288)
);

OAI211xp5_ASAP7_75t_SL g3289 ( 
.A1(n_3243),
.A2(n_3248),
.B(n_3244),
.C(n_3260),
.Y(n_3289)
);

INVx2_ASAP7_75t_SL g3290 ( 
.A(n_3271),
.Y(n_3290)
);

OAI22xp5_ASAP7_75t_L g3291 ( 
.A1(n_3271),
.A2(n_626),
.B1(n_624),
.B2(n_625),
.Y(n_3291)
);

AOI221xp5_ASAP7_75t_L g3292 ( 
.A1(n_3251),
.A2(n_633),
.B1(n_628),
.B2(n_629),
.C(n_634),
.Y(n_3292)
);

OAI22xp5_ASAP7_75t_L g3293 ( 
.A1(n_3256),
.A2(n_637),
.B1(n_635),
.B2(n_636),
.Y(n_3293)
);

NAND3xp33_ASAP7_75t_SL g3294 ( 
.A(n_3257),
.B(n_638),
.C(n_639),
.Y(n_3294)
);

INVx1_ASAP7_75t_L g3295 ( 
.A(n_3261),
.Y(n_3295)
);

INVx2_ASAP7_75t_L g3296 ( 
.A(n_3259),
.Y(n_3296)
);

AND2x4_ASAP7_75t_L g3297 ( 
.A(n_3250),
.B(n_641),
.Y(n_3297)
);

OAI22xp33_ASAP7_75t_L g3298 ( 
.A1(n_3245),
.A2(n_645),
.B1(n_642),
.B2(n_643),
.Y(n_3298)
);

AOI222xp33_ASAP7_75t_L g3299 ( 
.A1(n_3254),
.A2(n_652),
.B1(n_654),
.B2(n_649),
.C1(n_650),
.C2(n_653),
.Y(n_3299)
);

AO22x2_ASAP7_75t_L g3300 ( 
.A1(n_3286),
.A2(n_657),
.B1(n_655),
.B2(n_656),
.Y(n_3300)
);

AOI322xp5_ASAP7_75t_L g3301 ( 
.A1(n_3255),
.A2(n_665),
.A3(n_664),
.B1(n_661),
.B2(n_659),
.C1(n_660),
.C2(n_662),
.Y(n_3301)
);

XOR2xp5_ASAP7_75t_L g3302 ( 
.A(n_3262),
.B(n_666),
.Y(n_3302)
);

NAND4xp75_ASAP7_75t_L g3303 ( 
.A(n_3268),
.B(n_669),
.C(n_667),
.D(n_668),
.Y(n_3303)
);

NAND3xp33_ASAP7_75t_L g3304 ( 
.A(n_3272),
.B(n_670),
.C(n_671),
.Y(n_3304)
);

AOI22xp5_ASAP7_75t_L g3305 ( 
.A1(n_3284),
.A2(n_678),
.B1(n_675),
.B2(n_677),
.Y(n_3305)
);

OAI22xp5_ASAP7_75t_L g3306 ( 
.A1(n_3288),
.A2(n_3277),
.B1(n_3274),
.B2(n_3266),
.Y(n_3306)
);

AOI22xp5_ASAP7_75t_L g3307 ( 
.A1(n_3289),
.A2(n_3247),
.B1(n_3246),
.B2(n_3275),
.Y(n_3307)
);

OAI221xp5_ASAP7_75t_L g3308 ( 
.A1(n_3290),
.A2(n_3283),
.B1(n_3269),
.B2(n_3282),
.C(n_3285),
.Y(n_3308)
);

XNOR2xp5_ASAP7_75t_L g3309 ( 
.A(n_3305),
.B(n_3265),
.Y(n_3309)
);

NAND2xp5_ASAP7_75t_L g3310 ( 
.A(n_3295),
.B(n_3276),
.Y(n_3310)
);

NOR3xp33_ASAP7_75t_L g3311 ( 
.A(n_3296),
.B(n_3253),
.C(n_3279),
.Y(n_3311)
);

A2O1A1Ixp33_ASAP7_75t_L g3312 ( 
.A1(n_3304),
.A2(n_3273),
.B(n_3249),
.C(n_3263),
.Y(n_3312)
);

INVx1_ASAP7_75t_L g3313 ( 
.A(n_3302),
.Y(n_3313)
);

NOR3xp33_ASAP7_75t_L g3314 ( 
.A(n_3294),
.B(n_3270),
.C(n_3278),
.Y(n_3314)
);

OAI22xp5_ASAP7_75t_SL g3315 ( 
.A1(n_3293),
.A2(n_3267),
.B1(n_3252),
.B2(n_3280),
.Y(n_3315)
);

OAI221xp5_ASAP7_75t_L g3316 ( 
.A1(n_3299),
.A2(n_3252),
.B1(n_3281),
.B2(n_3264),
.C(n_681),
.Y(n_3316)
);

NOR4xp25_ASAP7_75t_L g3317 ( 
.A(n_3298),
.B(n_682),
.C(n_679),
.D(n_680),
.Y(n_3317)
);

AOI21xp33_ASAP7_75t_L g3318 ( 
.A1(n_3291),
.A2(n_683),
.B(n_684),
.Y(n_3318)
);

AND3x1_ASAP7_75t_L g3319 ( 
.A(n_3292),
.B(n_685),
.C(n_686),
.Y(n_3319)
);

NAND2xp5_ASAP7_75t_L g3320 ( 
.A(n_3297),
.B(n_687),
.Y(n_3320)
);

AOI21xp5_ASAP7_75t_L g3321 ( 
.A1(n_3308),
.A2(n_3300),
.B(n_3287),
.Y(n_3321)
);

AO22x2_ASAP7_75t_L g3322 ( 
.A1(n_3306),
.A2(n_3303),
.B1(n_3300),
.B2(n_3301),
.Y(n_3322)
);

OR2x6_ASAP7_75t_L g3323 ( 
.A(n_3310),
.B(n_3313),
.Y(n_3323)
);

INVx2_ASAP7_75t_L g3324 ( 
.A(n_3320),
.Y(n_3324)
);

INVx2_ASAP7_75t_L g3325 ( 
.A(n_3319),
.Y(n_3325)
);

AOI221xp5_ASAP7_75t_L g3326 ( 
.A1(n_3317),
.A2(n_3316),
.B1(n_3318),
.B2(n_3311),
.C(n_3315),
.Y(n_3326)
);

OAI32xp33_ASAP7_75t_L g3327 ( 
.A1(n_3314),
.A2(n_692),
.A3(n_689),
.B1(n_690),
.B2(n_696),
.Y(n_3327)
);

NAND2xp5_ASAP7_75t_L g3328 ( 
.A(n_3307),
.B(n_698),
.Y(n_3328)
);

AND2x2_ASAP7_75t_L g3329 ( 
.A(n_3312),
.B(n_700),
.Y(n_3329)
);

INVx4_ASAP7_75t_L g3330 ( 
.A(n_3309),
.Y(n_3330)
);

INVx1_ASAP7_75t_L g3331 ( 
.A(n_3320),
.Y(n_3331)
);

AOI211xp5_ASAP7_75t_L g3332 ( 
.A1(n_3308),
.A2(n_707),
.B(n_702),
.C(n_704),
.Y(n_3332)
);

OAI22xp5_ASAP7_75t_L g3333 ( 
.A1(n_3307),
.A2(n_710),
.B1(n_708),
.B2(n_709),
.Y(n_3333)
);

NAND4xp75_ASAP7_75t_L g3334 ( 
.A(n_3329),
.B(n_714),
.C(n_712),
.D(n_713),
.Y(n_3334)
);

XNOR2xp5_ASAP7_75t_L g3335 ( 
.A(n_3322),
.B(n_715),
.Y(n_3335)
);

OAI22xp5_ASAP7_75t_L g3336 ( 
.A1(n_3328),
.A2(n_719),
.B1(n_716),
.B2(n_718),
.Y(n_3336)
);

INVx2_ASAP7_75t_L g3337 ( 
.A(n_3325),
.Y(n_3337)
);

NOR2xp67_ASAP7_75t_L g3338 ( 
.A(n_3321),
.B(n_722),
.Y(n_3338)
);

INVx4_ASAP7_75t_L g3339 ( 
.A(n_3323),
.Y(n_3339)
);

AOI22xp5_ASAP7_75t_L g3340 ( 
.A1(n_3333),
.A2(n_725),
.B1(n_723),
.B2(n_724),
.Y(n_3340)
);

NAND2xp5_ASAP7_75t_L g3341 ( 
.A(n_3332),
.B(n_726),
.Y(n_3341)
);

XOR2xp5_ASAP7_75t_L g3342 ( 
.A(n_3331),
.B(n_907),
.Y(n_3342)
);

OR2x6_ASAP7_75t_L g3343 ( 
.A(n_3330),
.B(n_728),
.Y(n_3343)
);

NAND3xp33_ASAP7_75t_L g3344 ( 
.A(n_3326),
.B(n_729),
.C(n_730),
.Y(n_3344)
);

INVx1_ASAP7_75t_L g3345 ( 
.A(n_3324),
.Y(n_3345)
);

OAI22xp5_ASAP7_75t_L g3346 ( 
.A1(n_3339),
.A2(n_3327),
.B1(n_733),
.B2(n_731),
.Y(n_3346)
);

OAI22x1_ASAP7_75t_L g3347 ( 
.A1(n_3335),
.A2(n_735),
.B1(n_732),
.B2(n_734),
.Y(n_3347)
);

AOI21xp33_ASAP7_75t_L g3348 ( 
.A1(n_3345),
.A2(n_736),
.B(n_739),
.Y(n_3348)
);

AOI22xp5_ASAP7_75t_L g3349 ( 
.A1(n_3338),
.A2(n_744),
.B1(n_741),
.B2(n_743),
.Y(n_3349)
);

OR2x2_ASAP7_75t_L g3350 ( 
.A(n_3344),
.B(n_746),
.Y(n_3350)
);

OAI22xp5_ASAP7_75t_SL g3351 ( 
.A1(n_3343),
.A2(n_751),
.B1(n_747),
.B2(n_749),
.Y(n_3351)
);

AOI22xp5_ASAP7_75t_L g3352 ( 
.A1(n_3337),
.A2(n_755),
.B1(n_752),
.B2(n_754),
.Y(n_3352)
);

NAND2xp5_ASAP7_75t_SL g3353 ( 
.A(n_3349),
.B(n_3340),
.Y(n_3353)
);

AOI22xp33_ASAP7_75t_SL g3354 ( 
.A1(n_3346),
.A2(n_3341),
.B1(n_3336),
.B2(n_3343),
.Y(n_3354)
);

NAND3xp33_ASAP7_75t_L g3355 ( 
.A(n_3350),
.B(n_3334),
.C(n_3342),
.Y(n_3355)
);

AOI22xp33_ASAP7_75t_SL g3356 ( 
.A1(n_3351),
.A2(n_758),
.B1(n_756),
.B2(n_757),
.Y(n_3356)
);

OAI21xp5_ASAP7_75t_L g3357 ( 
.A1(n_3355),
.A2(n_3348),
.B(n_3347),
.Y(n_3357)
);

NAND3xp33_ASAP7_75t_L g3358 ( 
.A(n_3354),
.B(n_3352),
.C(n_759),
.Y(n_3358)
);

XNOR2xp5_ASAP7_75t_L g3359 ( 
.A(n_3353),
.B(n_761),
.Y(n_3359)
);

INVx1_ASAP7_75t_L g3360 ( 
.A(n_3358),
.Y(n_3360)
);

INVx1_ASAP7_75t_SL g3361 ( 
.A(n_3359),
.Y(n_3361)
);

OA21x2_ASAP7_75t_L g3362 ( 
.A1(n_3360),
.A2(n_3357),
.B(n_3356),
.Y(n_3362)
);

AOI221xp5_ASAP7_75t_L g3363 ( 
.A1(n_3362),
.A2(n_3361),
.B1(n_766),
.B2(n_762),
.C(n_763),
.Y(n_3363)
);

AOI211xp5_ASAP7_75t_L g3364 ( 
.A1(n_3363),
.A2(n_772),
.B(n_770),
.C(n_771),
.Y(n_3364)
);


endmodule