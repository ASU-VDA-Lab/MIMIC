module fake_ibex_236_n_977 (n_151, n_147, n_85, n_167, n_128, n_84, n_64, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_177, n_148, n_2, n_76, n_8, n_118, n_183, n_67, n_9, n_164, n_38, n_124, n_37, n_110, n_47, n_169, n_108, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_180, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_172, n_49, n_40, n_66, n_17, n_74, n_90, n_176, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_166, n_163, n_26, n_188, n_114, n_34, n_97, n_102, n_181, n_15, n_131, n_123, n_24, n_52, n_189, n_99, n_135, n_105, n_156, n_126, n_187, n_1, n_154, n_182, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_186, n_50, n_11, n_92, n_144, n_170, n_101, n_113, n_138, n_96, n_185, n_68, n_117, n_79, n_81, n_35, n_159, n_158, n_132, n_174, n_157, n_160, n_184, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_977);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_177;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_183;
input n_67;
input n_9;
input n_164;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_169;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_180;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_172;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_176;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_166;
input n_163;
input n_26;
input n_188;
input n_114;
input n_34;
input n_97;
input n_102;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_189;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_187;
input n_1;
input n_154;
input n_182;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_186;
input n_50;
input n_11;
input n_92;
input n_144;
input n_170;
input n_101;
input n_113;
input n_138;
input n_96;
input n_185;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_159;
input n_158;
input n_132;
input n_174;
input n_157;
input n_160;
input n_184;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_977;

wire n_599;
wire n_778;
wire n_822;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_946;
wire n_707;
wire n_273;
wire n_330;
wire n_309;
wire n_926;
wire n_328;
wire n_293;
wire n_341;
wire n_372;
wire n_256;
wire n_418;
wire n_193;
wire n_510;
wire n_845;
wire n_947;
wire n_972;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_956;
wire n_790;
wire n_920;
wire n_452;
wire n_664;
wire n_255;
wire n_586;
wire n_773;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_191;
wire n_873;
wire n_962;
wire n_593;
wire n_862;
wire n_545;
wire n_909;
wire n_583;
wire n_887;
wire n_957;
wire n_678;
wire n_663;
wire n_969;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_961;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_974;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_357;
wire n_412;
wire n_457;
wire n_494;
wire n_226;
wire n_930;
wire n_336;
wire n_959;
wire n_258;
wire n_861;
wire n_449;
wire n_547;
wire n_727;
wire n_216;
wire n_915;
wire n_911;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_963;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_498;
wire n_708;
wire n_280;
wire n_375;
wire n_340;
wire n_317;
wire n_698;
wire n_901;
wire n_667;
wire n_884;
wire n_682;
wire n_850;
wire n_196;
wire n_327;
wire n_326;
wire n_879;
wire n_723;
wire n_270;
wire n_383;
wire n_346;
wire n_886;
wire n_840;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_948;
wire n_859;
wire n_259;
wire n_339;
wire n_276;
wire n_470;
wire n_770;
wire n_965;
wire n_210;
wire n_348;
wire n_220;
wire n_875;
wire n_941;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_671;
wire n_228;
wire n_711;
wire n_876;
wire n_552;
wire n_384;
wire n_251;
wire n_632;
wire n_373;
wire n_854;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_936;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_533;
wire n_508;
wire n_939;
wire n_453;
wire n_591;
wire n_898;
wire n_655;
wire n_333;
wire n_928;
wire n_967;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_673;
wire n_732;
wire n_798;
wire n_832;
wire n_242;
wire n_278;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_914;
wire n_835;
wire n_526;
wire n_785;
wire n_824;
wire n_929;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_923;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_933;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_938;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_281;
wire n_758;
wire n_594;
wire n_636;
wire n_720;
wire n_710;
wire n_407;
wire n_490;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_944;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_543;
wire n_580;
wire n_483;
wire n_420;
wire n_769;
wire n_487;
wire n_222;
wire n_660;
wire n_524;
wire n_349;
wire n_765;
wire n_849;
wire n_857;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_917;
wire n_388;
wire n_953;
wire n_625;
wire n_968;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_931;
wire n_666;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_858;
wire n_207;
wire n_922;
wire n_438;
wire n_851;
wire n_689;
wire n_960;
wire n_793;
wire n_676;
wire n_937;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_973;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_514;
wire n_488;
wire n_705;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_635;
wire n_844;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_847;
wire n_830;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_966;
wire n_359;
wire n_826;
wire n_262;
wire n_299;
wire n_439;
wire n_433;
wire n_704;
wire n_949;
wire n_924;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_696;
wire n_796;
wire n_837;
wire n_797;
wire n_477;
wire n_640;
wire n_954;
wire n_363;
wire n_402;
wire n_725;
wire n_369;
wire n_976;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_935;
wire n_869;
wire n_925;
wire n_718;
wire n_801;
wire n_918;
wire n_672;
wire n_722;
wire n_401;
wire n_553;
wire n_554;
wire n_735;
wire n_305;
wire n_882;
wire n_942;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_605;
wire n_539;
wire n_354;
wire n_206;
wire n_630;
wire n_392;
wire n_516;
wire n_567;
wire n_548;
wire n_943;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_940;
wire n_200;
wire n_444;
wire n_506;
wire n_562;
wire n_564;
wire n_868;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_975;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_927;
wire n_934;
wire n_658;
wire n_512;
wire n_615;
wire n_950;
wire n_685;
wire n_283;
wire n_397;
wire n_366;
wire n_803;
wire n_894;
wire n_692;
wire n_627;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_757;
wire n_248;
wire n_712;
wire n_451;
wire n_702;
wire n_971;
wire n_190;
wire n_906;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_818;
wire n_653;
wire n_214;
wire n_238;
wire n_579;
wire n_843;
wire n_899;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_951;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_919;
wire n_780;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_597;
wire n_415;
wire n_288;
wire n_320;
wire n_247;
wire n_379;
wire n_285;
wire n_551;
wire n_612;
wire n_318;
wire n_291;
wire n_819;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_955;
wire n_385;
wire n_233;
wire n_414;
wire n_342;
wire n_430;
wire n_741;
wire n_729;
wire n_603;
wire n_378;
wire n_486;
wire n_952;
wire n_422;
wire n_264;
wire n_198;
wire n_616;
wire n_782;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_805;
wire n_670;
wire n_820;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_958;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_808;
wire n_250;
wire n_945;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_903;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_885;
wire n_513;
wire n_212;
wire n_588;
wire n_877;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_896;
wire n_197;
wire n_528;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_794;
wire n_836;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_572;
wire n_867;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_897;
wire n_889;
wire n_436;
wire n_428;
wire n_970;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_396;
wire n_252;
wire n_697;
wire n_816;
wire n_890;
wire n_874;
wire n_912;
wire n_921;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_213;
wire n_964;
wire n_424;
wire n_565;
wire n_916;
wire n_823;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_394;
wire n_364;
wire n_687;
wire n_895;
wire n_202;
wire n_298;
wire n_231;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_932;
wire n_657;
wire n_764;
wire n_492;
wire n_649;
wire n_855;
wire n_812;
wire n_232;
wire n_380;
wire n_749;
wire n_866;
wire n_559;
wire n_425;

INVx1_ASAP7_75t_L g190 ( 
.A(n_5),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_167),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_129),
.Y(n_192)
);

INVxp67_ASAP7_75t_SL g193 ( 
.A(n_141),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_182),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_35),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_71),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_105),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_151),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_159),
.Y(n_199)
);

BUFx5_ASAP7_75t_L g200 ( 
.A(n_177),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_64),
.Y(n_201)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_27),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_115),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_13),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_137),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_25),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_59),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_88),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_150),
.Y(n_209)
);

BUFx5_ASAP7_75t_L g210 ( 
.A(n_55),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_50),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_153),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_106),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_49),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_187),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_48),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_112),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_45),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_26),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_176),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_46),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_20),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_8),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_53),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_180),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_83),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_124),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_173),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_73),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_104),
.Y(n_230)
);

INVxp33_ASAP7_75t_SL g231 ( 
.A(n_12),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_128),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_60),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_122),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_15),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_27),
.Y(n_236)
);

INVxp67_ASAP7_75t_SL g237 ( 
.A(n_114),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_107),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_183),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_108),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_161),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_174),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_118),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_188),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_4),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_148),
.B(n_72),
.Y(n_246)
);

CKINVDCx14_ASAP7_75t_R g247 ( 
.A(n_132),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_68),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_6),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_4),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_47),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_85),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_125),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_184),
.B(n_146),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_163),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_157),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_91),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_13),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_29),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_172),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_123),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_15),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_109),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_21),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_149),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_169),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_93),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_74),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_43),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_31),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_144),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_111),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_22),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_103),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_98),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_66),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_37),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_11),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_62),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_28),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_131),
.Y(n_281)
);

INVxp67_ASAP7_75t_SL g282 ( 
.A(n_162),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_22),
.Y(n_283)
);

INVx2_ASAP7_75t_SL g284 ( 
.A(n_97),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_143),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_133),
.Y(n_286)
);

INVx2_ASAP7_75t_SL g287 ( 
.A(n_152),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_119),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_154),
.Y(n_289)
);

NOR2xp67_ASAP7_75t_L g290 ( 
.A(n_36),
.B(n_41),
.Y(n_290)
);

INVx1_ASAP7_75t_SL g291 ( 
.A(n_35),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_79),
.B(n_126),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_175),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_54),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_41),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_142),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_40),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_127),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_16),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_8),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_52),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_70),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_86),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_18),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_145),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_87),
.Y(n_306)
);

INVx2_ASAP7_75t_SL g307 ( 
.A(n_11),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_140),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_136),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g310 ( 
.A(n_96),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_94),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_7),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_138),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_171),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_67),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_147),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_120),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_42),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_158),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_170),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_116),
.Y(n_321)
);

BUFx5_ASAP7_75t_L g322 ( 
.A(n_139),
.Y(n_322)
);

INVx1_ASAP7_75t_SL g323 ( 
.A(n_168),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_89),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_240),
.B(n_0),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_307),
.B(n_0),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_202),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_217),
.A2(n_257),
.B1(n_279),
.B2(n_242),
.Y(n_328)
);

AND2x4_ASAP7_75t_L g329 ( 
.A(n_202),
.B(n_1),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_200),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_274),
.Y(n_331)
);

OA21x2_ASAP7_75t_L g332 ( 
.A1(n_191),
.A2(n_90),
.B(n_186),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_284),
.B(n_1),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_274),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_298),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_200),
.Y(n_336)
);

CKINVDCx8_ASAP7_75t_R g337 ( 
.A(n_195),
.Y(n_337)
);

AND2x2_ASAP7_75t_SL g338 ( 
.A(n_194),
.B(n_44),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_219),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_219),
.Y(n_340)
);

BUFx2_ASAP7_75t_L g341 ( 
.A(n_204),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_274),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_247),
.Y(n_343)
);

INVx6_ASAP7_75t_L g344 ( 
.A(n_200),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_245),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_287),
.B(n_2),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_274),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_245),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_310),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_200),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_247),
.B(n_2),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_190),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_206),
.Y(n_353)
);

BUFx2_ASAP7_75t_L g354 ( 
.A(n_250),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_310),
.B(n_3),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_200),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_191),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_222),
.B(n_3),
.Y(n_358)
);

INVx2_ASAP7_75t_SL g359 ( 
.A(n_293),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_235),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_223),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_258),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_259),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_262),
.B(n_9),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_200),
.Y(n_365)
);

OA21x2_ASAP7_75t_L g366 ( 
.A1(n_293),
.A2(n_99),
.B(n_185),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_231),
.A2(n_10),
.B1(n_14),
.B2(n_16),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_270),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_223),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_273),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_213),
.Y(n_371)
);

BUFx2_ASAP7_75t_L g372 ( 
.A(n_264),
.Y(n_372)
);

AND2x4_ASAP7_75t_L g373 ( 
.A(n_296),
.B(n_14),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_277),
.Y(n_374)
);

INVx5_ASAP7_75t_L g375 ( 
.A(n_246),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_278),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_295),
.Y(n_377)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_300),
.Y(n_378)
);

AND2x4_ASAP7_75t_L g379 ( 
.A(n_296),
.B(n_17),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_210),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_318),
.B(n_197),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_210),
.Y(n_382)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_324),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_198),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_199),
.Y(n_385)
);

OA21x2_ASAP7_75t_L g386 ( 
.A1(n_201),
.A2(n_101),
.B(n_181),
.Y(n_386)
);

INVx3_ASAP7_75t_L g387 ( 
.A(n_208),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_210),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_210),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_213),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_209),
.Y(n_391)
);

CKINVDCx16_ASAP7_75t_R g392 ( 
.A(n_236),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_313),
.B(n_18),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_210),
.Y(n_394)
);

HB1xp67_ASAP7_75t_L g395 ( 
.A(n_280),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_322),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_215),
.Y(n_397)
);

CKINVDCx6p67_ASAP7_75t_R g398 ( 
.A(n_322),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_322),
.Y(n_399)
);

BUFx12f_ASAP7_75t_L g400 ( 
.A(n_192),
.Y(n_400)
);

NOR2x1_ASAP7_75t_L g401 ( 
.A(n_216),
.B(n_220),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_224),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_225),
.B(n_19),
.Y(n_403)
);

INVx1_ASAP7_75t_SL g404 ( 
.A(n_341),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_329),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_371),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_384),
.B(n_227),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_357),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_357),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_373),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_373),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_402),
.B(n_228),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_373),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_327),
.B(n_232),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_331),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_357),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_357),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_379),
.B(n_375),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_341),
.B(n_283),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_357),
.Y(n_420)
);

INVx3_ASAP7_75t_L g421 ( 
.A(n_379),
.Y(n_421)
);

NAND3xp33_ASAP7_75t_L g422 ( 
.A(n_352),
.B(n_299),
.C(n_297),
.Y(n_422)
);

BUFx6f_ASAP7_75t_SL g423 ( 
.A(n_338),
.Y(n_423)
);

NAND3xp33_ASAP7_75t_L g424 ( 
.A(n_353),
.B(n_312),
.C(n_304),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_355),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_355),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_378),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_378),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_371),
.Y(n_429)
);

BUFx6f_ASAP7_75t_SL g430 ( 
.A(n_338),
.Y(n_430)
);

BUFx3_ASAP7_75t_L g431 ( 
.A(n_349),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_330),
.Y(n_432)
);

INVx5_ASAP7_75t_L g433 ( 
.A(n_344),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_378),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_383),
.B(n_234),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_326),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_354),
.B(n_291),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_354),
.B(n_196),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_372),
.B(n_203),
.Y(n_439)
);

NAND3xp33_ASAP7_75t_L g440 ( 
.A(n_325),
.B(n_243),
.C(n_241),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_364),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_364),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_L g443 ( 
.A1(n_335),
.A2(n_311),
.B1(n_244),
.B2(n_288),
.Y(n_443)
);

INVx1_ASAP7_75t_SL g444 ( 
.A(n_372),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_390),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_330),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_383),
.B(n_205),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_336),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_383),
.B(n_387),
.Y(n_449)
);

AND2x4_ASAP7_75t_L g450 ( 
.A(n_401),
.B(n_290),
.Y(n_450)
);

BUFx6f_ASAP7_75t_SL g451 ( 
.A(n_360),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_387),
.B(n_248),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_387),
.B(n_207),
.Y(n_453)
);

NAND2xp33_ASAP7_75t_L g454 ( 
.A(n_343),
.B(n_322),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_398),
.B(n_251),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_SL g456 ( 
.A(n_351),
.B(n_244),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_375),
.B(n_322),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_390),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_328),
.A2(n_311),
.B1(n_288),
.B2(n_236),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_375),
.B(n_322),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_359),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_398),
.B(n_212),
.Y(n_462)
);

INVx3_ASAP7_75t_L g463 ( 
.A(n_385),
.Y(n_463)
);

NAND3xp33_ASAP7_75t_L g464 ( 
.A(n_393),
.B(n_255),
.C(n_253),
.Y(n_464)
);

AND2x4_ASAP7_75t_L g465 ( 
.A(n_359),
.B(n_256),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_385),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_350),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_350),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_356),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_356),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_395),
.B(n_214),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_365),
.Y(n_472)
);

INVx4_ASAP7_75t_L g473 ( 
.A(n_344),
.Y(n_473)
);

AND2x6_ASAP7_75t_L g474 ( 
.A(n_351),
.B(n_393),
.Y(n_474)
);

AOI22xp33_ASAP7_75t_L g475 ( 
.A1(n_363),
.A2(n_272),
.B1(n_321),
.B2(n_320),
.Y(n_475)
);

AOI22xp33_ASAP7_75t_L g476 ( 
.A1(n_368),
.A2(n_308),
.B1(n_319),
.B2(n_285),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_385),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_335),
.B(n_218),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_375),
.B(n_221),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_365),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_385),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_380),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_380),
.Y(n_483)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_391),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_391),
.Y(n_485)
);

INVxp33_ASAP7_75t_L g486 ( 
.A(n_381),
.Y(n_486)
);

INVxp33_ASAP7_75t_L g487 ( 
.A(n_333),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_382),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_391),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_382),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_400),
.A2(n_263),
.B1(n_301),
.B2(n_249),
.Y(n_491)
);

AND2x6_ASAP7_75t_L g492 ( 
.A(n_388),
.B(n_260),
.Y(n_492)
);

OR2x6_ASAP7_75t_L g493 ( 
.A(n_400),
.B(n_265),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_331),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_391),
.Y(n_495)
);

INVx2_ASAP7_75t_SL g496 ( 
.A(n_344),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_391),
.B(n_267),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_388),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_389),
.Y(n_499)
);

AOI22xp33_ASAP7_75t_L g500 ( 
.A1(n_370),
.A2(n_314),
.B1(n_306),
.B2(n_309),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_397),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_389),
.Y(n_502)
);

INVx4_ASAP7_75t_L g503 ( 
.A(n_344),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_397),
.B(n_286),
.Y(n_504)
);

INVx4_ASAP7_75t_L g505 ( 
.A(n_349),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_394),
.Y(n_506)
);

INVxp67_ASAP7_75t_SL g507 ( 
.A(n_374),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_394),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_376),
.B(n_226),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_396),
.Y(n_510)
);

INVx3_ASAP7_75t_L g511 ( 
.A(n_397),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_396),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_399),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_486),
.B(n_377),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_486),
.B(n_337),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_436),
.B(n_403),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_427),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_487),
.B(n_337),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_507),
.B(n_346),
.Y(n_519)
);

AND2x4_ASAP7_75t_SL g520 ( 
.A(n_493),
.B(n_369),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_428),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_423),
.A2(n_367),
.B1(n_358),
.B2(n_362),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_487),
.B(n_229),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_438),
.B(n_339),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_431),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_455),
.B(n_230),
.Y(n_526)
);

INVx2_ASAP7_75t_SL g527 ( 
.A(n_404),
.Y(n_527)
);

INVx2_ASAP7_75t_SL g528 ( 
.A(n_444),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_465),
.B(n_340),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_434),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_455),
.B(n_233),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_439),
.B(n_345),
.Y(n_532)
);

AOI22xp33_ASAP7_75t_SL g533 ( 
.A1(n_423),
.A2(n_361),
.B1(n_348),
.B2(n_369),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_465),
.B(n_509),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_461),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_465),
.B(n_238),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_474),
.B(n_239),
.Y(n_537)
);

AOI22xp33_ASAP7_75t_L g538 ( 
.A1(n_421),
.A2(n_397),
.B1(n_349),
.B2(n_366),
.Y(n_538)
);

AOI22xp5_ASAP7_75t_L g539 ( 
.A1(n_430),
.A2(n_193),
.B1(n_282),
.B2(n_237),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_464),
.B(n_302),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_441),
.B(n_442),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_474),
.B(n_252),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_405),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_410),
.Y(n_544)
);

AOI21xp5_ASAP7_75t_L g545 ( 
.A1(n_418),
.A2(n_366),
.B(n_332),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_505),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_474),
.B(n_261),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_411),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_437),
.B(n_332),
.Y(n_549)
);

AND2x2_ASAP7_75t_L g550 ( 
.A(n_478),
.B(n_332),
.Y(n_550)
);

OAI22xp5_ASAP7_75t_SL g551 ( 
.A1(n_459),
.A2(n_386),
.B1(n_366),
.B2(n_323),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_425),
.B(n_211),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_471),
.B(n_266),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_426),
.B(n_268),
.Y(n_554)
);

AND2x6_ASAP7_75t_SL g555 ( 
.A(n_493),
.B(n_254),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_413),
.Y(n_556)
);

INVxp67_ASAP7_75t_L g557 ( 
.A(n_456),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_505),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_462),
.B(n_269),
.Y(n_559)
);

INVx2_ASAP7_75t_SL g560 ( 
.A(n_419),
.Y(n_560)
);

INVx5_ASAP7_75t_L g561 ( 
.A(n_463),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_449),
.B(n_271),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_440),
.B(n_275),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_422),
.B(n_276),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_492),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_492),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_R g567 ( 
.A(n_406),
.B(n_429),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_424),
.B(n_281),
.Y(n_568)
);

OR2x2_ASAP7_75t_L g569 ( 
.A(n_443),
.B(n_19),
.Y(n_569)
);

NAND2xp33_ASAP7_75t_L g570 ( 
.A(n_492),
.B(n_289),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_447),
.B(n_294),
.Y(n_571)
);

BUFx8_ASAP7_75t_L g572 ( 
.A(n_451),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_449),
.B(n_453),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_435),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_452),
.Y(n_575)
);

A2O1A1Ixp33_ASAP7_75t_L g576 ( 
.A1(n_452),
.A2(n_254),
.B(n_292),
.C(n_349),
.Y(n_576)
);

INVx3_ASAP7_75t_L g577 ( 
.A(n_492),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_450),
.B(n_303),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_473),
.B(n_305),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_414),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_407),
.B(n_315),
.Y(n_581)
);

NOR2xp67_ASAP7_75t_L g582 ( 
.A(n_491),
.B(n_20),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_407),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_412),
.B(n_316),
.Y(n_584)
);

AOI22xp33_ASAP7_75t_L g585 ( 
.A1(n_430),
.A2(n_386),
.B1(n_292),
.B2(n_342),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_412),
.B(n_317),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_475),
.B(n_331),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_454),
.B(n_51),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_475),
.B(n_331),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_476),
.B(n_331),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_484),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_476),
.B(n_334),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_473),
.B(n_334),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_500),
.B(n_334),
.Y(n_594)
);

AO221x1_ASAP7_75t_L g595 ( 
.A1(n_445),
.A2(n_347),
.B1(n_342),
.B2(n_334),
.C(n_25),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_503),
.B(n_334),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_457),
.Y(n_597)
);

NAND3xp33_ASAP7_75t_L g598 ( 
.A(n_500),
.B(n_347),
.C(n_342),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_493),
.B(n_21),
.Y(n_599)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_492),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_503),
.B(n_342),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_479),
.B(n_342),
.Y(n_602)
);

AOI22xp33_ASAP7_75t_L g603 ( 
.A1(n_432),
.A2(n_347),
.B1(n_24),
.B2(n_26),
.Y(n_603)
);

AOI22xp33_ASAP7_75t_L g604 ( 
.A1(n_432),
.A2(n_347),
.B1(n_24),
.B2(n_28),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_458),
.B(n_23),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_516),
.B(n_513),
.Y(n_606)
);

NAND3xp33_ASAP7_75t_L g607 ( 
.A(n_515),
.B(n_528),
.C(n_533),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_514),
.B(n_513),
.Y(n_608)
);

AOI21xp5_ASAP7_75t_L g609 ( 
.A1(n_545),
.A2(n_460),
.B(n_496),
.Y(n_609)
);

AOI21xp5_ASAP7_75t_L g610 ( 
.A1(n_545),
.A2(n_497),
.B(n_504),
.Y(n_610)
);

A2O1A1Ixp33_ASAP7_75t_L g611 ( 
.A1(n_574),
.A2(n_512),
.B(n_446),
.C(n_510),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_519),
.B(n_560),
.Y(n_612)
);

OAI22xp5_ASAP7_75t_L g613 ( 
.A1(n_583),
.A2(n_490),
.B1(n_510),
.B2(n_508),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_524),
.B(n_448),
.Y(n_614)
);

INVx2_ASAP7_75t_SL g615 ( 
.A(n_572),
.Y(n_615)
);

OAI22xp5_ASAP7_75t_L g616 ( 
.A1(n_580),
.A2(n_490),
.B1(n_508),
.B2(n_506),
.Y(n_616)
);

NOR3xp33_ASAP7_75t_L g617 ( 
.A(n_533),
.B(n_518),
.C(n_557),
.Y(n_617)
);

AOI21xp5_ASAP7_75t_L g618 ( 
.A1(n_573),
.A2(n_497),
.B(n_504),
.Y(n_618)
);

CKINVDCx10_ASAP7_75t_R g619 ( 
.A(n_520),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_524),
.B(n_448),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_532),
.B(n_467),
.Y(n_621)
);

AOI21xp5_ASAP7_75t_L g622 ( 
.A1(n_550),
.A2(n_534),
.B(n_549),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_575),
.B(n_467),
.Y(n_623)
);

AND2x4_ASAP7_75t_L g624 ( 
.A(n_541),
.B(n_433),
.Y(n_624)
);

A2O1A1Ixp33_ASAP7_75t_L g625 ( 
.A1(n_543),
.A2(n_480),
.B(n_506),
.C(n_502),
.Y(n_625)
);

AOI21xp5_ASAP7_75t_L g626 ( 
.A1(n_538),
.A2(n_480),
.B(n_502),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_546),
.Y(n_627)
);

BUFx8_ASAP7_75t_L g628 ( 
.A(n_599),
.Y(n_628)
);

AOI22xp5_ASAP7_75t_L g629 ( 
.A1(n_522),
.A2(n_470),
.B1(n_468),
.B2(n_499),
.Y(n_629)
);

AOI21xp5_ASAP7_75t_L g630 ( 
.A1(n_538),
.A2(n_472),
.B(n_468),
.Y(n_630)
);

O2A1O1Ixp33_ASAP7_75t_L g631 ( 
.A1(n_569),
.A2(n_483),
.B(n_470),
.C(n_498),
.Y(n_631)
);

NAND2x1_ASAP7_75t_L g632 ( 
.A(n_577),
.B(n_469),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_565),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_540),
.B(n_472),
.Y(n_634)
);

O2A1O1Ixp33_ASAP7_75t_L g635 ( 
.A1(n_557),
.A2(n_482),
.B(n_483),
.C(n_498),
.Y(n_635)
);

AOI21xp5_ASAP7_75t_L g636 ( 
.A1(n_602),
.A2(n_488),
.B(n_433),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_567),
.B(n_488),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_535),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_540),
.B(n_511),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_578),
.B(n_29),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_605),
.B(n_30),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_552),
.B(n_582),
.Y(n_642)
);

OAI21xp33_ASAP7_75t_L g643 ( 
.A1(n_552),
.A2(n_477),
.B(n_501),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_SL g644 ( 
.A(n_551),
.B(n_466),
.Y(n_644)
);

OAI21xp5_ASAP7_75t_L g645 ( 
.A1(n_587),
.A2(n_481),
.B(n_495),
.Y(n_645)
);

AOI21xp33_ASAP7_75t_L g646 ( 
.A1(n_537),
.A2(n_489),
.B(n_485),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_544),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_548),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_523),
.B(n_30),
.Y(n_649)
);

AOI21xp5_ASAP7_75t_L g650 ( 
.A1(n_562),
.A2(n_420),
.B(n_417),
.Y(n_650)
);

AOI21xp5_ASAP7_75t_L g651 ( 
.A1(n_597),
.A2(n_417),
.B(n_416),
.Y(n_651)
);

OAI22xp5_ASAP7_75t_L g652 ( 
.A1(n_556),
.A2(n_408),
.B1(n_409),
.B2(n_33),
.Y(n_652)
);

OAI21xp5_ASAP7_75t_L g653 ( 
.A1(n_589),
.A2(n_494),
.B(n_415),
.Y(n_653)
);

AOI22xp5_ASAP7_75t_L g654 ( 
.A1(n_539),
.A2(n_494),
.B1(n_415),
.B2(n_33),
.Y(n_654)
);

NOR2xp67_ASAP7_75t_L g655 ( 
.A(n_577),
.B(n_56),
.Y(n_655)
);

AND2x4_ASAP7_75t_L g656 ( 
.A(n_553),
.B(n_31),
.Y(n_656)
);

OAI21xp33_ASAP7_75t_SL g657 ( 
.A1(n_517),
.A2(n_32),
.B(n_34),
.Y(n_657)
);

OAI21xp5_ASAP7_75t_L g658 ( 
.A1(n_590),
.A2(n_594),
.B(n_592),
.Y(n_658)
);

INVxp33_ASAP7_75t_SL g659 ( 
.A(n_571),
.Y(n_659)
);

CKINVDCx12_ASAP7_75t_R g660 ( 
.A(n_555),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_521),
.Y(n_661)
);

AOI21xp5_ASAP7_75t_L g662 ( 
.A1(n_536),
.A2(n_117),
.B(n_179),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_584),
.B(n_32),
.Y(n_663)
);

AOI21xp5_ASAP7_75t_L g664 ( 
.A1(n_530),
.A2(n_121),
.B(n_178),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_529),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_554),
.B(n_34),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_554),
.B(n_36),
.Y(n_667)
);

AOI22xp5_ASAP7_75t_L g668 ( 
.A1(n_563),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_668)
);

BUFx6f_ASAP7_75t_L g669 ( 
.A(n_566),
.Y(n_669)
);

BUFx6f_ASAP7_75t_L g670 ( 
.A(n_566),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_571),
.B(n_38),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_581),
.B(n_39),
.Y(n_672)
);

OAI21xp5_ASAP7_75t_L g673 ( 
.A1(n_585),
.A2(n_113),
.B(n_166),
.Y(n_673)
);

AOI21xp5_ASAP7_75t_L g674 ( 
.A1(n_601),
.A2(n_110),
.B(n_165),
.Y(n_674)
);

OAI22xp5_ASAP7_75t_L g675 ( 
.A1(n_542),
.A2(n_40),
.B1(n_42),
.B2(n_57),
.Y(n_675)
);

AND2x2_ASAP7_75t_SL g676 ( 
.A(n_566),
.B(n_58),
.Y(n_676)
);

OA22x2_ASAP7_75t_L g677 ( 
.A1(n_595),
.A2(n_568),
.B1(n_531),
.B2(n_526),
.Y(n_677)
);

BUFx8_ASAP7_75t_L g678 ( 
.A(n_558),
.Y(n_678)
);

BUFx3_ASAP7_75t_L g679 ( 
.A(n_525),
.Y(n_679)
);

A2O1A1Ixp33_ASAP7_75t_L g680 ( 
.A1(n_576),
.A2(n_61),
.B(n_63),
.C(n_65),
.Y(n_680)
);

INVx3_ASAP7_75t_L g681 ( 
.A(n_600),
.Y(n_681)
);

OAI21xp33_ASAP7_75t_L g682 ( 
.A1(n_586),
.A2(n_69),
.B(n_75),
.Y(n_682)
);

OAI21xp33_ASAP7_75t_L g683 ( 
.A1(n_563),
.A2(n_76),
.B(n_77),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_547),
.B(n_600),
.Y(n_684)
);

OAI22xp5_ASAP7_75t_L g685 ( 
.A1(n_585),
.A2(n_78),
.B1(n_80),
.B2(n_81),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_564),
.B(n_82),
.Y(n_686)
);

NAND2x1p5_ASAP7_75t_L g687 ( 
.A(n_559),
.B(n_84),
.Y(n_687)
);

AOI21xp5_ASAP7_75t_L g688 ( 
.A1(n_579),
.A2(n_596),
.B(n_593),
.Y(n_688)
);

AOI21xp33_ASAP7_75t_L g689 ( 
.A1(n_570),
.A2(n_92),
.B(n_95),
.Y(n_689)
);

O2A1O1Ixp33_ASAP7_75t_L g690 ( 
.A1(n_603),
.A2(n_100),
.B(n_102),
.C(n_130),
.Y(n_690)
);

O2A1O1Ixp33_ASAP7_75t_L g691 ( 
.A1(n_603),
.A2(n_189),
.B(n_134),
.C(n_135),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_598),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_525),
.B(n_155),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_604),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_588),
.B(n_164),
.Y(n_695)
);

OA21x2_ASAP7_75t_L g696 ( 
.A1(n_653),
.A2(n_604),
.B(n_591),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_638),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_661),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_665),
.B(n_606),
.Y(n_699)
);

A2O1A1Ixp33_ASAP7_75t_L g700 ( 
.A1(n_631),
.A2(n_561),
.B(n_156),
.C(n_160),
.Y(n_700)
);

AND2x4_ASAP7_75t_L g701 ( 
.A(n_647),
.B(n_561),
.Y(n_701)
);

INVx2_ASAP7_75t_SL g702 ( 
.A(n_619),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_648),
.Y(n_703)
);

AOI21xp5_ASAP7_75t_L g704 ( 
.A1(n_610),
.A2(n_626),
.B(n_630),
.Y(n_704)
);

AOI21xp5_ASAP7_75t_L g705 ( 
.A1(n_618),
.A2(n_658),
.B(n_650),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_642),
.B(n_637),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_617),
.B(n_608),
.Y(n_707)
);

AOI21xp5_ASAP7_75t_L g708 ( 
.A1(n_623),
.A2(n_695),
.B(n_620),
.Y(n_708)
);

OAI22x1_ASAP7_75t_L g709 ( 
.A1(n_607),
.A2(n_656),
.B1(n_668),
.B2(n_615),
.Y(n_709)
);

OAI22xp5_ASAP7_75t_L g710 ( 
.A1(n_614),
.A2(n_621),
.B1(n_629),
.B2(n_616),
.Y(n_710)
);

AOI21xp5_ASAP7_75t_L g711 ( 
.A1(n_645),
.A2(n_611),
.B(n_651),
.Y(n_711)
);

A2O1A1Ixp33_ASAP7_75t_L g712 ( 
.A1(n_671),
.A2(n_667),
.B(n_666),
.C(n_657),
.Y(n_712)
);

BUFx3_ASAP7_75t_L g713 ( 
.A(n_678),
.Y(n_713)
);

AOI21xp5_ASAP7_75t_L g714 ( 
.A1(n_684),
.A2(n_646),
.B(n_634),
.Y(n_714)
);

OAI22xp5_ASAP7_75t_L g715 ( 
.A1(n_613),
.A2(n_694),
.B1(n_641),
.B2(n_663),
.Y(n_715)
);

NOR4xp25_ASAP7_75t_L g716 ( 
.A(n_680),
.B(n_683),
.C(n_675),
.D(n_672),
.Y(n_716)
);

AOI21xp5_ASAP7_75t_SL g717 ( 
.A1(n_673),
.A2(n_685),
.B(n_633),
.Y(n_717)
);

A2O1A1Ixp33_ASAP7_75t_L g718 ( 
.A1(n_635),
.A2(n_649),
.B(n_640),
.C(n_643),
.Y(n_718)
);

AO21x1_ASAP7_75t_L g719 ( 
.A1(n_686),
.A2(n_691),
.B(n_690),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_656),
.B(n_678),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_654),
.B(n_624),
.Y(n_721)
);

AO21x1_ASAP7_75t_L g722 ( 
.A1(n_662),
.A2(n_664),
.B(n_692),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_624),
.B(n_627),
.Y(n_723)
);

OAI21xp5_ASAP7_75t_SL g724 ( 
.A1(n_652),
.A2(n_687),
.B(n_689),
.Y(n_724)
);

OAI21xp5_ASAP7_75t_L g725 ( 
.A1(n_625),
.A2(n_639),
.B(n_636),
.Y(n_725)
);

CKINVDCx20_ASAP7_75t_R g726 ( 
.A(n_628),
.Y(n_726)
);

A2O1A1Ixp33_ASAP7_75t_L g727 ( 
.A1(n_688),
.A2(n_682),
.B(n_693),
.C(n_655),
.Y(n_727)
);

OAI22xp5_ASAP7_75t_L g728 ( 
.A1(n_677),
.A2(n_670),
.B1(n_669),
.B2(n_679),
.Y(n_728)
);

BUFx2_ASAP7_75t_R g729 ( 
.A(n_660),
.Y(n_729)
);

A2O1A1Ixp33_ASAP7_75t_L g730 ( 
.A1(n_655),
.A2(n_674),
.B(n_681),
.C(n_632),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_628),
.B(n_681),
.Y(n_731)
);

OAI22x1_ASAP7_75t_L g732 ( 
.A1(n_607),
.A2(n_459),
.B1(n_390),
.B2(n_371),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_612),
.B(n_486),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_612),
.B(n_486),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_612),
.Y(n_735)
);

OAI21xp5_ASAP7_75t_L g736 ( 
.A1(n_622),
.A2(n_630),
.B(n_626),
.Y(n_736)
);

OAI21xp5_ASAP7_75t_L g737 ( 
.A1(n_622),
.A2(n_630),
.B(n_626),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_612),
.B(n_486),
.Y(n_738)
);

OR2x2_ASAP7_75t_L g739 ( 
.A(n_612),
.B(n_527),
.Y(n_739)
);

BUFx2_ASAP7_75t_L g740 ( 
.A(n_678),
.Y(n_740)
);

NOR2xp67_ASAP7_75t_SL g741 ( 
.A(n_615),
.B(n_527),
.Y(n_741)
);

INVxp67_ASAP7_75t_SL g742 ( 
.A(n_678),
.Y(n_742)
);

NOR2xp67_ASAP7_75t_L g743 ( 
.A(n_612),
.B(n_606),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_612),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_612),
.B(n_486),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_612),
.B(n_486),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_659),
.B(n_527),
.Y(n_747)
);

A2O1A1Ixp33_ASAP7_75t_L g748 ( 
.A1(n_631),
.A2(n_574),
.B(n_575),
.C(n_622),
.Y(n_748)
);

AOI22xp5_ASAP7_75t_L g749 ( 
.A1(n_617),
.A2(n_430),
.B1(n_423),
.B2(n_474),
.Y(n_749)
);

A2O1A1Ixp33_ASAP7_75t_L g750 ( 
.A1(n_631),
.A2(n_574),
.B(n_575),
.C(n_622),
.Y(n_750)
);

OAI21xp5_ASAP7_75t_L g751 ( 
.A1(n_622),
.A2(n_630),
.B(n_626),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_612),
.B(n_486),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_612),
.B(n_486),
.Y(n_753)
);

NAND3x1_ASAP7_75t_L g754 ( 
.A(n_617),
.B(n_459),
.C(n_367),
.Y(n_754)
);

CKINVDCx20_ASAP7_75t_R g755 ( 
.A(n_678),
.Y(n_755)
);

AOI21xp5_ASAP7_75t_L g756 ( 
.A1(n_610),
.A2(n_545),
.B(n_609),
.Y(n_756)
);

AOI21xp5_ASAP7_75t_SL g757 ( 
.A1(n_673),
.A2(n_685),
.B(n_622),
.Y(n_757)
);

AO21x1_ASAP7_75t_L g758 ( 
.A1(n_644),
.A2(n_673),
.B(n_685),
.Y(n_758)
);

AO31x2_ASAP7_75t_L g759 ( 
.A1(n_680),
.A2(n_545),
.A3(n_622),
.B(n_685),
.Y(n_759)
);

BUFx6f_ASAP7_75t_L g760 ( 
.A(n_633),
.Y(n_760)
);

BUFx6f_ASAP7_75t_L g761 ( 
.A(n_633),
.Y(n_761)
);

INVx3_ASAP7_75t_L g762 ( 
.A(n_678),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_619),
.Y(n_763)
);

OAI22xp5_ASAP7_75t_L g764 ( 
.A1(n_614),
.A2(n_620),
.B1(n_621),
.B2(n_606),
.Y(n_764)
);

OAI22xp5_ASAP7_75t_L g765 ( 
.A1(n_614),
.A2(n_620),
.B1(n_621),
.B2(n_606),
.Y(n_765)
);

AOI21xp5_ASAP7_75t_L g766 ( 
.A1(n_610),
.A2(n_545),
.B(n_609),
.Y(n_766)
);

OAI21xp5_ASAP7_75t_L g767 ( 
.A1(n_622),
.A2(n_545),
.B(n_658),
.Y(n_767)
);

OAI22x1_ASAP7_75t_L g768 ( 
.A1(n_607),
.A2(n_459),
.B1(n_390),
.B2(n_371),
.Y(n_768)
);

AO31x2_ASAP7_75t_L g769 ( 
.A1(n_680),
.A2(n_545),
.A3(n_622),
.B(n_685),
.Y(n_769)
);

AOI21xp5_ASAP7_75t_L g770 ( 
.A1(n_610),
.A2(n_545),
.B(n_609),
.Y(n_770)
);

OAI21xp5_ASAP7_75t_L g771 ( 
.A1(n_622),
.A2(n_545),
.B(n_658),
.Y(n_771)
);

BUFx4f_ASAP7_75t_L g772 ( 
.A(n_615),
.Y(n_772)
);

A2O1A1Ixp33_ASAP7_75t_L g773 ( 
.A1(n_631),
.A2(n_574),
.B(n_575),
.C(n_622),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_612),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_612),
.Y(n_775)
);

NOR4xp25_ASAP7_75t_L g776 ( 
.A(n_657),
.B(n_631),
.C(n_576),
.D(n_569),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_612),
.B(n_486),
.Y(n_777)
);

NOR2x1_ASAP7_75t_L g778 ( 
.A(n_612),
.B(n_607),
.Y(n_778)
);

CKINVDCx11_ASAP7_75t_R g779 ( 
.A(n_619),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_638),
.Y(n_780)
);

AND2x2_ASAP7_75t_SL g781 ( 
.A(n_676),
.B(n_520),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_612),
.Y(n_782)
);

BUFx2_ASAP7_75t_L g783 ( 
.A(n_678),
.Y(n_783)
);

OAI22xp5_ASAP7_75t_L g784 ( 
.A1(n_614),
.A2(n_620),
.B1(n_621),
.B2(n_606),
.Y(n_784)
);

INVx1_ASAP7_75t_SL g785 ( 
.A(n_612),
.Y(n_785)
);

INVx3_ASAP7_75t_SL g786 ( 
.A(n_615),
.Y(n_786)
);

OAI21xp5_ASAP7_75t_L g787 ( 
.A1(n_748),
.A2(n_773),
.B(n_750),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_733),
.Y(n_788)
);

OAI21x1_ASAP7_75t_SL g789 ( 
.A1(n_764),
.A2(n_784),
.B(n_765),
.Y(n_789)
);

INVx6_ASAP7_75t_L g790 ( 
.A(n_713),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_738),
.B(n_753),
.Y(n_791)
);

BUFx2_ASAP7_75t_L g792 ( 
.A(n_755),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_735),
.Y(n_793)
);

AOI21xp5_ASAP7_75t_L g794 ( 
.A1(n_757),
.A2(n_708),
.B(n_704),
.Y(n_794)
);

INVx2_ASAP7_75t_SL g795 ( 
.A(n_740),
.Y(n_795)
);

AOI21xp5_ASAP7_75t_L g796 ( 
.A1(n_766),
.A2(n_770),
.B(n_751),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_744),
.Y(n_797)
);

OAI21xp5_ASAP7_75t_L g798 ( 
.A1(n_767),
.A2(n_771),
.B(n_712),
.Y(n_798)
);

INVx8_ASAP7_75t_L g799 ( 
.A(n_763),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_699),
.B(n_743),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_720),
.B(n_747),
.Y(n_801)
);

BUFx2_ASAP7_75t_R g802 ( 
.A(n_783),
.Y(n_802)
);

OAI21x1_ASAP7_75t_SL g803 ( 
.A1(n_728),
.A2(n_749),
.B(n_707),
.Y(n_803)
);

OA21x2_ASAP7_75t_L g804 ( 
.A1(n_705),
.A2(n_727),
.B(n_725),
.Y(n_804)
);

AOI21xp5_ASAP7_75t_L g805 ( 
.A1(n_717),
.A2(n_711),
.B(n_715),
.Y(n_805)
);

AND2x2_ASAP7_75t_L g806 ( 
.A(n_785),
.B(n_734),
.Y(n_806)
);

BUFx10_ASAP7_75t_L g807 ( 
.A(n_702),
.Y(n_807)
);

OAI21x1_ASAP7_75t_SL g808 ( 
.A1(n_749),
.A2(n_758),
.B(n_778),
.Y(n_808)
);

NAND3xp33_ASAP7_75t_L g809 ( 
.A(n_776),
.B(n_718),
.C(n_724),
.Y(n_809)
);

OAI21xp5_ASAP7_75t_L g810 ( 
.A1(n_776),
.A2(n_710),
.B(n_714),
.Y(n_810)
);

HB1xp67_ASAP7_75t_L g811 ( 
.A(n_774),
.Y(n_811)
);

AO31x2_ASAP7_75t_L g812 ( 
.A1(n_719),
.A2(n_700),
.A3(n_730),
.B(n_709),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_775),
.B(n_782),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_716),
.A2(n_724),
.B(n_696),
.Y(n_814)
);

AND2x2_ASAP7_75t_L g815 ( 
.A(n_745),
.B(n_746),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_752),
.Y(n_816)
);

OAI21xp5_ASAP7_75t_SL g817 ( 
.A1(n_739),
.A2(n_762),
.B(n_777),
.Y(n_817)
);

BUFx2_ASAP7_75t_L g818 ( 
.A(n_742),
.Y(n_818)
);

A2O1A1Ixp33_ASAP7_75t_L g819 ( 
.A1(n_706),
.A2(n_697),
.B(n_698),
.C(n_703),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_716),
.A2(n_721),
.B(n_723),
.Y(n_820)
);

OA21x2_ASAP7_75t_L g821 ( 
.A1(n_759),
.A2(n_769),
.B(n_780),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_731),
.Y(n_822)
);

OA21x2_ASAP7_75t_L g823 ( 
.A1(n_701),
.A2(n_760),
.B(n_761),
.Y(n_823)
);

AOI21x1_ASAP7_75t_L g824 ( 
.A1(n_741),
.A2(n_768),
.B(n_732),
.Y(n_824)
);

OAI21xp5_ASAP7_75t_L g825 ( 
.A1(n_754),
.A2(n_781),
.B(n_772),
.Y(n_825)
);

OAI21xp5_ASAP7_75t_L g826 ( 
.A1(n_772),
.A2(n_726),
.B(n_786),
.Y(n_826)
);

OA21x2_ASAP7_75t_L g827 ( 
.A1(n_729),
.A2(n_737),
.B(n_736),
.Y(n_827)
);

AND2x4_ASAP7_75t_L g828 ( 
.A(n_779),
.B(n_743),
.Y(n_828)
);

INVx4_ASAP7_75t_L g829 ( 
.A(n_713),
.Y(n_829)
);

AO31x2_ASAP7_75t_L g830 ( 
.A1(n_758),
.A2(n_704),
.A3(n_722),
.B(n_756),
.Y(n_830)
);

AOI21xp5_ASAP7_75t_L g831 ( 
.A1(n_764),
.A2(n_784),
.B(n_765),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_733),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_699),
.B(n_743),
.Y(n_833)
);

AO31x2_ASAP7_75t_L g834 ( 
.A1(n_758),
.A2(n_704),
.A3(n_722),
.B(n_756),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_733),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_781),
.B(n_527),
.Y(n_836)
);

BUFx10_ASAP7_75t_L g837 ( 
.A(n_763),
.Y(n_837)
);

OAI21xp5_ASAP7_75t_L g838 ( 
.A1(n_748),
.A2(n_622),
.B(n_750),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_779),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_733),
.Y(n_840)
);

AO31x2_ASAP7_75t_L g841 ( 
.A1(n_758),
.A2(n_704),
.A3(n_722),
.B(n_756),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_781),
.B(n_527),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_764),
.A2(n_784),
.B(n_765),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_L g844 ( 
.A(n_720),
.B(n_392),
.Y(n_844)
);

BUFx3_ASAP7_75t_L g845 ( 
.A(n_755),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_811),
.B(n_806),
.Y(n_846)
);

AOI22xp33_ASAP7_75t_L g847 ( 
.A1(n_789),
.A2(n_843),
.B1(n_831),
.B2(n_825),
.Y(n_847)
);

AO21x2_ASAP7_75t_L g848 ( 
.A1(n_814),
.A2(n_794),
.B(n_805),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_811),
.B(n_800),
.Y(n_849)
);

AO21x2_ASAP7_75t_L g850 ( 
.A1(n_796),
.A2(n_810),
.B(n_787),
.Y(n_850)
);

BUFx3_ASAP7_75t_L g851 ( 
.A(n_823),
.Y(n_851)
);

INVx2_ASAP7_75t_SL g852 ( 
.A(n_790),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_821),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_798),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_800),
.B(n_833),
.Y(n_855)
);

BUFx2_ASAP7_75t_R g856 ( 
.A(n_845),
.Y(n_856)
);

BUFx12f_ASAP7_75t_L g857 ( 
.A(n_837),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_793),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_815),
.B(n_813),
.Y(n_859)
);

OR2x2_ASAP7_75t_L g860 ( 
.A(n_817),
.B(n_813),
.Y(n_860)
);

OR2x2_ASAP7_75t_L g861 ( 
.A(n_817),
.B(n_809),
.Y(n_861)
);

INVx2_ASAP7_75t_SL g862 ( 
.A(n_790),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_797),
.Y(n_863)
);

HB1xp67_ASAP7_75t_L g864 ( 
.A(n_818),
.Y(n_864)
);

OR2x2_ASAP7_75t_L g865 ( 
.A(n_791),
.B(n_816),
.Y(n_865)
);

OA21x2_ASAP7_75t_L g866 ( 
.A1(n_810),
.A2(n_820),
.B(n_838),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_830),
.Y(n_867)
);

AND2x2_ASAP7_75t_L g868 ( 
.A(n_819),
.B(n_788),
.Y(n_868)
);

INVx8_ASAP7_75t_L g869 ( 
.A(n_828),
.Y(n_869)
);

BUFx2_ASAP7_75t_L g870 ( 
.A(n_851),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_853),
.Y(n_871)
);

AND2x2_ASAP7_75t_L g872 ( 
.A(n_854),
.B(n_827),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_859),
.B(n_840),
.Y(n_873)
);

HB1xp67_ASAP7_75t_L g874 ( 
.A(n_864),
.Y(n_874)
);

BUFx3_ASAP7_75t_L g875 ( 
.A(n_851),
.Y(n_875)
);

OR2x2_ASAP7_75t_L g876 ( 
.A(n_860),
.B(n_830),
.Y(n_876)
);

AOI221xp5_ASAP7_75t_L g877 ( 
.A1(n_847),
.A2(n_835),
.B1(n_832),
.B2(n_825),
.C(n_801),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_859),
.B(n_822),
.Y(n_878)
);

AOI22xp33_ASAP7_75t_L g879 ( 
.A1(n_860),
.A2(n_828),
.B1(n_808),
.B2(n_803),
.Y(n_879)
);

OR2x2_ASAP7_75t_L g880 ( 
.A(n_861),
.B(n_841),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_846),
.B(n_834),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_855),
.B(n_804),
.Y(n_882)
);

BUFx3_ASAP7_75t_L g883 ( 
.A(n_869),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_850),
.B(n_804),
.Y(n_884)
);

OR2x2_ASAP7_75t_L g885 ( 
.A(n_861),
.B(n_812),
.Y(n_885)
);

AOI22xp33_ASAP7_75t_L g886 ( 
.A1(n_868),
.A2(n_795),
.B1(n_844),
.B2(n_842),
.Y(n_886)
);

BUFx3_ASAP7_75t_L g887 ( 
.A(n_869),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_850),
.B(n_849),
.Y(n_888)
);

INVxp67_ASAP7_75t_L g889 ( 
.A(n_865),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_849),
.B(n_812),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_888),
.B(n_882),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_871),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_871),
.Y(n_893)
);

OR2x2_ASAP7_75t_L g894 ( 
.A(n_888),
.B(n_866),
.Y(n_894)
);

BUFx3_ASAP7_75t_L g895 ( 
.A(n_875),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_884),
.B(n_866),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_881),
.B(n_866),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_881),
.B(n_848),
.Y(n_898)
);

INVx1_ASAP7_75t_SL g899 ( 
.A(n_870),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_878),
.B(n_792),
.Y(n_900)
);

HB1xp67_ASAP7_75t_L g901 ( 
.A(n_870),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_890),
.B(n_867),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_890),
.B(n_867),
.Y(n_903)
);

OR2x2_ASAP7_75t_L g904 ( 
.A(n_894),
.B(n_880),
.Y(n_904)
);

BUFx3_ASAP7_75t_L g905 ( 
.A(n_895),
.Y(n_905)
);

OR2x2_ASAP7_75t_L g906 ( 
.A(n_894),
.B(n_880),
.Y(n_906)
);

OR2x2_ASAP7_75t_L g907 ( 
.A(n_891),
.B(n_876),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_891),
.B(n_897),
.Y(n_908)
);

INVxp67_ASAP7_75t_SL g909 ( 
.A(n_901),
.Y(n_909)
);

AND2x2_ASAP7_75t_L g910 ( 
.A(n_897),
.B(n_898),
.Y(n_910)
);

INVxp67_ASAP7_75t_SL g911 ( 
.A(n_901),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_892),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_893),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_897),
.B(n_872),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_902),
.B(n_874),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_902),
.B(n_889),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_893),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_SL g918 ( 
.A(n_899),
.B(n_883),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_L g919 ( 
.A(n_915),
.B(n_900),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_912),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_L g921 ( 
.A(n_916),
.B(n_907),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_912),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_908),
.B(n_896),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_910),
.B(n_898),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_913),
.Y(n_925)
);

INVx1_ASAP7_75t_SL g926 ( 
.A(n_905),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_913),
.Y(n_927)
);

OR2x2_ASAP7_75t_L g928 ( 
.A(n_907),
.B(n_903),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_917),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_920),
.Y(n_930)
);

AOI21xp33_ASAP7_75t_L g931 ( 
.A1(n_919),
.A2(n_865),
.B(n_862),
.Y(n_931)
);

NAND4xp25_ASAP7_75t_L g932 ( 
.A(n_919),
.B(n_879),
.C(n_877),
.D(n_886),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_922),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_923),
.B(n_908),
.Y(n_934)
);

INVxp67_ASAP7_75t_SL g935 ( 
.A(n_926),
.Y(n_935)
);

OAI22x1_ASAP7_75t_L g936 ( 
.A1(n_921),
.A2(n_918),
.B1(n_911),
.B2(n_909),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_925),
.B(n_910),
.Y(n_937)
);

OR2x2_ASAP7_75t_L g938 ( 
.A(n_928),
.B(n_904),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_927),
.Y(n_939)
);

OR2x2_ASAP7_75t_L g940 ( 
.A(n_924),
.B(n_904),
.Y(n_940)
);

NAND3xp33_ASAP7_75t_L g941 ( 
.A(n_929),
.B(n_906),
.C(n_885),
.Y(n_941)
);

AOI211xp5_ASAP7_75t_L g942 ( 
.A1(n_931),
.A2(n_826),
.B(n_921),
.C(n_906),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_938),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_937),
.B(n_923),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_934),
.B(n_914),
.Y(n_945)
);

OAI22xp33_ASAP7_75t_R g946 ( 
.A1(n_935),
.A2(n_856),
.B1(n_802),
.B2(n_857),
.Y(n_946)
);

AOI22xp33_ASAP7_75t_L g947 ( 
.A1(n_932),
.A2(n_931),
.B1(n_936),
.B2(n_869),
.Y(n_947)
);

OAI221xp5_ASAP7_75t_L g948 ( 
.A1(n_947),
.A2(n_942),
.B1(n_943),
.B2(n_946),
.C(n_941),
.Y(n_948)
);

A2O1A1Ixp33_ASAP7_75t_L g949 ( 
.A1(n_947),
.A2(n_869),
.B(n_887),
.C(n_883),
.Y(n_949)
);

AOI211x1_ASAP7_75t_L g950 ( 
.A1(n_944),
.A2(n_937),
.B(n_826),
.C(n_824),
.Y(n_950)
);

NOR3xp33_ASAP7_75t_L g951 ( 
.A(n_948),
.B(n_829),
.C(n_839),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_949),
.A2(n_799),
.B(n_930),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_951),
.B(n_950),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_952),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_954),
.Y(n_955)
);

HB1xp67_ASAP7_75t_L g956 ( 
.A(n_953),
.Y(n_956)
);

INVx2_ASAP7_75t_SL g957 ( 
.A(n_955),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_955),
.Y(n_958)
);

INVxp33_ASAP7_75t_L g959 ( 
.A(n_958),
.Y(n_959)
);

AOI22xp5_ASAP7_75t_L g960 ( 
.A1(n_957),
.A2(n_956),
.B1(n_857),
.B2(n_799),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_957),
.Y(n_961)
);

OA21x2_ASAP7_75t_L g962 ( 
.A1(n_961),
.A2(n_837),
.B(n_807),
.Y(n_962)
);

OAI21xp5_ASAP7_75t_L g963 ( 
.A1(n_960),
.A2(n_829),
.B(n_852),
.Y(n_963)
);

NOR4xp75_ASAP7_75t_L g964 ( 
.A(n_959),
.B(n_799),
.C(n_807),
.D(n_857),
.Y(n_964)
);

AOI22x1_ASAP7_75t_L g965 ( 
.A1(n_961),
.A2(n_856),
.B1(n_802),
.B2(n_862),
.Y(n_965)
);

XNOR2xp5_ASAP7_75t_L g966 ( 
.A(n_964),
.B(n_852),
.Y(n_966)
);

OAI22xp5_ASAP7_75t_L g967 ( 
.A1(n_965),
.A2(n_790),
.B1(n_945),
.B2(n_940),
.Y(n_967)
);

OA21x2_ASAP7_75t_L g968 ( 
.A1(n_963),
.A2(n_836),
.B(n_933),
.Y(n_968)
);

XNOR2xp5_ASAP7_75t_L g969 ( 
.A(n_962),
.B(n_873),
.Y(n_969)
);

OAI22x1_ASAP7_75t_L g970 ( 
.A1(n_962),
.A2(n_939),
.B1(n_858),
.B2(n_863),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_969),
.Y(n_971)
);

INVxp67_ASAP7_75t_SL g972 ( 
.A(n_966),
.Y(n_972)
);

OAI21xp33_ASAP7_75t_L g973 ( 
.A1(n_967),
.A2(n_905),
.B(n_887),
.Y(n_973)
);

INVxp67_ASAP7_75t_SL g974 ( 
.A(n_972),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_973),
.B(n_968),
.Y(n_975)
);

OR2x2_ASAP7_75t_L g976 ( 
.A(n_974),
.B(n_971),
.Y(n_976)
);

AOI21xp33_ASAP7_75t_L g977 ( 
.A1(n_976),
.A2(n_975),
.B(n_970),
.Y(n_977)
);


endmodule