module fake_jpeg_210_n_448 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_448);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_448;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_4),
.B(n_0),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx8_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_11),
.Y(n_41)
);

CKINVDCx11_ASAP7_75t_R g42 ( 
.A(n_4),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_6),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_12),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_21),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_48),
.B(n_50),
.Y(n_126)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_49),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_21),
.B(n_7),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_51),
.Y(n_101)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

BUFx4f_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_53),
.Y(n_108)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_54),
.Y(n_129)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_55),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_29),
.B(n_7),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_56),
.B(n_68),
.Y(n_127)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_57),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_16),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_58),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_59),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_60),
.Y(n_102)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_61),
.Y(n_112)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_16),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_62),
.Y(n_107)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_63),
.Y(n_128)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_64),
.Y(n_122)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_65),
.Y(n_130)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_66),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_16),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_67),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_34),
.B(n_7),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_69),
.Y(n_116)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_70),
.Y(n_131)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_26),
.Y(n_71)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_71),
.Y(n_109)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_72),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_73),
.Y(n_144)
);

BUFx24_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_74),
.Y(n_120)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_27),
.Y(n_75)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_75),
.Y(n_123)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_76),
.Y(n_136)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_22),
.Y(n_77)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_77),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_35),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_78),
.Y(n_147)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_26),
.Y(n_79)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_79),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_35),
.Y(n_80)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_80),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_29),
.B(n_8),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_81),
.B(n_83),
.Y(n_137)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_34),
.Y(n_82)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_82),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_41),
.B(n_42),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_37),
.Y(n_84)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_84),
.Y(n_134)
);

INVx2_ASAP7_75t_SL g85 ( 
.A(n_22),
.Y(n_85)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_85),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_35),
.Y(n_86)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_86),
.Y(n_145)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_22),
.Y(n_87)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_87),
.Y(n_140)
);

INVx4_ASAP7_75t_SL g88 ( 
.A(n_23),
.Y(n_88)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_88),
.Y(n_155)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_37),
.Y(n_89)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_89),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_25),
.Y(n_90)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_90),
.Y(n_139)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_23),
.Y(n_91)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_91),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_25),
.Y(n_92)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_92),
.Y(n_146)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_25),
.Y(n_93)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_93),
.Y(n_148)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_41),
.Y(n_94)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_94),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_23),
.A2(n_8),
.B1(n_2),
.B2(n_3),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_95),
.A2(n_17),
.B1(n_46),
.B2(n_43),
.Y(n_132)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_27),
.Y(n_96)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_96),
.Y(n_154)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_27),
.Y(n_97)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_97),
.Y(n_152)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_38),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_98),
.B(n_45),
.Y(n_100)
);

BUFx5_ASAP7_75t_L g99 ( 
.A(n_40),
.Y(n_99)
);

AND2x2_ASAP7_75t_SL g114 ( 
.A(n_99),
.B(n_44),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g184 ( 
.A(n_100),
.B(n_15),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_50),
.B(n_45),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_106),
.B(n_143),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_53),
.A2(n_44),
.B1(n_23),
.B2(n_19),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_110),
.A2(n_118),
.B1(n_149),
.B2(n_153),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_114),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_88),
.A2(n_44),
.B1(n_23),
.B2(n_19),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_48),
.B(n_47),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_124),
.B(n_68),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_132),
.A2(n_40),
.B1(n_80),
.B2(n_58),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_83),
.B(n_18),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_56),
.A2(n_44),
.B1(n_17),
.B2(n_38),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_81),
.A2(n_18),
.B1(n_46),
.B2(n_43),
.Y(n_153)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_148),
.Y(n_156)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_156),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_157),
.B(n_168),
.Y(n_216)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_108),
.Y(n_158)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_158),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_137),
.B(n_60),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_159),
.Y(n_199)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_135),
.Y(n_160)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_160),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_119),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_161),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_137),
.A2(n_47),
.B1(n_31),
.B2(n_85),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_162),
.A2(n_179),
.B1(n_188),
.B2(n_192),
.Y(n_207)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_131),
.Y(n_163)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_163),
.Y(n_209)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_104),
.Y(n_164)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_164),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_104),
.Y(n_165)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_165),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_120),
.Y(n_166)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_166),
.Y(n_212)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_116),
.Y(n_167)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_167),
.Y(n_230)
);

A2O1A1Ixp33_ASAP7_75t_L g168 ( 
.A1(n_126),
.A2(n_33),
.B(n_30),
.C(n_20),
.Y(n_168)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_115),
.Y(n_169)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_169),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_124),
.B(n_126),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_170),
.Y(n_205)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_133),
.Y(n_171)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_171),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_127),
.B(n_31),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_172),
.B(n_182),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_141),
.Y(n_173)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_173),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_149),
.A2(n_95),
.B1(n_90),
.B2(n_51),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_174),
.A2(n_141),
.B1(n_147),
.B2(n_144),
.Y(n_226)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_129),
.Y(n_175)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_175),
.Y(n_219)
);

INVx2_ASAP7_75t_SL g176 ( 
.A(n_155),
.Y(n_176)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_176),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_114),
.B(n_66),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_177),
.B(n_181),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_127),
.A2(n_33),
.B1(n_30),
.B2(n_20),
.Y(n_179)
);

AO22x2_ASAP7_75t_L g181 ( 
.A1(n_118),
.A2(n_74),
.B1(n_93),
.B2(n_62),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_130),
.B(n_44),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_150),
.Y(n_183)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_183),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_184),
.B(n_187),
.Y(n_203)
);

INVx13_ASAP7_75t_L g185 ( 
.A(n_102),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_185),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_103),
.B(n_15),
.Y(n_186)
);

OAI211xp5_ASAP7_75t_L g201 ( 
.A1(n_186),
.A2(n_191),
.B(n_180),
.C(n_151),
.Y(n_201)
);

AND2x2_ASAP7_75t_SL g187 ( 
.A(n_105),
.B(n_86),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_134),
.Y(n_188)
);

OAI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_110),
.A2(n_78),
.B1(n_73),
.B2(n_67),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_189),
.A2(n_147),
.B1(n_144),
.B2(n_101),
.Y(n_229)
);

BUFx12_ASAP7_75t_L g190 ( 
.A(n_121),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_190),
.Y(n_228)
);

BUFx12f_ASAP7_75t_L g192 ( 
.A(n_136),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_139),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_193),
.A2(n_194),
.B1(n_196),
.B2(n_197),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_121),
.Y(n_194)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_146),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_112),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_109),
.A2(n_40),
.B1(n_2),
.B2(n_3),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_198),
.A2(n_138),
.B1(n_111),
.B2(n_123),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_201),
.B(n_177),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_168),
.A2(n_122),
.B(n_117),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_206),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_178),
.A2(n_125),
.B1(n_145),
.B2(n_101),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_213),
.A2(n_165),
.B1(n_173),
.B2(n_182),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_186),
.A2(n_181),
.B1(n_191),
.B2(n_128),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_223),
.A2(n_226),
.B1(n_229),
.B2(n_177),
.Y(n_234)
);

BUFx2_ASAP7_75t_L g256 ( 
.A(n_225),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_174),
.A2(n_142),
.B1(n_140),
.B2(n_113),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_SL g251 ( 
.A(n_227),
.B(n_197),
.C(n_185),
.Y(n_251)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_221),
.Y(n_232)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_232),
.Y(n_263)
);

BUFx24_ASAP7_75t_SL g233 ( 
.A(n_205),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_233),
.B(n_255),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_L g268 ( 
.A1(n_234),
.A2(n_220),
.B1(n_224),
.B2(n_218),
.Y(n_268)
);

MAJx2_ASAP7_75t_L g235 ( 
.A(n_204),
.B(n_157),
.C(n_172),
.Y(n_235)
);

MAJx2_ASAP7_75t_L g264 ( 
.A(n_235),
.B(n_222),
.C(n_208),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_236),
.A2(n_251),
.B1(n_217),
.B2(n_212),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_237),
.A2(n_239),
.B1(n_208),
.B2(n_215),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_202),
.A2(n_223),
.B1(n_213),
.B2(n_226),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_205),
.B(n_195),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_240),
.B(n_245),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_203),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_241),
.B(n_242),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_217),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_202),
.A2(n_181),
.B1(n_160),
.B2(n_188),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_243),
.A2(n_246),
.B1(n_254),
.B2(n_237),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_204),
.B(n_176),
.C(n_187),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_244),
.B(n_241),
.C(n_258),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_206),
.B(n_187),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_202),
.A2(n_181),
.B1(n_184),
.B2(n_193),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_216),
.B(n_171),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_247),
.B(n_253),
.Y(n_269)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_221),
.Y(n_248)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_248),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_201),
.B(n_176),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_249),
.Y(n_271)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_210),
.Y(n_250)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_250),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_199),
.B(n_158),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_252),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_216),
.B(n_163),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_203),
.A2(n_196),
.B1(n_107),
.B2(n_156),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_219),
.B(n_169),
.Y(n_255)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_210),
.Y(n_257)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_257),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_203),
.B(n_167),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_258),
.B(n_215),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_246),
.A2(n_229),
.B1(n_207),
.B2(n_219),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_259),
.B(n_273),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_235),
.B(n_222),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_260),
.B(n_282),
.C(n_284),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_255),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_262),
.B(n_209),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_264),
.B(n_244),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_249),
.Y(n_267)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_267),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_268),
.A2(n_254),
.B1(n_232),
.B2(n_248),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_238),
.A2(n_249),
.B(n_236),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_270),
.B(n_272),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_243),
.A2(n_214),
.B1(n_164),
.B2(n_218),
.Y(n_273)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_274),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_236),
.A2(n_224),
.B1(n_145),
.B2(n_125),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_276),
.B(n_281),
.Y(n_290)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_250),
.Y(n_279)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_279),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_245),
.A2(n_228),
.B(n_230),
.Y(n_283)
);

OAI21xp33_ASAP7_75t_SL g310 ( 
.A1(n_283),
.A2(n_271),
.B(n_281),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_235),
.B(n_209),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_285),
.B(n_234),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_278),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_286),
.B(n_296),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_263),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_289),
.Y(n_315)
);

INVxp33_ASAP7_75t_L g319 ( 
.A(n_292),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_262),
.B(n_242),
.Y(n_293)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_293),
.Y(n_312)
);

INVxp33_ASAP7_75t_L g294 ( 
.A(n_280),
.Y(n_294)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_294),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_266),
.B(n_240),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_295),
.B(n_298),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_278),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_297),
.B(n_269),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_266),
.B(n_211),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_261),
.B(n_211),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_299),
.B(n_301),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_260),
.B(n_253),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_264),
.B(n_247),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_302),
.B(n_311),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_284),
.B(n_257),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_303),
.B(n_264),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_282),
.B(n_239),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_304),
.B(n_270),
.C(n_267),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_307),
.A2(n_309),
.B1(n_285),
.B2(n_273),
.Y(n_333)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_308),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_274),
.A2(n_256),
.B1(n_220),
.B2(n_251),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_310),
.A2(n_283),
.B(n_272),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_275),
.B(n_228),
.Y(n_311)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_293),
.Y(n_314)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_314),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_318),
.B(n_324),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_286),
.B(n_230),
.Y(n_320)
);

CKINVDCx16_ASAP7_75t_R g342 ( 
.A(n_320),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_321),
.B(n_325),
.C(n_231),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_322),
.A2(n_336),
.B1(n_288),
.B2(n_308),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_296),
.B(n_269),
.Y(n_323)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_323),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_305),
.B(n_263),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_304),
.B(n_231),
.Y(n_327)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_327),
.Y(n_340)
);

BUFx5_ASAP7_75t_L g329 ( 
.A(n_300),
.Y(n_329)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_329),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_300),
.A2(n_259),
.B(n_265),
.Y(n_330)
);

INVxp33_ASAP7_75t_L g346 ( 
.A(n_330),
.Y(n_346)
);

BUFx24_ASAP7_75t_SL g331 ( 
.A(n_288),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_331),
.B(n_212),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_307),
.A2(n_287),
.B1(n_291),
.B2(n_300),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_332),
.A2(n_334),
.B1(n_337),
.B2(n_292),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_333),
.A2(n_200),
.B1(n_107),
.B2(n_192),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_307),
.A2(n_256),
.B1(n_265),
.B2(n_275),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_291),
.A2(n_287),
.B1(n_309),
.B2(n_290),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_290),
.A2(n_256),
.B1(n_277),
.B2(n_279),
.Y(n_337)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_313),
.Y(n_341)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_341),
.Y(n_364)
);

BUFx3_ASAP7_75t_L g343 ( 
.A(n_326),
.Y(n_343)
);

HB1xp67_ASAP7_75t_L g378 ( 
.A(n_343),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_344),
.B(n_356),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_323),
.B(n_306),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_347),
.B(n_348),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_313),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_349),
.A2(n_352),
.B1(n_353),
.B2(n_336),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_SL g375 ( 
.A(n_350),
.B(n_359),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_SL g351 ( 
.A(n_318),
.B(n_297),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_351),
.B(n_357),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_332),
.A2(n_276),
.B1(n_306),
.B2(n_277),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_319),
.A2(n_303),
.B1(n_305),
.B2(n_289),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_312),
.Y(n_354)
);

INVxp67_ASAP7_75t_SL g376 ( 
.A(n_354),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_325),
.B(n_289),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_321),
.B(n_200),
.C(n_220),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_358),
.B(n_324),
.C(n_319),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_315),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_360),
.A2(n_334),
.B1(n_337),
.B2(n_312),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_362),
.B(n_374),
.C(n_367),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_363),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_365),
.A2(n_352),
.B1(n_355),
.B2(n_340),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_339),
.B(n_322),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_SL g387 ( 
.A(n_366),
.B(n_367),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_339),
.B(n_330),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_357),
.B(n_314),
.C(n_335),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_369),
.B(n_379),
.Y(n_384)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_346),
.A2(n_333),
.B(n_329),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_SL g382 ( 
.A1(n_371),
.A2(n_346),
.B(n_355),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_349),
.A2(n_317),
.B1(n_328),
.B2(n_316),
.Y(n_372)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_372),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_345),
.A2(n_315),
.B1(n_166),
.B2(n_192),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_373),
.B(n_377),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_353),
.B(n_152),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_348),
.B(n_11),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_SL g379 ( 
.A(n_343),
.B(n_154),
.Y(n_379)
);

CKINVDCx16_ASAP7_75t_R g380 ( 
.A(n_347),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_380),
.B(n_342),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_L g405 ( 
.A1(n_382),
.A2(n_366),
.B(n_190),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_383),
.B(n_374),
.Y(n_400)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_364),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_385),
.B(n_392),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_370),
.A2(n_364),
.B1(n_338),
.B2(n_345),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_386),
.A2(n_389),
.B1(n_190),
.B2(n_3),
.Y(n_406)
);

AOI22xp33_ASAP7_75t_SL g404 ( 
.A1(n_391),
.A2(n_397),
.B1(n_377),
.B2(n_365),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_362),
.B(n_356),
.C(n_358),
.Y(n_392)
);

BUFx4f_ASAP7_75t_SL g393 ( 
.A(n_378),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_393),
.B(n_395),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_SL g394 ( 
.A1(n_371),
.A2(n_360),
.B(n_351),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_SL g408 ( 
.A1(n_394),
.A2(n_5),
.B(n_6),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_375),
.B(n_9),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_370),
.B(n_9),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_396),
.B(n_3),
.Y(n_407)
);

INVx11_ASAP7_75t_L g397 ( 
.A(n_376),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_393),
.B(n_369),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_398),
.B(n_399),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_392),
.B(n_368),
.C(n_361),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_400),
.B(n_410),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_383),
.B(n_368),
.C(n_361),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_403),
.B(n_407),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_L g415 ( 
.A1(n_404),
.A2(n_381),
.B(n_389),
.Y(n_415)
);

OR2x2_ASAP7_75t_L g420 ( 
.A(n_405),
.B(n_406),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_L g422 ( 
.A1(n_408),
.A2(n_396),
.B(n_386),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_384),
.B(n_5),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_409),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_387),
.B(n_14),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_393),
.B(n_5),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_411),
.A2(n_412),
.B1(n_385),
.B2(n_13),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_390),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_412)
);

NAND3xp33_ASAP7_75t_SL g413 ( 
.A(n_405),
.B(n_382),
.C(n_394),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g431 ( 
.A1(n_413),
.A2(n_13),
.B(n_1),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_415),
.A2(n_406),
.B1(n_412),
.B2(n_410),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_401),
.B(n_388),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_418),
.B(n_419),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_399),
.B(n_390),
.C(n_387),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_422),
.B(n_424),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_400),
.B(n_381),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_423),
.B(n_397),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_414),
.B(n_403),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_426),
.B(n_427),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_421),
.B(n_402),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_428),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_429),
.B(n_433),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_416),
.B(n_13),
.Y(n_430)
);

AOI21xp33_ASAP7_75t_L g438 ( 
.A1(n_430),
.A2(n_431),
.B(n_1),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_423),
.B(n_1),
.C(n_419),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_425),
.B(n_417),
.C(n_420),
.Y(n_436)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_436),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_433),
.B(n_420),
.C(n_413),
.Y(n_437)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_437),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_SL g440 ( 
.A1(n_438),
.A2(n_432),
.B(n_429),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_440),
.B(n_439),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_442),
.Y(n_443)
);

FAx1_ASAP7_75t_R g445 ( 
.A(n_443),
.B(n_444),
.CI(n_441),
.CON(n_445),
.SN(n_445)
);

BUFx24_ASAP7_75t_SL g446 ( 
.A(n_445),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_SL g447 ( 
.A1(n_446),
.A2(n_435),
.B(n_434),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_447),
.B(n_435),
.Y(n_448)
);


endmodule