module fake_jpeg_923_n_74 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_74);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_74;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_73;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_48;
wire n_35;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_36;
wire n_11;
wire n_62;
wire n_25;
wire n_17;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

BUFx12_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_8),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_4),
.B(n_3),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_0),
.B(n_2),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_22),
.B(n_23),
.Y(n_40)
);

OR2x4_ASAP7_75t_L g23 ( 
.A(n_16),
.B(n_2),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_16),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_27),
.B(n_28),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_14),
.B(n_3),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_17),
.B(n_15),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_30),
.A2(n_15),
.B1(n_17),
.B2(n_19),
.Y(n_33)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_30),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_32),
.B(n_26),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_33),
.A2(n_37),
.B1(n_31),
.B2(n_24),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_23),
.A2(n_15),
.B1(n_19),
.B2(n_12),
.Y(n_37)
);

CKINVDCx12_ASAP7_75t_R g41 ( 
.A(n_26),
.Y(n_41)
);

OAI21xp33_ASAP7_75t_L g50 ( 
.A1(n_41),
.A2(n_21),
.B(n_18),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_37),
.A2(n_29),
.B1(n_25),
.B2(n_12),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_45),
.Y(n_52)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_46),
.Y(n_56)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_47),
.A2(n_49),
.B1(n_50),
.B2(n_51),
.Y(n_54)
);

AOI21xp33_ASAP7_75t_L g48 ( 
.A1(n_40),
.A2(n_21),
.B(n_18),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_33),
.C(n_38),
.Y(n_57)
);

AND2x6_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_35),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_57),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_52),
.A2(n_45),
.B1(n_44),
.B2(n_47),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_58),
.A2(n_61),
.B1(n_54),
.B2(n_57),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_55),
.A2(n_34),
.B1(n_39),
.B2(n_38),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_59),
.B(n_56),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_62),
.B(n_63),
.Y(n_66)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_60),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_64),
.B(n_65),
.C(n_34),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_59),
.B(n_53),
.Y(n_65)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_67),
.Y(n_69)
);

OAI22x1_ASAP7_75t_L g68 ( 
.A1(n_66),
.A2(n_64),
.B1(n_5),
.B2(n_7),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_68),
.B(n_4),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_70),
.B(n_7),
.Y(n_71)
);

AOI322xp5_ASAP7_75t_L g72 ( 
.A1(n_71),
.A2(n_9),
.A3(n_10),
.B1(n_11),
.B2(n_39),
.C1(n_69),
.C2(n_70),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_9),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_11),
.Y(n_74)
);


endmodule