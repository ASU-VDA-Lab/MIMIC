module fake_jpeg_28103_n_172 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_172);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_172;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_26),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_19),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_31),
.Y(n_56)
);

BUFx4f_ASAP7_75t_L g57 ( 
.A(n_8),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_2),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_11),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_34),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_15),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_0),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_43),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_1),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_0),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_2),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_13),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_10),
.Y(n_71)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_8),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_16),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_1),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_74),
.B(n_78),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_70),
.Y(n_75)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_61),
.Y(n_78)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_50),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_80),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_79),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_81),
.Y(n_112)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_82),
.B(n_71),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_76),
.Y(n_83)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_83),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_75),
.A2(n_72),
.B1(n_59),
.B2(n_63),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_85),
.A2(n_91),
.B1(n_62),
.B2(n_55),
.Y(n_102)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_75),
.A2(n_53),
.B1(n_66),
.B2(n_57),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_94),
.Y(n_96)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_93),
.Y(n_97)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_84),
.A2(n_73),
.B1(n_65),
.B2(n_78),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_99),
.A2(n_101),
.B1(n_102),
.B2(n_107),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_95),
.B(n_56),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_104),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_91),
.A2(n_62),
.B1(n_51),
.B2(n_56),
.Y(n_101)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_81),
.Y(n_103)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_103),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_67),
.Y(n_104)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_89),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_106),
.A2(n_113),
.B1(n_88),
.B2(n_92),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_88),
.A2(n_51),
.B1(n_54),
.B2(n_69),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_111),
.A2(n_71),
.B1(n_69),
.B2(n_68),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_86),
.B(n_52),
.Y(n_113)
);

BUFx5_ASAP7_75t_L g114 ( 
.A(n_108),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_114),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_116),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_117),
.A2(n_123),
.B1(n_4),
.B2(n_5),
.Y(n_135)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_110),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_119),
.Y(n_133)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_109),
.Y(n_121)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_121),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_98),
.A2(n_58),
.B1(n_4),
.B2(n_5),
.Y(n_123)
);

O2A1O1Ixp33_ASAP7_75t_L g125 ( 
.A1(n_124),
.A2(n_112),
.B(n_105),
.C(n_100),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_125),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_120),
.B(n_113),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_126),
.B(n_127),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_118),
.B(n_3),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_122),
.B(n_104),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_130),
.B(n_132),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_115),
.B(n_112),
.Y(n_132)
);

OAI32xp33_ASAP7_75t_L g134 ( 
.A1(n_117),
.A2(n_25),
.A3(n_48),
.B1(n_45),
.B2(n_42),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_134),
.B(n_123),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_135),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_136),
.B(n_137),
.Y(n_153)
);

OR2x2_ASAP7_75t_L g137 ( 
.A(n_125),
.B(n_121),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_133),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_138),
.B(n_141),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_133),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_140),
.Y(n_154)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_143),
.Y(n_151)
);

OAI22x1_ASAP7_75t_SL g144 ( 
.A1(n_134),
.A2(n_28),
.B1(n_41),
.B2(n_12),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_144),
.Y(n_149)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_128),
.Y(n_145)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_145),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_128),
.B(n_10),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_146),
.B(n_147),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_131),
.A2(n_11),
.B1(n_14),
.B2(n_17),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_129),
.B(n_49),
.Y(n_148)
);

MAJx2_ASAP7_75t_L g150 ( 
.A(n_148),
.B(n_18),
.C(n_20),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_150),
.A2(n_146),
.B1(n_156),
.B2(n_139),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_153),
.B(n_142),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_157),
.B(n_158),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_154),
.A2(n_137),
.B(n_144),
.Y(n_158)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_159),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_160),
.Y(n_162)
);

INVxp33_ASAP7_75t_L g163 ( 
.A(n_162),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_163),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_164),
.A2(n_161),
.B1(n_151),
.B2(n_155),
.Y(n_165)
);

OAI21x1_ASAP7_75t_SL g166 ( 
.A1(n_165),
.A2(n_149),
.B(n_152),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_166),
.A2(n_149),
.B(n_157),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_167),
.A2(n_150),
.B(n_23),
.Y(n_168)
);

A2O1A1O1Ixp25_ASAP7_75t_L g169 ( 
.A1(n_168),
.A2(n_22),
.B(n_27),
.C(n_29),
.D(n_30),
.Y(n_169)
);

A2O1A1Ixp33_ASAP7_75t_SL g170 ( 
.A1(n_169),
.A2(n_32),
.B(n_35),
.C(n_36),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_170),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_171),
.A2(n_39),
.B(n_40),
.Y(n_172)
);


endmodule