module real_aes_6367_n_222 (n_17, n_28, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_165, n_51, n_195, n_176, n_27, n_163, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_84, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_16, n_116, n_94, n_39, n_5, n_45, n_60, n_38, n_155, n_118, n_143, n_139, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_222);
input n_17;
input n_28;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_84;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_16;
input n_116;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_222;
wire n_480;
wire n_476;
wire n_599;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_673;
wire n_386;
wire n_518;
wire n_254;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_461;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_271;
wire n_489;
wire n_548;
wire n_678;
wire n_427;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_578;
wire n_372;
wire n_528;
wire n_495;
wire n_370;
wire n_384;
wire n_352;
wire n_467;
wire n_327;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_693;
wire n_281;
wire n_496;
wire n_468;
wire n_234;
wire n_284;
wire n_532;
wire n_316;
wire n_656;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_310;
wire n_455;
wire n_504;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_565;
wire n_443;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_331;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_527;
wire n_434;
wire n_502;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_246;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_269;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_498;
wire n_691;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_472;
wire n_452;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_266;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_705;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_541;
wire n_224;
wire n_546;
wire n_587;
wire n_639;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_228;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_241;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
CKINVDCx20_ASAP7_75t_R g666 ( .A(n_0), .Y(n_666) );
CKINVDCx20_ASAP7_75t_R g271 ( .A(n_1), .Y(n_271) );
XOR2x2_ASAP7_75t_L g416 ( .A(n_2), .B(n_417), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g298 ( .A1(n_3), .A2(n_14), .B1(n_299), .B2(n_304), .Y(n_298) );
AOI22xp33_ASAP7_75t_L g395 ( .A1(n_4), .A2(n_144), .B1(n_360), .B2(n_363), .Y(n_395) );
CKINVDCx20_ASAP7_75t_R g569 ( .A(n_5), .Y(n_569) );
INVx1_ASAP7_75t_L g386 ( .A(n_6), .Y(n_386) );
AOI22xp5_ASAP7_75t_L g239 ( .A1(n_7), .A2(n_240), .B1(n_333), .B2(n_334), .Y(n_239) );
INVx1_ASAP7_75t_L g333 ( .A(n_7), .Y(n_333) );
AOI222xp33_ASAP7_75t_L g434 ( .A1(n_8), .A2(n_23), .B1(n_178), .B2(n_266), .C1(n_435), .C2(n_437), .Y(n_434) );
AOI22xp5_ASAP7_75t_L g509 ( .A1(n_9), .A2(n_192), .B1(n_274), .B2(n_422), .Y(n_509) );
CKINVDCx20_ASAP7_75t_R g516 ( .A(n_10), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_11), .B(n_392), .Y(n_391) );
AOI22xp33_ASAP7_75t_L g425 ( .A1(n_12), .A2(n_62), .B1(n_426), .B2(n_428), .Y(n_425) );
AOI22xp33_ASAP7_75t_SL g487 ( .A1(n_13), .A2(n_82), .B1(n_363), .B2(n_422), .Y(n_487) );
AOI22xp33_ASAP7_75t_SL g370 ( .A1(n_15), .A2(n_52), .B1(n_325), .B2(n_329), .Y(n_370) );
AOI22xp33_ASAP7_75t_SL g542 ( .A1(n_16), .A2(n_181), .B1(n_543), .B2(n_544), .Y(n_542) );
CKINVDCx20_ASAP7_75t_R g665 ( .A(n_17), .Y(n_665) );
XOR2x2_ASAP7_75t_L g440 ( .A(n_18), .B(n_441), .Y(n_440) );
AOI22xp33_ASAP7_75t_L g358 ( .A1(n_19), .A2(n_164), .B1(n_359), .B2(n_362), .Y(n_358) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_20), .A2(n_74), .B1(n_437), .B2(n_599), .Y(n_598) );
AO22x2_ASAP7_75t_L g248 ( .A1(n_21), .A2(n_69), .B1(n_249), .B2(n_250), .Y(n_248) );
INVx1_ASAP7_75t_L g653 ( .A(n_21), .Y(n_653) );
AOI22xp33_ASAP7_75t_L g714 ( .A1(n_22), .A2(n_63), .B1(n_319), .B2(n_609), .Y(n_714) );
AOI222xp33_ASAP7_75t_L g494 ( .A1(n_24), .A2(n_81), .B1(n_104), .B2(n_273), .C1(n_342), .C2(n_435), .Y(n_494) );
CKINVDCx20_ASAP7_75t_R g412 ( .A(n_25), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_26), .A2(n_128), .B1(n_326), .B2(n_505), .Y(n_504) );
AOI22xp33_ASAP7_75t_SL g534 ( .A1(n_27), .A2(n_29), .B1(n_299), .B2(n_432), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g489 ( .A1(n_28), .A2(n_186), .B1(n_490), .B2(n_491), .Y(n_489) );
INVx1_ASAP7_75t_L g632 ( .A(n_30), .Y(n_632) );
AOI222xp33_ASAP7_75t_L g514 ( .A1(n_31), .A2(n_73), .B1(n_201), .B2(n_385), .C1(n_389), .C2(n_515), .Y(n_514) );
CKINVDCx20_ASAP7_75t_R g701 ( .A(n_32), .Y(n_701) );
AOI22xp33_ASAP7_75t_SL g529 ( .A1(n_33), .A2(n_53), .B1(n_362), .B2(n_530), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g419 ( .A1(n_34), .A2(n_35), .B1(n_392), .B2(n_420), .Y(n_419) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_36), .A2(n_133), .B1(n_300), .B2(n_478), .Y(n_477) );
AO22x2_ASAP7_75t_L g252 ( .A1(n_37), .A2(n_70), .B1(n_249), .B2(n_253), .Y(n_252) );
INVx1_ASAP7_75t_L g654 ( .A(n_37), .Y(n_654) );
CKINVDCx20_ASAP7_75t_R g573 ( .A(n_38), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g409 ( .A1(n_39), .A2(n_110), .B1(n_322), .B2(n_410), .Y(n_409) );
AOI22xp33_ASAP7_75t_SL g606 ( .A1(n_40), .A2(n_42), .B1(n_463), .B2(n_607), .Y(n_606) );
AOI22xp33_ASAP7_75t_SL g602 ( .A1(n_41), .A2(n_95), .B1(n_426), .B2(n_490), .Y(n_602) );
AOI22xp33_ASAP7_75t_SL g594 ( .A1(n_43), .A2(n_213), .B1(n_273), .B2(n_435), .Y(n_594) );
CKINVDCx20_ASAP7_75t_R g678 ( .A(n_44), .Y(n_678) );
AOI22xp33_ASAP7_75t_L g324 ( .A1(n_45), .A2(n_123), .B1(n_325), .B2(n_329), .Y(n_324) );
AOI22xp33_ASAP7_75t_L g471 ( .A1(n_46), .A2(n_187), .B1(n_472), .B2(n_473), .Y(n_471) );
CKINVDCx20_ASAP7_75t_R g553 ( .A(n_47), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g318 ( .A1(n_48), .A2(n_96), .B1(n_319), .B2(n_322), .Y(n_318) );
AOI22xp33_ASAP7_75t_SL g603 ( .A1(n_49), .A2(n_163), .B1(n_329), .B2(n_604), .Y(n_603) );
XOR2x2_ASAP7_75t_L g589 ( .A(n_50), .B(n_590), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g662 ( .A1(n_51), .A2(n_172), .B1(n_402), .B2(n_663), .Y(n_662) );
CKINVDCx20_ASAP7_75t_R g558 ( .A(n_54), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_55), .B(n_456), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g309 ( .A1(n_56), .A2(n_71), .B1(n_310), .B2(n_314), .Y(n_309) );
AOI22xp33_ASAP7_75t_SL g387 ( .A1(n_57), .A2(n_211), .B1(n_388), .B2(n_389), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_58), .B(n_394), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g433 ( .A1(n_59), .A2(n_169), .B1(n_320), .B2(n_402), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_60), .B(n_351), .Y(n_350) );
AOI22xp33_ASAP7_75t_L g492 ( .A1(n_61), .A2(n_135), .B1(n_368), .B2(n_493), .Y(n_492) );
CKINVDCx20_ASAP7_75t_R g680 ( .A(n_64), .Y(n_680) );
AOI22xp33_ASAP7_75t_SL g365 ( .A1(n_65), .A2(n_94), .B1(n_366), .B2(n_369), .Y(n_365) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_66), .A2(n_205), .B1(n_394), .B2(n_532), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_67), .A2(n_214), .B1(n_353), .B2(n_454), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g715 ( .A1(n_68), .A2(n_132), .B1(n_304), .B2(n_323), .Y(n_715) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_72), .A2(n_208), .B1(n_369), .B2(n_403), .Y(n_506) );
INVx1_ASAP7_75t_L g230 ( .A(n_75), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_76), .B(n_453), .Y(n_452) );
AOI22xp5_ASAP7_75t_L g661 ( .A1(n_77), .A2(n_105), .B1(n_490), .B2(n_541), .Y(n_661) );
CKINVDCx20_ASAP7_75t_R g527 ( .A(n_78), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_79), .B(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g228 ( .A(n_80), .Y(n_228) );
AOI22xp33_ASAP7_75t_SL g540 ( .A1(n_83), .A2(n_212), .B1(n_512), .B2(n_541), .Y(n_540) );
CKINVDCx20_ASAP7_75t_R g561 ( .A(n_84), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g405 ( .A1(n_85), .A2(n_124), .B1(n_406), .B2(n_408), .Y(n_405) );
AOI22xp33_ASAP7_75t_L g424 ( .A1(n_86), .A2(n_188), .B1(n_330), .B2(n_376), .Y(n_424) );
CKINVDCx20_ASAP7_75t_R g445 ( .A(n_87), .Y(n_445) );
AOI22xp33_ASAP7_75t_L g461 ( .A1(n_88), .A2(n_156), .B1(n_368), .B2(n_462), .Y(n_461) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_89), .A2(n_143), .B1(n_312), .B2(n_320), .Y(n_513) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_90), .A2(n_98), .B1(n_376), .B2(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g634 ( .A(n_91), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_92), .B(n_282), .Y(n_281) );
AOI222xp33_ASAP7_75t_L g581 ( .A1(n_93), .A2(n_109), .B1(n_175), .B2(n_458), .C1(n_582), .C2(n_584), .Y(n_581) );
CKINVDCx20_ASAP7_75t_R g565 ( .A(n_97), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_99), .B(n_282), .Y(n_708) );
CKINVDCx20_ASAP7_75t_R g711 ( .A(n_100), .Y(n_711) );
AOI22xp33_ASAP7_75t_L g421 ( .A1(n_101), .A2(n_106), .B1(n_274), .B2(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g627 ( .A(n_102), .Y(n_627) );
CKINVDCx20_ASAP7_75t_R g673 ( .A(n_103), .Y(n_673) );
AOI22xp33_ASAP7_75t_L g431 ( .A1(n_107), .A2(n_217), .B1(n_406), .B2(n_432), .Y(n_431) );
AO22x2_ASAP7_75t_L g549 ( .A1(n_108), .A2(n_550), .B1(n_585), .B2(n_586), .Y(n_549) );
CKINVDCx20_ASAP7_75t_R g585 ( .A(n_108), .Y(n_585) );
XNOR2xp5_ASAP7_75t_L g656 ( .A(n_111), .B(n_657), .Y(n_656) );
AOI22xp33_ASAP7_75t_SL g535 ( .A1(n_112), .A2(n_200), .B1(n_536), .B2(n_538), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g615 ( .A1(n_113), .A2(n_116), .B1(n_616), .B2(n_617), .Y(n_615) );
INVx1_ASAP7_75t_L g630 ( .A(n_114), .Y(n_630) );
CKINVDCx20_ASAP7_75t_R g523 ( .A(n_115), .Y(n_523) );
AOI222xp33_ASAP7_75t_L g636 ( .A1(n_117), .A2(n_150), .B1(n_154), .B2(n_267), .C1(n_274), .C2(n_282), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_118), .B(n_458), .Y(n_681) );
CKINVDCx20_ASAP7_75t_R g704 ( .A(n_119), .Y(n_704) );
AOI221xp5_ASAP7_75t_L g575 ( .A1(n_120), .A2(n_221), .B1(n_532), .B2(n_576), .C(n_577), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g457 ( .A1(n_121), .A2(n_198), .B1(n_359), .B2(n_458), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_122), .A2(n_161), .B1(n_465), .B2(n_466), .Y(n_464) );
AOI22xp33_ASAP7_75t_SL g377 ( .A1(n_125), .A2(n_153), .B1(n_378), .B2(n_379), .Y(n_377) );
INVx2_ASAP7_75t_L g231 ( .A(n_126), .Y(n_231) );
AOI22xp33_ASAP7_75t_L g446 ( .A1(n_127), .A2(n_193), .B1(n_447), .B2(n_448), .Y(n_446) );
CKINVDCx20_ASAP7_75t_R g707 ( .A(n_129), .Y(n_707) );
CKINVDCx20_ASAP7_75t_R g259 ( .A(n_130), .Y(n_259) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_131), .A2(n_203), .B1(n_480), .B2(n_481), .Y(n_479) );
AOI22xp5_ASAP7_75t_L g468 ( .A1(n_134), .A2(n_177), .B1(n_314), .B2(n_469), .Y(n_468) );
AND2x6_ASAP7_75t_L g227 ( .A(n_136), .B(n_228), .Y(n_227) );
HB1xp67_ASAP7_75t_L g647 ( .A(n_136), .Y(n_647) );
AO22x2_ASAP7_75t_L g258 ( .A1(n_137), .A2(n_185), .B1(n_249), .B2(n_253), .Y(n_258) );
AOI22xp33_ASAP7_75t_L g619 ( .A1(n_138), .A2(n_209), .B1(n_469), .B2(n_473), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g717 ( .A1(n_139), .A2(n_170), .B1(n_299), .B2(n_432), .Y(n_717) );
AOI211xp5_ASAP7_75t_L g222 ( .A1(n_140), .A2(n_223), .B(n_232), .C(n_655), .Y(n_222) );
AOI22xp33_ASAP7_75t_SL g345 ( .A1(n_141), .A2(n_167), .B1(n_282), .B2(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_142), .B(n_454), .Y(n_486) );
AOI22xp33_ASAP7_75t_SL g372 ( .A1(n_145), .A2(n_219), .B1(n_373), .B2(n_374), .Y(n_372) );
CKINVDCx20_ASAP7_75t_R g580 ( .A(n_146), .Y(n_580) );
CKINVDCx20_ASAP7_75t_R g685 ( .A(n_147), .Y(n_685) );
INVx1_ASAP7_75t_L g621 ( .A(n_148), .Y(n_621) );
AOI22xp33_ASAP7_75t_L g718 ( .A1(n_149), .A2(n_191), .B1(n_604), .B2(n_719), .Y(n_718) );
CKINVDCx20_ASAP7_75t_R g495 ( .A(n_151), .Y(n_495) );
INVx1_ASAP7_75t_L g637 ( .A(n_152), .Y(n_637) );
AO22x2_ASAP7_75t_L g256 ( .A1(n_155), .A2(n_194), .B1(n_249), .B2(n_250), .Y(n_256) );
CKINVDCx20_ASAP7_75t_R g676 ( .A(n_157), .Y(n_676) );
AOI22xp33_ASAP7_75t_SL g398 ( .A1(n_158), .A2(n_196), .B1(n_399), .B2(n_400), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_159), .B(n_351), .Y(n_596) );
CKINVDCx20_ASAP7_75t_R g286 ( .A(n_160), .Y(n_286) );
AOI22xp33_ASAP7_75t_SL g401 ( .A1(n_162), .A2(n_165), .B1(n_402), .B2(n_403), .Y(n_401) );
CKINVDCx20_ASAP7_75t_R g289 ( .A(n_166), .Y(n_289) );
AOI22xp33_ASAP7_75t_L g624 ( .A1(n_168), .A2(n_199), .B1(n_515), .B2(n_599), .Y(n_624) );
CKINVDCx20_ASAP7_75t_R g280 ( .A(n_171), .Y(n_280) );
CKINVDCx20_ASAP7_75t_R g669 ( .A(n_173), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_174), .B(n_623), .Y(n_622) );
AOI22xp33_ASAP7_75t_SL g608 ( .A1(n_176), .A2(n_215), .B1(n_505), .B2(n_609), .Y(n_608) );
CKINVDCx20_ASAP7_75t_R g566 ( .A(n_179), .Y(n_566) );
CKINVDCx20_ASAP7_75t_R g668 ( .A(n_180), .Y(n_668) );
CKINVDCx20_ASAP7_75t_R g683 ( .A(n_182), .Y(n_683) );
CKINVDCx20_ASAP7_75t_R g710 ( .A(n_183), .Y(n_710) );
XOR2x2_ASAP7_75t_L g337 ( .A(n_184), .B(n_338), .Y(n_337) );
NOR2xp33_ASAP7_75t_L g651 ( .A(n_185), .B(n_652), .Y(n_651) );
CKINVDCx20_ASAP7_75t_R g483 ( .A(n_189), .Y(n_483) );
CKINVDCx20_ASAP7_75t_R g578 ( .A(n_190), .Y(n_578) );
INVx1_ASAP7_75t_L g650 ( .A(n_194), .Y(n_650) );
INVx1_ASAP7_75t_L g344 ( .A(n_195), .Y(n_344) );
OA22x2_ASAP7_75t_L g518 ( .A1(n_197), .A2(n_519), .B1(n_520), .B2(n_546), .Y(n_518) );
CKINVDCx20_ASAP7_75t_R g519 ( .A(n_197), .Y(n_519) );
CKINVDCx20_ASAP7_75t_R g593 ( .A(n_202), .Y(n_593) );
CKINVDCx20_ASAP7_75t_R g525 ( .A(n_204), .Y(n_525) );
CKINVDCx20_ASAP7_75t_R g243 ( .A(n_206), .Y(n_243) );
INVx1_ASAP7_75t_L g249 ( .A(n_207), .Y(n_249) );
INVx1_ASAP7_75t_L g251 ( .A(n_207), .Y(n_251) );
CKINVDCx20_ASAP7_75t_R g706 ( .A(n_210), .Y(n_706) );
INVx1_ASAP7_75t_L g694 ( .A(n_216), .Y(n_694) );
AOI22x1_ASAP7_75t_L g697 ( .A1(n_216), .A2(n_694), .B1(n_698), .B2(n_720), .Y(n_697) );
CKINVDCx20_ASAP7_75t_R g554 ( .A(n_218), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_220), .B(n_454), .Y(n_597) );
CKINVDCx20_ASAP7_75t_R g223 ( .A(n_224), .Y(n_223) );
CKINVDCx20_ASAP7_75t_R g224 ( .A(n_225), .Y(n_224) );
HB1xp67_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
AND2x4_ASAP7_75t_L g226 ( .A(n_227), .B(n_229), .Y(n_226) );
HB1xp67_ASAP7_75t_L g646 ( .A(n_228), .Y(n_646) );
OAI21xp5_ASAP7_75t_L g692 ( .A1(n_229), .A2(n_645), .B(n_693), .Y(n_692) );
AND2x2_ASAP7_75t_L g229 ( .A(n_230), .B(n_231), .Y(n_229) );
AOI221xp5_ASAP7_75t_L g232 ( .A1(n_233), .A2(n_548), .B1(n_640), .B2(n_641), .C(n_642), .Y(n_232) );
INVx1_ASAP7_75t_L g640 ( .A(n_233), .Y(n_640) );
AOI22xp5_ASAP7_75t_SL g233 ( .A1(n_234), .A2(n_235), .B1(n_499), .B2(n_500), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
XNOR2xp5_ASAP7_75t_SL g235 ( .A(n_236), .B(n_413), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
AOI22xp5_ASAP7_75t_L g237 ( .A1(n_238), .A2(n_239), .B1(n_335), .B2(n_336), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
INVx1_ASAP7_75t_L g334 ( .A(n_240), .Y(n_334) );
AND2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_296), .Y(n_240) );
NOR3xp33_ASAP7_75t_L g241 ( .A(n_242), .B(n_264), .C(n_285), .Y(n_241) );
OAI22xp5_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_244), .B1(n_259), .B2(n_260), .Y(n_242) );
BUFx6f_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
BUFx3_ASAP7_75t_L g684 ( .A(n_245), .Y(n_684) );
INVx2_ASAP7_75t_L g703 ( .A(n_245), .Y(n_703) );
OR2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_254), .Y(n_245) );
INVx2_ASAP7_75t_L g313 ( .A(n_246), .Y(n_313) );
OR2x2_ASAP7_75t_L g246 ( .A(n_247), .B(n_252), .Y(n_246) );
AND2x2_ASAP7_75t_L g263 ( .A(n_247), .B(n_252), .Y(n_263) );
AND2x2_ASAP7_75t_L g303 ( .A(n_247), .B(n_278), .Y(n_303) );
INVx2_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g268 ( .A(n_248), .B(n_252), .Y(n_268) );
AND2x2_ASAP7_75t_L g279 ( .A(n_248), .B(n_258), .Y(n_279) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
INVx1_ASAP7_75t_L g253 ( .A(n_251), .Y(n_253) );
INVx2_ASAP7_75t_L g278 ( .A(n_252), .Y(n_278) );
INVx1_ASAP7_75t_L g332 ( .A(n_252), .Y(n_332) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
NAND2x1p5_ASAP7_75t_L g262 ( .A(n_255), .B(n_263), .Y(n_262) );
AND2x4_ASAP7_75t_L g323 ( .A(n_255), .B(n_303), .Y(n_323) );
AND2x6_ASAP7_75t_L g353 ( .A(n_255), .B(n_263), .Y(n_353) );
AND2x4_ASAP7_75t_L g357 ( .A(n_255), .B(n_313), .Y(n_357) );
AND2x2_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .Y(n_255) );
INVx1_ASAP7_75t_L g270 ( .A(n_256), .Y(n_270) );
INVx1_ASAP7_75t_L g277 ( .A(n_256), .Y(n_277) );
INVx1_ASAP7_75t_L g295 ( .A(n_256), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_256), .B(n_258), .Y(n_308) );
AND2x2_ASAP7_75t_L g269 ( .A(n_257), .B(n_270), .Y(n_269) );
INVx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g302 ( .A(n_258), .B(n_295), .Y(n_302) );
INVx1_ASAP7_75t_SL g260 ( .A(n_261), .Y(n_260) );
INVx1_ASAP7_75t_L g686 ( .A(n_261), .Y(n_686) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
BUFx3_ASAP7_75t_L g485 ( .A(n_262), .Y(n_485) );
AND2x4_ASAP7_75t_L g316 ( .A(n_263), .B(n_269), .Y(n_316) );
AND2x2_ASAP7_75t_L g328 ( .A(n_263), .B(n_302), .Y(n_328) );
NAND2xp5_ASAP7_75t_SL g560 ( .A(n_263), .B(n_302), .Y(n_560) );
OAI221xp5_ASAP7_75t_L g264 ( .A1(n_265), .A2(n_271), .B1(n_272), .B2(n_280), .C(n_281), .Y(n_264) );
OAI21xp5_ASAP7_75t_SL g592 ( .A1(n_265), .A2(n_593), .B(n_594), .Y(n_592) );
OAI221xp5_ASAP7_75t_SL g705 ( .A1(n_265), .A2(n_524), .B1(n_706), .B2(n_707), .C(n_708), .Y(n_705) );
INVx2_ASAP7_75t_SL g265 ( .A(n_266), .Y(n_265) );
BUFx6f_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVx4_ASAP7_75t_L g343 ( .A(n_267), .Y(n_343) );
BUFx3_ASAP7_75t_L g385 ( .A(n_267), .Y(n_385) );
INVx2_ASAP7_75t_SL g444 ( .A(n_267), .Y(n_444) );
AND2x6_ASAP7_75t_L g267 ( .A(n_268), .B(n_269), .Y(n_267) );
INVx1_ASAP7_75t_L g292 ( .A(n_268), .Y(n_292) );
AND2x4_ASAP7_75t_L g363 ( .A(n_268), .B(n_294), .Y(n_363) );
AND2x6_ASAP7_75t_L g312 ( .A(n_269), .B(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g321 ( .A(n_269), .B(n_303), .Y(n_321) );
INVx2_ASAP7_75t_SL g272 ( .A(n_273), .Y(n_272) );
BUFx6f_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
BUFx6f_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
BUFx6f_ASAP7_75t_L g348 ( .A(n_275), .Y(n_348) );
BUFx4f_ASAP7_75t_SL g388 ( .A(n_275), .Y(n_388) );
BUFx6f_ASAP7_75t_L g458 ( .A(n_275), .Y(n_458) );
AND2x4_ASAP7_75t_L g275 ( .A(n_276), .B(n_279), .Y(n_275) );
AND2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
INVx1_ASAP7_75t_L g284 ( .A(n_277), .Y(n_284) );
INVx1_ASAP7_75t_L g288 ( .A(n_278), .Y(n_288) );
AND2x4_ASAP7_75t_L g283 ( .A(n_279), .B(n_284), .Y(n_283) );
NAND2x1p5_ASAP7_75t_L g287 ( .A(n_279), .B(n_288), .Y(n_287) );
AND2x4_ASAP7_75t_L g360 ( .A(n_279), .B(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g526 ( .A(n_282), .Y(n_526) );
BUFx6f_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
BUFx12f_ASAP7_75t_L g389 ( .A(n_283), .Y(n_389) );
BUFx6f_ASAP7_75t_L g447 ( .A(n_283), .Y(n_447) );
OAI22xp5_ASAP7_75t_L g285 ( .A1(n_286), .A2(n_287), .B1(n_289), .B2(n_290), .Y(n_285) );
BUFx3_ASAP7_75t_L g579 ( .A(n_287), .Y(n_579) );
INVx4_ASAP7_75t_L g675 ( .A(n_287), .Y(n_675) );
AND2x2_ASAP7_75t_L g403 ( .A(n_288), .B(n_307), .Y(n_403) );
OAI22xp5_ASAP7_75t_L g577 ( .A1(n_290), .A2(n_578), .B1(n_579), .B2(n_580), .Y(n_577) );
OAI22xp5_ASAP7_75t_L g709 ( .A1(n_290), .A2(n_579), .B1(n_710), .B2(n_711), .Y(n_709) );
BUFx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
OAI22xp5_ASAP7_75t_L g672 ( .A1(n_291), .A2(n_673), .B1(n_674), .B2(n_676), .Y(n_672) );
OR2x6_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
NOR2xp33_ASAP7_75t_L g296 ( .A(n_297), .B(n_317), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_298), .B(n_309), .Y(n_297) );
BUFx3_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
BUFx3_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
BUFx3_ASAP7_75t_L g376 ( .A(n_301), .Y(n_376) );
BUFx3_ASAP7_75t_L g399 ( .A(n_301), .Y(n_399) );
BUFx3_ASAP7_75t_L g463 ( .A(n_301), .Y(n_463) );
AND2x2_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_302), .B(n_303), .Y(n_572) );
AND2x4_ASAP7_75t_L g306 ( .A(n_303), .B(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g574 ( .A(n_304), .Y(n_574) );
BUFx2_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
BUFx3_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
BUFx2_ASAP7_75t_SL g379 ( .A(n_306), .Y(n_379) );
BUFx2_ASAP7_75t_L g400 ( .A(n_306), .Y(n_400) );
INVx1_ASAP7_75t_L g429 ( .A(n_306), .Y(n_429) );
BUFx3_ASAP7_75t_L g466 ( .A(n_306), .Y(n_466) );
BUFx3_ASAP7_75t_L g478 ( .A(n_306), .Y(n_478) );
BUFx3_ASAP7_75t_L g512 ( .A(n_306), .Y(n_512) );
BUFx2_ASAP7_75t_SL g607 ( .A(n_306), .Y(n_607) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
OR2x6_ASAP7_75t_L g331 ( .A(n_308), .B(n_332), .Y(n_331) );
INVx4_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx2_ASAP7_75t_SL g368 ( .A(n_311), .Y(n_368) );
INVx11_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx11_ASAP7_75t_L g407 ( .A(n_312), .Y(n_407) );
INVx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx2_ASAP7_75t_L g378 ( .A(n_315), .Y(n_378) );
INVx3_ASAP7_75t_L g408 ( .A(n_315), .Y(n_408) );
INVx6_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
BUFx3_ASAP7_75t_L g432 ( .A(n_316), .Y(n_432) );
BUFx3_ASAP7_75t_L g493 ( .A(n_316), .Y(n_493) );
BUFx3_ASAP7_75t_L g505 ( .A(n_316), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_318), .B(n_324), .Y(n_317) );
BUFx3_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
BUFx6f_ASAP7_75t_L g373 ( .A(n_320), .Y(n_373) );
BUFx3_ASAP7_75t_L g543 ( .A(n_320), .Y(n_543) );
BUFx6f_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx2_ASAP7_75t_L g411 ( .A(n_321), .Y(n_411) );
BUFx2_ASAP7_75t_SL g490 ( .A(n_321), .Y(n_490) );
BUFx2_ASAP7_75t_SL g616 ( .A(n_321), .Y(n_616) );
INVx1_ASAP7_75t_L g545 ( .A(n_322), .Y(n_545) );
BUFx3_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
BUFx6f_ASAP7_75t_L g369 ( .A(n_323), .Y(n_369) );
INVx2_ASAP7_75t_L g427 ( .A(n_323), .Y(n_427) );
BUFx3_ASAP7_75t_L g472 ( .A(n_323), .Y(n_472) );
BUFx3_ASAP7_75t_L g491 ( .A(n_323), .Y(n_491) );
BUFx2_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
BUFx6f_ASAP7_75t_L g604 ( .A(n_326), .Y(n_604) );
INVx5_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx2_ASAP7_75t_L g402 ( .A(n_327), .Y(n_402) );
BUFx3_ASAP7_75t_L g470 ( .A(n_327), .Y(n_470) );
INVx3_ASAP7_75t_L g480 ( .A(n_327), .Y(n_480) );
INVx1_ASAP7_75t_L g537 ( .A(n_327), .Y(n_537) );
INVx8_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
BUFx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
BUFx2_ASAP7_75t_L g473 ( .A(n_330), .Y(n_473) );
BUFx2_ASAP7_75t_L g481 ( .A(n_330), .Y(n_481) );
BUFx2_ASAP7_75t_L g538 ( .A(n_330), .Y(n_538) );
BUFx4f_ASAP7_75t_SL g719 ( .A(n_330), .Y(n_719) );
INVx6_ASAP7_75t_SL g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g663 ( .A(n_331), .Y(n_663) );
INVx1_ASAP7_75t_L g361 ( .A(n_332), .Y(n_361) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
XNOR2xp5_ASAP7_75t_L g336 ( .A(n_337), .B(n_380), .Y(n_336) );
NAND3x2_ASAP7_75t_L g338 ( .A(n_339), .B(n_364), .C(n_371), .Y(n_338) );
NOR2x1_ASAP7_75t_SL g339 ( .A(n_340), .B(n_349), .Y(n_339) );
OAI21xp5_ASAP7_75t_SL g340 ( .A1(n_341), .A2(n_344), .B(n_345), .Y(n_340) );
OAI222xp33_ASAP7_75t_L g522 ( .A1(n_341), .A2(n_523), .B1(n_524), .B2(n_525), .C1(n_526), .C2(n_527), .Y(n_522) );
INVx2_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx4_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
BUFx2_ASAP7_75t_L g583 ( .A(n_343), .Y(n_583) );
OAI221xp5_ASAP7_75t_L g677 ( .A1(n_343), .A2(n_678), .B1(n_679), .B2(n_680), .C(n_681), .Y(n_677) );
INVx3_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx4_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
NAND3xp33_ASAP7_75t_L g349 ( .A(n_350), .B(n_354), .C(n_358), .Y(n_349) );
INVx1_ASAP7_75t_SL g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_SL g352 ( .A(n_353), .Y(n_352) );
BUFx4f_ASAP7_75t_L g392 ( .A(n_353), .Y(n_392) );
BUFx2_ASAP7_75t_L g456 ( .A(n_353), .Y(n_456) );
BUFx2_ASAP7_75t_L g532 ( .A(n_353), .Y(n_532) );
INVx2_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx2_ASAP7_75t_L g394 ( .A(n_356), .Y(n_394) );
INVx2_ASAP7_75t_L g420 ( .A(n_356), .Y(n_420) );
INVx5_ASAP7_75t_L g454 ( .A(n_356), .Y(n_454) );
INVx4_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
BUFx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
BUFx3_ASAP7_75t_L g422 ( .A(n_360), .Y(n_422) );
BUFx2_ASAP7_75t_L g530 ( .A(n_360), .Y(n_530) );
INVx1_ASAP7_75t_L g600 ( .A(n_360), .Y(n_600) );
BUFx2_ASAP7_75t_SL g362 ( .A(n_363), .Y(n_362) );
BUFx2_ASAP7_75t_SL g437 ( .A(n_363), .Y(n_437) );
BUFx6f_ASAP7_75t_L g450 ( .A(n_363), .Y(n_450) );
BUFx3_ASAP7_75t_L g515 ( .A(n_363), .Y(n_515) );
AND2x2_ASAP7_75t_L g364 ( .A(n_365), .B(n_370), .Y(n_364) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx4_ASAP7_75t_L g618 ( .A(n_369), .Y(n_618) );
AND2x2_ASAP7_75t_L g371 ( .A(n_372), .B(n_377), .Y(n_371) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
XOR2x2_ASAP7_75t_L g380 ( .A(n_381), .B(n_412), .Y(n_380) );
NAND2xp5_ASAP7_75t_SL g381 ( .A(n_382), .B(n_396), .Y(n_381) );
NOR2xp33_ASAP7_75t_L g382 ( .A(n_383), .B(n_390), .Y(n_382) );
OAI21xp5_ASAP7_75t_SL g383 ( .A1(n_384), .A2(n_386), .B(n_387), .Y(n_383) );
INVx3_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g524 ( .A(n_388), .Y(n_524) );
INVx2_ASAP7_75t_L g436 ( .A(n_389), .Y(n_436) );
NAND3xp33_ASAP7_75t_L g390 ( .A(n_391), .B(n_393), .C(n_395), .Y(n_390) );
BUFx2_ASAP7_75t_L g623 ( .A(n_394), .Y(n_623) );
NOR2xp33_ASAP7_75t_L g396 ( .A(n_397), .B(n_404), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_398), .B(n_401), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_405), .B(n_409), .Y(n_404) );
INVx4_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx3_ASAP7_75t_L g541 ( .A(n_407), .Y(n_541) );
OAI22xp5_ASAP7_75t_L g564 ( .A1(n_407), .A2(n_565), .B1(n_566), .B2(n_567), .Y(n_564) );
INVx2_ASAP7_75t_SL g609 ( .A(n_407), .Y(n_609) );
INVx1_ASAP7_75t_L g635 ( .A(n_408), .Y(n_635) );
INVx3_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx3_ASAP7_75t_L g465 ( .A(n_411), .Y(n_465) );
OAI22xp5_ASAP7_75t_L g552 ( .A1(n_411), .A2(n_553), .B1(n_554), .B2(n_555), .Y(n_552) );
AOI22xp5_ASAP7_75t_L g413 ( .A1(n_414), .A2(n_415), .B1(n_438), .B2(n_498), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
NAND4xp75_ASAP7_75t_L g417 ( .A(n_418), .B(n_423), .C(n_430), .D(n_434), .Y(n_417) );
AND2x2_ASAP7_75t_SL g418 ( .A(n_419), .B(n_421), .Y(n_418) );
AND2x2_ASAP7_75t_L g423 ( .A(n_424), .B(n_425), .Y(n_423) );
INVx2_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
AND2x2_ASAP7_75t_L g430 ( .A(n_431), .B(n_433), .Y(n_430) );
INVx3_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g498 ( .A(n_438), .Y(n_498) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
AO22x2_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_474), .B1(n_496), .B2(n_497), .Y(n_439) );
INVx2_ASAP7_75t_L g496 ( .A(n_440), .Y(n_496) );
NAND2xp5_ASAP7_75t_SL g441 ( .A(n_442), .B(n_459), .Y(n_441) );
NOR2xp33_ASAP7_75t_SL g442 ( .A(n_443), .B(n_451), .Y(n_442) );
OAI21xp5_ASAP7_75t_SL g443 ( .A1(n_444), .A2(n_445), .B(n_446), .Y(n_443) );
BUFx3_ASAP7_75t_L g584 ( .A(n_447), .Y(n_584) );
INVx2_ASAP7_75t_L g679 ( .A(n_447), .Y(n_679) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_SL g449 ( .A(n_450), .Y(n_449) );
NAND3xp33_ASAP7_75t_L g451 ( .A(n_452), .B(n_455), .C(n_457), .Y(n_451) );
HB1xp67_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
BUFx6f_ASAP7_75t_L g576 ( .A(n_454), .Y(n_576) );
NOR2x1_ASAP7_75t_L g459 ( .A(n_460), .B(n_467), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_461), .B(n_464), .Y(n_460) );
BUFx4f_ASAP7_75t_SL g462 ( .A(n_463), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_468), .B(n_471), .Y(n_467) );
INVx3_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx3_ASAP7_75t_SL g497 ( .A(n_474), .Y(n_497) );
XOR2x2_ASAP7_75t_L g474 ( .A(n_475), .B(n_495), .Y(n_474) );
NAND4xp75_ASAP7_75t_L g475 ( .A(n_476), .B(n_482), .C(n_488), .D(n_494), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_477), .B(n_479), .Y(n_476) );
INVxp67_ASAP7_75t_L g629 ( .A(n_478), .Y(n_629) );
OA211x2_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_484), .B(n_486), .C(n_487), .Y(n_482) );
OA211x2_ASAP7_75t_L g620 ( .A1(n_484), .A2(n_621), .B(n_622), .C(n_624), .Y(n_620) );
BUFx3_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
AND2x2_ASAP7_75t_L g488 ( .A(n_489), .B(n_492), .Y(n_488) );
BUFx2_ASAP7_75t_L g556 ( .A(n_491), .Y(n_556) );
INVx1_ASAP7_75t_L g567 ( .A(n_493), .Y(n_567) );
CKINVDCx16_ASAP7_75t_R g499 ( .A(n_500), .Y(n_499) );
AOI22xp5_ASAP7_75t_L g500 ( .A1(n_501), .A2(n_517), .B1(n_518), .B2(n_547), .Y(n_500) );
INVx2_ASAP7_75t_SL g547 ( .A(n_501), .Y(n_547) );
XOR2x2_ASAP7_75t_L g501 ( .A(n_502), .B(n_516), .Y(n_501) );
NAND4xp75_ASAP7_75t_L g502 ( .A(n_503), .B(n_507), .C(n_510), .D(n_514), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_504), .B(n_506), .Y(n_503) );
AND2x2_ASAP7_75t_SL g507 ( .A(n_508), .B(n_509), .Y(n_507) );
AND2x2_ASAP7_75t_L g510 ( .A(n_511), .B(n_513), .Y(n_510) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx2_ASAP7_75t_L g546 ( .A(n_520), .Y(n_546) );
NAND3x1_ASAP7_75t_L g520 ( .A(n_521), .B(n_533), .C(n_539), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_522), .B(n_528), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_529), .B(n_531), .Y(n_528) );
AND2x2_ASAP7_75t_L g533 ( .A(n_534), .B(n_535), .Y(n_533) );
HB1xp67_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVxp67_ASAP7_75t_L g562 ( .A(n_538), .Y(n_562) );
AND2x2_ASAP7_75t_L g539 ( .A(n_540), .B(n_542), .Y(n_539) );
INVx1_ASAP7_75t_L g633 ( .A(n_541), .Y(n_633) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g641 ( .A(n_548), .Y(n_641) );
AOI22xp5_ASAP7_75t_L g548 ( .A1(n_549), .A2(n_587), .B1(n_588), .B2(n_639), .Y(n_548) );
INVx1_ASAP7_75t_L g639 ( .A(n_549), .Y(n_639) );
INVx1_ASAP7_75t_L g586 ( .A(n_550), .Y(n_586) );
AND4x1_ASAP7_75t_L g550 ( .A(n_551), .B(n_563), .C(n_575), .D(n_581), .Y(n_550) );
NOR2xp33_ASAP7_75t_SL g551 ( .A(n_552), .B(n_557), .Y(n_551) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
OAI22xp5_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_559), .B1(n_561), .B2(n_562), .Y(n_557) );
BUFx2_ASAP7_75t_R g559 ( .A(n_560), .Y(n_559) );
NOR2xp33_ASAP7_75t_SL g563 ( .A(n_564), .B(n_568), .Y(n_563) );
OAI22xp5_ASAP7_75t_L g568 ( .A1(n_569), .A2(n_570), .B1(n_573), .B2(n_574), .Y(n_568) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g628 ( .A(n_571), .Y(n_628) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
OAI22xp5_ASAP7_75t_SL g588 ( .A1(n_589), .A2(n_610), .B1(n_611), .B2(n_638), .Y(n_588) );
INVx1_ASAP7_75t_L g638 ( .A(n_589), .Y(n_638) );
NAND3xp33_ASAP7_75t_L g590 ( .A(n_591), .B(n_601), .C(n_605), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g591 ( .A(n_592), .B(n_595), .Y(n_591) );
NAND3xp33_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .C(n_598), .Y(n_595) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .Y(n_601) );
AND2x2_ASAP7_75t_L g605 ( .A(n_606), .B(n_608), .Y(n_605) );
INVx1_ASAP7_75t_SL g670 ( .A(n_607), .Y(n_670) );
INVx1_ASAP7_75t_SL g610 ( .A(n_611), .Y(n_610) );
INVx2_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
XOR2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_637), .Y(n_612) );
NAND4xp75_ASAP7_75t_L g613 ( .A(n_614), .B(n_620), .C(n_625), .D(n_636), .Y(n_613) );
AND2x2_ASAP7_75t_L g614 ( .A(n_615), .B(n_619), .Y(n_614) );
INVx3_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
OAI22xp5_ASAP7_75t_L g667 ( .A1(n_618), .A2(n_668), .B1(n_669), .B2(n_670), .Y(n_667) );
NOR2xp33_ASAP7_75t_L g625 ( .A(n_626), .B(n_631), .Y(n_625) );
OAI22xp5_ASAP7_75t_L g626 ( .A1(n_627), .A2(n_628), .B1(n_629), .B2(n_630), .Y(n_626) );
OAI22xp5_ASAP7_75t_L g664 ( .A1(n_628), .A2(n_635), .B1(n_665), .B2(n_666), .Y(n_664) );
OAI22xp5_ASAP7_75t_L g631 ( .A1(n_632), .A2(n_633), .B1(n_634), .B2(n_635), .Y(n_631) );
INVx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
NOR2x1_ASAP7_75t_L g643 ( .A(n_644), .B(n_648), .Y(n_643) );
OR2x2_ASAP7_75t_SL g723 ( .A(n_644), .B(n_649), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_645), .B(n_647), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
HB1xp67_ASAP7_75t_L g687 ( .A(n_646), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_646), .B(n_690), .Y(n_693) );
CKINVDCx16_ASAP7_75t_R g690 ( .A(n_647), .Y(n_690) );
CKINVDCx20_ASAP7_75t_R g648 ( .A(n_649), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_650), .B(n_651), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_653), .B(n_654), .Y(n_652) );
OAI322xp33_ASAP7_75t_L g655 ( .A1(n_656), .A2(n_687), .A3(n_688), .B1(n_691), .B2(n_694), .C1(n_695), .C2(n_721), .Y(n_655) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
AND2x2_ASAP7_75t_L g658 ( .A(n_659), .B(n_671), .Y(n_658) );
NOR3xp33_ASAP7_75t_L g659 ( .A(n_660), .B(n_664), .C(n_667), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_661), .B(n_662), .Y(n_660) );
NOR3xp33_ASAP7_75t_L g671 ( .A(n_672), .B(n_677), .C(n_682), .Y(n_671) );
INVx3_ASAP7_75t_SL g674 ( .A(n_675), .Y(n_674) );
OAI22xp5_ASAP7_75t_L g682 ( .A1(n_683), .A2(n_684), .B1(n_685), .B2(n_686), .Y(n_682) );
OAI22xp5_ASAP7_75t_L g700 ( .A1(n_686), .A2(n_701), .B1(n_702), .B2(n_704), .Y(n_700) );
HB1xp67_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
CKINVDCx20_ASAP7_75t_R g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx2_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx2_ASAP7_75t_SL g720 ( .A(n_698), .Y(n_720) );
AND2x2_ASAP7_75t_L g698 ( .A(n_699), .B(n_712), .Y(n_698) );
NOR3xp33_ASAP7_75t_L g699 ( .A(n_700), .B(n_705), .C(n_709), .Y(n_699) );
INVx2_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
NOR2xp33_ASAP7_75t_L g712 ( .A(n_713), .B(n_716), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_714), .B(n_715), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_717), .B(n_718), .Y(n_716) );
CKINVDCx20_ASAP7_75t_R g721 ( .A(n_722), .Y(n_721) );
CKINVDCx20_ASAP7_75t_R g722 ( .A(n_723), .Y(n_722) );
endmodule