module fake_netlist_6_2299_n_1731 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1731);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1731;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_701;
wire n_295;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1373;
wire n_1292;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_8),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_62),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_80),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_133),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_66),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_24),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_41),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_115),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_2),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_105),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_27),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_147),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_96),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_108),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_100),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_17),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_151),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_94),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_111),
.Y(n_173)
);

INVx2_ASAP7_75t_SL g174 ( 
.A(n_73),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_50),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_114),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_95),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_77),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_124),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_20),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_118),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_137),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_28),
.Y(n_183)
);

BUFx8_ASAP7_75t_SL g184 ( 
.A(n_54),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_72),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_13),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_101),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_79),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_36),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_13),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_42),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_12),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_84),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_87),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_3),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_9),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_55),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_93),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_78),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_117),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_122),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_30),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_6),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_17),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_20),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_37),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_126),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_71),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_145),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_40),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_63),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_35),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_132),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_16),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_68),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_113),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_120),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_107),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_50),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_55),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_24),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_18),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_148),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_37),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_82),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_144),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_67),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_47),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_59),
.Y(n_229)
);

BUFx10_ASAP7_75t_L g230 ( 
.A(n_57),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_5),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_146),
.Y(n_232)
);

BUFx2_ASAP7_75t_L g233 ( 
.A(n_23),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_47),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_49),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_112),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_154),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_56),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_31),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_106),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_41),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_29),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_44),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_83),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_38),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_65),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_74),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_29),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_7),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_44),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_31),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_152),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_5),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_8),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_28),
.Y(n_255)
);

BUFx10_ASAP7_75t_L g256 ( 
.A(n_60),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_102),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_0),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_35),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_89),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_48),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_92),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_30),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_116),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_136),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_138),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_121),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_103),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_0),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_129),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_21),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_27),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_42),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_58),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_56),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_15),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_85),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_32),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_64),
.Y(n_279)
);

INVx1_ASAP7_75t_SL g280 ( 
.A(n_109),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_49),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_10),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_25),
.Y(n_283)
);

BUFx10_ASAP7_75t_L g284 ( 
.A(n_134),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_149),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_38),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_125),
.Y(n_287)
);

INVxp67_ASAP7_75t_SL g288 ( 
.A(n_104),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_139),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_86),
.Y(n_290)
);

INVx1_ASAP7_75t_SL g291 ( 
.A(n_39),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_127),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_88),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_153),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_15),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_4),
.Y(n_296)
);

CKINVDCx14_ASAP7_75t_R g297 ( 
.A(n_97),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_48),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_16),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_14),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_46),
.Y(n_301)
);

BUFx5_ASAP7_75t_L g302 ( 
.A(n_22),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_130),
.Y(n_303)
);

BUFx10_ASAP7_75t_L g304 ( 
.A(n_19),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_12),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_33),
.Y(n_306)
);

BUFx3_ASAP7_75t_L g307 ( 
.A(n_36),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_150),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_14),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_184),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_156),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_302),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_157),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_166),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_287),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_198),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_158),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_182),
.B(n_1),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_302),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_302),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_159),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_287),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_297),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_302),
.Y(n_324)
);

INVxp67_ASAP7_75t_SL g325 ( 
.A(n_200),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_162),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_164),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_233),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_211),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_167),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_168),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_302),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_244),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_173),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_302),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_302),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_302),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_265),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_302),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_176),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_270),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_196),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_196),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_178),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_228),
.Y(n_345)
);

HB1xp67_ASAP7_75t_L g346 ( 
.A(n_233),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_228),
.Y(n_347)
);

INVxp67_ASAP7_75t_SL g348 ( 
.A(n_200),
.Y(n_348)
);

INVxp67_ASAP7_75t_SL g349 ( 
.A(n_273),
.Y(n_349)
);

INVx3_ASAP7_75t_L g350 ( 
.A(n_169),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_179),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_235),
.Y(n_352)
);

NOR2xp67_ASAP7_75t_L g353 ( 
.A(n_235),
.B(n_1),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_186),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_174),
.B(n_2),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_181),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_186),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_185),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_188),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_171),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_190),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_190),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_193),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_203),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_174),
.B(n_3),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_169),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_203),
.Y(n_367)
);

INVxp33_ASAP7_75t_L g368 ( 
.A(n_204),
.Y(n_368)
);

CKINVDCx16_ASAP7_75t_R g369 ( 
.A(n_230),
.Y(n_369)
);

BUFx2_ASAP7_75t_L g370 ( 
.A(n_273),
.Y(n_370)
);

CKINVDCx16_ASAP7_75t_R g371 ( 
.A(n_230),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_204),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_194),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_199),
.Y(n_374)
);

INVxp67_ASAP7_75t_SL g375 ( 
.A(n_307),
.Y(n_375)
);

BUFx2_ASAP7_75t_L g376 ( 
.A(n_307),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_205),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_201),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_207),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_208),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_205),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_213),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_206),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_215),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_217),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_366),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_312),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_366),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_312),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_319),
.B(n_267),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_319),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_320),
.B(n_267),
.Y(n_392)
);

OA21x2_ASAP7_75t_L g393 ( 
.A1(n_360),
.A2(n_221),
.B(n_206),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_320),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_324),
.Y(n_395)
);

AND2x4_ASAP7_75t_L g396 ( 
.A(n_350),
.B(n_171),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_355),
.B(n_280),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_366),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_324),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_350),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_325),
.B(n_348),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_332),
.B(n_172),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_332),
.Y(n_403)
);

HB1xp67_ASAP7_75t_L g404 ( 
.A(n_370),
.Y(n_404)
);

AND2x4_ASAP7_75t_L g405 ( 
.A(n_350),
.B(n_172),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_335),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_335),
.Y(n_407)
);

INVx4_ASAP7_75t_L g408 ( 
.A(n_350),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_336),
.Y(n_409)
);

INVx3_ASAP7_75t_L g410 ( 
.A(n_336),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_337),
.B(n_177),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_337),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_339),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_339),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_365),
.B(n_177),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_360),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_342),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_342),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_343),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_343),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_349),
.B(n_375),
.Y(n_421)
);

BUFx2_ASAP7_75t_L g422 ( 
.A(n_370),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_345),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_345),
.Y(n_424)
);

AND2x4_ASAP7_75t_L g425 ( 
.A(n_353),
.B(n_187),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_347),
.Y(n_426)
);

AND2x6_ASAP7_75t_L g427 ( 
.A(n_347),
.B(n_169),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_352),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_352),
.Y(n_429)
);

NAND2xp33_ASAP7_75t_SL g430 ( 
.A(n_368),
.B(n_191),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_354),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_376),
.B(n_187),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_354),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_357),
.Y(n_434)
);

CKINVDCx6p67_ASAP7_75t_R g435 ( 
.A(n_315),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_357),
.Y(n_436)
);

BUFx2_ASAP7_75t_L g437 ( 
.A(n_376),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_361),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_361),
.B(n_216),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_L g440 ( 
.A1(n_328),
.A2(n_255),
.B1(n_286),
.B2(n_160),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_362),
.Y(n_441)
);

AND2x4_ASAP7_75t_L g442 ( 
.A(n_353),
.B(n_216),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_362),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_364),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_364),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_367),
.B(n_218),
.Y(n_446)
);

INVx3_ASAP7_75t_L g447 ( 
.A(n_367),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_372),
.B(n_218),
.Y(n_448)
);

NAND2xp33_ASAP7_75t_R g449 ( 
.A(n_310),
.B(n_155),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_372),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_377),
.Y(n_451)
);

OA21x2_ASAP7_75t_L g452 ( 
.A1(n_377),
.A2(n_234),
.B(n_221),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_381),
.B(n_223),
.Y(n_453)
);

HB1xp67_ASAP7_75t_L g454 ( 
.A(n_346),
.Y(n_454)
);

OR2x2_ASAP7_75t_L g455 ( 
.A(n_422),
.B(n_315),
.Y(n_455)
);

NOR3xp33_ASAP7_75t_L g456 ( 
.A(n_440),
.B(n_322),
.C(n_318),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_409),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_397),
.B(n_311),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_397),
.B(n_313),
.Y(n_459)
);

INVxp67_ASAP7_75t_SL g460 ( 
.A(n_410),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_394),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_394),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_394),
.Y(n_463)
);

INVx1_ASAP7_75t_SL g464 ( 
.A(n_430),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_394),
.Y(n_465)
);

BUFx10_ASAP7_75t_L g466 ( 
.A(n_415),
.Y(n_466)
);

BUFx3_ASAP7_75t_L g467 ( 
.A(n_393),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_401),
.B(n_317),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_401),
.B(n_321),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_415),
.B(n_326),
.Y(n_470)
);

INVx4_ASAP7_75t_L g471 ( 
.A(n_389),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_393),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_394),
.Y(n_473)
);

NAND2xp33_ASAP7_75t_R g474 ( 
.A(n_422),
.B(n_327),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_449),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_421),
.B(n_322),
.Y(n_476)
);

INVx3_ASAP7_75t_L g477 ( 
.A(n_408),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_393),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_401),
.B(n_330),
.Y(n_479)
);

NOR3xp33_ASAP7_75t_L g480 ( 
.A(n_440),
.B(n_371),
.C(n_369),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_393),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_393),
.Y(n_482)
);

BUFx3_ASAP7_75t_L g483 ( 
.A(n_393),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_387),
.Y(n_484)
);

BUFx10_ASAP7_75t_L g485 ( 
.A(n_425),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_387),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_401),
.B(n_331),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_421),
.B(n_323),
.Y(n_488)
);

AND2x6_ASAP7_75t_L g489 ( 
.A(n_425),
.B(n_223),
.Y(n_489)
);

INVx1_ASAP7_75t_SL g490 ( 
.A(n_430),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_387),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_421),
.B(n_334),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_393),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_421),
.B(n_340),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_422),
.B(n_351),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_409),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_437),
.B(n_358),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_387),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_409),
.Y(n_499)
);

AOI22xp33_ASAP7_75t_L g500 ( 
.A1(n_425),
.A2(n_275),
.B1(n_271),
.B2(n_269),
.Y(n_500)
);

AND2x2_ASAP7_75t_SL g501 ( 
.A(n_425),
.B(n_225),
.Y(n_501)
);

INVx5_ASAP7_75t_L g502 ( 
.A(n_427),
.Y(n_502)
);

INVx1_ASAP7_75t_SL g503 ( 
.A(n_437),
.Y(n_503)
);

AND2x2_ASAP7_75t_SL g504 ( 
.A(n_425),
.B(n_225),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_449),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_439),
.B(n_381),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_412),
.B(n_413),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_403),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g509 ( 
.A(n_389),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_412),
.Y(n_510)
);

INVx2_ASAP7_75t_SL g511 ( 
.A(n_404),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_412),
.Y(n_512)
);

NOR2x1p5_ASAP7_75t_L g513 ( 
.A(n_435),
.B(n_161),
.Y(n_513)
);

AOI22xp33_ASAP7_75t_L g514 ( 
.A1(n_425),
.A2(n_243),
.B1(n_242),
.B2(n_239),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_437),
.B(n_363),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_439),
.B(n_383),
.Y(n_516)
);

NAND2xp33_ASAP7_75t_SL g517 ( 
.A(n_432),
.B(n_165),
.Y(n_517)
);

BUFx3_ASAP7_75t_L g518 ( 
.A(n_452),
.Y(n_518)
);

INVx4_ASAP7_75t_L g519 ( 
.A(n_389),
.Y(n_519)
);

INVxp67_ASAP7_75t_SL g520 ( 
.A(n_410),
.Y(n_520)
);

AOI22xp33_ASAP7_75t_L g521 ( 
.A1(n_425),
.A2(n_242),
.B1(n_243),
.B2(n_239),
.Y(n_521)
);

INVx4_ASAP7_75t_L g522 ( 
.A(n_389),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_403),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_413),
.Y(n_524)
);

INVx4_ASAP7_75t_L g525 ( 
.A(n_389),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_404),
.B(n_378),
.Y(n_526)
);

INVx5_ASAP7_75t_L g527 ( 
.A(n_427),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_439),
.B(n_383),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_403),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_413),
.Y(n_530)
);

BUFx2_ASAP7_75t_L g531 ( 
.A(n_454),
.Y(n_531)
);

OR2x6_ASAP7_75t_L g532 ( 
.A(n_432),
.B(n_163),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_414),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_414),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_432),
.A2(n_359),
.B1(n_344),
.B2(n_373),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_408),
.Y(n_536)
);

AOI22xp33_ASAP7_75t_SL g537 ( 
.A1(n_440),
.A2(n_369),
.B1(n_371),
.B2(n_341),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_414),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_403),
.Y(n_539)
);

NAND2xp33_ASAP7_75t_L g540 ( 
.A(n_402),
.B(n_169),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_408),
.B(n_379),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_407),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_432),
.B(n_323),
.Y(n_543)
);

INVxp33_ASAP7_75t_L g544 ( 
.A(n_454),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_410),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_408),
.B(n_380),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_407),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_408),
.B(n_382),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_407),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_407),
.Y(n_550)
);

AND2x6_ASAP7_75t_L g551 ( 
.A(n_442),
.B(n_227),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_410),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_439),
.B(n_384),
.Y(n_553)
);

AOI22xp33_ASAP7_75t_L g554 ( 
.A1(n_442),
.A2(n_446),
.B1(n_448),
.B2(n_452),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_408),
.B(n_385),
.Y(n_555)
);

AOI22xp5_ASAP7_75t_L g556 ( 
.A1(n_435),
.A2(n_356),
.B1(n_374),
.B2(n_442),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_408),
.B(n_226),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_410),
.Y(n_558)
);

CKINVDCx20_ASAP7_75t_R g559 ( 
.A(n_435),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_410),
.Y(n_560)
);

OR2x6_ASAP7_75t_L g561 ( 
.A(n_442),
.B(n_189),
.Y(n_561)
);

AOI22xp33_ASAP7_75t_L g562 ( 
.A1(n_442),
.A2(n_446),
.B1(n_448),
.B2(n_452),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_442),
.B(n_256),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_441),
.B(n_338),
.Y(n_564)
);

AO21x2_ASAP7_75t_L g565 ( 
.A1(n_402),
.A2(n_236),
.B(n_227),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g566 ( 
.A(n_446),
.B(n_236),
.Y(n_566)
);

OAI22xp33_ASAP7_75t_L g567 ( 
.A1(n_435),
.A2(n_214),
.B1(n_291),
.B2(n_306),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_442),
.B(n_256),
.Y(n_568)
);

AND2x6_ASAP7_75t_L g569 ( 
.A(n_446),
.B(n_262),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_448),
.B(n_262),
.Y(n_570)
);

OAI22xp33_ASAP7_75t_L g571 ( 
.A1(n_453),
.A2(n_276),
.B1(n_309),
.B2(n_231),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_389),
.B(n_229),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_SL g573 ( 
.A(n_448),
.B(n_314),
.Y(n_573)
);

OR2x2_ASAP7_75t_L g574 ( 
.A(n_452),
.B(n_170),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_396),
.B(n_256),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_396),
.B(n_256),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_452),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_389),
.B(n_232),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_441),
.B(n_316),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_396),
.B(n_284),
.Y(n_580)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_389),
.Y(n_581)
);

AND2x6_ASAP7_75t_L g582 ( 
.A(n_396),
.B(n_264),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_452),
.Y(n_583)
);

CKINVDCx20_ASAP7_75t_R g584 ( 
.A(n_452),
.Y(n_584)
);

INVx1_ASAP7_75t_SL g585 ( 
.A(n_453),
.Y(n_585)
);

AOI22xp33_ASAP7_75t_L g586 ( 
.A1(n_396),
.A2(n_234),
.B1(n_283),
.B2(n_296),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_441),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_443),
.Y(n_588)
);

BUFx6f_ASAP7_75t_L g589 ( 
.A(n_389),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_416),
.Y(n_590)
);

OAI22xp5_ASAP7_75t_L g591 ( 
.A1(n_402),
.A2(n_219),
.B1(n_305),
.B2(n_301),
.Y(n_591)
);

AOI22xp33_ASAP7_75t_L g592 ( 
.A1(n_396),
.A2(n_296),
.B1(n_283),
.B2(n_275),
.Y(n_592)
);

AOI22xp33_ASAP7_75t_L g593 ( 
.A1(n_396),
.A2(n_269),
.B1(n_271),
.B2(n_289),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_389),
.B(n_237),
.Y(n_594)
);

BUFx10_ASAP7_75t_L g595 ( 
.A(n_405),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_443),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_391),
.B(n_240),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_443),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_405),
.Y(n_599)
);

INVx2_ASAP7_75t_SL g600 ( 
.A(n_405),
.Y(n_600)
);

AND2x2_ASAP7_75t_SL g601 ( 
.A(n_405),
.B(n_264),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_416),
.Y(n_602)
);

BUFx3_ASAP7_75t_L g603 ( 
.A(n_405),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_391),
.B(n_246),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_467),
.Y(n_605)
);

NOR3xp33_ASAP7_75t_L g606 ( 
.A(n_459),
.B(n_453),
.C(n_288),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_585),
.B(n_447),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_467),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_599),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_483),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_470),
.B(n_329),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_468),
.B(n_411),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_479),
.B(n_447),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_492),
.B(n_447),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_501),
.B(n_447),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_466),
.B(n_333),
.Y(n_616)
);

AOI221xp5_ASAP7_75t_L g617 ( 
.A1(n_456),
.A2(n_249),
.B1(n_212),
.B2(n_210),
.C(n_222),
.Y(n_617)
);

INVxp67_ASAP7_75t_L g618 ( 
.A(n_495),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_501),
.B(n_447),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_504),
.B(n_447),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_469),
.B(n_411),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_466),
.B(n_247),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_487),
.B(n_411),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_504),
.B(n_391),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_494),
.B(n_175),
.Y(n_625)
);

INVx3_ASAP7_75t_L g626 ( 
.A(n_603),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_554),
.B(n_391),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_599),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_466),
.B(n_252),
.Y(n_629)
);

NAND2xp33_ASAP7_75t_L g630 ( 
.A(n_584),
.B(n_257),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_562),
.B(n_391),
.Y(n_631)
);

INVxp67_ASAP7_75t_L g632 ( 
.A(n_497),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_511),
.B(n_230),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_458),
.B(n_391),
.Y(n_634)
);

NOR2xp67_ASAP7_75t_SL g635 ( 
.A(n_477),
.B(n_169),
.Y(n_635)
);

AOI22xp5_ASAP7_75t_L g636 ( 
.A1(n_584),
.A2(n_405),
.B1(n_260),
.B2(n_308),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_603),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_476),
.B(n_180),
.Y(n_638)
);

BUFx6f_ASAP7_75t_L g639 ( 
.A(n_518),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_506),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_506),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_516),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_516),
.B(n_391),
.Y(n_643)
);

BUFx6f_ASAP7_75t_SL g644 ( 
.A(n_511),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_483),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_528),
.B(n_391),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_518),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_601),
.B(n_391),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_528),
.B(n_391),
.Y(n_649)
);

NAND3xp33_ASAP7_75t_L g650 ( 
.A(n_517),
.B(n_248),
.C(n_183),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_587),
.Y(n_651)
);

NOR3xp33_ASAP7_75t_L g652 ( 
.A(n_564),
.B(n_250),
.C(n_195),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_488),
.B(n_192),
.Y(n_653)
);

AOI22xp33_ASAP7_75t_L g654 ( 
.A1(n_577),
.A2(n_289),
.B1(n_293),
.B2(n_392),
.Y(n_654)
);

NAND2xp33_ASAP7_75t_L g655 ( 
.A(n_489),
.B(n_266),
.Y(n_655)
);

INVx3_ASAP7_75t_L g656 ( 
.A(n_595),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_596),
.Y(n_657)
);

OR2x6_ASAP7_75t_L g658 ( 
.A(n_531),
.B(n_455),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_553),
.B(n_197),
.Y(n_659)
);

BUFx2_ASAP7_75t_L g660 ( 
.A(n_531),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_596),
.Y(n_661)
);

INVx2_ASAP7_75t_SL g662 ( 
.A(n_455),
.Y(n_662)
);

BUFx6f_ASAP7_75t_L g663 ( 
.A(n_595),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_598),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_598),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_510),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_477),
.B(n_395),
.Y(n_667)
);

AOI22xp33_ASAP7_75t_L g668 ( 
.A1(n_577),
.A2(n_293),
.B1(n_392),
.B2(n_390),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_510),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_553),
.B(n_268),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_472),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_477),
.B(n_395),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_536),
.B(n_395),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_512),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_536),
.B(n_395),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_475),
.B(n_274),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_543),
.B(n_202),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_536),
.B(n_395),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_526),
.B(n_220),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_515),
.B(n_224),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_457),
.B(n_395),
.Y(n_681)
);

BUFx8_ASAP7_75t_L g682 ( 
.A(n_574),
.Y(n_682)
);

OAI221xp5_ASAP7_75t_L g683 ( 
.A1(n_500),
.A2(n_390),
.B1(n_392),
.B2(n_429),
.C(n_424),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_475),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_464),
.B(n_238),
.Y(n_685)
);

NAND2xp33_ASAP7_75t_L g686 ( 
.A(n_489),
.B(n_277),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_472),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_496),
.B(n_395),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_499),
.B(n_395),
.Y(n_689)
);

AOI22xp33_ASAP7_75t_L g690 ( 
.A1(n_583),
.A2(n_565),
.B1(n_478),
.B2(n_482),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_524),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_505),
.B(n_279),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_478),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_524),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_530),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_460),
.B(n_395),
.Y(n_696)
);

AOI22xp33_ASAP7_75t_L g697 ( 
.A1(n_583),
.A2(n_390),
.B1(n_405),
.B2(n_451),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_505),
.B(n_285),
.Y(n_698)
);

BUFx6f_ASAP7_75t_L g699 ( 
.A(n_595),
.Y(n_699)
);

INVxp67_ASAP7_75t_L g700 ( 
.A(n_474),
.Y(n_700)
);

INVxp67_ASAP7_75t_L g701 ( 
.A(n_579),
.Y(n_701)
);

NOR2xp67_ASAP7_75t_L g702 ( 
.A(n_535),
.B(n_417),
.Y(n_702)
);

O2A1O1Ixp5_ASAP7_75t_L g703 ( 
.A1(n_481),
.A2(n_400),
.B(n_434),
.C(n_445),
.Y(n_703)
);

INVx3_ASAP7_75t_L g704 ( 
.A(n_600),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_490),
.B(n_241),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_503),
.B(n_230),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_530),
.Y(n_707)
);

BUFx10_ASAP7_75t_L g708 ( 
.A(n_513),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_533),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_532),
.B(n_574),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_533),
.Y(n_711)
);

OAI21xp5_ASAP7_75t_L g712 ( 
.A1(n_481),
.A2(n_400),
.B(n_416),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_520),
.B(n_395),
.Y(n_713)
);

BUFx8_ASAP7_75t_L g714 ( 
.A(n_566),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_532),
.B(n_245),
.Y(n_715)
);

OAI22xp5_ASAP7_75t_L g716 ( 
.A1(n_601),
.A2(n_303),
.B1(n_294),
.B2(n_292),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_588),
.B(n_566),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_534),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_600),
.B(n_399),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_570),
.B(n_399),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_570),
.B(n_399),
.Y(n_721)
);

O2A1O1Ixp5_ASAP7_75t_L g722 ( 
.A1(n_482),
.A2(n_493),
.B(n_534),
.C(n_538),
.Y(n_722)
);

AND2x2_ASAP7_75t_SL g723 ( 
.A(n_480),
.B(n_209),
.Y(n_723)
);

AOI22xp5_ASAP7_75t_L g724 ( 
.A1(n_573),
.A2(n_290),
.B1(n_438),
.B2(n_445),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_493),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_538),
.B(n_399),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_545),
.B(n_399),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_545),
.B(n_399),
.Y(n_728)
);

BUFx6f_ASAP7_75t_SL g729 ( 
.A(n_532),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_590),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_552),
.B(n_558),
.Y(n_731)
);

NAND2xp33_ASAP7_75t_SL g732 ( 
.A(n_544),
.B(n_251),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_552),
.B(n_399),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_532),
.B(n_253),
.Y(n_734)
);

NOR3xp33_ASAP7_75t_L g735 ( 
.A(n_537),
.B(n_254),
.C(n_258),
.Y(n_735)
);

BUFx6f_ASAP7_75t_L g736 ( 
.A(n_485),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_558),
.B(n_399),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_485),
.B(n_399),
.Y(n_738)
);

AOI22xp33_ASAP7_75t_SL g739 ( 
.A1(n_559),
.A2(n_569),
.B1(n_591),
.B2(n_561),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_560),
.B(n_399),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_507),
.B(n_406),
.Y(n_741)
);

AOI22xp5_ASAP7_75t_L g742 ( 
.A1(n_561),
.A2(n_431),
.B1(n_433),
.B2(n_445),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_569),
.B(n_541),
.Y(n_743)
);

INVxp67_ASAP7_75t_L g744 ( 
.A(n_517),
.Y(n_744)
);

INVxp67_ASAP7_75t_L g745 ( 
.A(n_567),
.Y(n_745)
);

NAND2xp33_ASAP7_75t_L g746 ( 
.A(n_489),
.B(n_551),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_590),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_602),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_602),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_569),
.B(n_406),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_571),
.B(n_284),
.Y(n_751)
);

NOR2x1p5_ASAP7_75t_L g752 ( 
.A(n_559),
.B(n_259),
.Y(n_752)
);

AO22x2_ASAP7_75t_L g753 ( 
.A1(n_563),
.A2(n_429),
.B1(n_417),
.B2(n_419),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_569),
.B(n_406),
.Y(n_754)
);

OR2x2_ASAP7_75t_L g755 ( 
.A(n_561),
.B(n_261),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_485),
.B(n_284),
.Y(n_756)
);

INVxp67_ASAP7_75t_L g757 ( 
.A(n_556),
.Y(n_757)
);

NOR3xp33_ASAP7_75t_L g758 ( 
.A(n_568),
.B(n_263),
.C(n_272),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_569),
.B(n_406),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_514),
.B(n_284),
.Y(n_760)
);

NAND2x1_ASAP7_75t_L g761 ( 
.A(n_471),
.B(n_400),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_561),
.B(n_278),
.Y(n_762)
);

AOI22xp33_ASAP7_75t_L g763 ( 
.A1(n_565),
.A2(n_451),
.B1(n_431),
.B2(n_445),
.Y(n_763)
);

AOI22xp33_ASAP7_75t_L g764 ( 
.A1(n_565),
.A2(n_451),
.B1(n_431),
.B2(n_433),
.Y(n_764)
);

AOI22xp5_ASAP7_75t_L g765 ( 
.A1(n_569),
.A2(n_431),
.B1(n_438),
.B2(n_436),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_521),
.B(n_209),
.Y(n_766)
);

AOI22xp33_ASAP7_75t_L g767 ( 
.A1(n_489),
.A2(n_551),
.B1(n_582),
.B2(n_593),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_484),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_486),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_546),
.B(n_406),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_548),
.B(n_406),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_555),
.B(n_209),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_575),
.B(n_576),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_486),
.Y(n_774)
);

INVx2_ASAP7_75t_SL g775 ( 
.A(n_580),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_612),
.B(n_489),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_612),
.B(n_489),
.Y(n_777)
);

NOR2xp67_ASAP7_75t_L g778 ( 
.A(n_701),
.B(n_604),
.Y(n_778)
);

AOI21xp5_ASAP7_75t_L g779 ( 
.A1(n_712),
.A2(n_557),
.B(n_594),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_618),
.B(n_572),
.Y(n_780)
);

AOI33xp33_ASAP7_75t_L g781 ( 
.A1(n_662),
.A2(n_586),
.A3(n_592),
.B1(n_429),
.B2(n_428),
.B3(n_417),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_651),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_621),
.B(n_551),
.Y(n_783)
);

AOI22xp33_ASAP7_75t_L g784 ( 
.A1(n_654),
.A2(n_551),
.B1(n_582),
.B2(n_540),
.Y(n_784)
);

AOI21x1_ASAP7_75t_L g785 ( 
.A1(n_635),
.A2(n_597),
.B(n_578),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_621),
.B(n_551),
.Y(n_786)
);

OAI21xp5_ASAP7_75t_L g787 ( 
.A1(n_627),
.A2(n_631),
.B(n_722),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_632),
.B(n_471),
.Y(n_788)
);

A2O1A1Ixp33_ASAP7_75t_L g789 ( 
.A1(n_623),
.A2(n_540),
.B(n_581),
.C(n_550),
.Y(n_789)
);

BUFx12f_ASAP7_75t_L g790 ( 
.A(n_708),
.Y(n_790)
);

BUFx2_ASAP7_75t_L g791 ( 
.A(n_658),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_607),
.B(n_581),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_625),
.B(n_581),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_625),
.B(n_491),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_613),
.B(n_491),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_651),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_614),
.B(n_498),
.Y(n_797)
);

BUFx6f_ASAP7_75t_L g798 ( 
.A(n_639),
.Y(n_798)
);

AOI21xp5_ASAP7_75t_L g799 ( 
.A1(n_743),
.A2(n_471),
.B(n_519),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_661),
.Y(n_800)
);

AOI21xp5_ASAP7_75t_L g801 ( 
.A1(n_667),
.A2(n_519),
.B(n_522),
.Y(n_801)
);

INVx2_ASAP7_75t_SL g802 ( 
.A(n_660),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_680),
.B(n_498),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_639),
.B(n_509),
.Y(n_804)
);

AND2x4_ASAP7_75t_L g805 ( 
.A(n_640),
.B(n_582),
.Y(n_805)
);

INVx11_ASAP7_75t_L g806 ( 
.A(n_714),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_700),
.B(n_519),
.Y(n_807)
);

OAI21xp5_ASAP7_75t_L g808 ( 
.A1(n_703),
.A2(n_523),
.B(n_508),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_680),
.B(n_508),
.Y(n_809)
);

AOI21xp33_ASAP7_75t_L g810 ( 
.A1(n_679),
.A2(n_281),
.B(n_300),
.Y(n_810)
);

OAI21xp5_ASAP7_75t_L g811 ( 
.A1(n_615),
.A2(n_539),
.B(n_523),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_633),
.B(n_304),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_639),
.B(n_509),
.Y(n_813)
);

INVx3_ASAP7_75t_L g814 ( 
.A(n_639),
.Y(n_814)
);

BUFx2_ASAP7_75t_L g815 ( 
.A(n_658),
.Y(n_815)
);

NOR3xp33_ASAP7_75t_L g816 ( 
.A(n_679),
.B(n_282),
.C(n_295),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_654),
.B(n_529),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_664),
.Y(n_818)
);

OAI21xp5_ASAP7_75t_L g819 ( 
.A1(n_619),
.A2(n_620),
.B(n_624),
.Y(n_819)
);

OAI22xp5_ASAP7_75t_L g820 ( 
.A1(n_690),
.A2(n_529),
.B1(n_539),
.B2(n_550),
.Y(n_820)
);

BUFx6f_ASAP7_75t_L g821 ( 
.A(n_663),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_665),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_672),
.A2(n_522),
.B(n_525),
.Y(n_823)
);

OAI21xp5_ASAP7_75t_L g824 ( 
.A1(n_690),
.A2(n_542),
.B(n_547),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_671),
.B(n_687),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_671),
.B(n_542),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_687),
.B(n_547),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_665),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_609),
.Y(n_829)
);

NOR2x1p5_ASAP7_75t_SL g830 ( 
.A(n_693),
.B(n_461),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_628),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_605),
.B(n_509),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_693),
.B(n_549),
.Y(n_833)
);

INVx2_ASAP7_75t_SL g834 ( 
.A(n_658),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_725),
.B(n_461),
.Y(n_835)
);

AOI21xp5_ASAP7_75t_L g836 ( 
.A1(n_673),
.A2(n_522),
.B(n_525),
.Y(n_836)
);

AOI21xp5_ASAP7_75t_L g837 ( 
.A1(n_675),
.A2(n_525),
.B(n_589),
.Y(n_837)
);

OR2x6_ASAP7_75t_L g838 ( 
.A(n_616),
.B(n_209),
.Y(n_838)
);

O2A1O1Ixp33_ASAP7_75t_L g839 ( 
.A1(n_744),
.A2(n_473),
.B(n_463),
.C(n_462),
.Y(n_839)
);

INVx11_ASAP7_75t_L g840 ( 
.A(n_714),
.Y(n_840)
);

INVx11_ASAP7_75t_L g841 ( 
.A(n_682),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_745),
.B(n_462),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_678),
.A2(n_509),
.B(n_589),
.Y(n_843)
);

OAI22xp5_ASAP7_75t_L g844 ( 
.A1(n_668),
.A2(n_463),
.B1(n_465),
.B2(n_589),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_605),
.B(n_509),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_657),
.Y(n_846)
);

AOI22xp5_ASAP7_75t_L g847 ( 
.A1(n_710),
.A2(n_582),
.B1(n_465),
.B2(n_589),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_710),
.B(n_589),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_738),
.A2(n_527),
.B(n_502),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_725),
.B(n_582),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_666),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_608),
.B(n_582),
.Y(n_852)
);

BUFx4f_ASAP7_75t_L g853 ( 
.A(n_755),
.Y(n_853)
);

BUFx6f_ASAP7_75t_L g854 ( 
.A(n_663),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_738),
.A2(n_527),
.B(n_502),
.Y(n_855)
);

INVx4_ASAP7_75t_L g856 ( 
.A(n_663),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_768),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_611),
.B(n_298),
.Y(n_858)
);

OAI21xp5_ASAP7_75t_L g859 ( 
.A1(n_648),
.A2(n_416),
.B(n_398),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_720),
.A2(n_527),
.B(n_502),
.Y(n_860)
);

HB1xp67_ASAP7_75t_L g861 ( 
.A(n_608),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_610),
.B(n_406),
.Y(n_862)
);

OAI321xp33_ASAP7_75t_L g863 ( 
.A1(n_751),
.A2(n_424),
.A3(n_428),
.B1(n_420),
.B2(n_419),
.C(n_304),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_721),
.A2(n_527),
.B(n_502),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_610),
.B(n_406),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_768),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_769),
.Y(n_867)
);

INVx3_ASAP7_75t_L g868 ( 
.A(n_626),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_645),
.B(n_717),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_697),
.A2(n_527),
.B(n_502),
.Y(n_870)
);

NOR2x1_ASAP7_75t_L g871 ( 
.A(n_676),
.B(n_433),
.Y(n_871)
);

AND2x4_ASAP7_75t_L g872 ( 
.A(n_641),
.B(n_419),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_645),
.B(n_406),
.Y(n_873)
);

AOI21x1_ASAP7_75t_L g874 ( 
.A1(n_719),
.A2(n_398),
.B(n_386),
.Y(n_874)
);

O2A1O1Ixp33_ASAP7_75t_L g875 ( 
.A1(n_630),
.A2(n_451),
.B(n_438),
.C(n_436),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_SL g876 ( 
.A(n_684),
.B(n_304),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_647),
.B(n_406),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_606),
.B(n_450),
.Y(n_878)
);

OAI22xp5_ASAP7_75t_L g879 ( 
.A1(n_668),
.A2(n_209),
.B1(n_444),
.B2(n_450),
.Y(n_879)
);

BUFx2_ASAP7_75t_L g880 ( 
.A(n_682),
.Y(n_880)
);

OAI22xp5_ASAP7_75t_L g881 ( 
.A1(n_647),
.A2(n_450),
.B1(n_444),
.B2(n_299),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_704),
.B(n_450),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_697),
.A2(n_771),
.B(n_770),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_704),
.B(n_450),
.Y(n_884)
);

OR2x2_ASAP7_75t_L g885 ( 
.A(n_706),
.B(n_659),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_634),
.A2(n_438),
.B(n_436),
.Y(n_886)
);

OAI21xp5_ASAP7_75t_L g887 ( 
.A1(n_643),
.A2(n_649),
.B(n_646),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_642),
.B(n_444),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_669),
.B(n_444),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_730),
.Y(n_890)
);

INVx2_ASAP7_75t_SL g891 ( 
.A(n_752),
.Y(n_891)
);

INVx1_ASAP7_75t_SL g892 ( 
.A(n_732),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_674),
.B(n_444),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_773),
.A2(n_436),
.B(n_434),
.Y(n_894)
);

A2O1A1Ixp33_ASAP7_75t_L g895 ( 
.A1(n_638),
.A2(n_428),
.B(n_424),
.C(n_420),
.Y(n_895)
);

OAI22xp5_ASAP7_75t_L g896 ( 
.A1(n_775),
.A2(n_450),
.B1(n_444),
.B2(n_434),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_663),
.B(n_450),
.Y(n_897)
);

OAI22xp5_ASAP7_75t_L g898 ( 
.A1(n_626),
.A2(n_450),
.B1(n_444),
.B2(n_434),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_741),
.A2(n_433),
.B(n_388),
.Y(n_899)
);

AOI21xp33_ASAP7_75t_L g900 ( 
.A1(n_638),
.A2(n_420),
.B(n_6),
.Y(n_900)
);

NOR3xp33_ASAP7_75t_L g901 ( 
.A(n_757),
.B(n_423),
.C(n_418),
.Y(n_901)
);

A2O1A1Ixp33_ASAP7_75t_L g902 ( 
.A1(n_653),
.A2(n_418),
.B(n_426),
.C(n_423),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_SL g903 ( 
.A(n_699),
.B(n_450),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_691),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_747),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_694),
.B(n_444),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_695),
.Y(n_907)
);

BUFx6f_ASAP7_75t_L g908 ( 
.A(n_699),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_746),
.A2(n_386),
.B(n_388),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_747),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_L g911 ( 
.A(n_659),
.B(n_4),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_L g912 ( 
.A(n_685),
.B(n_7),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_707),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_709),
.Y(n_914)
);

AOI21x1_ASAP7_75t_L g915 ( 
.A1(n_719),
.A2(n_386),
.B(n_388),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_699),
.B(n_444),
.Y(n_916)
);

A2O1A1Ixp33_ASAP7_75t_L g917 ( 
.A1(n_653),
.A2(n_426),
.B(n_418),
.C(n_423),
.Y(n_917)
);

AND2x4_ASAP7_75t_L g918 ( 
.A(n_637),
.B(n_423),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_L g919 ( 
.A(n_685),
.B(n_9),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_SL g920 ( 
.A(n_699),
.B(n_444),
.Y(n_920)
);

NOR3xp33_ASAP7_75t_L g921 ( 
.A(n_617),
.B(n_418),
.C(n_426),
.Y(n_921)
);

OR2x2_ASAP7_75t_L g922 ( 
.A(n_705),
.B(n_418),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_705),
.B(n_304),
.Y(n_923)
);

INVx11_ASAP7_75t_L g924 ( 
.A(n_644),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_711),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_736),
.B(n_426),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_718),
.B(n_656),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_L g928 ( 
.A(n_692),
.B(n_10),
.Y(n_928)
);

INVx3_ASAP7_75t_L g929 ( 
.A(n_656),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_696),
.A2(n_398),
.B(n_426),
.Y(n_930)
);

OR2x2_ASAP7_75t_L g931 ( 
.A(n_698),
.B(n_11),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_736),
.B(n_427),
.Y(n_932)
);

AO21x1_ASAP7_75t_L g933 ( 
.A1(n_772),
.A2(n_11),
.B(n_18),
.Y(n_933)
);

INVxp67_ASAP7_75t_R g934 ( 
.A(n_644),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_677),
.B(n_19),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_774),
.Y(n_936)
);

A2O1A1Ixp33_ASAP7_75t_L g937 ( 
.A1(n_677),
.A2(n_723),
.B(n_762),
.C(n_734),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_713),
.A2(n_427),
.B(n_70),
.Y(n_938)
);

AOI21xp33_ASAP7_75t_L g939 ( 
.A1(n_715),
.A2(n_21),
.B(n_22),
.Y(n_939)
);

INVx3_ASAP7_75t_L g940 ( 
.A(n_736),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_736),
.B(n_427),
.Y(n_941)
);

AND2x4_ASAP7_75t_L g942 ( 
.A(n_702),
.B(n_650),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_731),
.B(n_427),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_748),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_750),
.A2(n_427),
.B(n_76),
.Y(n_945)
);

OAI22xp33_ASAP7_75t_L g946 ( 
.A1(n_683),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_946)
);

AOI21xp33_ASAP7_75t_L g947 ( 
.A1(n_715),
.A2(n_26),
.B(n_32),
.Y(n_947)
);

AOI21xp33_ASAP7_75t_L g948 ( 
.A1(n_734),
.A2(n_33),
.B(n_34),
.Y(n_948)
);

BUFx6f_ASAP7_75t_L g949 ( 
.A(n_761),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_754),
.A2(n_427),
.B(n_91),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_723),
.B(n_427),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_652),
.B(n_34),
.Y(n_952)
);

NOR3xp33_ASAP7_75t_L g953 ( 
.A(n_762),
.B(n_735),
.C(n_670),
.Y(n_953)
);

BUFx6f_ASAP7_75t_L g954 ( 
.A(n_759),
.Y(n_954)
);

INVx11_ASAP7_75t_L g955 ( 
.A(n_708),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_767),
.A2(n_427),
.B(n_98),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_782),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_SL g958 ( 
.A(n_937),
.B(n_739),
.Y(n_958)
);

BUFx6f_ASAP7_75t_L g959 ( 
.A(n_798),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_937),
.B(n_767),
.Y(n_960)
);

NOR3xp33_ASAP7_75t_SL g961 ( 
.A(n_935),
.B(n_622),
.C(n_629),
.Y(n_961)
);

OAI22xp5_ASAP7_75t_L g962 ( 
.A1(n_776),
.A2(n_636),
.B1(n_753),
.B2(n_724),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_780),
.B(n_753),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_923),
.B(n_753),
.Y(n_964)
);

OAI21x1_ASAP7_75t_L g965 ( 
.A1(n_808),
.A2(n_726),
.B(n_727),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_SL g966 ( 
.A(n_954),
.B(n_742),
.Y(n_966)
);

AOI22xp33_ASAP7_75t_L g967 ( 
.A1(n_946),
.A2(n_935),
.B1(n_911),
.B2(n_919),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_861),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_883),
.A2(n_655),
.B(n_686),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_779),
.A2(n_756),
.B(n_763),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_885),
.B(n_729),
.Y(n_971)
);

HB1xp67_ASAP7_75t_L g972 ( 
.A(n_861),
.Y(n_972)
);

CKINVDCx20_ASAP7_75t_R g973 ( 
.A(n_790),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_796),
.Y(n_974)
);

O2A1O1Ixp33_ASAP7_75t_L g975 ( 
.A1(n_912),
.A2(n_919),
.B(n_911),
.C(n_900),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_800),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_777),
.A2(n_764),
.B(n_763),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_780),
.B(n_758),
.Y(n_978)
);

NAND3xp33_ASAP7_75t_SL g979 ( 
.A(n_816),
.B(n_760),
.C(n_716),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_857),
.Y(n_980)
);

AOI22xp33_ASAP7_75t_L g981 ( 
.A1(n_946),
.A2(n_766),
.B1(n_729),
.B2(n_764),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_SL g982 ( 
.A(n_954),
.B(n_783),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_866),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_867),
.Y(n_984)
);

AOI22xp33_ASAP7_75t_L g985 ( 
.A1(n_912),
.A2(n_749),
.B1(n_688),
.B2(n_689),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_786),
.A2(n_681),
.B(n_737),
.Y(n_986)
);

BUFx12f_ASAP7_75t_L g987 ( 
.A(n_880),
.Y(n_987)
);

INVx2_ASAP7_75t_SL g988 ( 
.A(n_802),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_SL g989 ( 
.A(n_954),
.B(n_765),
.Y(n_989)
);

AO22x1_ASAP7_75t_L g990 ( 
.A1(n_816),
.A2(n_733),
.B1(n_728),
.B2(n_740),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_812),
.B(n_858),
.Y(n_991)
);

AOI21x1_ASAP7_75t_L g992 ( 
.A1(n_785),
.A2(n_427),
.B(n_90),
.Y(n_992)
);

OAI21xp33_ASAP7_75t_SL g993 ( 
.A1(n_784),
.A2(n_39),
.B(n_40),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_842),
.B(n_43),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_L g995 ( 
.A(n_810),
.B(n_43),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_818),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_822),
.Y(n_997)
);

HB1xp67_ASAP7_75t_L g998 ( 
.A(n_798),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_SL g999 ( 
.A(n_954),
.B(n_99),
.Y(n_999)
);

NOR2xp33_ASAP7_75t_R g1000 ( 
.A(n_853),
.B(n_110),
.Y(n_1000)
);

AOI211xp5_ASAP7_75t_L g1001 ( 
.A1(n_858),
.A2(n_45),
.B(n_46),
.C(n_51),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_887),
.A2(n_119),
.B(n_143),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_842),
.B(n_45),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_793),
.A2(n_81),
.B(n_142),
.Y(n_1004)
);

INVx5_ASAP7_75t_L g1005 ( 
.A(n_798),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_828),
.Y(n_1006)
);

AOI221xp5_ASAP7_75t_L g1007 ( 
.A1(n_939),
.A2(n_51),
.B1(n_52),
.B2(n_53),
.C(n_54),
.Y(n_1007)
);

AOI22xp33_ASAP7_75t_L g1008 ( 
.A1(n_947),
.A2(n_427),
.B1(n_53),
.B2(n_57),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_890),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_829),
.Y(n_1010)
);

OAI22xp5_ASAP7_75t_SL g1011 ( 
.A1(n_838),
.A2(n_52),
.B1(n_61),
.B2(n_69),
.Y(n_1011)
);

NOR2xp33_ASAP7_75t_SL g1012 ( 
.A(n_791),
.B(n_427),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_869),
.A2(n_75),
.B(n_123),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_SL g1014 ( 
.A(n_819),
.B(n_128),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_SL g1015 ( 
.A(n_778),
.B(n_131),
.Y(n_1015)
);

A2O1A1Ixp33_ASAP7_75t_L g1016 ( 
.A1(n_928),
.A2(n_135),
.B(n_140),
.C(n_141),
.Y(n_1016)
);

CKINVDCx14_ASAP7_75t_R g1017 ( 
.A(n_815),
.Y(n_1017)
);

A2O1A1Ixp33_ASAP7_75t_L g1018 ( 
.A1(n_928),
.A2(n_953),
.B(n_848),
.C(n_831),
.Y(n_1018)
);

HB1xp67_ASAP7_75t_L g1019 ( 
.A(n_798),
.Y(n_1019)
);

O2A1O1Ixp5_ASAP7_75t_SL g1020 ( 
.A1(n_948),
.A2(n_926),
.B(n_879),
.C(n_896),
.Y(n_1020)
);

OAI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_784),
.A2(n_922),
.B1(n_848),
.B2(n_809),
.Y(n_1021)
);

INVx4_ASAP7_75t_L g1022 ( 
.A(n_821),
.Y(n_1022)
);

INVx3_ASAP7_75t_L g1023 ( 
.A(n_821),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_L g1024 ( 
.A(n_913),
.B(n_914),
.Y(n_1024)
);

AO21x1_ASAP7_75t_L g1025 ( 
.A1(n_803),
.A2(n_953),
.B(n_794),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_846),
.B(n_851),
.Y(n_1026)
);

INVx2_ASAP7_75t_SL g1027 ( 
.A(n_834),
.Y(n_1027)
);

INVx4_ASAP7_75t_L g1028 ( 
.A(n_821),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_904),
.B(n_907),
.Y(n_1029)
);

BUFx2_ASAP7_75t_L g1030 ( 
.A(n_853),
.Y(n_1030)
);

A2O1A1Ixp33_ASAP7_75t_L g1031 ( 
.A1(n_942),
.A2(n_925),
.B(n_787),
.C(n_956),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_L g1032 ( 
.A(n_892),
.B(n_931),
.Y(n_1032)
);

A2O1A1Ixp33_ASAP7_75t_L g1033 ( 
.A1(n_942),
.A2(n_788),
.B(n_807),
.C(n_781),
.Y(n_1033)
);

AND2x4_ASAP7_75t_L g1034 ( 
.A(n_872),
.B(n_856),
.Y(n_1034)
);

OR2x2_ASAP7_75t_L g1035 ( 
.A(n_872),
.B(n_838),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_SL g1036 ( 
.A(n_821),
.B(n_854),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_L g1037 ( 
.A(n_838),
.B(n_788),
.Y(n_1037)
);

BUFx6f_ASAP7_75t_L g1038 ( 
.A(n_854),
.Y(n_1038)
);

NOR3xp33_ASAP7_75t_SL g1039 ( 
.A(n_863),
.B(n_807),
.C(n_951),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_SL g1040 ( 
.A(n_854),
.B(n_908),
.Y(n_1040)
);

OAI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_868),
.A2(n_817),
.B1(n_825),
.B2(n_927),
.Y(n_1041)
);

BUFx6f_ASAP7_75t_L g1042 ( 
.A(n_854),
.Y(n_1042)
);

OAI21x1_ASAP7_75t_L g1043 ( 
.A1(n_843),
.A2(n_837),
.B(n_799),
.Y(n_1043)
);

OAI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_868),
.A2(n_850),
.B1(n_814),
.B2(n_847),
.Y(n_1044)
);

AND2x2_ASAP7_75t_L g1045 ( 
.A(n_952),
.B(n_876),
.Y(n_1045)
);

AND2x2_ASAP7_75t_SL g1046 ( 
.A(n_908),
.B(n_856),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_795),
.B(n_797),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_944),
.B(n_792),
.Y(n_1048)
);

AND2x4_ASAP7_75t_L g1049 ( 
.A(n_805),
.B(n_940),
.Y(n_1049)
);

NOR2xp67_ASAP7_75t_SL g1050 ( 
.A(n_908),
.B(n_940),
.Y(n_1050)
);

AOI22xp33_ASAP7_75t_L g1051 ( 
.A1(n_933),
.A2(n_901),
.B1(n_921),
.B2(n_936),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_L g1052 ( 
.A(n_878),
.B(n_814),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_870),
.A2(n_804),
.B(n_813),
.Y(n_1053)
);

OAI22xp5_ASAP7_75t_L g1054 ( 
.A1(n_929),
.A2(n_908),
.B1(n_852),
.B2(n_804),
.Y(n_1054)
);

OAI22x1_ASAP7_75t_L g1055 ( 
.A1(n_891),
.A2(n_918),
.B1(n_813),
.B2(n_929),
.Y(n_1055)
);

INVx2_ASAP7_75t_SL g1056 ( 
.A(n_924),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_901),
.B(n_905),
.Y(n_1057)
);

BUFx6f_ASAP7_75t_L g1058 ( 
.A(n_805),
.Y(n_1058)
);

A2O1A1Ixp33_ASAP7_75t_L g1059 ( 
.A1(n_895),
.A2(n_894),
.B(n_830),
.C(n_871),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_910),
.B(n_918),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_897),
.A2(n_920),
.B(n_916),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_897),
.A2(n_920),
.B(n_916),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_903),
.A2(n_836),
.B(n_801),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_934),
.B(n_921),
.Y(n_1064)
);

A2O1A1Ixp33_ASAP7_75t_L g1065 ( 
.A1(n_839),
.A2(n_888),
.B(n_875),
.C(n_789),
.Y(n_1065)
);

NOR2xp67_ASAP7_75t_L g1066 ( 
.A(n_932),
.B(n_941),
.Y(n_1066)
);

AND2x4_ASAP7_75t_L g1067 ( 
.A(n_949),
.B(n_926),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_826),
.B(n_827),
.Y(n_1068)
);

O2A1O1Ixp33_ASAP7_75t_L g1069 ( 
.A1(n_902),
.A2(n_917),
.B(n_881),
.C(n_889),
.Y(n_1069)
);

INVxp67_ASAP7_75t_L g1070 ( 
.A(n_893),
.Y(n_1070)
);

AND2x2_ASAP7_75t_L g1071 ( 
.A(n_824),
.B(n_859),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_903),
.A2(n_823),
.B(n_873),
.Y(n_1072)
);

INVx3_ASAP7_75t_L g1073 ( 
.A(n_949),
.Y(n_1073)
);

CKINVDCx10_ASAP7_75t_R g1074 ( 
.A(n_806),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_833),
.Y(n_1075)
);

OR2x6_ASAP7_75t_L g1076 ( 
.A(n_840),
.B(n_949),
.Y(n_1076)
);

OAI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_832),
.A2(n_845),
.B1(n_835),
.B2(n_949),
.Y(n_1077)
);

HB1xp67_ASAP7_75t_L g1078 ( 
.A(n_906),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_862),
.A2(n_865),
.B(n_832),
.Y(n_1079)
);

NOR2xp33_ASAP7_75t_L g1080 ( 
.A(n_845),
.B(n_877),
.Y(n_1080)
);

A2O1A1Ixp33_ASAP7_75t_L g1081 ( 
.A1(n_943),
.A2(n_917),
.B(n_886),
.C(n_811),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_820),
.B(n_877),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_882),
.A2(n_884),
.B(n_844),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_L g1084 ( 
.A(n_955),
.B(n_915),
.Y(n_1084)
);

BUFx3_ASAP7_75t_L g1085 ( 
.A(n_841),
.Y(n_1085)
);

AOI21x1_ASAP7_75t_L g1086 ( 
.A1(n_874),
.A2(n_899),
.B(n_930),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_L g1087 ( 
.A(n_898),
.B(n_909),
.Y(n_1087)
);

AND2x2_ASAP7_75t_L g1088 ( 
.A(n_945),
.B(n_950),
.Y(n_1088)
);

AND2x2_ASAP7_75t_L g1089 ( 
.A(n_938),
.B(n_849),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_SL g1090 ( 
.A(n_860),
.B(n_864),
.Y(n_1090)
);

O2A1O1Ixp5_ASAP7_75t_L g1091 ( 
.A1(n_855),
.A2(n_935),
.B(n_911),
.C(n_937),
.Y(n_1091)
);

O2A1O1Ixp33_ASAP7_75t_SL g1092 ( 
.A1(n_937),
.A2(n_946),
.B(n_900),
.C(n_935),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_861),
.Y(n_1093)
);

BUFx3_ASAP7_75t_L g1094 ( 
.A(n_802),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_L g1095 ( 
.A(n_885),
.B(n_701),
.Y(n_1095)
);

OAI22xp5_ASAP7_75t_L g1096 ( 
.A1(n_937),
.A2(n_777),
.B1(n_783),
.B2(n_776),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_861),
.Y(n_1097)
);

BUFx3_ASAP7_75t_L g1098 ( 
.A(n_802),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_883),
.A2(n_536),
.B(n_477),
.Y(n_1099)
);

OA21x2_ASAP7_75t_L g1100 ( 
.A1(n_970),
.A2(n_1091),
.B(n_1065),
.Y(n_1100)
);

AOI21x1_ASAP7_75t_L g1101 ( 
.A1(n_990),
.A2(n_969),
.B(n_1090),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_1099),
.A2(n_1047),
.B(n_1063),
.Y(n_1102)
);

BUFx3_ASAP7_75t_L g1103 ( 
.A(n_1094),
.Y(n_1103)
);

AOI22xp5_ASAP7_75t_L g1104 ( 
.A1(n_995),
.A2(n_967),
.B1(n_1095),
.B2(n_958),
.Y(n_1104)
);

AOI221xp5_ASAP7_75t_SL g1105 ( 
.A1(n_967),
.A2(n_975),
.B1(n_1007),
.B2(n_995),
.C(n_1008),
.Y(n_1105)
);

NAND3xp33_ASAP7_75t_L g1106 ( 
.A(n_961),
.B(n_1018),
.C(n_1001),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_1095),
.B(n_991),
.Y(n_1107)
);

INVx3_ASAP7_75t_L g1108 ( 
.A(n_1058),
.Y(n_1108)
);

AO31x2_ASAP7_75t_L g1109 ( 
.A1(n_1025),
.A2(n_1096),
.A3(n_1081),
.B(n_962),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_978),
.B(n_1024),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_977),
.A2(n_1031),
.B(n_1021),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_1024),
.B(n_1032),
.Y(n_1112)
);

INVxp67_ASAP7_75t_L g1113 ( 
.A(n_1098),
.Y(n_1113)
);

AOI22xp5_ASAP7_75t_L g1114 ( 
.A1(n_958),
.A2(n_1032),
.B1(n_964),
.B2(n_1045),
.Y(n_1114)
);

OAI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_1033),
.A2(n_1052),
.B(n_1092),
.Y(n_1115)
);

OAI21x1_ASAP7_75t_L g1116 ( 
.A1(n_1043),
.A2(n_1072),
.B(n_1086),
.Y(n_1116)
);

INVx2_ASAP7_75t_SL g1117 ( 
.A(n_988),
.Y(n_1117)
);

O2A1O1Ixp33_ASAP7_75t_SL g1118 ( 
.A1(n_960),
.A2(n_1016),
.B(n_1014),
.C(n_979),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_1083),
.A2(n_1068),
.B(n_1071),
.Y(n_1119)
);

NOR2xp33_ASAP7_75t_L g1120 ( 
.A(n_1030),
.B(n_972),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_1075),
.B(n_972),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_1048),
.B(n_968),
.Y(n_1122)
);

NOR2xp33_ASAP7_75t_SL g1123 ( 
.A(n_1046),
.B(n_1011),
.Y(n_1123)
);

NOR4xp25_ASAP7_75t_L g1124 ( 
.A(n_994),
.B(n_1003),
.C(n_1008),
.D(n_960),
.Y(n_1124)
);

AOI221x1_ASAP7_75t_L g1125 ( 
.A1(n_1002),
.A2(n_963),
.B1(n_1037),
.B2(n_1053),
.C(n_1059),
.Y(n_1125)
);

OAI21x1_ASAP7_75t_L g1126 ( 
.A1(n_1079),
.A2(n_1090),
.B(n_965),
.Y(n_1126)
);

O2A1O1Ixp33_ASAP7_75t_L g1127 ( 
.A1(n_961),
.A2(n_1037),
.B(n_1014),
.C(n_1064),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1026),
.Y(n_1128)
);

CKINVDCx20_ASAP7_75t_R g1129 ( 
.A(n_973),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_1087),
.A2(n_986),
.B(n_982),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_1087),
.A2(n_982),
.B(n_966),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_1093),
.B(n_1097),
.Y(n_1132)
);

OR2x2_ASAP7_75t_L g1133 ( 
.A(n_1029),
.B(n_1035),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_974),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1052),
.B(n_1034),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_966),
.A2(n_1082),
.B(n_989),
.Y(n_1136)
);

BUFx3_ASAP7_75t_L g1137 ( 
.A(n_1085),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_1034),
.B(n_1070),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_976),
.Y(n_1139)
);

O2A1O1Ixp33_ASAP7_75t_SL g1140 ( 
.A1(n_1015),
.A2(n_999),
.B(n_989),
.C(n_1057),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_SL g1141 ( 
.A(n_1046),
.B(n_971),
.Y(n_1141)
);

AO32x2_ASAP7_75t_L g1142 ( 
.A1(n_1041),
.A2(n_1044),
.A3(n_1077),
.B1(n_1054),
.B2(n_1020),
.Y(n_1142)
);

OAI21x1_ASAP7_75t_L g1143 ( 
.A1(n_992),
.A2(n_1062),
.B(n_1061),
.Y(n_1143)
);

INVx2_ASAP7_75t_SL g1144 ( 
.A(n_1027),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_1089),
.A2(n_1088),
.B(n_1069),
.Y(n_1145)
);

OR2x6_ASAP7_75t_L g1146 ( 
.A(n_1076),
.B(n_1058),
.Y(n_1146)
);

AO31x2_ASAP7_75t_L g1147 ( 
.A1(n_1080),
.A2(n_1055),
.A3(n_1004),
.B(n_1013),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1078),
.B(n_981),
.Y(n_1148)
);

NAND2xp33_ASAP7_75t_L g1149 ( 
.A(n_1058),
.B(n_1000),
.Y(n_1149)
);

O2A1O1Ixp33_ASAP7_75t_L g1150 ( 
.A1(n_1015),
.A2(n_993),
.B(n_971),
.C(n_999),
.Y(n_1150)
);

AO31x2_ASAP7_75t_L g1151 ( 
.A1(n_1080),
.A2(n_997),
.A3(n_996),
.B(n_1006),
.Y(n_1151)
);

NOR2xp33_ASAP7_75t_L g1152 ( 
.A(n_1017),
.B(n_1058),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_1074),
.Y(n_1153)
);

OAI21x1_ASAP7_75t_L g1154 ( 
.A1(n_1051),
.A2(n_1036),
.B(n_1040),
.Y(n_1154)
);

OR2x2_ASAP7_75t_L g1155 ( 
.A(n_1060),
.B(n_957),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1078),
.B(n_981),
.Y(n_1156)
);

OAI21x1_ASAP7_75t_L g1157 ( 
.A1(n_1051),
.A2(n_1040),
.B(n_1036),
.Y(n_1157)
);

BUFx3_ASAP7_75t_L g1158 ( 
.A(n_1056),
.Y(n_1158)
);

OAI21x1_ASAP7_75t_L g1159 ( 
.A1(n_1073),
.A2(n_985),
.B(n_1066),
.Y(n_1159)
);

OR2x6_ASAP7_75t_L g1160 ( 
.A(n_1076),
.B(n_1049),
.Y(n_1160)
);

BUFx3_ASAP7_75t_L g1161 ( 
.A(n_987),
.Y(n_1161)
);

O2A1O1Ixp33_ASAP7_75t_L g1162 ( 
.A1(n_1084),
.A2(n_1039),
.B(n_1076),
.C(n_980),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1005),
.A2(n_985),
.B(n_1067),
.Y(n_1163)
);

BUFx6f_ASAP7_75t_L g1164 ( 
.A(n_1038),
.Y(n_1164)
);

O2A1O1Ixp5_ASAP7_75t_L g1165 ( 
.A1(n_1084),
.A2(n_1067),
.B(n_1050),
.C(n_1023),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1005),
.A2(n_1049),
.B(n_1019),
.Y(n_1166)
);

A2O1A1Ixp33_ASAP7_75t_L g1167 ( 
.A1(n_1039),
.A2(n_983),
.B(n_984),
.C(n_1009),
.Y(n_1167)
);

BUFx6f_ASAP7_75t_L g1168 ( 
.A(n_1038),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_998),
.B(n_1019),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_998),
.B(n_1022),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_959),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_959),
.Y(n_1172)
);

BUFx8_ASAP7_75t_L g1173 ( 
.A(n_1038),
.Y(n_1173)
);

AOI21x1_ASAP7_75t_L g1174 ( 
.A1(n_1005),
.A2(n_959),
.B(n_1042),
.Y(n_1174)
);

AND2x6_ASAP7_75t_L g1175 ( 
.A(n_1042),
.B(n_1000),
.Y(n_1175)
);

AOI31xp67_ASAP7_75t_L g1176 ( 
.A1(n_1012),
.A2(n_1005),
.A3(n_1042),
.B(n_1028),
.Y(n_1176)
);

AOI221x1_ASAP7_75t_L g1177 ( 
.A1(n_1028),
.A2(n_937),
.B1(n_935),
.B2(n_911),
.C(n_912),
.Y(n_1177)
);

BUFx6f_ASAP7_75t_L g1178 ( 
.A(n_1038),
.Y(n_1178)
);

INVx3_ASAP7_75t_L g1179 ( 
.A(n_1058),
.Y(n_1179)
);

OA21x2_ASAP7_75t_L g1180 ( 
.A1(n_970),
.A2(n_1091),
.B(n_1065),
.Y(n_1180)
);

CKINVDCx20_ASAP7_75t_R g1181 ( 
.A(n_973),
.Y(n_1181)
);

O2A1O1Ixp33_ASAP7_75t_SL g1182 ( 
.A1(n_975),
.A2(n_937),
.B(n_1033),
.C(n_958),
.Y(n_1182)
);

INVx1_ASAP7_75t_SL g1183 ( 
.A(n_1094),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_SL g1184 ( 
.A(n_991),
.B(n_475),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_1074),
.Y(n_1185)
);

AOI21x1_ASAP7_75t_L g1186 ( 
.A1(n_990),
.A2(n_970),
.B(n_969),
.Y(n_1186)
);

BUFx10_ASAP7_75t_L g1187 ( 
.A(n_995),
.Y(n_1187)
);

BUFx6f_ASAP7_75t_L g1188 ( 
.A(n_1038),
.Y(n_1188)
);

OR2x6_ASAP7_75t_L g1189 ( 
.A(n_1076),
.B(n_1030),
.Y(n_1189)
);

OR2x6_ASAP7_75t_L g1190 ( 
.A(n_1076),
.B(n_1030),
.Y(n_1190)
);

INVx2_ASAP7_75t_SL g1191 ( 
.A(n_1094),
.Y(n_1191)
);

BUFx2_ASAP7_75t_L g1192 ( 
.A(n_1094),
.Y(n_1192)
);

AOI22xp5_ASAP7_75t_L g1193 ( 
.A1(n_995),
.A2(n_911),
.B1(n_935),
.B2(n_919),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1095),
.B(n_585),
.Y(n_1194)
);

O2A1O1Ixp33_ASAP7_75t_SL g1195 ( 
.A1(n_975),
.A2(n_937),
.B(n_1033),
.C(n_958),
.Y(n_1195)
);

O2A1O1Ixp33_ASAP7_75t_SL g1196 ( 
.A1(n_975),
.A2(n_937),
.B(n_1033),
.C(n_958),
.Y(n_1196)
);

O2A1O1Ixp33_ASAP7_75t_L g1197 ( 
.A1(n_975),
.A2(n_937),
.B(n_701),
.C(n_919),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_970),
.A2(n_969),
.B(n_883),
.Y(n_1198)
);

INVx2_ASAP7_75t_SL g1199 ( 
.A(n_1094),
.Y(n_1199)
);

NAND3xp33_ASAP7_75t_L g1200 ( 
.A(n_975),
.B(n_967),
.C(n_995),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_970),
.A2(n_969),
.B(n_883),
.Y(n_1201)
);

AO31x2_ASAP7_75t_L g1202 ( 
.A1(n_1025),
.A2(n_1096),
.A3(n_1065),
.B(n_1081),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1095),
.B(n_585),
.Y(n_1203)
);

OAI21x1_ASAP7_75t_L g1204 ( 
.A1(n_1043),
.A2(n_1063),
.B(n_1072),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_970),
.A2(n_969),
.B(n_883),
.Y(n_1205)
);

INVx3_ASAP7_75t_L g1206 ( 
.A(n_1058),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1095),
.B(n_585),
.Y(n_1207)
);

NOR2xp33_ASAP7_75t_L g1208 ( 
.A(n_1095),
.B(n_701),
.Y(n_1208)
);

OAI21x1_ASAP7_75t_L g1209 ( 
.A1(n_1043),
.A2(n_1063),
.B(n_1072),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_970),
.A2(n_969),
.B(n_883),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_970),
.A2(n_969),
.B(n_883),
.Y(n_1211)
);

NAND2xp33_ASAP7_75t_SL g1212 ( 
.A(n_961),
.B(n_1000),
.Y(n_1212)
);

O2A1O1Ixp5_ASAP7_75t_L g1213 ( 
.A1(n_958),
.A2(n_935),
.B(n_911),
.C(n_919),
.Y(n_1213)
);

OAI21x1_ASAP7_75t_L g1214 ( 
.A1(n_1043),
.A2(n_1063),
.B(n_1072),
.Y(n_1214)
);

NOR2xp33_ASAP7_75t_L g1215 ( 
.A(n_1095),
.B(n_701),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_970),
.A2(n_969),
.B(n_883),
.Y(n_1216)
);

AOI22xp5_ASAP7_75t_L g1217 ( 
.A1(n_995),
.A2(n_911),
.B1(n_935),
.B2(n_919),
.Y(n_1217)
);

AOI22xp33_ASAP7_75t_L g1218 ( 
.A1(n_967),
.A2(n_935),
.B1(n_911),
.B2(n_995),
.Y(n_1218)
);

OAI21x1_ASAP7_75t_L g1219 ( 
.A1(n_1043),
.A2(n_1063),
.B(n_1072),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_970),
.A2(n_969),
.B(n_883),
.Y(n_1220)
);

AO31x2_ASAP7_75t_L g1221 ( 
.A1(n_1025),
.A2(n_1096),
.A3(n_1065),
.B(n_1081),
.Y(n_1221)
);

OA21x2_ASAP7_75t_L g1222 ( 
.A1(n_970),
.A2(n_1091),
.B(n_1065),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1095),
.B(n_585),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1095),
.B(n_585),
.Y(n_1224)
);

O2A1O1Ixp33_ASAP7_75t_SL g1225 ( 
.A1(n_975),
.A2(n_937),
.B(n_1033),
.C(n_958),
.Y(n_1225)
);

AND2x2_ASAP7_75t_L g1226 ( 
.A(n_1095),
.B(n_585),
.Y(n_1226)
);

OAI22xp33_ASAP7_75t_L g1227 ( 
.A1(n_978),
.A2(n_701),
.B1(n_573),
.B2(n_505),
.Y(n_1227)
);

AOI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_995),
.A2(n_911),
.B1(n_935),
.B2(n_919),
.Y(n_1228)
);

AO31x2_ASAP7_75t_L g1229 ( 
.A1(n_1025),
.A2(n_1096),
.A3(n_1065),
.B(n_1081),
.Y(n_1229)
);

OAI21xp33_ASAP7_75t_L g1230 ( 
.A1(n_967),
.A2(n_680),
.B(n_911),
.Y(n_1230)
);

INVx4_ASAP7_75t_L g1231 ( 
.A(n_1005),
.Y(n_1231)
);

AND2x2_ASAP7_75t_L g1232 ( 
.A(n_1095),
.B(n_585),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1095),
.B(n_585),
.Y(n_1233)
);

NOR2xp33_ASAP7_75t_L g1234 ( 
.A(n_1095),
.B(n_701),
.Y(n_1234)
);

OAI22x1_ASAP7_75t_L g1235 ( 
.A1(n_995),
.A2(n_935),
.B1(n_919),
.B2(n_912),
.Y(n_1235)
);

CKINVDCx11_ASAP7_75t_R g1236 ( 
.A(n_973),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1010),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_970),
.A2(n_969),
.B(n_883),
.Y(n_1238)
);

OAI21x1_ASAP7_75t_L g1239 ( 
.A1(n_1043),
.A2(n_1063),
.B(n_1072),
.Y(n_1239)
);

OAI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_975),
.A2(n_967),
.B(n_1091),
.Y(n_1240)
);

O2A1O1Ixp33_ASAP7_75t_SL g1241 ( 
.A1(n_975),
.A2(n_937),
.B(n_1033),
.C(n_958),
.Y(n_1241)
);

AOI22xp33_ASAP7_75t_L g1242 ( 
.A1(n_1230),
.A2(n_1200),
.B1(n_1218),
.B2(n_1228),
.Y(n_1242)
);

INVx3_ASAP7_75t_SL g1243 ( 
.A(n_1153),
.Y(n_1243)
);

CKINVDCx11_ASAP7_75t_R g1244 ( 
.A(n_1236),
.Y(n_1244)
);

CKINVDCx11_ASAP7_75t_R g1245 ( 
.A(n_1129),
.Y(n_1245)
);

OR2x2_ASAP7_75t_L g1246 ( 
.A(n_1107),
.B(n_1112),
.Y(n_1246)
);

BUFx3_ASAP7_75t_L g1247 ( 
.A(n_1103),
.Y(n_1247)
);

INVx4_ASAP7_75t_SL g1248 ( 
.A(n_1175),
.Y(n_1248)
);

BUFx8_ASAP7_75t_L g1249 ( 
.A(n_1192),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1110),
.B(n_1226),
.Y(n_1250)
);

BUFx6f_ASAP7_75t_SL g1251 ( 
.A(n_1137),
.Y(n_1251)
);

AOI22xp33_ASAP7_75t_SL g1252 ( 
.A1(n_1123),
.A2(n_1200),
.B1(n_1106),
.B2(n_1240),
.Y(n_1252)
);

AOI22xp33_ASAP7_75t_SL g1253 ( 
.A1(n_1123),
.A2(n_1106),
.B1(n_1187),
.B2(n_1234),
.Y(n_1253)
);

CKINVDCx20_ASAP7_75t_R g1254 ( 
.A(n_1181),
.Y(n_1254)
);

AOI22xp33_ASAP7_75t_L g1255 ( 
.A1(n_1230),
.A2(n_1217),
.B1(n_1193),
.B2(n_1228),
.Y(n_1255)
);

BUFx12f_ASAP7_75t_L g1256 ( 
.A(n_1185),
.Y(n_1256)
);

INVx8_ASAP7_75t_L g1257 ( 
.A(n_1175),
.Y(n_1257)
);

AOI22xp33_ASAP7_75t_L g1258 ( 
.A1(n_1193),
.A2(n_1217),
.B1(n_1235),
.B2(n_1104),
.Y(n_1258)
);

OR2x2_ASAP7_75t_L g1259 ( 
.A(n_1133),
.B(n_1194),
.Y(n_1259)
);

BUFx3_ASAP7_75t_L g1260 ( 
.A(n_1173),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_1183),
.Y(n_1261)
);

INVx1_ASAP7_75t_SL g1262 ( 
.A(n_1117),
.Y(n_1262)
);

AOI22xp33_ASAP7_75t_SL g1263 ( 
.A1(n_1187),
.A2(n_1208),
.B1(n_1215),
.B2(n_1115),
.Y(n_1263)
);

BUFx3_ASAP7_75t_L g1264 ( 
.A(n_1158),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_L g1265 ( 
.A1(n_1104),
.A2(n_1212),
.B1(n_1227),
.B2(n_1114),
.Y(n_1265)
);

BUFx12f_ASAP7_75t_L g1266 ( 
.A(n_1191),
.Y(n_1266)
);

OAI22xp5_ASAP7_75t_L g1267 ( 
.A1(n_1203),
.A2(n_1224),
.B1(n_1207),
.B2(n_1233),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1232),
.B(n_1114),
.Y(n_1268)
);

AOI22xp33_ASAP7_75t_L g1269 ( 
.A1(n_1111),
.A2(n_1136),
.B1(n_1128),
.B2(n_1156),
.Y(n_1269)
);

BUFx3_ASAP7_75t_L g1270 ( 
.A(n_1199),
.Y(n_1270)
);

INVx3_ASAP7_75t_SL g1271 ( 
.A(n_1189),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1223),
.B(n_1122),
.Y(n_1272)
);

AND2x4_ASAP7_75t_SL g1273 ( 
.A(n_1189),
.B(n_1190),
.Y(n_1273)
);

NAND2x1p5_ASAP7_75t_L g1274 ( 
.A(n_1141),
.B(n_1159),
.Y(n_1274)
);

OAI22xp5_ASAP7_75t_L g1275 ( 
.A1(n_1148),
.A2(n_1135),
.B1(n_1138),
.B2(n_1120),
.Y(n_1275)
);

CKINVDCx11_ASAP7_75t_R g1276 ( 
.A(n_1161),
.Y(n_1276)
);

OAI22xp5_ASAP7_75t_L g1277 ( 
.A1(n_1184),
.A2(n_1190),
.B1(n_1189),
.B2(n_1127),
.Y(n_1277)
);

NAND2x1p5_ASAP7_75t_L g1278 ( 
.A(n_1174),
.B(n_1163),
.Y(n_1278)
);

OR2x2_ASAP7_75t_L g1279 ( 
.A(n_1121),
.B(n_1132),
.Y(n_1279)
);

NAND2x1p5_ASAP7_75t_L g1280 ( 
.A(n_1108),
.B(n_1179),
.Y(n_1280)
);

BUFx6f_ASAP7_75t_L g1281 ( 
.A(n_1164),
.Y(n_1281)
);

OAI22xp5_ASAP7_75t_L g1282 ( 
.A1(n_1190),
.A2(n_1197),
.B1(n_1162),
.B2(n_1146),
.Y(n_1282)
);

INVx2_ASAP7_75t_R g1283 ( 
.A(n_1172),
.Y(n_1283)
);

HB1xp67_ASAP7_75t_L g1284 ( 
.A(n_1151),
.Y(n_1284)
);

NAND2xp33_ASAP7_75t_SL g1285 ( 
.A(n_1144),
.B(n_1237),
.Y(n_1285)
);

BUFx6f_ASAP7_75t_L g1286 ( 
.A(n_1164),
.Y(n_1286)
);

BUFx4_ASAP7_75t_R g1287 ( 
.A(n_1171),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1134),
.Y(n_1288)
);

BUFx6f_ASAP7_75t_L g1289 ( 
.A(n_1168),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1139),
.Y(n_1290)
);

BUFx12f_ASAP7_75t_L g1291 ( 
.A(n_1173),
.Y(n_1291)
);

BUFx6f_ASAP7_75t_L g1292 ( 
.A(n_1168),
.Y(n_1292)
);

CKINVDCx20_ASAP7_75t_R g1293 ( 
.A(n_1152),
.Y(n_1293)
);

OAI22xp5_ASAP7_75t_L g1294 ( 
.A1(n_1146),
.A2(n_1160),
.B1(n_1150),
.B2(n_1145),
.Y(n_1294)
);

INVxp67_ASAP7_75t_SL g1295 ( 
.A(n_1154),
.Y(n_1295)
);

OAI22xp5_ASAP7_75t_L g1296 ( 
.A1(n_1146),
.A2(n_1160),
.B1(n_1167),
.B2(n_1155),
.Y(n_1296)
);

INVx4_ASAP7_75t_L g1297 ( 
.A(n_1175),
.Y(n_1297)
);

BUFx2_ASAP7_75t_L g1298 ( 
.A(n_1113),
.Y(n_1298)
);

AOI22xp33_ASAP7_75t_L g1299 ( 
.A1(n_1105),
.A2(n_1100),
.B1(n_1222),
.B2(n_1180),
.Y(n_1299)
);

BUFx10_ASAP7_75t_L g1300 ( 
.A(n_1175),
.Y(n_1300)
);

OAI22x1_ASAP7_75t_L g1301 ( 
.A1(n_1105),
.A2(n_1100),
.B1(n_1222),
.B2(n_1180),
.Y(n_1301)
);

AOI22xp33_ASAP7_75t_L g1302 ( 
.A1(n_1131),
.A2(n_1119),
.B1(n_1213),
.B2(n_1130),
.Y(n_1302)
);

OAI22xp5_ASAP7_75t_L g1303 ( 
.A1(n_1160),
.A2(n_1170),
.B1(n_1206),
.B2(n_1108),
.Y(n_1303)
);

AOI22xp33_ASAP7_75t_L g1304 ( 
.A1(n_1182),
.A2(n_1241),
.B1(n_1195),
.B2(n_1225),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1151),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1151),
.Y(n_1306)
);

BUFx2_ASAP7_75t_L g1307 ( 
.A(n_1169),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1178),
.Y(n_1308)
);

AOI22xp33_ASAP7_75t_SL g1309 ( 
.A1(n_1196),
.A2(n_1149),
.B1(n_1124),
.B2(n_1177),
.Y(n_1309)
);

INVx4_ASAP7_75t_L g1310 ( 
.A(n_1188),
.Y(n_1310)
);

BUFx2_ASAP7_75t_SL g1311 ( 
.A(n_1188),
.Y(n_1311)
);

BUFx8_ASAP7_75t_L g1312 ( 
.A(n_1188),
.Y(n_1312)
);

AO22x1_ASAP7_75t_L g1313 ( 
.A1(n_1179),
.A2(n_1206),
.B1(n_1165),
.B2(n_1118),
.Y(n_1313)
);

BUFx12f_ASAP7_75t_L g1314 ( 
.A(n_1166),
.Y(n_1314)
);

AOI22xp33_ASAP7_75t_L g1315 ( 
.A1(n_1124),
.A2(n_1198),
.B1(n_1201),
.B2(n_1210),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_SL g1316 ( 
.A1(n_1157),
.A2(n_1205),
.B1(n_1211),
.B2(n_1220),
.Y(n_1316)
);

CKINVDCx11_ASAP7_75t_R g1317 ( 
.A(n_1176),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_1102),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1202),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1202),
.Y(n_1320)
);

AOI22xp5_ASAP7_75t_SL g1321 ( 
.A1(n_1216),
.A2(n_1238),
.B1(n_1140),
.B2(n_1125),
.Y(n_1321)
);

AOI22xp33_ASAP7_75t_L g1322 ( 
.A1(n_1126),
.A2(n_1109),
.B1(n_1143),
.B2(n_1229),
.Y(n_1322)
);

BUFx12f_ASAP7_75t_L g1323 ( 
.A(n_1147),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1202),
.B(n_1229),
.Y(n_1324)
);

OAI22xp5_ASAP7_75t_L g1325 ( 
.A1(n_1186),
.A2(n_1101),
.B1(n_1229),
.B2(n_1221),
.Y(n_1325)
);

CKINVDCx11_ASAP7_75t_R g1326 ( 
.A(n_1147),
.Y(n_1326)
);

INVx4_ASAP7_75t_L g1327 ( 
.A(n_1221),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1109),
.A2(n_1221),
.B1(n_1116),
.B2(n_1204),
.Y(n_1328)
);

AOI21xp33_ASAP7_75t_L g1329 ( 
.A1(n_1209),
.A2(n_1214),
.B(n_1219),
.Y(n_1329)
);

INVxp67_ASAP7_75t_L g1330 ( 
.A(n_1239),
.Y(n_1330)
);

AOI22xp33_ASAP7_75t_L g1331 ( 
.A1(n_1142),
.A2(n_1230),
.B1(n_1200),
.B2(n_1218),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1142),
.Y(n_1332)
);

BUFx4f_ASAP7_75t_SL g1333 ( 
.A(n_1129),
.Y(n_1333)
);

AOI22xp33_ASAP7_75t_L g1334 ( 
.A1(n_1230),
.A2(n_1200),
.B1(n_1218),
.B2(n_1217),
.Y(n_1334)
);

AOI22xp33_ASAP7_75t_L g1335 ( 
.A1(n_1230),
.A2(n_1200),
.B1(n_1218),
.B2(n_1217),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1230),
.A2(n_1200),
.B1(n_1218),
.B2(n_1217),
.Y(n_1336)
);

AOI22xp33_ASAP7_75t_L g1337 ( 
.A1(n_1230),
.A2(n_1200),
.B1(n_1218),
.B2(n_1217),
.Y(n_1337)
);

BUFx3_ASAP7_75t_L g1338 ( 
.A(n_1103),
.Y(n_1338)
);

OAI22xp5_ASAP7_75t_L g1339 ( 
.A1(n_1193),
.A2(n_1228),
.B1(n_1217),
.B2(n_967),
.Y(n_1339)
);

OAI22xp5_ASAP7_75t_L g1340 ( 
.A1(n_1193),
.A2(n_1228),
.B1(n_1217),
.B2(n_967),
.Y(n_1340)
);

INVx1_ASAP7_75t_SL g1341 ( 
.A(n_1183),
.Y(n_1341)
);

CKINVDCx16_ASAP7_75t_R g1342 ( 
.A(n_1129),
.Y(n_1342)
);

AOI22xp33_ASAP7_75t_L g1343 ( 
.A1(n_1230),
.A2(n_1200),
.B1(n_1218),
.B2(n_1217),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_L g1344 ( 
.A1(n_1230),
.A2(n_1200),
.B1(n_1218),
.B2(n_1217),
.Y(n_1344)
);

INVx5_ASAP7_75t_L g1345 ( 
.A(n_1175),
.Y(n_1345)
);

OAI22xp5_ASAP7_75t_SL g1346 ( 
.A1(n_1218),
.A2(n_537),
.B1(n_559),
.B2(n_701),
.Y(n_1346)
);

BUFx6f_ASAP7_75t_L g1347 ( 
.A(n_1164),
.Y(n_1347)
);

INVx4_ASAP7_75t_L g1348 ( 
.A(n_1231),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1230),
.A2(n_1200),
.B1(n_1218),
.B2(n_1217),
.Y(n_1349)
);

OAI21xp5_ASAP7_75t_SL g1350 ( 
.A1(n_1193),
.A2(n_537),
.B(n_1217),
.Y(n_1350)
);

BUFx3_ASAP7_75t_L g1351 ( 
.A(n_1103),
.Y(n_1351)
);

AOI22xp33_ASAP7_75t_L g1352 ( 
.A1(n_1230),
.A2(n_1200),
.B1(n_1218),
.B2(n_1217),
.Y(n_1352)
);

BUFx3_ASAP7_75t_L g1353 ( 
.A(n_1103),
.Y(n_1353)
);

BUFx12f_ASAP7_75t_L g1354 ( 
.A(n_1236),
.Y(n_1354)
);

BUFx3_ASAP7_75t_L g1355 ( 
.A(n_1103),
.Y(n_1355)
);

INVx6_ASAP7_75t_L g1356 ( 
.A(n_1173),
.Y(n_1356)
);

OAI22xp33_ASAP7_75t_L g1357 ( 
.A1(n_1193),
.A2(n_1228),
.B1(n_1217),
.B2(n_1104),
.Y(n_1357)
);

AOI22xp33_ASAP7_75t_L g1358 ( 
.A1(n_1230),
.A2(n_1200),
.B1(n_1218),
.B2(n_1217),
.Y(n_1358)
);

NAND2x1p5_ASAP7_75t_L g1359 ( 
.A(n_1231),
.B(n_1046),
.Y(n_1359)
);

AOI22xp5_ASAP7_75t_L g1360 ( 
.A1(n_1193),
.A2(n_1228),
.B1(n_1217),
.B2(n_505),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1252),
.B(n_1268),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1252),
.B(n_1258),
.Y(n_1362)
);

AOI21x1_ASAP7_75t_L g1363 ( 
.A1(n_1313),
.A2(n_1325),
.B(n_1301),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1305),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1306),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1284),
.Y(n_1366)
);

CKINVDCx20_ASAP7_75t_R g1367 ( 
.A(n_1245),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1284),
.Y(n_1368)
);

OR2x2_ASAP7_75t_L g1369 ( 
.A(n_1324),
.B(n_1319),
.Y(n_1369)
);

HB1xp67_ASAP7_75t_L g1370 ( 
.A(n_1307),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1320),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1295),
.Y(n_1372)
);

AOI22xp33_ASAP7_75t_L g1373 ( 
.A1(n_1339),
.A2(n_1340),
.B1(n_1357),
.B2(n_1346),
.Y(n_1373)
);

OR2x2_ASAP7_75t_L g1374 ( 
.A(n_1259),
.B(n_1258),
.Y(n_1374)
);

OR2x6_ASAP7_75t_L g1375 ( 
.A(n_1294),
.B(n_1323),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1295),
.Y(n_1376)
);

HB1xp67_ASAP7_75t_L g1377 ( 
.A(n_1279),
.Y(n_1377)
);

HB1xp67_ASAP7_75t_L g1378 ( 
.A(n_1275),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1288),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1290),
.Y(n_1380)
);

NOR2xp33_ASAP7_75t_L g1381 ( 
.A(n_1261),
.B(n_1250),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1255),
.B(n_1331),
.Y(n_1382)
);

BUFx6f_ASAP7_75t_L g1383 ( 
.A(n_1345),
.Y(n_1383)
);

OA21x2_ASAP7_75t_L g1384 ( 
.A1(n_1315),
.A2(n_1302),
.B(n_1299),
.Y(n_1384)
);

OAI21x1_ASAP7_75t_L g1385 ( 
.A1(n_1315),
.A2(n_1302),
.B(n_1328),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1255),
.B(n_1331),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1242),
.B(n_1334),
.Y(n_1387)
);

BUFx3_ASAP7_75t_L g1388 ( 
.A(n_1249),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1327),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1332),
.Y(n_1390)
);

OR2x2_ASAP7_75t_L g1391 ( 
.A(n_1274),
.B(n_1357),
.Y(n_1391)
);

NOR2xp67_ASAP7_75t_SL g1392 ( 
.A(n_1350),
.B(n_1314),
.Y(n_1392)
);

HB1xp67_ASAP7_75t_L g1393 ( 
.A(n_1303),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1242),
.B(n_1334),
.Y(n_1394)
);

AOI21xp5_ASAP7_75t_L g1395 ( 
.A1(n_1318),
.A2(n_1321),
.B(n_1304),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1278),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1335),
.B(n_1336),
.Y(n_1397)
);

NAND3xp33_ASAP7_75t_L g1398 ( 
.A(n_1253),
.B(n_1360),
.C(n_1263),
.Y(n_1398)
);

OAI211xp5_ASAP7_75t_L g1399 ( 
.A1(n_1263),
.A2(n_1253),
.B(n_1358),
.C(n_1352),
.Y(n_1399)
);

OAI21x1_ASAP7_75t_L g1400 ( 
.A1(n_1328),
.A2(n_1322),
.B(n_1299),
.Y(n_1400)
);

AOI21x1_ASAP7_75t_L g1401 ( 
.A1(n_1277),
.A2(n_1282),
.B(n_1296),
.Y(n_1401)
);

BUFx2_ASAP7_75t_L g1402 ( 
.A(n_1285),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1326),
.Y(n_1403)
);

INVx4_ASAP7_75t_SL g1404 ( 
.A(n_1271),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_L g1405 ( 
.A1(n_1322),
.A2(n_1304),
.B(n_1269),
.Y(n_1405)
);

AND2x4_ASAP7_75t_L g1406 ( 
.A(n_1248),
.B(n_1297),
.Y(n_1406)
);

HB1xp67_ASAP7_75t_L g1407 ( 
.A(n_1287),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1330),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1317),
.Y(n_1409)
);

BUFx2_ASAP7_75t_L g1410 ( 
.A(n_1359),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1283),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1283),
.Y(n_1412)
);

AO31x2_ASAP7_75t_L g1413 ( 
.A1(n_1267),
.A2(n_1309),
.A3(n_1316),
.B(n_1352),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1269),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1272),
.B(n_1246),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1316),
.Y(n_1416)
);

INVx2_ASAP7_75t_SL g1417 ( 
.A(n_1273),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1309),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1280),
.Y(n_1419)
);

HB1xp67_ASAP7_75t_L g1420 ( 
.A(n_1287),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1308),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1335),
.Y(n_1422)
);

OAI21x1_ASAP7_75t_L g1423 ( 
.A1(n_1265),
.A2(n_1359),
.B(n_1358),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1336),
.B(n_1349),
.Y(n_1424)
);

INVx1_ASAP7_75t_SL g1425 ( 
.A(n_1341),
.Y(n_1425)
);

OAI22xp5_ASAP7_75t_L g1426 ( 
.A1(n_1337),
.A2(n_1349),
.B1(n_1344),
.B2(n_1343),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1337),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1343),
.Y(n_1428)
);

OAI21xp5_ASAP7_75t_L g1429 ( 
.A1(n_1344),
.A2(n_1265),
.B(n_1262),
.Y(n_1429)
);

INVx2_ASAP7_75t_SL g1430 ( 
.A(n_1312),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1298),
.B(n_1342),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1329),
.Y(n_1432)
);

AOI22xp33_ASAP7_75t_SL g1433 ( 
.A1(n_1257),
.A2(n_1356),
.B1(n_1333),
.B2(n_1260),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1293),
.B(n_1254),
.Y(n_1434)
);

AOI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1251),
.A2(n_1356),
.B1(n_1291),
.B2(n_1249),
.Y(n_1435)
);

OAI211xp5_ASAP7_75t_L g1436 ( 
.A1(n_1399),
.A2(n_1244),
.B(n_1276),
.C(n_1270),
.Y(n_1436)
);

OR2x2_ASAP7_75t_L g1437 ( 
.A(n_1416),
.B(n_1260),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1377),
.B(n_1333),
.Y(n_1438)
);

NAND4xp25_ASAP7_75t_L g1439 ( 
.A(n_1373),
.B(n_1398),
.C(n_1415),
.D(n_1429),
.Y(n_1439)
);

OA21x2_ASAP7_75t_L g1440 ( 
.A1(n_1400),
.A2(n_1300),
.B(n_1311),
.Y(n_1440)
);

OA21x2_ASAP7_75t_L g1441 ( 
.A1(n_1400),
.A2(n_1385),
.B(n_1405),
.Y(n_1441)
);

NAND3xp33_ASAP7_75t_L g1442 ( 
.A(n_1426),
.B(n_1312),
.C(n_1348),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1361),
.B(n_1292),
.Y(n_1443)
);

OAI21xp5_ASAP7_75t_L g1444 ( 
.A1(n_1395),
.A2(n_1353),
.B(n_1338),
.Y(n_1444)
);

NOR2xp33_ASAP7_75t_L g1445 ( 
.A(n_1381),
.B(n_1247),
.Y(n_1445)
);

CKINVDCx8_ASAP7_75t_R g1446 ( 
.A(n_1406),
.Y(n_1446)
);

NAND3xp33_ASAP7_75t_L g1447 ( 
.A(n_1392),
.B(n_1353),
.C(n_1338),
.Y(n_1447)
);

AOI221xp5_ASAP7_75t_L g1448 ( 
.A1(n_1362),
.A2(n_1251),
.B1(n_1264),
.B2(n_1355),
.C(n_1351),
.Y(n_1448)
);

OAI21xp5_ASAP7_75t_L g1449 ( 
.A1(n_1424),
.A2(n_1310),
.B(n_1266),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1378),
.B(n_1289),
.Y(n_1450)
);

OA21x2_ASAP7_75t_L g1451 ( 
.A1(n_1385),
.A2(n_1281),
.B(n_1286),
.Y(n_1451)
);

A2O1A1Ixp33_ASAP7_75t_L g1452 ( 
.A1(n_1362),
.A2(n_1286),
.B(n_1347),
.C(n_1356),
.Y(n_1452)
);

NOR2xp33_ASAP7_75t_SL g1453 ( 
.A(n_1367),
.B(n_1354),
.Y(n_1453)
);

O2A1O1Ixp33_ASAP7_75t_SL g1454 ( 
.A1(n_1430),
.A2(n_1243),
.B(n_1256),
.C(n_1347),
.Y(n_1454)
);

OAI22xp5_ASAP7_75t_L g1455 ( 
.A1(n_1409),
.A2(n_1243),
.B1(n_1347),
.B2(n_1407),
.Y(n_1455)
);

NOR2xp33_ASAP7_75t_L g1456 ( 
.A(n_1425),
.B(n_1434),
.Y(n_1456)
);

NAND2xp33_ASAP7_75t_L g1457 ( 
.A(n_1383),
.B(n_1387),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1379),
.B(n_1380),
.Y(n_1458)
);

OAI21xp5_ASAP7_75t_L g1459 ( 
.A1(n_1387),
.A2(n_1394),
.B(n_1397),
.Y(n_1459)
);

AOI221xp5_ASAP7_75t_L g1460 ( 
.A1(n_1394),
.A2(n_1397),
.B1(n_1427),
.B2(n_1428),
.C(n_1422),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1370),
.B(n_1374),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1364),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1364),
.Y(n_1463)
);

OR2x2_ASAP7_75t_L g1464 ( 
.A(n_1372),
.B(n_1376),
.Y(n_1464)
);

OAI22xp5_ASAP7_75t_L g1465 ( 
.A1(n_1409),
.A2(n_1420),
.B1(n_1433),
.B2(n_1403),
.Y(n_1465)
);

CKINVDCx20_ASAP7_75t_R g1466 ( 
.A(n_1388),
.Y(n_1466)
);

OAI21xp33_ASAP7_75t_SL g1467 ( 
.A1(n_1382),
.A2(n_1386),
.B(n_1423),
.Y(n_1467)
);

AO21x2_ASAP7_75t_L g1468 ( 
.A1(n_1432),
.A2(n_1363),
.B(n_1376),
.Y(n_1468)
);

OR2x2_ASAP7_75t_L g1469 ( 
.A(n_1366),
.B(n_1368),
.Y(n_1469)
);

AO21x2_ASAP7_75t_L g1470 ( 
.A1(n_1432),
.A2(n_1363),
.B(n_1405),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1390),
.B(n_1413),
.Y(n_1471)
);

O2A1O1Ixp33_ASAP7_75t_L g1472 ( 
.A1(n_1422),
.A2(n_1428),
.B(n_1427),
.C(n_1418),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1390),
.B(n_1413),
.Y(n_1473)
);

AND2x4_ASAP7_75t_L g1474 ( 
.A(n_1404),
.B(n_1411),
.Y(n_1474)
);

AND2x4_ASAP7_75t_L g1475 ( 
.A(n_1404),
.B(n_1411),
.Y(n_1475)
);

OR2x2_ASAP7_75t_L g1476 ( 
.A(n_1461),
.B(n_1366),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1471),
.B(n_1414),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1462),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1471),
.B(n_1412),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1473),
.B(n_1413),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1462),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1473),
.B(n_1412),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1463),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1443),
.B(n_1408),
.Y(n_1484)
);

AOI211x1_ASAP7_75t_SL g1485 ( 
.A1(n_1439),
.A2(n_1421),
.B(n_1431),
.C(n_1419),
.Y(n_1485)
);

AND2x4_ASAP7_75t_L g1486 ( 
.A(n_1474),
.B(n_1396),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1463),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1458),
.B(n_1413),
.Y(n_1488)
);

CKINVDCx16_ASAP7_75t_R g1489 ( 
.A(n_1453),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1469),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1469),
.Y(n_1491)
);

OR2x2_ASAP7_75t_L g1492 ( 
.A(n_1468),
.B(n_1368),
.Y(n_1492)
);

NOR2xp33_ASAP7_75t_L g1493 ( 
.A(n_1438),
.B(n_1403),
.Y(n_1493)
);

NOR2x1_ASAP7_75t_L g1494 ( 
.A(n_1447),
.B(n_1402),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1464),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1442),
.A2(n_1392),
.B1(n_1386),
.B2(n_1382),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1470),
.B(n_1391),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1470),
.B(n_1468),
.Y(n_1498)
);

AOI22xp33_ASAP7_75t_L g1499 ( 
.A1(n_1460),
.A2(n_1375),
.B1(n_1418),
.B2(n_1393),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1470),
.B(n_1391),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1468),
.B(n_1389),
.Y(n_1501)
);

INVx3_ASAP7_75t_L g1502 ( 
.A(n_1474),
.Y(n_1502)
);

NOR2xp33_ASAP7_75t_L g1503 ( 
.A(n_1445),
.B(n_1417),
.Y(n_1503)
);

AOI22xp5_ASAP7_75t_L g1504 ( 
.A1(n_1436),
.A2(n_1423),
.B1(n_1374),
.B2(n_1375),
.Y(n_1504)
);

AOI22xp33_ASAP7_75t_SL g1505 ( 
.A1(n_1457),
.A2(n_1402),
.B1(n_1375),
.B2(n_1410),
.Y(n_1505)
);

HB1xp67_ASAP7_75t_L g1506 ( 
.A(n_1487),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1479),
.B(n_1441),
.Y(n_1507)
);

INVx5_ASAP7_75t_L g1508 ( 
.A(n_1498),
.Y(n_1508)
);

OR2x2_ASAP7_75t_L g1509 ( 
.A(n_1488),
.B(n_1441),
.Y(n_1509)
);

AND2x4_ASAP7_75t_L g1510 ( 
.A(n_1502),
.B(n_1475),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1482),
.B(n_1440),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1495),
.B(n_1467),
.Y(n_1512)
);

NOR2xp33_ASAP7_75t_L g1513 ( 
.A(n_1489),
.B(n_1435),
.Y(n_1513)
);

NOR2x1_ASAP7_75t_L g1514 ( 
.A(n_1494),
.B(n_1457),
.Y(n_1514)
);

INVx1_ASAP7_75t_SL g1515 ( 
.A(n_1476),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1487),
.Y(n_1516)
);

OAI22xp5_ASAP7_75t_L g1517 ( 
.A1(n_1499),
.A2(n_1459),
.B1(n_1446),
.B2(n_1452),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1482),
.B(n_1440),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1478),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1495),
.B(n_1413),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1478),
.Y(n_1521)
);

INVxp67_ASAP7_75t_SL g1522 ( 
.A(n_1492),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1502),
.B(n_1440),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_SL g1524 ( 
.A(n_1489),
.B(n_1448),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1481),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1483),
.Y(n_1526)
);

AO21x2_ASAP7_75t_L g1527 ( 
.A1(n_1501),
.A2(n_1365),
.B(n_1371),
.Y(n_1527)
);

AOI22xp33_ASAP7_75t_SL g1528 ( 
.A1(n_1480),
.A2(n_1465),
.B1(n_1384),
.B2(n_1444),
.Y(n_1528)
);

BUFx2_ASAP7_75t_L g1529 ( 
.A(n_1494),
.Y(n_1529)
);

AND2x4_ASAP7_75t_L g1530 ( 
.A(n_1486),
.B(n_1475),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1497),
.B(n_1451),
.Y(n_1531)
);

OAI322xp33_ASAP7_75t_L g1532 ( 
.A1(n_1480),
.A2(n_1472),
.A3(n_1437),
.B1(n_1450),
.B2(n_1455),
.C1(n_1435),
.C2(n_1369),
.Y(n_1532)
);

OAI21xp5_ASAP7_75t_L g1533 ( 
.A1(n_1504),
.A2(n_1401),
.B(n_1449),
.Y(n_1533)
);

INVxp67_ASAP7_75t_SL g1534 ( 
.A(n_1514),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1527),
.Y(n_1535)
);

AND2x4_ASAP7_75t_L g1536 ( 
.A(n_1523),
.B(n_1501),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1519),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1519),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1521),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1511),
.B(n_1500),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1527),
.Y(n_1541)
);

OR2x2_ASAP7_75t_L g1542 ( 
.A(n_1509),
.B(n_1492),
.Y(n_1542)
);

NAND2x1_ASAP7_75t_SL g1543 ( 
.A(n_1514),
.B(n_1500),
.Y(n_1543)
);

BUFx3_ASAP7_75t_L g1544 ( 
.A(n_1529),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1515),
.B(n_1512),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1527),
.Y(n_1546)
);

HB1xp67_ASAP7_75t_L g1547 ( 
.A(n_1506),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1518),
.B(n_1531),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1527),
.Y(n_1549)
);

NOR2xp33_ASAP7_75t_L g1550 ( 
.A(n_1524),
.B(n_1493),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1518),
.B(n_1531),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1516),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1512),
.B(n_1490),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1516),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1518),
.B(n_1484),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1525),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1529),
.B(n_1491),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1531),
.B(n_1484),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1525),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1522),
.B(n_1491),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1522),
.B(n_1477),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1526),
.Y(n_1562)
);

OR2x2_ASAP7_75t_L g1563 ( 
.A(n_1509),
.B(n_1477),
.Y(n_1563)
);

CKINVDCx14_ASAP7_75t_R g1564 ( 
.A(n_1550),
.Y(n_1564)
);

OR2x2_ASAP7_75t_L g1565 ( 
.A(n_1545),
.B(n_1509),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1537),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1553),
.B(n_1507),
.Y(n_1567)
);

OR2x2_ASAP7_75t_L g1568 ( 
.A(n_1545),
.B(n_1520),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1537),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1538),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1538),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_1552),
.Y(n_1572)
);

OR2x6_ASAP7_75t_L g1573 ( 
.A(n_1544),
.B(n_1533),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1534),
.B(n_1510),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1539),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1534),
.B(n_1510),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1555),
.B(n_1510),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1539),
.Y(n_1578)
);

OR2x6_ASAP7_75t_L g1579 ( 
.A(n_1544),
.B(n_1533),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_1552),
.Y(n_1580)
);

INVx2_ASAP7_75t_SL g1581 ( 
.A(n_1543),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1552),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1553),
.B(n_1507),
.Y(n_1583)
);

INVxp67_ASAP7_75t_SL g1584 ( 
.A(n_1543),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1558),
.B(n_1530),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1552),
.Y(n_1586)
);

AND2x4_ASAP7_75t_L g1587 ( 
.A(n_1544),
.B(n_1530),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1554),
.Y(n_1588)
);

CKINVDCx5p33_ASAP7_75t_R g1589 ( 
.A(n_1550),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1556),
.Y(n_1590)
);

INVx1_ASAP7_75t_SL g1591 ( 
.A(n_1544),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1554),
.Y(n_1592)
);

NAND3xp33_ASAP7_75t_L g1593 ( 
.A(n_1542),
.B(n_1528),
.C(n_1517),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1556),
.B(n_1507),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1558),
.B(n_1548),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1559),
.Y(n_1596)
);

INVxp67_ASAP7_75t_L g1597 ( 
.A(n_1547),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1558),
.B(n_1530),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1559),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1562),
.Y(n_1600)
);

NOR2xp67_ASAP7_75t_L g1601 ( 
.A(n_1547),
.B(n_1508),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1564),
.B(n_1589),
.Y(n_1602)
);

AND2x2_ASAP7_75t_SL g1603 ( 
.A(n_1587),
.B(n_1513),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1572),
.Y(n_1604)
);

INVx1_ASAP7_75t_SL g1605 ( 
.A(n_1591),
.Y(n_1605)
);

NOR2xp33_ASAP7_75t_L g1606 ( 
.A(n_1593),
.B(n_1466),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1574),
.B(n_1540),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1593),
.B(n_1561),
.Y(n_1608)
);

NOR2xp33_ASAP7_75t_L g1609 ( 
.A(n_1573),
.B(n_1466),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1566),
.Y(n_1610)
);

OAI31xp33_ASAP7_75t_L g1611 ( 
.A1(n_1581),
.A2(n_1517),
.A3(n_1496),
.B(n_1454),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1574),
.B(n_1540),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_SL g1613 ( 
.A(n_1587),
.B(n_1528),
.Y(n_1613)
);

INVx1_ASAP7_75t_SL g1614 ( 
.A(n_1591),
.Y(n_1614)
);

AND2x4_ASAP7_75t_L g1615 ( 
.A(n_1601),
.B(n_1508),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1572),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1597),
.B(n_1557),
.Y(n_1617)
);

OR2x2_ASAP7_75t_L g1618 ( 
.A(n_1568),
.B(n_1565),
.Y(n_1618)
);

OR2x2_ASAP7_75t_L g1619 ( 
.A(n_1568),
.B(n_1563),
.Y(n_1619)
);

INVx2_ASAP7_75t_SL g1620 ( 
.A(n_1587),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1566),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1572),
.Y(n_1622)
);

AND2x4_ASAP7_75t_L g1623 ( 
.A(n_1601),
.B(n_1508),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1597),
.B(n_1557),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1569),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1569),
.Y(n_1626)
);

NOR2xp33_ASAP7_75t_L g1627 ( 
.A(n_1573),
.B(n_1388),
.Y(n_1627)
);

OR2x2_ASAP7_75t_L g1628 ( 
.A(n_1565),
.B(n_1563),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1576),
.B(n_1540),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1570),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1576),
.B(n_1548),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1570),
.Y(n_1632)
);

INVx3_ASAP7_75t_L g1633 ( 
.A(n_1581),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1587),
.B(n_1548),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1580),
.Y(n_1635)
);

OR2x2_ASAP7_75t_L g1636 ( 
.A(n_1567),
.B(n_1563),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1610),
.Y(n_1637)
);

OAI21xp33_ASAP7_75t_L g1638 ( 
.A1(n_1608),
.A2(n_1579),
.B(n_1573),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1610),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1603),
.B(n_1585),
.Y(n_1640)
);

NOR2xp33_ASAP7_75t_SL g1641 ( 
.A(n_1603),
.B(n_1532),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1633),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1606),
.B(n_1595),
.Y(n_1643)
);

NOR2x1_ASAP7_75t_L g1644 ( 
.A(n_1602),
.B(n_1573),
.Y(n_1644)
);

OR2x2_ASAP7_75t_L g1645 ( 
.A(n_1605),
.B(n_1567),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1633),
.Y(n_1646)
);

NAND3xp33_ASAP7_75t_L g1647 ( 
.A(n_1611),
.B(n_1579),
.C(n_1573),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1621),
.Y(n_1648)
);

AOI32xp33_ASAP7_75t_L g1649 ( 
.A1(n_1609),
.A2(n_1584),
.A3(n_1581),
.B1(n_1595),
.B2(n_1585),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1621),
.Y(n_1650)
);

NOR3xp33_ASAP7_75t_L g1651 ( 
.A(n_1613),
.B(n_1614),
.C(n_1605),
.Y(n_1651)
);

INVxp67_ASAP7_75t_L g1652 ( 
.A(n_1614),
.Y(n_1652)
);

AOI22xp5_ASAP7_75t_L g1653 ( 
.A1(n_1603),
.A2(n_1579),
.B1(n_1505),
.B2(n_1504),
.Y(n_1653)
);

OR2x2_ASAP7_75t_L g1654 ( 
.A(n_1617),
.B(n_1583),
.Y(n_1654)
);

INVx2_ASAP7_75t_SL g1655 ( 
.A(n_1633),
.Y(n_1655)
);

AOI21xp33_ASAP7_75t_L g1656 ( 
.A1(n_1611),
.A2(n_1579),
.B(n_1575),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1625),
.Y(n_1657)
);

INVxp67_ASAP7_75t_SL g1658 ( 
.A(n_1633),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1625),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1634),
.B(n_1598),
.Y(n_1660)
);

OAI21xp33_ASAP7_75t_L g1661 ( 
.A1(n_1627),
.A2(n_1579),
.B(n_1543),
.Y(n_1661)
);

AOI222xp33_ASAP7_75t_L g1662 ( 
.A1(n_1641),
.A2(n_1624),
.B1(n_1617),
.B2(n_1631),
.C1(n_1607),
.C2(n_1612),
.Y(n_1662)
);

INVxp67_ASAP7_75t_L g1663 ( 
.A(n_1658),
.Y(n_1663)
);

NAND3x2_ASAP7_75t_L g1664 ( 
.A(n_1640),
.B(n_1618),
.C(n_1628),
.Y(n_1664)
);

HB1xp67_ASAP7_75t_L g1665 ( 
.A(n_1652),
.Y(n_1665)
);

OAI211xp5_ASAP7_75t_L g1666 ( 
.A1(n_1651),
.A2(n_1624),
.B(n_1620),
.C(n_1630),
.Y(n_1666)
);

NOR2xp33_ASAP7_75t_SL g1667 ( 
.A(n_1644),
.B(n_1532),
.Y(n_1667)
);

NOR2xp33_ASAP7_75t_L g1668 ( 
.A(n_1652),
.B(n_1620),
.Y(n_1668)
);

BUFx2_ASAP7_75t_SL g1669 ( 
.A(n_1655),
.Y(n_1669)
);

AOI211x1_ASAP7_75t_SL g1670 ( 
.A1(n_1656),
.A2(n_1622),
.B(n_1635),
.C(n_1616),
.Y(n_1670)
);

OAI22xp5_ASAP7_75t_L g1671 ( 
.A1(n_1647),
.A2(n_1631),
.B1(n_1607),
.B2(n_1612),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1655),
.Y(n_1672)
);

AOI322xp5_ASAP7_75t_L g1673 ( 
.A1(n_1651),
.A2(n_1629),
.A3(n_1634),
.B1(n_1551),
.B2(n_1583),
.C1(n_1536),
.C2(n_1630),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1643),
.B(n_1629),
.Y(n_1674)
);

OAI32xp33_ASAP7_75t_L g1675 ( 
.A1(n_1638),
.A2(n_1618),
.A3(n_1619),
.B1(n_1628),
.B2(n_1636),
.Y(n_1675)
);

OAI21xp5_ASAP7_75t_L g1676 ( 
.A1(n_1653),
.A2(n_1623),
.B(n_1615),
.Y(n_1676)
);

AOI22xp5_ASAP7_75t_L g1677 ( 
.A1(n_1661),
.A2(n_1615),
.B1(n_1623),
.B2(n_1632),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_1660),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1658),
.Y(n_1679)
);

NOR2x1_ASAP7_75t_L g1680 ( 
.A(n_1642),
.B(n_1626),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1680),
.Y(n_1681)
);

AOI222xp33_ASAP7_75t_L g1682 ( 
.A1(n_1665),
.A2(n_1659),
.B1(n_1657),
.B2(n_1637),
.C1(n_1650),
.C2(n_1639),
.Y(n_1682)
);

AOI322xp5_ASAP7_75t_L g1683 ( 
.A1(n_1665),
.A2(n_1648),
.A3(n_1642),
.B1(n_1646),
.B2(n_1551),
.C1(n_1626),
.C2(n_1632),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1668),
.B(n_1649),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1668),
.B(n_1645),
.Y(n_1685)
);

HB1xp67_ASAP7_75t_L g1686 ( 
.A(n_1663),
.Y(n_1686)
);

OR2x2_ASAP7_75t_L g1687 ( 
.A(n_1664),
.B(n_1654),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1663),
.Y(n_1688)
);

AOI21xp33_ASAP7_75t_SL g1689 ( 
.A1(n_1671),
.A2(n_1646),
.B(n_1623),
.Y(n_1689)
);

OAI222xp33_ASAP7_75t_L g1690 ( 
.A1(n_1677),
.A2(n_1619),
.B1(n_1636),
.B2(n_1623),
.C1(n_1615),
.C2(n_1508),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1686),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1688),
.B(n_1678),
.Y(n_1692)
);

NOR2x1_ASAP7_75t_L g1693 ( 
.A(n_1681),
.B(n_1679),
.Y(n_1693)
);

AOI22xp33_ASAP7_75t_L g1694 ( 
.A1(n_1684),
.A2(n_1667),
.B1(n_1662),
.B2(n_1676),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1685),
.B(n_1672),
.Y(n_1695)
);

NOR4xp25_ASAP7_75t_L g1696 ( 
.A(n_1687),
.B(n_1666),
.C(n_1674),
.D(n_1670),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1682),
.Y(n_1697)
);

NOR3x1_ASAP7_75t_L g1698 ( 
.A(n_1689),
.B(n_1430),
.C(n_1675),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1682),
.Y(n_1699)
);

AOI222xp33_ASAP7_75t_L g1700 ( 
.A1(n_1697),
.A2(n_1690),
.B1(n_1673),
.B2(n_1683),
.C1(n_1615),
.C2(n_1669),
.Y(n_1700)
);

AOI221xp5_ASAP7_75t_L g1701 ( 
.A1(n_1696),
.A2(n_1635),
.B1(n_1622),
.B2(n_1616),
.C(n_1604),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1694),
.B(n_1598),
.Y(n_1702)
);

AOI321xp33_ASAP7_75t_L g1703 ( 
.A1(n_1694),
.A2(n_1635),
.A3(n_1622),
.B1(n_1616),
.B2(n_1604),
.C(n_1456),
.Y(n_1703)
);

OAI21xp5_ASAP7_75t_SL g1704 ( 
.A1(n_1699),
.A2(n_1503),
.B(n_1485),
.Y(n_1704)
);

OAI22xp5_ASAP7_75t_L g1705 ( 
.A1(n_1702),
.A2(n_1695),
.B1(n_1691),
.B2(n_1692),
.Y(n_1705)
);

NAND4xp25_ASAP7_75t_L g1706 ( 
.A(n_1703),
.B(n_1698),
.C(n_1693),
.D(n_1604),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1700),
.B(n_1577),
.Y(n_1707)
);

AOI221xp5_ASAP7_75t_L g1708 ( 
.A1(n_1704),
.A2(n_1535),
.B1(n_1549),
.B2(n_1546),
.C(n_1541),
.Y(n_1708)
);

AOI211xp5_ASAP7_75t_L g1709 ( 
.A1(n_1701),
.A2(n_1600),
.B(n_1599),
.C(n_1596),
.Y(n_1709)
);

NAND3xp33_ASAP7_75t_SL g1710 ( 
.A(n_1703),
.B(n_1485),
.C(n_1542),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1705),
.B(n_1577),
.Y(n_1711)
);

NOR2xp67_ASAP7_75t_L g1712 ( 
.A(n_1706),
.B(n_1571),
.Y(n_1712)
);

NOR4xp75_ASAP7_75t_L g1713 ( 
.A(n_1707),
.B(n_1594),
.C(n_1561),
.D(n_1560),
.Y(n_1713)
);

NOR2x1_ASAP7_75t_L g1714 ( 
.A(n_1710),
.B(n_1571),
.Y(n_1714)
);

OR2x2_ASAP7_75t_L g1715 ( 
.A(n_1709),
.B(n_1594),
.Y(n_1715)
);

INVxp67_ASAP7_75t_L g1716 ( 
.A(n_1711),
.Y(n_1716)
);

AOI21xp33_ASAP7_75t_SL g1717 ( 
.A1(n_1715),
.A2(n_1578),
.B(n_1575),
.Y(n_1717)
);

NOR2x1_ASAP7_75t_L g1718 ( 
.A(n_1712),
.B(n_1714),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1718),
.Y(n_1719)
);

AOI22xp5_ASAP7_75t_SL g1720 ( 
.A1(n_1719),
.A2(n_1716),
.B1(n_1713),
.B2(n_1717),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1720),
.B(n_1708),
.Y(n_1721)
);

OAI22xp5_ASAP7_75t_L g1722 ( 
.A1(n_1720),
.A2(n_1580),
.B1(n_1582),
.B2(n_1586),
.Y(n_1722)
);

XNOR2xp5_ASAP7_75t_L g1723 ( 
.A(n_1721),
.B(n_1406),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1722),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_SL g1725 ( 
.A(n_1723),
.B(n_1580),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1724),
.Y(n_1726)
);

AOI22xp33_ASAP7_75t_L g1727 ( 
.A1(n_1726),
.A2(n_1582),
.B1(n_1586),
.B2(n_1588),
.Y(n_1727)
);

AOI21xp5_ASAP7_75t_L g1728 ( 
.A1(n_1727),
.A2(n_1725),
.B(n_1586),
.Y(n_1728)
);

OAI21x1_ASAP7_75t_SL g1729 ( 
.A1(n_1728),
.A2(n_1588),
.B(n_1582),
.Y(n_1729)
);

OAI221xp5_ASAP7_75t_R g1730 ( 
.A1(n_1729),
.A2(n_1588),
.B1(n_1592),
.B2(n_1596),
.C(n_1599),
.Y(n_1730)
);

AOI211xp5_ASAP7_75t_L g1731 ( 
.A1(n_1730),
.A2(n_1592),
.B(n_1600),
.C(n_1590),
.Y(n_1731)
);


endmodule