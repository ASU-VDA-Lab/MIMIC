module fake_jpeg_1829_n_635 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_635);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_635;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

OR2x2_ASAP7_75t_L g20 ( 
.A(n_15),
.B(n_7),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_17),
.B(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_3),
.B(n_11),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_17),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_19),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_12),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_12),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_10),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_6),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_7),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_26),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_58),
.B(n_61),
.Y(n_140)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g135 ( 
.A(n_59),
.Y(n_135)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_60),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_21),
.B(n_19),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_62),
.Y(n_132)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_63),
.Y(n_165)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_64),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_21),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_65),
.B(n_67),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g179 ( 
.A(n_66),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_32),
.B(n_0),
.Y(n_67)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g184 ( 
.A(n_68),
.Y(n_184)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g207 ( 
.A(n_69),
.Y(n_207)
);

BUFx4f_ASAP7_75t_SL g70 ( 
.A(n_47),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_70),
.Y(n_188)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_71),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_54),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_72),
.B(n_76),
.Y(n_154)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_33),
.Y(n_73)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_73),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_74),
.Y(n_156)
);

INVx6_ASAP7_75t_SL g75 ( 
.A(n_56),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g194 ( 
.A(n_75),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_32),
.B(n_0),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_25),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_77),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_54),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_78),
.B(n_79),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_29),
.Y(n_79)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

INVx5_ASAP7_75t_L g195 ( 
.A(n_80),
.Y(n_195)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

INVx5_ASAP7_75t_L g225 ( 
.A(n_81),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_82),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_83),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_26),
.B(n_0),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_84),
.B(n_97),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_85),
.Y(n_150)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_86),
.Y(n_147)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_87),
.Y(n_171)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_88),
.Y(n_186)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_89),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_45),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_90),
.Y(n_205)
);

INVx11_ASAP7_75t_SL g91 ( 
.A(n_24),
.Y(n_91)
);

INVx8_ASAP7_75t_L g185 ( 
.A(n_91),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_92),
.Y(n_224)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_93),
.Y(n_200)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_94),
.Y(n_133)
);

BUFx12f_ASAP7_75t_SL g95 ( 
.A(n_43),
.Y(n_95)
);

OR2x4_ASAP7_75t_L g148 ( 
.A(n_95),
.B(n_91),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_20),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_96),
.A2(n_37),
.B1(n_36),
.B2(n_34),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_54),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_48),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_98),
.B(n_100),
.Y(n_192)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_40),
.Y(n_99)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_99),
.Y(n_142)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_40),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_48),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_101),
.B(n_107),
.Y(n_198)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_47),
.Y(n_102)
);

INVx8_ASAP7_75t_L g191 ( 
.A(n_102),
.Y(n_191)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_40),
.Y(n_103)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_103),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_20),
.B(n_1),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_104),
.B(n_119),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_53),
.Y(n_105)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_105),
.Y(n_134)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_38),
.Y(n_106)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_106),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_22),
.B(n_2),
.Y(n_107)
);

INVx6_ASAP7_75t_SL g108 ( 
.A(n_29),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g223 ( 
.A(n_108),
.Y(n_223)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_47),
.Y(n_109)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_109),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_35),
.B(n_2),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_110),
.B(n_116),
.Y(n_216)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_43),
.Y(n_111)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_111),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_53),
.Y(n_112)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_112),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_53),
.Y(n_113)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_113),
.Y(n_160)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_57),
.Y(n_114)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_114),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_28),
.Y(n_115)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_115),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_48),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_28),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_117),
.B(n_126),
.Y(n_219)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_43),
.Y(n_118)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_118),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_20),
.B(n_5),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g120 ( 
.A(n_47),
.Y(n_120)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_120),
.Y(n_174)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_57),
.Y(n_121)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_121),
.Y(n_217)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_28),
.Y(n_122)
);

INVx3_ASAP7_75t_SL g170 ( 
.A(n_122),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_39),
.Y(n_123)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_123),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_30),
.B(n_5),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_124),
.B(n_130),
.Y(n_145)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_43),
.Y(n_125)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_125),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_39),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_39),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_127),
.B(n_128),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_42),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_42),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_129),
.B(n_35),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_42),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g136 ( 
.A(n_75),
.Y(n_136)
);

BUFx5_ASAP7_75t_L g247 ( 
.A(n_136),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_108),
.A2(n_27),
.B1(n_49),
.B2(n_30),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_138),
.A2(n_141),
.B1(n_169),
.B2(n_175),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_95),
.A2(n_27),
.B1(n_49),
.B2(n_30),
.Y(n_141)
);

OR2x4_ASAP7_75t_L g249 ( 
.A(n_148),
.B(n_70),
.Y(n_249)
);

AOI21xp33_ASAP7_75t_L g149 ( 
.A1(n_104),
.A2(n_22),
.B(n_44),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_149),
.B(n_204),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_152),
.B(n_15),
.Y(n_274)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_86),
.Y(n_158)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_158),
.Y(n_258)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_87),
.Y(n_161)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_161),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_58),
.A2(n_44),
.B1(n_24),
.B2(n_52),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g229 ( 
.A(n_162),
.B(n_172),
.Y(n_229)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_88),
.Y(n_163)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_163),
.Y(n_265)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_62),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_167),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_130),
.A2(n_49),
.B1(n_27),
.B2(n_52),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_119),
.A2(n_51),
.B1(n_23),
.B2(n_41),
.Y(n_172)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_100),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_173),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_124),
.A2(n_51),
.B1(n_23),
.B2(n_41),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_93),
.Y(n_176)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_176),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_177),
.A2(n_183),
.B1(n_193),
.B2(n_70),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_106),
.A2(n_37),
.B1(n_36),
.B2(n_34),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_180),
.A2(n_120),
.B1(n_7),
.B2(n_8),
.Y(n_252)
);

INVx3_ASAP7_75t_SL g181 ( 
.A(n_59),
.Y(n_181)
);

BUFx2_ASAP7_75t_L g228 ( 
.A(n_181),
.Y(n_228)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_73),
.Y(n_182)
);

INVx4_ASAP7_75t_L g254 ( 
.A(n_182),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_96),
.A2(n_29),
.B1(n_38),
.B2(n_47),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_122),
.A2(n_71),
.B1(n_123),
.B2(n_115),
.Y(n_193)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_64),
.Y(n_196)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_196),
.Y(n_256)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_66),
.Y(n_197)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_197),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_60),
.B(n_38),
.C(n_6),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_202),
.B(n_118),
.C(n_112),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_114),
.B(n_121),
.Y(n_204)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_99),
.Y(n_206)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_206),
.Y(n_296)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_102),
.Y(n_208)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_208),
.Y(n_277)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_103),
.Y(n_209)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_209),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_94),
.B(n_5),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_210),
.B(n_6),
.Y(n_253)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_102),
.Y(n_211)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_211),
.Y(n_281)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_74),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_212),
.Y(n_291)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_109),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g305 ( 
.A(n_213),
.Y(n_305)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_111),
.Y(n_214)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_214),
.Y(n_300)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_69),
.Y(n_215)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_215),
.Y(n_237)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_89),
.Y(n_218)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_218),
.Y(n_250)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_63),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_220),
.Y(n_243)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_109),
.Y(n_221)
);

INVx5_ASAP7_75t_L g266 ( 
.A(n_221),
.Y(n_266)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_68),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_227),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_145),
.B(n_192),
.Y(n_231)
);

CKINVDCx14_ASAP7_75t_R g316 ( 
.A(n_231),
.Y(n_316)
);

XNOR2x1_ASAP7_75t_L g355 ( 
.A(n_233),
.B(n_282),
.Y(n_355)
);

OAI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_175),
.A2(n_198),
.B1(n_216),
.B2(n_190),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_L g367 ( 
.A1(n_234),
.A2(n_270),
.B1(n_260),
.B2(n_262),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_192),
.B(n_125),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g318 ( 
.A(n_235),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_168),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_236),
.B(n_238),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_219),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_239),
.A2(n_242),
.B1(n_245),
.B2(n_311),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_203),
.A2(n_85),
.B1(n_82),
.B2(n_105),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_240),
.A2(n_272),
.B1(n_132),
.B2(n_199),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_219),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_241),
.B(n_244),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_198),
.A2(n_92),
.B1(n_90),
.B2(n_83),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_222),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_190),
.A2(n_77),
.B1(n_113),
.B2(n_80),
.Y(n_245)
);

INVx11_ASAP7_75t_L g248 ( 
.A(n_223),
.Y(n_248)
);

INVx4_ASAP7_75t_L g365 ( 
.A(n_248),
.Y(n_365)
);

OR2x2_ASAP7_75t_L g336 ( 
.A(n_249),
.B(n_267),
.Y(n_336)
);

O2A1O1Ixp33_ASAP7_75t_L g251 ( 
.A1(n_141),
.A2(n_81),
.B(n_120),
.C(n_8),
.Y(n_251)
);

OA22x2_ASAP7_75t_L g349 ( 
.A1(n_251),
.A2(n_199),
.B1(n_308),
.B2(n_245),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_252),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_253),
.B(n_137),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_203),
.B(n_216),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_255),
.B(n_261),
.Y(n_315)
);

AND2x2_ASAP7_75t_SL g257 ( 
.A(n_147),
.B(n_8),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_257),
.Y(n_323)
);

AND2x2_ASAP7_75t_SL g259 ( 
.A(n_171),
.B(n_8),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_259),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_140),
.B(n_9),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_260),
.B(n_187),
.C(n_160),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_154),
.B(n_9),
.Y(n_261)
);

CKINVDCx6p67_ASAP7_75t_R g262 ( 
.A(n_223),
.Y(n_262)
);

INVx5_ASAP7_75t_SL g337 ( 
.A(n_262),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_154),
.B(n_10),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_264),
.B(n_269),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_140),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_186),
.B(n_11),
.Y(n_269)
);

OAI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_180),
.A2(n_11),
.B1(n_12),
.B2(n_14),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_169),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_200),
.B(n_14),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_273),
.B(n_280),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_274),
.B(n_276),
.Y(n_338)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_222),
.Y(n_275)
);

HB1xp67_ASAP7_75t_L g341 ( 
.A(n_275),
.Y(n_341)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_168),
.Y(n_276)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_201),
.Y(n_279)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_279),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_217),
.B(n_15),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_207),
.B(n_139),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_153),
.B(n_194),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_283),
.B(n_286),
.Y(n_343)
);

AOI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_153),
.A2(n_151),
.B1(n_207),
.B2(n_179),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_284),
.A2(n_225),
.B1(n_195),
.B2(n_164),
.Y(n_320)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_142),
.Y(n_285)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_285),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_178),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_155),
.B(n_144),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_287),
.B(n_293),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_135),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_288),
.B(n_289),
.Y(n_348)
);

CKINVDCx14_ASAP7_75t_R g289 ( 
.A(n_179),
.Y(n_289)
);

INVx8_ASAP7_75t_L g292 ( 
.A(n_194),
.Y(n_292)
);

INVx3_ASAP7_75t_SL g333 ( 
.A(n_292),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_131),
.B(n_133),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_166),
.Y(n_294)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_294),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_188),
.B(n_185),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_295),
.B(n_302),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_146),
.B(n_170),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_298),
.B(n_304),
.Y(n_362)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_181),
.Y(n_299)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_299),
.Y(n_334)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_170),
.Y(n_301)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_301),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_189),
.B(n_174),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_143),
.B(n_184),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g335 ( 
.A(n_303),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_178),
.B(n_184),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_135),
.B(n_165),
.Y(n_306)
);

AND2x2_ASAP7_75t_SL g328 ( 
.A(n_306),
.B(n_156),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_165),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_307),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_138),
.Y(n_308)
);

BUFx2_ASAP7_75t_L g352 ( 
.A(n_308),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_191),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_309),
.Y(n_364)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_159),
.Y(n_310)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_310),
.Y(n_346)
);

AOI22xp33_ASAP7_75t_L g311 ( 
.A1(n_150),
.A2(n_224),
.B1(n_205),
.B2(n_226),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g373 ( 
.A(n_312),
.B(n_282),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_314),
.A2(n_332),
.B1(n_351),
.B2(n_361),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_246),
.A2(n_146),
.B1(n_226),
.B2(n_132),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_317),
.A2(n_363),
.B1(n_296),
.B2(n_228),
.Y(n_387)
);

INVx13_ASAP7_75t_L g319 ( 
.A(n_262),
.Y(n_319)
);

INVx1_ASAP7_75t_SL g395 ( 
.A(n_319),
.Y(n_395)
);

OAI21xp33_ASAP7_75t_L g375 ( 
.A1(n_320),
.A2(n_340),
.B(n_369),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_324),
.B(n_358),
.Y(n_389)
);

INVx5_ASAP7_75t_L g325 ( 
.A(n_292),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_325),
.Y(n_401)
);

CKINVDCx16_ASAP7_75t_R g411 ( 
.A(n_328),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_239),
.A2(n_134),
.B1(n_156),
.B2(n_157),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g340 ( 
.A(n_235),
.B(n_249),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_231),
.B(n_157),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_342),
.B(n_344),
.C(n_306),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_231),
.B(n_255),
.C(n_233),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_299),
.Y(n_345)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_345),
.Y(n_390)
);

AOI21xp33_ASAP7_75t_L g407 ( 
.A1(n_349),
.A2(n_230),
.B(n_330),
.Y(n_407)
);

INVx3_ASAP7_75t_L g350 ( 
.A(n_262),
.Y(n_350)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_350),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_242),
.A2(n_229),
.B1(n_269),
.B2(n_273),
.Y(n_351)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_293),
.Y(n_356)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_356),
.Y(n_403)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_287),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_228),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_359),
.B(n_368),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_229),
.A2(n_280),
.B1(n_290),
.B2(n_261),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_240),
.A2(n_272),
.B1(n_235),
.B2(n_298),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_257),
.A2(n_259),
.B1(n_267),
.B2(n_264),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_366),
.A2(n_271),
.B1(n_243),
.B2(n_278),
.Y(n_391)
);

OAI22xp33_ASAP7_75t_SL g398 ( 
.A1(n_367),
.A2(n_277),
.B1(n_281),
.B2(n_256),
.Y(n_398)
);

INVx4_ASAP7_75t_L g368 ( 
.A(n_248),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_282),
.B(n_306),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_258),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_370),
.B(n_334),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_363),
.A2(n_257),
.B1(n_259),
.B2(n_232),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_371),
.A2(n_372),
.B1(n_382),
.B2(n_383),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_356),
.A2(n_291),
.B1(n_232),
.B2(n_251),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_373),
.Y(n_429)
);

AOI22xp33_ASAP7_75t_L g376 ( 
.A1(n_322),
.A2(n_268),
.B1(n_265),
.B2(n_263),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_376),
.A2(n_404),
.B1(n_406),
.B2(n_334),
.Y(n_436)
);

OA22x2_ASAP7_75t_L g377 ( 
.A1(n_314),
.A2(n_268),
.B1(n_265),
.B2(n_263),
.Y(n_377)
);

AO21x2_ASAP7_75t_L g444 ( 
.A1(n_377),
.A2(n_321),
.B(n_345),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_326),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_378),
.B(n_381),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_379),
.B(n_386),
.C(n_400),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_325),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_358),
.A2(n_291),
.B1(n_258),
.B2(n_285),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_316),
.A2(n_297),
.B1(n_296),
.B2(n_271),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_357),
.B(n_300),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_384),
.B(n_392),
.Y(n_426)
);

NOR4xp25_ASAP7_75t_L g385 ( 
.A(n_315),
.B(n_237),
.C(n_250),
.D(n_278),
.Y(n_385)
);

MAJx2_ASAP7_75t_L g438 ( 
.A(n_385),
.B(n_328),
.C(n_364),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_344),
.B(n_300),
.C(n_297),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_387),
.A2(n_398),
.B1(n_383),
.B2(n_411),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g388 ( 
.A1(n_340),
.A2(n_309),
.B(n_243),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g418 ( 
.A1(n_388),
.A2(n_407),
.B(n_369),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_391),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_357),
.B(n_254),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_360),
.B(n_254),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_394),
.B(n_414),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_335),
.B(n_230),
.Y(n_396)
);

CKINVDCx14_ASAP7_75t_R g441 ( 
.A(n_396),
.Y(n_441)
);

AO21x1_ASAP7_75t_L g397 ( 
.A1(n_340),
.A2(n_305),
.B(n_247),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_SL g430 ( 
.A1(n_397),
.A2(n_410),
.B(n_347),
.Y(n_430)
);

INVx6_ASAP7_75t_L g399 ( 
.A(n_337),
.Y(n_399)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_399),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_355),
.B(n_277),
.C(n_281),
.Y(n_400)
);

AND2x6_ASAP7_75t_L g402 ( 
.A(n_355),
.B(n_247),
.Y(n_402)
);

AND2x6_ASAP7_75t_L g427 ( 
.A(n_402),
.B(n_349),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_317),
.A2(n_360),
.B1(n_362),
.B2(n_336),
.Y(n_404)
);

NOR2x1_ASAP7_75t_L g405 ( 
.A(n_343),
.B(n_266),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_SL g421 ( 
.A(n_405),
.B(n_415),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_362),
.A2(n_256),
.B1(n_266),
.B2(n_305),
.Y(n_406)
);

INVx6_ASAP7_75t_L g408 ( 
.A(n_337),
.Y(n_408)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_408),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_SL g409 ( 
.A(n_315),
.B(n_338),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_409),
.B(n_346),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_L g410 ( 
.A1(n_336),
.A2(n_318),
.B(n_323),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_342),
.B(n_324),
.C(n_331),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_412),
.B(n_416),
.C(n_312),
.Y(n_437)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_413),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_353),
.B(n_366),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_341),
.B(n_353),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_329),
.B(n_354),
.C(n_369),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_SL g463 ( 
.A1(n_418),
.A2(n_428),
.B(n_430),
.Y(n_463)
);

INVx1_ASAP7_75t_SL g419 ( 
.A(n_397),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_419),
.B(n_391),
.Y(n_458)
);

CKINVDCx16_ASAP7_75t_R g423 ( 
.A(n_374),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_423),
.B(n_438),
.Y(n_478)
);

BUFx5_ASAP7_75t_L g476 ( 
.A(n_427),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_L g428 ( 
.A1(n_410),
.A2(n_375),
.B(n_388),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_L g432 ( 
.A1(n_405),
.A2(n_397),
.B(n_414),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_SL g477 ( 
.A1(n_432),
.A2(n_446),
.B(n_455),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_379),
.B(n_312),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_433),
.B(n_437),
.C(n_386),
.Y(n_457)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_390),
.Y(n_435)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_435),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_436),
.B(n_440),
.Y(n_464)
);

MAJx2_ASAP7_75t_L g439 ( 
.A(n_412),
.B(n_328),
.C(n_313),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_SL g493 ( 
.A(n_439),
.B(n_365),
.Y(n_493)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_390),
.Y(n_442)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_442),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_378),
.B(n_364),
.Y(n_443)
);

INVxp33_ASAP7_75t_L g490 ( 
.A(n_443),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_444),
.A2(n_448),
.B1(n_451),
.B2(n_382),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_389),
.B(n_313),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_SL g480 ( 
.A(n_445),
.B(n_377),
.Y(n_480)
);

AOI21xp5_ASAP7_75t_L g446 ( 
.A1(n_402),
.A2(n_352),
.B(n_330),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_380),
.A2(n_349),
.B1(n_352),
.B2(n_347),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_404),
.A2(n_349),
.B1(n_321),
.B2(n_339),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_L g472 ( 
.A1(n_449),
.A2(n_452),
.B1(n_454),
.B2(n_456),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_SL g479 ( 
.A(n_450),
.B(n_453),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_380),
.A2(n_339),
.B1(n_327),
.B2(n_346),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_387),
.A2(n_327),
.B1(n_333),
.B2(n_348),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_409),
.B(n_350),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_371),
.A2(n_403),
.B1(n_372),
.B2(n_392),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_L g455 ( 
.A1(n_394),
.A2(n_333),
.B(n_370),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_403),
.A2(n_333),
.B1(n_359),
.B2(n_368),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_457),
.B(n_466),
.C(n_492),
.Y(n_498)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_458),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_421),
.B(n_384),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_459),
.B(n_465),
.Y(n_502)
);

CKINVDCx16_ASAP7_75t_R g461 ( 
.A(n_424),
.Y(n_461)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_461),
.Y(n_501)
);

OAI21xp5_ASAP7_75t_L g462 ( 
.A1(n_430),
.A2(n_385),
.B(n_400),
.Y(n_462)
);

OAI21xp5_ASAP7_75t_SL g497 ( 
.A1(n_462),
.A2(n_467),
.B(n_473),
.Y(n_497)
);

OA21x2_ASAP7_75t_L g465 ( 
.A1(n_432),
.A2(n_377),
.B(n_406),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_431),
.B(n_416),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_L g467 ( 
.A1(n_418),
.A2(n_373),
.B(n_381),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_L g515 ( 
.A1(n_469),
.A2(n_482),
.B1(n_491),
.B2(n_444),
.Y(n_515)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_435),
.Y(n_470)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_470),
.Y(n_513)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_442),
.Y(n_471)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_471),
.Y(n_518)
);

OAI21xp5_ASAP7_75t_L g473 ( 
.A1(n_428),
.A2(n_429),
.B(n_419),
.Y(n_473)
);

FAx1_ASAP7_75t_SL g474 ( 
.A(n_438),
.B(n_377),
.CI(n_399),
.CON(n_474),
.SN(n_474)
);

NOR2xp33_ASAP7_75t_SL g514 ( 
.A(n_474),
.B(n_481),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_421),
.B(n_393),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_475),
.B(n_486),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_480),
.B(n_485),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_425),
.B(n_393),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_L g482 ( 
.A1(n_454),
.A2(n_408),
.B1(n_401),
.B2(n_395),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_417),
.Y(n_483)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_483),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_425),
.B(n_441),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_SL g525 ( 
.A(n_484),
.B(n_487),
.Y(n_525)
);

OAI21xp5_ASAP7_75t_SL g485 ( 
.A1(n_446),
.A2(n_395),
.B(n_401),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_451),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_445),
.B(n_401),
.Y(n_487)
);

OAI21xp5_ASAP7_75t_L g488 ( 
.A1(n_429),
.A2(n_447),
.B(n_426),
.Y(n_488)
);

CKINVDCx16_ASAP7_75t_R g509 ( 
.A(n_488),
.Y(n_509)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_417),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_489),
.B(n_420),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_L g491 ( 
.A1(n_449),
.A2(n_422),
.B1(n_447),
.B2(n_426),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_431),
.B(n_319),
.Y(n_492)
);

XNOR2x1_ASAP7_75t_L g512 ( 
.A(n_493),
.B(n_480),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_481),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_494),
.B(n_519),
.Y(n_538)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_466),
.B(n_433),
.Y(n_499)
);

XOR2xp5_ASAP7_75t_L g530 ( 
.A(n_499),
.B(n_510),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_491),
.A2(n_448),
.B1(n_422),
.B2(n_434),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_SL g550 ( 
.A1(n_500),
.A2(n_505),
.B1(n_506),
.B2(n_521),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_457),
.B(n_437),
.C(n_439),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_504),
.B(n_507),
.C(n_526),
.Y(n_549)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_472),
.A2(n_434),
.B1(n_444),
.B2(n_455),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_472),
.A2(n_486),
.B1(n_464),
.B2(n_469),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_492),
.B(n_420),
.C(n_427),
.Y(n_507)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_508),
.Y(n_532)
);

XOR2xp5_ASAP7_75t_L g510 ( 
.A(n_493),
.B(n_452),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_464),
.A2(n_444),
.B1(n_440),
.B2(n_456),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_511),
.A2(n_515),
.B1(n_522),
.B2(n_474),
.Y(n_534)
);

XNOR2x1_ASAP7_75t_L g537 ( 
.A(n_512),
.B(n_476),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_484),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_516),
.B(n_517),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_479),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_479),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_519),
.B(n_468),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_L g520 ( 
.A1(n_461),
.A2(n_488),
.B1(n_464),
.B2(n_478),
.Y(n_520)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_520),
.Y(n_535)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_465),
.A2(n_365),
.B1(n_444),
.B2(n_462),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_465),
.A2(n_459),
.B1(n_473),
.B2(n_458),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_L g523 ( 
.A1(n_475),
.A2(n_465),
.B1(n_482),
.B2(n_490),
.Y(n_523)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_523),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_483),
.B(n_489),
.Y(n_524)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_524),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_467),
.B(n_463),
.C(n_477),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_517),
.B(n_477),
.Y(n_528)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_528),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_516),
.B(n_460),
.Y(n_531)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_531),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_524),
.B(n_460),
.Y(n_533)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_533),
.Y(n_573)
);

AOI22xp5_ASAP7_75t_L g574 ( 
.A1(n_534),
.A2(n_536),
.B1(n_550),
.B2(n_543),
.Y(n_574)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_500),
.A2(n_474),
.B1(n_463),
.B2(n_476),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_SL g562 ( 
.A(n_537),
.B(n_539),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_SL g555 ( 
.A(n_538),
.B(n_501),
.Y(n_555)
);

XOR2xp5_ASAP7_75t_L g539 ( 
.A(n_499),
.B(n_485),
.Y(n_539)
);

XOR2xp5_ASAP7_75t_L g559 ( 
.A(n_539),
.B(n_540),
.Y(n_559)
);

XOR2xp5_ASAP7_75t_L g540 ( 
.A(n_498),
.B(n_471),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g561 ( 
.A(n_541),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_508),
.B(n_468),
.Y(n_542)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_542),
.Y(n_571)
);

OAI21xp5_ASAP7_75t_SL g544 ( 
.A1(n_521),
.A2(n_470),
.B(n_497),
.Y(n_544)
);

AOI21xp5_ASAP7_75t_L g567 ( 
.A1(n_544),
.A2(n_553),
.B(n_512),
.Y(n_567)
);

INVx2_ASAP7_75t_SL g545 ( 
.A(n_527),
.Y(n_545)
);

INVxp67_ASAP7_75t_L g563 ( 
.A(n_545),
.Y(n_563)
);

AOI21xp5_ASAP7_75t_L g546 ( 
.A1(n_497),
.A2(n_526),
.B(n_502),
.Y(n_546)
);

OAI21xp5_ASAP7_75t_L g566 ( 
.A1(n_546),
.A2(n_547),
.B(n_525),
.Y(n_566)
);

AOI21xp5_ASAP7_75t_L g547 ( 
.A1(n_502),
.A2(n_522),
.B(n_496),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_527),
.B(n_496),
.Y(n_548)
);

XNOR2xp5_ASAP7_75t_L g572 ( 
.A(n_548),
.B(n_552),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_503),
.B(n_509),
.Y(n_552)
);

XOR2x2_ASAP7_75t_L g553 ( 
.A(n_510),
.B(n_495),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_513),
.Y(n_554)
);

BUFx2_ASAP7_75t_L g568 ( 
.A(n_554),
.Y(n_568)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_555),
.Y(n_579)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_540),
.B(n_498),
.C(n_504),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_558),
.B(n_566),
.Y(n_589)
);

A2O1A1Ixp33_ASAP7_75t_SL g560 ( 
.A1(n_550),
.A2(n_511),
.B(n_503),
.C(n_505),
.Y(n_560)
);

INVxp67_ASAP7_75t_L g583 ( 
.A(n_560),
.Y(n_583)
);

XNOR2xp5_ASAP7_75t_SL g588 ( 
.A(n_562),
.B(n_567),
.Y(n_588)
);

XOR2xp5_ASAP7_75t_L g564 ( 
.A(n_530),
.B(n_507),
.Y(n_564)
);

XNOR2xp5_ASAP7_75t_L g580 ( 
.A(n_564),
.B(n_565),
.Y(n_580)
);

XOR2xp5_ASAP7_75t_L g565 ( 
.A(n_530),
.B(n_495),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_535),
.B(n_501),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_569),
.B(n_576),
.Y(n_590)
);

AOI321xp33_ASAP7_75t_L g570 ( 
.A1(n_529),
.A2(n_506),
.A3(n_513),
.B1(n_514),
.B2(n_518),
.C(n_541),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_SL g584 ( 
.A(n_570),
.B(n_531),
.Y(n_584)
);

OAI22xp5_ASAP7_75t_SL g582 ( 
.A1(n_574),
.A2(n_534),
.B1(n_543),
.B2(n_532),
.Y(n_582)
);

NAND5xp2_ASAP7_75t_L g575 ( 
.A(n_544),
.B(n_518),
.C(n_552),
.D(n_529),
.E(n_547),
.Y(n_575)
);

XOR2xp5_ASAP7_75t_L g585 ( 
.A(n_575),
.B(n_542),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_549),
.B(n_546),
.C(n_553),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g577 ( 
.A(n_558),
.B(n_549),
.C(n_535),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_577),
.B(n_578),
.Y(n_600)
);

OAI21xp5_ASAP7_75t_SL g578 ( 
.A1(n_566),
.A2(n_528),
.B(n_536),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g581 ( 
.A(n_576),
.B(n_553),
.C(n_537),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g597 ( 
.A(n_581),
.B(n_587),
.C(n_592),
.Y(n_597)
);

AOI22xp5_ASAP7_75t_L g601 ( 
.A1(n_582),
.A2(n_571),
.B1(n_560),
.B2(n_563),
.Y(n_601)
);

NOR2xp67_ASAP7_75t_L g605 ( 
.A(n_584),
.B(n_560),
.Y(n_605)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_585),
.Y(n_607)
);

XNOR2xp5_ASAP7_75t_L g586 ( 
.A(n_556),
.B(n_548),
.Y(n_586)
);

XOR2xp5_ASAP7_75t_L g595 ( 
.A(n_586),
.B(n_572),
.Y(n_595)
);

MAJIxp5_ASAP7_75t_L g587 ( 
.A(n_559),
.B(n_545),
.C(n_532),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_561),
.B(n_551),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_SL g603 ( 
.A(n_591),
.B(n_568),
.Y(n_603)
);

MAJIxp5_ASAP7_75t_L g592 ( 
.A(n_559),
.B(n_545),
.C(n_551),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_564),
.B(n_554),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_SL g602 ( 
.A(n_593),
.B(n_594),
.Y(n_602)
);

MAJIxp5_ASAP7_75t_L g594 ( 
.A(n_565),
.B(n_533),
.C(n_562),
.Y(n_594)
);

XOR2xp5_ASAP7_75t_L g609 ( 
.A(n_595),
.B(n_598),
.Y(n_609)
);

AOI21xp5_ASAP7_75t_L g596 ( 
.A1(n_585),
.A2(n_557),
.B(n_574),
.Y(n_596)
);

AOI21xp5_ASAP7_75t_L g615 ( 
.A1(n_596),
.A2(n_605),
.B(n_606),
.Y(n_615)
);

XOR2xp5_ASAP7_75t_L g598 ( 
.A(n_594),
.B(n_572),
.Y(n_598)
);

OAI22xp5_ASAP7_75t_SL g599 ( 
.A1(n_583),
.A2(n_573),
.B1(n_560),
.B2(n_575),
.Y(n_599)
);

OAI22xp5_ASAP7_75t_SL g610 ( 
.A1(n_599),
.A2(n_601),
.B1(n_608),
.B2(n_588),
.Y(n_610)
);

OAI22xp5_ASAP7_75t_L g616 ( 
.A1(n_603),
.A2(n_607),
.B1(n_596),
.B2(n_595),
.Y(n_616)
);

XOR2xp5_ASAP7_75t_L g604 ( 
.A(n_581),
.B(n_587),
.Y(n_604)
);

MAJIxp5_ASAP7_75t_L g611 ( 
.A(n_604),
.B(n_577),
.C(n_597),
.Y(n_611)
);

NOR2x1_ASAP7_75t_L g606 ( 
.A(n_586),
.B(n_563),
.Y(n_606)
);

OAI22xp5_ASAP7_75t_SL g608 ( 
.A1(n_583),
.A2(n_568),
.B1(n_590),
.B2(n_589),
.Y(n_608)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_610),
.Y(n_624)
);

MAJIxp5_ASAP7_75t_L g625 ( 
.A(n_611),
.B(n_613),
.C(n_614),
.Y(n_625)
);

FAx1_ASAP7_75t_SL g612 ( 
.A(n_599),
.B(n_588),
.CI(n_592),
.CON(n_612),
.SN(n_612)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_612),
.B(n_616),
.Y(n_619)
);

MAJIxp5_ASAP7_75t_L g613 ( 
.A(n_597),
.B(n_580),
.C(n_579),
.Y(n_613)
);

MAJIxp5_ASAP7_75t_L g614 ( 
.A(n_604),
.B(n_598),
.C(n_600),
.Y(n_614)
);

NOR2xp67_ASAP7_75t_SL g617 ( 
.A(n_607),
.B(n_601),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_617),
.B(n_618),
.Y(n_621)
);

OAI22xp5_ASAP7_75t_L g618 ( 
.A1(n_603),
.A2(n_608),
.B1(n_602),
.B2(n_606),
.Y(n_618)
);

OAI21xp33_ASAP7_75t_L g620 ( 
.A1(n_615),
.A2(n_610),
.B(n_618),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_620),
.B(n_623),
.Y(n_626)
);

OAI21xp5_ASAP7_75t_SL g622 ( 
.A1(n_615),
.A2(n_614),
.B(n_613),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_622),
.B(n_609),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g623 ( 
.A(n_611),
.Y(n_623)
);

AOI21xp5_ASAP7_75t_L g631 ( 
.A1(n_627),
.A2(n_619),
.B(n_621),
.Y(n_631)
);

INVxp67_ASAP7_75t_L g628 ( 
.A(n_625),
.Y(n_628)
);

NAND3xp33_ASAP7_75t_L g630 ( 
.A(n_628),
.B(n_629),
.C(n_623),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_620),
.B(n_609),
.Y(n_629)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_630),
.Y(n_632)
);

OAI221xp5_ASAP7_75t_L g633 ( 
.A1(n_632),
.A2(n_626),
.B1(n_631),
.B2(n_624),
.C(n_617),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_633),
.B(n_612),
.Y(n_634)
);

XOR2xp5_ASAP7_75t_L g635 ( 
.A(n_634),
.B(n_612),
.Y(n_635)
);


endmodule