module real_jpeg_4733_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_464;
wire n_423;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_531;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g198 ( 
.A(n_0),
.Y(n_198)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_0),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_0),
.Y(n_233)
);

BUFx5_ASAP7_75t_L g286 ( 
.A(n_0),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_0),
.Y(n_417)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_1),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_1),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g329 ( 
.A(n_1),
.Y(n_329)
);

INVx3_ASAP7_75t_L g429 ( 
.A(n_1),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_1),
.Y(n_458)
);

AOI22xp33_ASAP7_75t_L g280 ( 
.A1(n_2),
.A2(n_281),
.B1(n_283),
.B2(n_284),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_2),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_SL g364 ( 
.A1(n_2),
.A2(n_283),
.B1(n_365),
.B2(n_367),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_2),
.A2(n_283),
.B1(n_288),
.B2(n_391),
.Y(n_390)
);

OAI22xp33_ASAP7_75t_L g455 ( 
.A1(n_2),
.A2(n_67),
.B1(n_283),
.B2(n_456),
.Y(n_455)
);

AOI22xp33_ASAP7_75t_L g211 ( 
.A1(n_3),
.A2(n_212),
.B1(n_216),
.B2(n_217),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_3),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_3),
.A2(n_204),
.B1(n_216),
.B2(n_238),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g306 ( 
.A1(n_3),
.A2(n_102),
.B1(n_216),
.B2(n_307),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_3),
.A2(n_216),
.B1(n_328),
.B2(n_428),
.Y(n_427)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_4),
.A2(n_44),
.B1(n_46),
.B2(n_47),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_4),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_4),
.A2(n_47),
.B1(n_107),
.B2(n_108),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_4),
.A2(n_47),
.B1(n_142),
.B2(n_143),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_4),
.A2(n_47),
.B1(n_381),
.B2(n_382),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_6),
.A2(n_142),
.B1(n_171),
.B2(n_172),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_6),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_6),
.A2(n_172),
.B1(n_204),
.B2(n_207),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_6),
.A2(n_172),
.B1(n_275),
.B2(n_276),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_6),
.A2(n_46),
.B1(n_172),
.B2(n_355),
.Y(n_354)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_7),
.Y(n_534)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_8),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_8),
.Y(n_123)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_8),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_8),
.Y(n_179)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_9),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_10),
.A2(n_163),
.B1(n_165),
.B2(n_168),
.Y(n_162)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_10),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_10),
.B(n_179),
.C(n_180),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_10),
.B(n_89),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_10),
.B(n_233),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_10),
.B(n_140),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_10),
.B(n_270),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_11),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_11),
.Y(n_134)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_11),
.Y(n_185)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_12),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_13),
.Y(n_537)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_14),
.A2(n_51),
.B1(n_56),
.B2(n_57),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_14),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_14),
.A2(n_57),
.B1(n_99),
.B2(n_102),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_SL g376 ( 
.A1(n_14),
.A2(n_57),
.B1(n_181),
.B2(n_377),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_14),
.A2(n_57),
.B1(n_406),
.B2(n_410),
.Y(n_405)
);

OAI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_15),
.A2(n_189),
.B1(n_191),
.B2(n_192),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_15),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_15),
.A2(n_142),
.B1(n_191),
.B2(n_213),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_L g360 ( 
.A1(n_15),
.A2(n_191),
.B1(n_288),
.B2(n_361),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_15),
.A2(n_70),
.B1(n_73),
.B2(n_191),
.Y(n_401)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_16),
.A2(n_67),
.B1(n_69),
.B2(n_71),
.Y(n_66)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_16),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g313 ( 
.A1(n_16),
.A2(n_71),
.B1(n_314),
.B2(n_315),
.Y(n_313)
);

OAI22xp33_ASAP7_75t_SL g385 ( 
.A1(n_16),
.A2(n_71),
.B1(n_212),
.B2(n_367),
.Y(n_385)
);

AOI22xp33_ASAP7_75t_SL g394 ( 
.A1(n_16),
.A2(n_71),
.B1(n_395),
.B2(n_397),
.Y(n_394)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_18),
.A2(n_44),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_18),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g340 ( 
.A1(n_18),
.A2(n_74),
.B1(n_341),
.B2(n_343),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_18),
.A2(n_74),
.B1(n_144),
.B2(n_387),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_18),
.A2(n_74),
.B1(n_391),
.B2(n_441),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_533),
.B(n_535),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_60),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_59),
.Y(n_21)
);

OR2x2_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_48),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_23),
.B(n_48),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_36),
.B(n_42),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_24),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_24),
.B(n_354),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_24),
.B(n_455),
.Y(n_454)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_37),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_29),
.B1(n_32),
.B2(n_34),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx4_ASAP7_75t_L g333 ( 
.A(n_28),
.Y(n_333)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_31),
.Y(n_83)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_31),
.Y(n_101)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_31),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_31),
.Y(n_272)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_33),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_33),
.Y(n_107)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g49 ( 
.A(n_36),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_36),
.A2(n_350),
.B(n_352),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_36),
.B(n_354),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_37)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_38),
.Y(n_331)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

INVx8_ASAP7_75t_L g351 ( 
.A(n_39),
.Y(n_351)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_43),
.A2(n_49),
.B1(n_50),
.B2(n_58),
.Y(n_48)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_48),
.B(n_62),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_48),
.B(n_62),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_49),
.A2(n_58),
.B1(n_66),
.B2(n_72),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_49),
.A2(n_50),
.B1(n_58),
.B2(n_72),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g400 ( 
.A1(n_49),
.A2(n_353),
.B(n_401),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g426 ( 
.A1(n_49),
.A2(n_58),
.B1(n_401),
.B2(n_427),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g504 ( 
.A1(n_49),
.A2(n_58),
.B1(n_66),
.B2(n_505),
.Y(n_504)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_52),
.B(n_168),
.Y(n_334)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_55),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_58),
.B(n_168),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g469 ( 
.A1(n_58),
.A2(n_427),
.B(n_459),
.Y(n_469)
);

AO21x1_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_152),
.B(n_532),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_148),
.C(n_149),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g527 ( 
.A1(n_63),
.A2(n_64),
.B1(n_528),
.B2(n_529),
.Y(n_527)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_75),
.C(n_111),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_SL g519 ( 
.A(n_65),
.B(n_520),
.Y(n_519)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_75),
.A2(n_111),
.B1(n_112),
.B2(n_521),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_75),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_76),
.A2(n_98),
.B1(n_105),
.B2(n_106),
.Y(n_75)
);

INVx2_ASAP7_75t_SL g150 ( 
.A(n_76),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_76),
.A2(n_105),
.B1(n_306),
.B2(n_360),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_76),
.A2(n_105),
.B1(n_390),
.B2(n_394),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g508 ( 
.A1(n_76),
.A2(n_98),
.B1(n_105),
.B2(n_509),
.Y(n_508)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_89),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_80),
.B1(n_84),
.B2(n_87),
.Y(n_77)
);

INVx6_ASAP7_75t_L g295 ( 
.A(n_78),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_79),
.Y(n_86)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_80),
.Y(n_275)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_83),
.Y(n_267)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_83),
.Y(n_327)
);

INVx3_ASAP7_75t_L g443 ( 
.A(n_83),
.Y(n_443)
);

AO22x2_ASAP7_75t_L g89 ( 
.A1(n_84),
.A2(n_90),
.B1(n_94),
.B2(n_96),
.Y(n_89)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_86),
.Y(n_293)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g399 ( 
.A(n_88),
.Y(n_399)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_89),
.A2(n_150),
.B(n_151),
.Y(n_149)
);

AOI22x1_ASAP7_75t_L g430 ( 
.A1(n_89),
.A2(n_150),
.B1(n_309),
.B2(n_431),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_89),
.A2(n_150),
.B1(n_439),
.B2(n_440),
.Y(n_438)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_93),
.Y(n_95)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_93),
.Y(n_117)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_93),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_93),
.Y(n_142)
);

INVx11_ASAP7_75t_L g147 ( 
.A(n_93),
.Y(n_147)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_93),
.Y(n_164)
);

BUFx5_ASAP7_75t_L g409 ( 
.A(n_93),
.Y(n_409)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_99),
.B(n_333),
.Y(n_332)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_101),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_101),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_101),
.Y(n_396)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx5_ASAP7_75t_L g276 ( 
.A(n_103),
.Y(n_276)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_105),
.B(n_274),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_105),
.A2(n_306),
.B(n_308),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_106),
.Y(n_151)
);

INVx4_ASAP7_75t_L g288 ( 
.A(n_107),
.Y(n_288)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_111),
.A2(n_112),
.B1(n_507),
.B2(n_508),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_111),
.B(n_504),
.C(n_507),
.Y(n_515)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_113),
.A2(n_139),
.B(n_141),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_113),
.A2(n_162),
.B(n_169),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_113),
.A2(n_139),
.B1(n_211),
.B2(n_263),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_113),
.A2(n_169),
.B(n_263),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_113),
.A2(n_139),
.B1(n_364),
.B2(n_422),
.Y(n_421)
);

INVx2_ASAP7_75t_SL g113 ( 
.A(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_114),
.B(n_170),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_114),
.A2(n_140),
.B1(n_385),
.B2(n_386),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_114),
.A2(n_140),
.B1(n_386),
.B2(n_405),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_114),
.A2(n_140),
.B1(n_405),
.B2(n_446),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_126),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_118),
.B1(n_121),
.B2(n_124),
.Y(n_115)
);

INVx4_ASAP7_75t_SL g367 ( 
.A(n_116),
.Y(n_367)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g387 ( 
.A(n_117),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_123),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_125),
.Y(n_291)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_126),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_126),
.A2(n_211),
.B(n_220),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_129),
.B1(n_133),
.B2(n_135),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_132),
.Y(n_200)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_132),
.Y(n_285)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_132),
.Y(n_314)
);

BUFx8_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_134),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_134),
.Y(n_240)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g363 ( 
.A1(n_139),
.A2(n_220),
.B(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_140),
.B(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_141),
.Y(n_446)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

NAND2xp33_ASAP7_75t_SL g294 ( 
.A(n_145),
.B(n_295),
.Y(n_294)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_146),
.Y(n_177)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_147),
.Y(n_167)
);

INVx5_ASAP7_75t_L g215 ( 
.A(n_147),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_147),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_147),
.Y(n_366)
);

INVx6_ASAP7_75t_L g413 ( 
.A(n_147),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g529 ( 
.A(n_148),
.B(n_149),
.Y(n_529)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_150),
.A2(n_266),
.B(n_273),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_150),
.B(n_309),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g471 ( 
.A1(n_150),
.A2(n_273),
.B(n_472),
.Y(n_471)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_526),
.B(n_531),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_498),
.B(n_523),
.Y(n_153)
);

OAI311xp33_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_370),
.A3(n_474),
.B1(n_492),
.C1(n_493),
.Y(n_154)
);

AOI21x1_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_320),
.B(n_369),
.Y(n_155)
);

AO21x1_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_297),
.B(n_319),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_257),
.B(n_296),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_223),
.B(n_256),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_186),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_160),
.B(n_186),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_161),
.B(n_173),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_161),
.A2(n_173),
.B1(n_174),
.B2(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_161),
.Y(n_254)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_163),
.Y(n_171)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_168),
.A2(n_195),
.B(n_201),
.Y(n_234)
);

OAI21xp33_ASAP7_75t_SL g266 ( 
.A1(n_168),
.A2(n_267),
.B(n_268),
.Y(n_266)
);

OAI21xp33_ASAP7_75t_SL g350 ( 
.A1(n_168),
.A2(n_334),
.B(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_178),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_183),
.Y(n_342)
);

INVx5_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_184),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_185),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_185),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_208),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_187),
.B(n_209),
.C(n_222),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_195),
.B(n_201),
.Y(n_187)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_188),
.Y(n_249)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_192),
.Y(n_315)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_194),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_195),
.A2(n_337),
.B1(n_338),
.B2(n_339),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_195),
.A2(n_251),
.B1(n_376),
.B2(n_380),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_SL g414 ( 
.A1(n_195),
.A2(n_380),
.B(n_415),
.Y(n_414)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_196),
.B(n_203),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_196),
.A2(n_248),
.B1(n_249),
.B2(n_250),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_196),
.A2(n_280),
.B1(n_313),
.B2(n_316),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_196),
.A2(n_316),
.B1(n_340),
.B2(n_424),
.Y(n_423)
);

OR2x2_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_199),
.Y(n_196)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_197),
.Y(n_242)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_198),
.Y(n_252)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_198),
.Y(n_317)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_199),
.Y(n_207)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx8_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx4_ASAP7_75t_L g343 ( 
.A(n_206),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_209),
.A2(n_210),
.B1(n_221),
.B2(n_222),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_213),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx11_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_246),
.B(n_255),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_235),
.B(n_245),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_234),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_232),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx6_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_231),
.Y(n_282)
);

INVx3_ASAP7_75t_L g379 ( 
.A(n_231),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_236),
.B(n_244),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_236),
.B(n_244),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_241),
.B(n_243),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_237),
.Y(n_248)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx5_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_243),
.A2(n_279),
.B(n_286),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_253),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_247),
.B(n_253),
.Y(n_255)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx8_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_258),
.B(n_259),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_277),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_262),
.B1(n_264),
.B2(n_265),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_262),
.B(n_264),
.C(n_277),
.Y(n_298)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVxp33_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

AOI32xp33_ASAP7_75t_L g287 ( 
.A1(n_269),
.A2(n_288),
.A3(n_289),
.B1(n_292),
.B2(n_294),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_271),
.Y(n_270)
);

INVx6_ASAP7_75t_SL g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_274),
.Y(n_309)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_276),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_287),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_278),
.B(n_287),
.Y(n_303)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx6_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx5_ASAP7_75t_SL g289 ( 
.A(n_290),
.Y(n_289)
);

INVx4_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx5_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_298),
.B(n_299),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_300),
.A2(n_301),
.B1(n_304),
.B2(n_318),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_SL g301 ( 
.A(n_302),
.B(n_303),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_302),
.B(n_303),
.C(n_318),
.Y(n_321)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_304),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_SL g304 ( 
.A(n_305),
.B(n_310),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_305),
.B(n_311),
.C(n_312),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_313),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_316),
.Y(n_338)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_322),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g369 ( 
.A(n_321),
.B(n_322),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_347),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_324),
.A2(n_344),
.B1(n_345),
.B2(n_346),
.Y(n_323)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_324),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_325),
.A2(n_326),
.B1(n_335),
.B2(n_336),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_326),
.B(n_335),
.Y(n_470)
);

OAI32xp33_ASAP7_75t_L g326 ( 
.A1(n_327),
.A2(n_328),
.A3(n_330),
.B1(n_332),
.B2(n_334),
.Y(n_326)
);

INVx3_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_SL g330 ( 
.A(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_341),
.Y(n_381)
);

INVx3_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_344),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_344),
.B(n_345),
.C(n_347),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_348),
.A2(n_349),
.B1(n_358),
.B2(n_368),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_348),
.B(n_359),
.C(n_363),
.Y(n_483)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx4_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_358),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_SL g358 ( 
.A(n_359),
.B(n_363),
.Y(n_358)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_360),
.Y(n_472)
);

INVx3_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx5_ASAP7_75t_L g393 ( 
.A(n_362),
.Y(n_393)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

NAND2xp33_ASAP7_75t_SL g370 ( 
.A(n_371),
.B(n_460),
.Y(n_370)
);

A2O1A1Ixp33_ASAP7_75t_SL g493 ( 
.A1(n_371),
.A2(n_460),
.B(n_494),
.C(n_497),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_432),
.Y(n_371)
);

OR2x2_ASAP7_75t_L g492 ( 
.A(n_372),
.B(n_432),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_402),
.C(n_419),
.Y(n_372)
);

FAx1_ASAP7_75t_L g473 ( 
.A(n_373),
.B(n_402),
.CI(n_419),
.CON(n_473),
.SN(n_473)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_388),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_374),
.B(n_389),
.C(n_400),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_384),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_375),
.B(n_384),
.Y(n_466)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_376),
.Y(n_424)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_SL g378 ( 
.A(n_379),
.Y(n_378)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_385),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_400),
.Y(n_388)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_390),
.Y(n_431)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx4_ASAP7_75t_SL g392 ( 
.A(n_393),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_394),
.Y(n_439)
);

INVx6_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_403),
.A2(n_404),
.B1(n_414),
.B2(n_418),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_404),
.B(n_414),
.Y(n_450)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx5_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

BUFx2_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx8_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_414),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_414),
.A2(n_418),
.B1(n_452),
.B2(n_453),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_L g501 ( 
.A1(n_414),
.A2(n_450),
.B(n_453),
.Y(n_501)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_420),
.B(n_425),
.C(n_430),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_420),
.B(n_464),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_421),
.B(n_423),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_421),
.B(n_423),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_425),
.A2(n_426),
.B1(n_430),
.B2(n_465),
.Y(n_464)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx6_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx1_ASAP7_75t_SL g465 ( 
.A(n_430),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_433),
.B(n_434),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_433),
.B(n_436),
.C(n_448),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_435),
.A2(n_436),
.B1(n_448),
.B2(n_449),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_L g436 ( 
.A1(n_437),
.A2(n_444),
.B(n_447),
.Y(n_436)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g447 ( 
.A(n_438),
.B(n_445),
.Y(n_447)
);

INVxp67_ASAP7_75t_L g509 ( 
.A(n_440),
.Y(n_509)
);

INVx5_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVx4_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

FAx1_ASAP7_75t_SL g500 ( 
.A(n_447),
.B(n_501),
.CI(n_502),
.CON(n_500),
.SN(n_500)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_447),
.B(n_501),
.C(n_502),
.Y(n_522)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_451),
.Y(n_449)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_459),
.Y(n_453)
);

INVxp67_ASAP7_75t_L g505 ( 
.A(n_455),
.Y(n_505)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_473),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_461),
.B(n_473),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_466),
.C(n_467),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_462),
.A2(n_463),
.B1(n_466),
.B2(n_486),
.Y(n_485)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_466),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_467),
.B(n_485),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_468),
.B(n_470),
.C(n_471),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_468),
.A2(n_469),
.B1(n_471),
.B2(n_480),
.Y(n_479)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_470),
.B(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_471),
.Y(n_480)
);

BUFx24_ASAP7_75t_SL g540 ( 
.A(n_473),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_475),
.B(n_487),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

OAI21xp5_ASAP7_75t_L g494 ( 
.A1(n_476),
.A2(n_495),
.B(n_496),
.Y(n_494)
);

NOR2x1_ASAP7_75t_L g476 ( 
.A(n_477),
.B(n_484),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_477),
.B(n_484),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_478),
.B(n_481),
.C(n_483),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_478),
.B(n_490),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_481),
.A2(n_482),
.B1(n_483),
.B2(n_491),
.Y(n_490)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_483),
.Y(n_491)
);

OR2x2_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_489),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_488),
.B(n_489),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_499),
.B(n_512),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_SL g499 ( 
.A(n_500),
.B(n_511),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_500),
.B(n_511),
.Y(n_524)
);

BUFx24_ASAP7_75t_SL g538 ( 
.A(n_500),
.Y(n_538)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_503),
.A2(n_504),
.B1(n_506),
.B2(n_510),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_503),
.A2(n_504),
.B1(n_518),
.B2(n_519),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_503),
.B(n_514),
.C(n_518),
.Y(n_530)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_506),
.Y(n_510)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_L g523 ( 
.A1(n_512),
.A2(n_524),
.B(n_525),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_SL g512 ( 
.A(n_513),
.B(n_522),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_513),
.B(n_522),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_L g513 ( 
.A1(n_514),
.A2(n_515),
.B1(n_516),
.B2(n_517),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_519),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_527),
.B(n_530),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_527),
.B(n_530),
.Y(n_531)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_529),
.Y(n_528)
);

INVx5_ASAP7_75t_L g533 ( 
.A(n_534),
.Y(n_533)
);

INVx8_ASAP7_75t_L g536 ( 
.A(n_534),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_536),
.B(n_537),
.Y(n_535)
);


endmodule