module fake_jpeg_31781_n_203 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_203);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_203;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx2_ASAP7_75t_SL g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_15),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_43),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_37),
.Y(n_79)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_15),
.B(n_19),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_41),
.B(n_25),
.Y(n_75)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_19),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

AOI21xp33_ASAP7_75t_L g45 ( 
.A1(n_17),
.A2(n_0),
.B(n_1),
.Y(n_45)
);

AND2x2_ASAP7_75t_SL g52 ( 
.A(n_45),
.B(n_0),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

BUFx16f_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_22),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_48),
.B(n_22),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_49),
.B(n_74),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

A2O1A1Ixp33_ASAP7_75t_L g93 ( 
.A1(n_52),
.A2(n_30),
.B(n_24),
.C(n_18),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_45),
.A2(n_21),
.B1(n_29),
.B2(n_31),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_55),
.A2(n_66),
.B1(n_70),
.B2(n_31),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_41),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_56),
.B(n_62),
.Y(n_83)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_36),
.B(n_25),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_34),
.A2(n_35),
.B1(n_37),
.B2(n_39),
.Y(n_66)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_35),
.A2(n_21),
.B1(n_29),
.B2(n_30),
.Y(n_70)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

INVx3_ASAP7_75t_SL g100 ( 
.A(n_71),
.Y(n_100)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_72),
.Y(n_96)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_73),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_75),
.B(n_76),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_43),
.B(n_33),
.Y(n_76)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_37),
.Y(n_78)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_78),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_50),
.A2(n_38),
.B1(n_40),
.B2(n_46),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_82),
.A2(n_66),
.B1(n_64),
.B2(n_78),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_85),
.A2(n_86),
.B1(n_67),
.B2(n_79),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_77),
.A2(n_20),
.B1(n_18),
.B2(n_17),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_61),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_90),
.B(n_91),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_70),
.B(n_48),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_32),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_94),
.B(n_95),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_69),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_52),
.B(n_24),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_102),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_68),
.B(n_79),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_59),
.Y(n_103)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_103),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_65),
.B(n_33),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_104),
.B(n_105),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_65),
.B(n_32),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_92),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_106),
.B(n_110),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_98),
.B(n_71),
.C(n_54),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_107),
.B(n_109),
.C(n_112),
.Y(n_130)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_108),
.Y(n_136)
);

AND2x2_ASAP7_75t_SL g109 ( 
.A(n_104),
.B(n_51),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_85),
.B(n_54),
.C(n_64),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_88),
.Y(n_113)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_113),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_114),
.A2(n_117),
.B1(n_118),
.B2(n_125),
.Y(n_138)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_97),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_115),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_93),
.B(n_26),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_116),
.B(n_89),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_91),
.A2(n_67),
.B1(n_53),
.B2(n_27),
.Y(n_118)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_84),
.Y(n_122)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_122),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_83),
.B(n_27),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_123),
.B(n_13),
.Y(n_144)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_84),
.Y(n_124)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_124),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_102),
.A2(n_53),
.B1(n_26),
.B2(n_20),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_96),
.Y(n_126)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_126),
.Y(n_141)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_96),
.Y(n_128)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_128),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_119),
.A2(n_105),
.B(n_94),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_129),
.A2(n_132),
.B(n_143),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_99),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_131),
.B(n_134),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_114),
.A2(n_100),
.B(n_89),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_133),
.B(n_127),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_112),
.A2(n_81),
.B1(n_103),
.B2(n_101),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_117),
.A2(n_81),
.B1(n_101),
.B2(n_100),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_135),
.B(n_134),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_107),
.A2(n_69),
.B(n_80),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_144),
.B(n_147),
.Y(n_153)
);

AND2x6_ASAP7_75t_L g147 ( 
.A(n_110),
.B(n_87),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_127),
.A2(n_80),
.B(n_87),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_148),
.A2(n_0),
.B(n_1),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_150),
.B(n_151),
.C(n_133),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_130),
.B(n_109),
.C(n_116),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_145),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_152),
.B(n_159),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_132),
.A2(n_120),
.B(n_109),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_155),
.A2(n_156),
.B(n_162),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_130),
.A2(n_118),
.B(n_125),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_138),
.A2(n_128),
.B1(n_121),
.B2(n_80),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_157),
.A2(n_158),
.B1(n_142),
.B2(n_146),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_131),
.A2(n_121),
.B1(n_1),
.B2(n_2),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_142),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_137),
.Y(n_160)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_160),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_161),
.A2(n_148),
.B1(n_135),
.B2(n_140),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_164),
.A2(n_174),
.B1(n_159),
.B2(n_157),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_155),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_165),
.A2(n_168),
.B1(n_161),
.B2(n_156),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_152),
.B(n_139),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_166),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_167),
.B(n_172),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_149),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_169),
.Y(n_181)
);

A2O1A1O1Ixp25_ASAP7_75t_L g170 ( 
.A1(n_154),
.A2(n_129),
.B(n_147),
.C(n_143),
.D(n_141),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_170),
.B(n_12),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_151),
.B(n_141),
.C(n_140),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_160),
.Y(n_174)
);

A2O1A1O1Ixp25_ASAP7_75t_L g175 ( 
.A1(n_169),
.A2(n_154),
.B(n_153),
.C(n_149),
.D(n_162),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_175),
.B(n_168),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_176),
.B(n_177),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_163),
.A2(n_137),
.B1(n_136),
.B2(n_150),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_178),
.B(n_182),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_163),
.A2(n_10),
.B(n_11),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_180),
.A2(n_3),
.B(n_4),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_179),
.B(n_172),
.C(n_167),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_184),
.B(n_186),
.C(n_4),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_179),
.B(n_173),
.C(n_170),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_188),
.A2(n_6),
.B(n_7),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_189),
.A2(n_183),
.B1(n_181),
.B2(n_182),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_190),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_187),
.A2(n_181),
.B1(n_175),
.B2(n_171),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_191),
.B(n_192),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_184),
.A2(n_3),
.B(n_4),
.Y(n_192)
);

OAI21xp33_ASAP7_75t_L g197 ( 
.A1(n_193),
.A2(n_194),
.B(n_6),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_197),
.B(n_185),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_195),
.B(n_193),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_198),
.B(n_199),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_200),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_201),
.B(n_196),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_202),
.B(n_188),
.Y(n_203)
);


endmodule