module fake_jpeg_18707_n_318 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_318);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_318;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx2_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_17),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx2_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

INVx5_ASAP7_75t_SL g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

HB1xp67_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

INVx3_ASAP7_75t_SL g91 ( 
.A(n_41),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_23),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_43),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_0),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_30),
.B(n_0),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_45),
.B(n_20),
.Y(n_83)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_30),
.B(n_0),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_37),
.C(n_20),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_23),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_55),
.Y(n_69)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_24),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_24),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_57),
.B(n_21),
.Y(n_97)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_58),
.Y(n_100)
);

BUFx10_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx13_ASAP7_75t_L g129 ( 
.A(n_59),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_28),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_60),
.B(n_64),
.Y(n_116)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_61),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_46),
.A2(n_18),
.B1(n_35),
.B2(n_29),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_62),
.A2(n_76),
.B1(n_78),
.B2(n_81),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_28),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_65),
.B(n_36),
.Y(n_108)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_71),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_72),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_51),
.B(n_18),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_73),
.A2(n_85),
.B1(n_93),
.B2(n_96),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_74),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_46),
.A2(n_35),
.B1(n_29),
.B2(n_31),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_43),
.A2(n_39),
.B1(n_31),
.B2(n_37),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_44),
.A2(n_31),
.B1(n_26),
.B2(n_39),
.Y(n_81)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_83),
.B(n_89),
.Y(n_112)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_51),
.B(n_34),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_49),
.A2(n_26),
.B1(n_27),
.B2(n_36),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_88),
.A2(n_41),
.B1(n_26),
.B2(n_53),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_42),
.B(n_19),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_90),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_51),
.A2(n_2),
.B(n_3),
.Y(n_92)
);

A2O1A1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_92),
.A2(n_41),
.B(n_27),
.C(n_32),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_51),
.B(n_34),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_94),
.Y(n_130)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_95),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_40),
.B(n_19),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_21),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_85),
.A2(n_48),
.B(n_47),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_99),
.A2(n_104),
.B(n_113),
.Y(n_167)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_86),
.Y(n_102)
);

INVx13_ASAP7_75t_L g139 ( 
.A(n_102),
.Y(n_139)
);

NAND2x1_ASAP7_75t_SL g104 ( 
.A(n_88),
.B(n_57),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_62),
.A2(n_57),
.B1(n_55),
.B2(n_53),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_105),
.A2(n_107),
.B1(n_117),
.B2(n_81),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_108),
.B(n_2),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_73),
.B(n_93),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_67),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_114),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_76),
.A2(n_55),
.B1(n_42),
.B2(n_41),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_69),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_128),
.Y(n_137)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_80),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_119),
.A2(n_126),
.B1(n_127),
.B2(n_79),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_120),
.B(n_122),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_121),
.B(n_123),
.Y(n_163)
);

OA22x2_ASAP7_75t_SL g122 ( 
.A1(n_68),
.A2(n_48),
.B1(n_52),
.B2(n_56),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_96),
.B(n_33),
.Y(n_123)
);

INVx11_ASAP7_75t_L g124 ( 
.A(n_90),
.Y(n_124)
);

INVx13_ASAP7_75t_L g152 ( 
.A(n_124),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_75),
.A2(n_32),
.B1(n_22),
.B2(n_33),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_125),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_87),
.A2(n_32),
.B1(n_22),
.B2(n_33),
.Y(n_126)
);

INVx11_ASAP7_75t_L g127 ( 
.A(n_59),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_59),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_63),
.B(n_32),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_52),
.Y(n_145)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_77),
.Y(n_134)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_134),
.Y(n_136)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_79),
.Y(n_135)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_135),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_140),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_141),
.A2(n_166),
.B1(n_110),
.B2(n_101),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_129),
.Y(n_142)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_142),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_113),
.B(n_67),
.C(n_70),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_144),
.B(n_154),
.C(n_99),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_145),
.Y(n_180)
);

CKINVDCx12_ASAP7_75t_R g146 ( 
.A(n_102),
.Y(n_146)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_146),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_98),
.B(n_56),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_147),
.B(n_103),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_116),
.B(n_86),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_148),
.B(n_151),
.Y(n_169)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_109),
.Y(n_149)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_149),
.Y(n_168)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_130),
.Y(n_150)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_150),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_112),
.B(n_82),
.Y(n_151)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_130),
.Y(n_153)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_153),
.Y(n_184)
);

AND2x2_ASAP7_75t_SL g154 ( 
.A(n_115),
.B(n_113),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_108),
.B(n_80),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_155),
.B(n_159),
.Y(n_170)
);

OAI21xp33_ASAP7_75t_L g193 ( 
.A1(n_157),
.A2(n_3),
.B(n_4),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_122),
.B(n_87),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_158),
.B(n_162),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_111),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_134),
.Y(n_160)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_160),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_122),
.B(n_70),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_108),
.B(n_91),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_164),
.B(n_165),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_109),
.B(n_100),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_115),
.A2(n_91),
.B1(n_66),
.B2(n_74),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_171),
.B(n_173),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_158),
.A2(n_104),
.B1(n_103),
.B2(n_114),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_172),
.A2(n_187),
.B1(n_189),
.B2(n_192),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_150),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_176),
.B(n_185),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_167),
.A2(n_120),
.B(n_131),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_177),
.A2(n_197),
.B(n_199),
.Y(n_211)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_153),
.Y(n_179)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_179),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_167),
.B(n_100),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_182),
.B(n_188),
.Y(n_205)
);

MAJx2_ASAP7_75t_L g183 ( 
.A(n_154),
.B(n_106),
.C(n_119),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_183),
.A2(n_147),
.B(n_163),
.Y(n_203)
);

NOR2x1_ASAP7_75t_L g185 ( 
.A(n_146),
.B(n_106),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_162),
.A2(n_110),
.B1(n_101),
.B2(n_66),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_154),
.B(n_135),
.Y(n_188)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_137),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_190),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_156),
.A2(n_154),
.B1(n_141),
.B2(n_166),
.Y(n_192)
);

BUFx24_ASAP7_75t_SL g209 ( 
.A(n_193),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_156),
.B(n_133),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_194),
.B(n_195),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_144),
.B(n_133),
.C(n_129),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_163),
.B(n_127),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_143),
.A2(n_124),
.B1(n_4),
.B2(n_5),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_198),
.A2(n_147),
.B1(n_7),
.B2(n_8),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_143),
.A2(n_3),
.B(n_4),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_186),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_SL g234 ( 
.A(n_201),
.B(n_202),
.C(n_212),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_179),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_203),
.B(n_222),
.Y(n_246)
);

INVx8_ASAP7_75t_L g207 ( 
.A(n_196),
.Y(n_207)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_207),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_181),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_178),
.B(n_159),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_213),
.B(n_220),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_215),
.A2(n_199),
.B1(n_180),
.B2(n_175),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_188),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_216),
.Y(n_236)
);

XOR2x2_ASAP7_75t_L g217 ( 
.A(n_183),
.B(n_157),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_217),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_192),
.A2(n_136),
.B1(n_160),
.B2(n_149),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_218),
.A2(n_219),
.B1(n_224),
.B2(n_196),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_172),
.A2(n_136),
.B1(n_138),
.B2(n_161),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_178),
.B(n_161),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_184),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_221),
.B(n_223),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_177),
.A2(n_139),
.B(n_142),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_194),
.A2(n_139),
.B(n_138),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_175),
.A2(n_161),
.B1(n_139),
.B2(n_152),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_168),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_225),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_168),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_226),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_200),
.B(n_169),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_228),
.B(n_235),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_208),
.B(n_171),
.C(n_182),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_229),
.B(n_232),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_231),
.A2(n_243),
.B1(n_247),
.B2(n_224),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_208),
.B(n_205),
.C(n_206),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_205),
.B(n_195),
.C(n_173),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_237),
.A2(n_215),
.B1(n_210),
.B2(n_219),
.Y(n_257)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_204),
.Y(n_238)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_238),
.Y(n_258)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_204),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_239),
.B(n_241),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_200),
.B(n_170),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_240),
.B(n_201),
.Y(n_264)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_220),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_214),
.A2(n_187),
.B1(n_191),
.B2(n_197),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_214),
.A2(n_197),
.B1(n_185),
.B2(n_198),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_206),
.B(n_203),
.C(n_217),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_248),
.B(n_211),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_248),
.B(n_217),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_249),
.B(n_250),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_252),
.A2(n_259),
.B1(n_261),
.B2(n_245),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_242),
.A2(n_222),
.B(n_211),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_253),
.B(n_262),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_238),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_256),
.B(n_264),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_257),
.B(n_246),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_231),
.A2(n_213),
.B1(n_218),
.B2(n_202),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_229),
.B(n_223),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_260),
.B(n_246),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_243),
.A2(n_221),
.B1(n_212),
.B2(n_226),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_242),
.A2(n_210),
.B(n_225),
.Y(n_262)
);

OR2x2_ASAP7_75t_L g263 ( 
.A(n_230),
.B(n_247),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_263),
.A2(n_245),
.B1(n_233),
.B2(n_241),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_239),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_265),
.B(n_227),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_266),
.A2(n_270),
.B1(n_277),
.B2(n_253),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_255),
.B(n_232),
.C(n_235),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_268),
.B(n_279),
.C(n_260),
.Y(n_280)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_269),
.Y(n_290)
);

AOI21xp33_ASAP7_75t_L g270 ( 
.A1(n_251),
.A2(n_236),
.B(n_234),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_271),
.B(n_273),
.Y(n_289)
);

BUFx12f_ASAP7_75t_SL g272 ( 
.A(n_263),
.Y(n_272)
);

XNOR2x1_ASAP7_75t_L g288 ( 
.A(n_272),
.B(n_6),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_262),
.B(n_233),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_275),
.B(n_244),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_252),
.A2(n_259),
.B1(n_261),
.B2(n_254),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_209),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_255),
.B(n_234),
.C(n_207),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_280),
.B(n_281),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_268),
.B(n_249),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_282),
.B(n_285),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_272),
.A2(n_254),
.B1(n_258),
.B2(n_250),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_283),
.A2(n_287),
.B1(n_275),
.B2(n_276),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_279),
.B(n_244),
.C(n_174),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_284),
.B(n_286),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_266),
.A2(n_152),
.B1(n_7),
.B2(n_9),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_288),
.A2(n_267),
.B(n_290),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_294),
.B(n_296),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_295),
.B(n_299),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_289),
.B(n_273),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_283),
.A2(n_277),
.B1(n_278),
.B2(n_274),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_297),
.B(n_298),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_288),
.A2(n_274),
.B1(n_152),
.B2(n_10),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_284),
.Y(n_299)
);

NOR2xp67_ASAP7_75t_SL g302 ( 
.A(n_291),
.B(n_280),
.Y(n_302)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_302),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_293),
.A2(n_282),
.B(n_285),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_303),
.B(n_305),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_297),
.A2(n_6),
.B(n_7),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_304),
.B(n_292),
.C(n_295),
.Y(n_306)
);

OR2x2_ASAP7_75t_L g311 ( 
.A(n_306),
.B(n_307),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_300),
.B(n_6),
.C(n_10),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_301),
.B(n_15),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_310),
.B(n_13),
.Y(n_313)
);

AOI322xp5_ASAP7_75t_L g312 ( 
.A1(n_309),
.A2(n_10),
.A3(n_11),
.B1(n_12),
.B2(n_13),
.C1(n_15),
.C2(n_308),
.Y(n_312)
);

AO21x2_ASAP7_75t_SL g315 ( 
.A1(n_312),
.A2(n_313),
.B(n_11),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_311),
.Y(n_314)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_314),
.Y(n_316)
);

FAx1_ASAP7_75t_SL g317 ( 
.A(n_316),
.B(n_315),
.CI(n_12),
.CON(n_317),
.SN(n_317)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_295),
.Y(n_318)
);


endmodule