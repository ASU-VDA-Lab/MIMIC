module fake_jpeg_18973_n_30 (n_3, n_2, n_1, n_0, n_4, n_30);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;

output n_30;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_5;
wire n_11;
wire n_17;
wire n_25;
wire n_29;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

INVx3_ASAP7_75t_L g5 ( 
.A(n_1),
.Y(n_5)
);

BUFx24_ASAP7_75t_L g6 ( 
.A(n_4),
.Y(n_6)
);

NAND2xp5_ASAP7_75t_L g7 ( 
.A(n_1),
.B(n_0),
.Y(n_7)
);

INVx2_ASAP7_75t_SL g8 ( 
.A(n_2),
.Y(n_8)
);

BUFx12_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

OAI22xp33_ASAP7_75t_L g10 ( 
.A1(n_5),
.A2(n_7),
.B1(n_8),
.B2(n_6),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_10),
.B(n_12),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

XNOR2xp5_ASAP7_75t_L g13 ( 
.A(n_7),
.B(n_0),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_13),
.B(n_14),
.Y(n_15)
);

INVx8_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_13),
.B(n_8),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_18),
.B(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_19),
.A2(n_11),
.B(n_9),
.Y(n_25)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_20),
.B(n_21),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_15),
.B(n_16),
.C(n_12),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_17),
.B(n_1),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_22),
.B(n_9),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_24),
.B(n_14),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_L g26 ( 
.A1(n_25),
.A2(n_21),
.B(n_9),
.Y(n_26)
);

OAI21xp33_ASAP7_75t_L g28 ( 
.A1(n_26),
.A2(n_27),
.B(n_23),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_28),
.B(n_2),
.C(n_3),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_29),
.B(n_3),
.C(n_4),
.Y(n_30)
);


endmodule