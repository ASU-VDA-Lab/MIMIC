module fake_jpeg_695_n_687 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_687);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_687;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_686;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

INVx2_ASAP7_75t_SL g22 ( 
.A(n_14),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx8_ASAP7_75t_SL g33 ( 
.A(n_2),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_12),
.Y(n_41)
);

BUFx8_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_9),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_12),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_12),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_9),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_7),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

BUFx10_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_15),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_6),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_13),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_59),
.Y(n_149)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g144 ( 
.A(n_60),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_61),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_31),
.B(n_8),
.C(n_18),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_62),
.B(n_65),
.Y(n_137)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_63),
.Y(n_134)
);

BUFx24_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g201 ( 
.A(n_64),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_28),
.B(n_8),
.Y(n_65)
);

BUFx12_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

CKINVDCx6p67_ASAP7_75t_R g157 ( 
.A(n_66),
.Y(n_157)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx8_ASAP7_75t_L g163 ( 
.A(n_67),
.Y(n_163)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_68),
.Y(n_133)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_69),
.Y(n_139)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_32),
.Y(n_70)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_70),
.Y(n_142)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_71),
.Y(n_141)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_72),
.Y(n_150)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_23),
.Y(n_73)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_73),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_74),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_26),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_75),
.Y(n_182)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_23),
.B(n_34),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_76),
.B(n_85),
.Y(n_138)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

INVx2_ASAP7_75t_SL g213 ( 
.A(n_77),
.Y(n_213)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_78),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_29),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_79),
.Y(n_208)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_32),
.Y(n_80)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_80),
.Y(n_151)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_34),
.Y(n_81)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_81),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_29),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_82),
.Y(n_214)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_27),
.Y(n_83)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_83),
.Y(n_162)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_27),
.Y(n_84)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_84),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_28),
.B(n_9),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_27),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g164 ( 
.A(n_86),
.Y(n_164)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_27),
.Y(n_87)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_87),
.Y(n_172)
);

AND2x6_ASAP7_75t_SL g88 ( 
.A(n_33),
.B(n_7),
.Y(n_88)
);

NAND2xp33_ASAP7_75t_SL g185 ( 
.A(n_88),
.B(n_126),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_30),
.B(n_10),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_89),
.B(n_90),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_30),
.B(n_10),
.Y(n_90)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_29),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_91),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_29),
.Y(n_92)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_92),
.Y(n_186)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_27),
.Y(n_93)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_93),
.Y(n_174)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_27),
.Y(n_94)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_94),
.Y(n_176)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_40),
.Y(n_95)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_95),
.Y(n_177)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_39),
.Y(n_96)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_96),
.Y(n_136)
);

BUFx8_ASAP7_75t_L g97 ( 
.A(n_39),
.Y(n_97)
);

BUFx2_ASAP7_75t_L g173 ( 
.A(n_97),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_38),
.Y(n_98)
);

INVx6_ASAP7_75t_L g215 ( 
.A(n_98),
.Y(n_215)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_36),
.Y(n_99)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_99),
.Y(n_168)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_40),
.Y(n_100)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_100),
.Y(n_148)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_38),
.Y(n_101)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_101),
.Y(n_158)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_37),
.Y(n_102)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_102),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_38),
.Y(n_103)
);

INVx6_ASAP7_75t_L g228 ( 
.A(n_103),
.Y(n_228)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_39),
.Y(n_104)
);

INVx6_ASAP7_75t_SL g171 ( 
.A(n_104),
.Y(n_171)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_36),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g187 ( 
.A(n_105),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_35),
.B(n_52),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_106),
.B(n_107),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_36),
.B(n_10),
.Y(n_107)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_40),
.Y(n_108)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_108),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_21),
.B(n_19),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_109),
.B(n_124),
.Y(n_140)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_58),
.Y(n_110)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_110),
.Y(n_167)
);

BUFx12f_ASAP7_75t_L g111 ( 
.A(n_38),
.Y(n_111)
);

INVx5_ASAP7_75t_L g211 ( 
.A(n_111),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_45),
.Y(n_112)
);

INVx6_ASAP7_75t_L g229 ( 
.A(n_112),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_35),
.B(n_6),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_113),
.B(n_128),
.Y(n_155)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_40),
.Y(n_114)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_114),
.Y(n_160)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_45),
.Y(n_115)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_115),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_45),
.Y(n_116)
);

INVx3_ASAP7_75t_SL g170 ( 
.A(n_116),
.Y(n_170)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_45),
.Y(n_117)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_117),
.Y(n_179)
);

INVx13_ASAP7_75t_L g118 ( 
.A(n_39),
.Y(n_118)
);

INVx6_ASAP7_75t_SL g198 ( 
.A(n_118),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_58),
.Y(n_119)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_119),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_58),
.A2(n_6),
.B1(n_18),
.B2(n_2),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_120),
.A2(n_55),
.B1(n_56),
.B2(n_24),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_58),
.Y(n_121)
);

INVx5_ASAP7_75t_L g218 ( 
.A(n_121),
.Y(n_218)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_22),
.Y(n_122)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_122),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_20),
.Y(n_123)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_123),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_21),
.B(n_11),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_22),
.Y(n_125)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_125),
.Y(n_194)
);

HAxp5_ASAP7_75t_SL g126 ( 
.A(n_54),
.B(n_0),
.CON(n_126),
.SN(n_126)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_20),
.Y(n_127)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_127),
.Y(n_195)
);

INVx4_ASAP7_75t_SL g128 ( 
.A(n_37),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_22),
.Y(n_129)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_129),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_20),
.Y(n_130)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_130),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_57),
.B(n_11),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_131),
.B(n_5),
.Y(n_145)
);

AOI21xp33_ASAP7_75t_L g132 ( 
.A1(n_24),
.A2(n_11),
.B(n_18),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_132),
.B(n_0),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_145),
.B(n_159),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_128),
.A2(n_22),
.B1(n_55),
.B2(n_44),
.Y(n_146)
);

OA22x2_ASAP7_75t_L g281 ( 
.A1(n_146),
.A2(n_197),
.B1(n_200),
.B2(n_206),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_107),
.B(n_57),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_61),
.A2(n_55),
.B1(n_44),
.B2(n_53),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_161),
.A2(n_169),
.B1(n_178),
.B2(n_204),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_165),
.B(n_0),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_76),
.A2(n_41),
.B1(n_52),
.B2(n_51),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_97),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_175),
.B(n_212),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_74),
.A2(n_55),
.B1(n_44),
.B2(n_53),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_67),
.B(n_50),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_181),
.B(n_189),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_184),
.A2(n_1),
.B1(n_14),
.B2(n_17),
.Y(n_313)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_78),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g299 ( 
.A(n_188),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_67),
.B(n_50),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_71),
.B(n_51),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_190),
.B(n_202),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_102),
.B(n_46),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_192),
.B(n_209),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_71),
.A2(n_25),
.B1(n_53),
.B2(n_49),
.Y(n_197)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_78),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g312 ( 
.A(n_199),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_126),
.A2(n_96),
.B1(n_86),
.B2(n_64),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_64),
.B(n_46),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_123),
.Y(n_203)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_203),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_59),
.A2(n_41),
.B1(n_56),
.B2(n_25),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_127),
.Y(n_205)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_205),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_101),
.A2(n_56),
.B1(n_25),
.B2(n_49),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_130),
.B(n_43),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_91),
.Y(n_212)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_104),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g317 ( 
.A(n_217),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_75),
.B(n_49),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_219),
.B(n_1),
.Y(n_298)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_79),
.Y(n_220)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_220),
.Y(n_234)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_118),
.Y(n_221)
);

INVx2_ASAP7_75t_SL g285 ( 
.A(n_221),
.Y(n_285)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_110),
.Y(n_222)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_222),
.Y(n_251)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_82),
.Y(n_223)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_223),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_101),
.A2(n_48),
.B1(n_43),
.B2(n_24),
.Y(n_224)
);

OA22x2_ASAP7_75t_L g311 ( 
.A1(n_224),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_311)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_92),
.Y(n_225)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_225),
.Y(n_252)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_98),
.Y(n_226)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_226),
.Y(n_257)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_103),
.Y(n_227)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_227),
.Y(n_259)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_112),
.Y(n_230)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_230),
.Y(n_269)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_116),
.Y(n_231)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_231),
.Y(n_284)
);

BUFx2_ASAP7_75t_L g233 ( 
.A(n_173),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g363 ( 
.A(n_233),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_171),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_235),
.B(n_238),
.Y(n_367)
);

INVx4_ASAP7_75t_SL g237 ( 
.A(n_198),
.Y(n_237)
);

INVx13_ASAP7_75t_L g321 ( 
.A(n_237),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_164),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_138),
.A2(n_111),
.B1(n_43),
.B2(n_48),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g322 ( 
.A1(n_240),
.A2(n_250),
.B1(n_253),
.B2(n_273),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_164),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_241),
.B(n_242),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_173),
.Y(n_242)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_201),
.Y(n_243)
);

INVx3_ASAP7_75t_L g343 ( 
.A(n_243),
.Y(n_343)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_201),
.Y(n_244)
);

INVx3_ASAP7_75t_L g359 ( 
.A(n_244),
.Y(n_359)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_141),
.Y(n_246)
);

INVx5_ASAP7_75t_L g352 ( 
.A(n_246),
.Y(n_352)
);

INVxp67_ASAP7_75t_SL g248 ( 
.A(n_157),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_248),
.Y(n_328)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_177),
.Y(n_249)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_249),
.Y(n_333)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_138),
.A2(n_155),
.B1(n_191),
.B2(n_195),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_155),
.A2(n_111),
.B1(n_48),
.B2(n_66),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g369 ( 
.A(n_254),
.B(n_279),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_157),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_255),
.B(n_258),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_157),
.Y(n_258)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_148),
.Y(n_260)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_260),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_181),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_261),
.B(n_263),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_189),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_179),
.Y(n_264)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_264),
.Y(n_341)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_196),
.Y(n_265)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_265),
.Y(n_345)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_135),
.Y(n_266)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_266),
.Y(n_329)
);

INVx6_ASAP7_75t_L g267 ( 
.A(n_152),
.Y(n_267)
);

INVx3_ASAP7_75t_L g366 ( 
.A(n_267),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_190),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_270),
.B(n_274),
.Y(n_379)
);

INVx5_ASAP7_75t_L g271 ( 
.A(n_163),
.Y(n_271)
);

INVx3_ASAP7_75t_L g373 ( 
.A(n_271),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_152),
.Y(n_272)
);

INVx6_ASAP7_75t_L g332 ( 
.A(n_272),
.Y(n_332)
);

AOI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_210),
.A2(n_121),
.B1(n_119),
.B2(n_47),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_187),
.Y(n_274)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_156),
.Y(n_276)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_276),
.Y(n_338)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_170),
.Y(n_277)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_277),
.Y(n_349)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_143),
.Y(n_278)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_278),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_187),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_153),
.Y(n_280)
);

INVx6_ASAP7_75t_L g350 ( 
.A(n_280),
.Y(n_350)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_183),
.Y(n_282)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_282),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_137),
.B(n_54),
.C(n_47),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_283),
.B(n_273),
.C(n_258),
.Y(n_380)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_167),
.Y(n_287)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_287),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_216),
.Y(n_288)
);

CKINVDCx14_ASAP7_75t_R g324 ( 
.A(n_288),
.Y(n_324)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_194),
.Y(n_289)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_289),
.Y(n_364)
);

BUFx3_ASAP7_75t_L g290 ( 
.A(n_158),
.Y(n_290)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_290),
.Y(n_365)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_202),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_291),
.B(n_296),
.Y(n_356)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_211),
.Y(n_292)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_292),
.Y(n_372)
);

OAI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_161),
.A2(n_54),
.B1(n_47),
.B2(n_37),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_293),
.A2(n_294),
.B1(n_310),
.B2(n_17),
.Y(n_355)
);

OAI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_178),
.A2(n_54),
.B1(n_1),
.B2(n_3),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_207),
.Y(n_295)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_295),
.Y(n_374)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_136),
.Y(n_296)
);

A2O1A1Ixp33_ASAP7_75t_L g297 ( 
.A1(n_165),
.A2(n_54),
.B(n_2),
.C(n_3),
.Y(n_297)
);

O2A1O1Ixp33_ASAP7_75t_L g331 ( 
.A1(n_297),
.A2(n_140),
.B(n_224),
.C(n_154),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_298),
.B(n_300),
.Y(n_375)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_180),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_154),
.B(n_13),
.Y(n_301)
);

OR2x2_ASAP7_75t_L g368 ( 
.A(n_301),
.B(n_302),
.Y(n_368)
);

NAND2x1_ASAP7_75t_L g302 ( 
.A(n_185),
.B(n_54),
.Y(n_302)
);

INVx4_ASAP7_75t_L g303 ( 
.A(n_160),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_303),
.Y(n_319)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_142),
.Y(n_304)
);

OR2x2_ASAP7_75t_L g376 ( 
.A(n_304),
.B(n_305),
.Y(n_376)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_150),
.Y(n_305)
);

AO22x2_ASAP7_75t_L g306 ( 
.A1(n_200),
.A2(n_218),
.B1(n_146),
.B2(n_168),
.Y(n_306)
);

AO22x1_ASAP7_75t_L g339 ( 
.A1(n_306),
.A2(n_182),
.B1(n_214),
.B2(n_208),
.Y(n_339)
);

AOI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_134),
.A2(n_13),
.B1(n_3),
.B2(n_4),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_SL g347 ( 
.A1(n_307),
.A2(n_311),
.B1(n_314),
.B2(n_315),
.Y(n_347)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_151),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_308),
.Y(n_326)
);

BUFx2_ASAP7_75t_L g309 ( 
.A(n_170),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_309),
.Y(n_342)
);

OAI22xp33_ASAP7_75t_SL g310 ( 
.A1(n_137),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_313),
.A2(n_147),
.B1(n_229),
.B2(n_228),
.Y(n_335)
);

INVx4_ASAP7_75t_L g314 ( 
.A(n_144),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_144),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_162),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_SL g370 ( 
.A1(n_316),
.A2(n_318),
.B1(n_233),
.B2(n_237),
.Y(n_370)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_193),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_302),
.A2(n_197),
.B(n_206),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g382 ( 
.A1(n_323),
.A2(n_334),
.B(n_340),
.Y(n_382)
);

AOI22xp33_ASAP7_75t_L g330 ( 
.A1(n_275),
.A2(n_213),
.B1(n_214),
.B2(n_208),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_330),
.A2(n_346),
.B1(n_348),
.B2(n_355),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_331),
.B(n_336),
.Y(n_388)
);

O2A1O1Ixp33_ASAP7_75t_L g334 ( 
.A1(n_297),
.A2(n_176),
.B(n_172),
.C(n_174),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_335),
.A2(n_351),
.B1(n_277),
.B2(n_309),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_310),
.B(n_147),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_283),
.B(n_133),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_337),
.B(n_377),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_339),
.B(n_361),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_250),
.A2(n_254),
.B(n_268),
.Y(n_340)
);

MAJx2_ASAP7_75t_L g344 ( 
.A(n_286),
.B(n_139),
.C(n_166),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_344),
.B(n_378),
.C(n_312),
.Y(n_426)
);

AOI22xp33_ASAP7_75t_L g346 ( 
.A1(n_293),
.A2(n_294),
.B1(n_239),
.B2(n_236),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_256),
.A2(n_215),
.B1(n_186),
.B2(n_182),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_313),
.A2(n_149),
.B1(n_232),
.B2(n_153),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_L g353 ( 
.A1(n_240),
.A2(n_213),
.B(n_149),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_L g411 ( 
.A1(n_353),
.A2(n_357),
.B(n_244),
.Y(n_411)
);

OAI22xp33_ASAP7_75t_SL g354 ( 
.A1(n_253),
.A2(n_232),
.B1(n_17),
.B2(n_19),
.Y(n_354)
);

AOI22xp33_ASAP7_75t_L g416 ( 
.A1(n_354),
.A2(n_353),
.B1(n_336),
.B2(n_324),
.Y(n_416)
);

O2A1O1Ixp33_ASAP7_75t_L g357 ( 
.A1(n_281),
.A2(n_19),
.B(n_306),
.C(n_311),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_306),
.A2(n_281),
.B1(n_301),
.B2(n_287),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_370),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_262),
.B(n_247),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_306),
.B(n_281),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_380),
.B(n_255),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_249),
.B(n_264),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_381),
.B(n_257),
.Y(n_390)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_320),
.Y(n_383)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_383),
.Y(n_447)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_320),
.Y(n_385)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_385),
.Y(n_453)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_381),
.Y(n_387)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_387),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_390),
.B(n_397),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_391),
.A2(n_404),
.B1(n_406),
.B2(n_407),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_367),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_393),
.B(n_405),
.Y(n_446)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_329),
.Y(n_394)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_394),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_339),
.A2(n_252),
.B1(n_265),
.B2(n_311),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_395),
.A2(n_425),
.B1(n_429),
.B2(n_430),
.Y(n_434)
);

INVx3_ASAP7_75t_L g396 ( 
.A(n_366),
.Y(n_396)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_396),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_337),
.B(n_234),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_344),
.B(n_251),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_398),
.B(n_409),
.C(n_427),
.Y(n_454)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_329),
.Y(n_399)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_399),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_331),
.B(n_284),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_400),
.B(n_410),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_327),
.Y(n_401)
);

INVxp33_ASAP7_75t_L g473 ( 
.A(n_401),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_356),
.B(n_243),
.Y(n_402)
);

AND2x2_ASAP7_75t_SL g458 ( 
.A(n_402),
.B(n_424),
.Y(n_458)
);

FAx1_ASAP7_75t_SL g403 ( 
.A(n_340),
.B(n_317),
.CI(n_307),
.CON(n_403),
.SN(n_403)
);

NOR2xp33_ASAP7_75t_SL g474 ( 
.A(n_403),
.B(n_352),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_361),
.A2(n_267),
.B1(n_272),
.B2(n_280),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_371),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_378),
.A2(n_259),
.B1(n_245),
.B2(n_269),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_322),
.A2(n_300),
.B1(n_318),
.B2(n_303),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_328),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_408),
.B(n_416),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_375),
.B(n_296),
.Y(n_410)
);

NAND2xp33_ASAP7_75t_SL g436 ( 
.A(n_411),
.B(n_413),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_L g412 ( 
.A1(n_355),
.A2(n_314),
.B1(n_292),
.B2(n_271),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_412),
.B(n_415),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_323),
.A2(n_285),
.B(n_299),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_332),
.Y(n_414)
);

INVxp67_ASAP7_75t_L g461 ( 
.A(n_414),
.Y(n_461)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_338),
.Y(n_415)
);

BUFx3_ASAP7_75t_L g417 ( 
.A(n_328),
.Y(n_417)
);

INVx11_ASAP7_75t_L g445 ( 
.A(n_417),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_377),
.B(n_285),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_SL g433 ( 
.A(n_418),
.B(n_319),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_375),
.B(n_278),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_419),
.B(n_420),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_375),
.B(n_246),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_379),
.B(n_290),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_421),
.B(n_343),
.Y(n_443)
);

AND2x2_ASAP7_75t_SL g422 ( 
.A(n_380),
.B(n_299),
.Y(n_422)
);

CKINVDCx14_ASAP7_75t_R g440 ( 
.A(n_422),
.Y(n_440)
);

INVx3_ASAP7_75t_L g423 ( 
.A(n_366),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_423),
.B(n_342),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_356),
.B(n_312),
.Y(n_424)
);

AOI22xp33_ASAP7_75t_L g425 ( 
.A1(n_339),
.A2(n_357),
.B1(n_326),
.B2(n_334),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_426),
.B(n_409),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_368),
.B(n_356),
.C(n_374),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_368),
.B(n_376),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_428),
.B(n_410),
.Y(n_450)
);

AOI22xp33_ASAP7_75t_L g429 ( 
.A1(n_326),
.A2(n_319),
.B1(n_342),
.B2(n_362),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_351),
.A2(n_325),
.B1(n_369),
.B2(n_347),
.Y(n_430)
);

O2A1O1Ixp33_ASAP7_75t_SL g431 ( 
.A1(n_369),
.A2(n_362),
.B(n_365),
.C(n_372),
.Y(n_431)
);

OA21x2_ASAP7_75t_L g459 ( 
.A1(n_431),
.A2(n_413),
.B(n_400),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_433),
.B(n_466),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_439),
.B(n_455),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_388),
.A2(n_376),
.B1(n_332),
.B2(n_350),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_441),
.A2(n_449),
.B1(n_468),
.B2(n_415),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_443),
.B(n_444),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_387),
.B(n_374),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_389),
.B(n_360),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_SL g505 ( 
.A(n_448),
.B(n_451),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_388),
.A2(n_350),
.B1(n_360),
.B2(n_338),
.Y(n_449)
);

INVx1_ASAP7_75t_SL g511 ( 
.A(n_450),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_389),
.B(n_364),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_390),
.Y(n_452)
);

INVx13_ASAP7_75t_L g500 ( 
.A(n_452),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_398),
.B(n_364),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_397),
.B(n_349),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_456),
.B(n_465),
.Y(n_499)
);

CKINVDCx16_ASAP7_75t_R g514 ( 
.A(n_459),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_408),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_462),
.B(n_436),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_L g463 ( 
.A1(n_411),
.A2(n_365),
.B(n_373),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_SL g506 ( 
.A1(n_463),
.A2(n_419),
.B(n_420),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_430),
.B(n_406),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_428),
.B(n_349),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_386),
.A2(n_373),
.B1(n_358),
.B2(n_372),
.Y(n_468)
);

XOR2x2_ASAP7_75t_L g469 ( 
.A(n_426),
.B(n_343),
.Y(n_469)
);

INVxp67_ASAP7_75t_L g487 ( 
.A(n_469),
.Y(n_487)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_470),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_401),
.B(n_358),
.Y(n_472)
);

NAND3xp33_ASAP7_75t_L g496 ( 
.A(n_472),
.B(n_427),
.C(n_424),
.Y(n_496)
);

OAI21xp5_ASAP7_75t_L g483 ( 
.A1(n_474),
.A2(n_382),
.B(n_428),
.Y(n_483)
);

BUFx5_ASAP7_75t_L g478 ( 
.A(n_445),
.Y(n_478)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_478),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_470),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_479),
.B(n_488),
.Y(n_547)
);

CKINVDCx16_ASAP7_75t_R g480 ( 
.A(n_472),
.Y(n_480)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_480),
.Y(n_526)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_447),
.Y(n_481)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_481),
.Y(n_515)
);

INVxp33_ASAP7_75t_L g482 ( 
.A(n_473),
.Y(n_482)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_482),
.Y(n_540)
);

OAI21xp5_ASAP7_75t_L g528 ( 
.A1(n_483),
.A2(n_495),
.B(n_497),
.Y(n_528)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_447),
.Y(n_484)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_484),
.Y(n_545)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_453),
.Y(n_485)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_485),
.Y(n_551)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_446),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_453),
.Y(n_489)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_489),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_462),
.B(n_421),
.Y(n_490)
);

CKINVDCx14_ASAP7_75t_R g522 ( 
.A(n_490),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_433),
.B(n_417),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_491),
.B(n_502),
.Y(n_538)
);

AND2x4_ASAP7_75t_L g530 ( 
.A(n_492),
.B(n_506),
.Y(n_530)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_460),
.Y(n_493)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_493),
.Y(n_536)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_460),
.Y(n_494)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_494),
.Y(n_537)
);

OAI21xp5_ASAP7_75t_L g495 ( 
.A1(n_436),
.A2(n_382),
.B(n_431),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_L g519 ( 
.A1(n_496),
.A2(n_507),
.B1(n_508),
.B2(n_464),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_L g497 ( 
.A1(n_474),
.A2(n_431),
.B(n_403),
.Y(n_497)
);

OAI21xp5_ASAP7_75t_L g498 ( 
.A1(n_459),
.A2(n_403),
.B(n_386),
.Y(n_498)
);

INVxp67_ASAP7_75t_L g517 ( 
.A(n_498),
.Y(n_517)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_471),
.Y(n_501)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_501),
.Y(n_543)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_444),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g503 ( 
.A(n_439),
.B(n_422),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_503),
.B(n_504),
.C(n_455),
.Y(n_531)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_454),
.B(n_422),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_L g507 ( 
.A1(n_434),
.A2(n_386),
.B1(n_395),
.B2(n_384),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_L g508 ( 
.A1(n_434),
.A2(n_391),
.B1(n_392),
.B2(n_407),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_509),
.B(n_512),
.Y(n_532)
);

OAI21xp5_ASAP7_75t_L g510 ( 
.A1(n_459),
.A2(n_392),
.B(n_402),
.Y(n_510)
);

INVxp67_ASAP7_75t_L g520 ( 
.A(n_510),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_L g512 ( 
.A1(n_459),
.A2(n_402),
.B(n_424),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_467),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_513),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_SL g516 ( 
.A1(n_514),
.A2(n_465),
.B1(n_464),
.B2(n_452),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_SL g582 ( 
.A1(n_516),
.A2(n_525),
.B1(n_529),
.B2(n_533),
.Y(n_582)
);

OAI22xp5_ASAP7_75t_L g568 ( 
.A1(n_519),
.A2(n_549),
.B1(n_438),
.B2(n_508),
.Y(n_568)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_504),
.B(n_454),
.Y(n_523)
);

XOR2xp5_ASAP7_75t_L g560 ( 
.A(n_523),
.B(n_531),
.Y(n_560)
);

CKINVDCx16_ASAP7_75t_R g524 ( 
.A(n_492),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_524),
.B(n_534),
.Y(n_578)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_507),
.A2(n_463),
.B1(n_457),
.B2(n_441),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_L g529 ( 
.A1(n_514),
.A2(n_457),
.B1(n_449),
.B2(n_437),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_SL g533 ( 
.A1(n_499),
.A2(n_432),
.B1(n_437),
.B2(n_435),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_500),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g535 ( 
.A(n_486),
.B(n_469),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g562 ( 
.A(n_535),
.B(n_539),
.Y(n_562)
);

XNOR2xp5_ASAP7_75t_L g539 ( 
.A(n_486),
.B(n_469),
.Y(n_539)
);

OAI22xp5_ASAP7_75t_SL g541 ( 
.A1(n_499),
.A2(n_432),
.B1(n_435),
.B2(n_438),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_SL g583 ( 
.A1(n_541),
.A2(n_542),
.B1(n_550),
.B2(n_493),
.Y(n_583)
);

AOI22xp5_ASAP7_75t_L g542 ( 
.A1(n_502),
.A2(n_438),
.B1(n_468),
.B2(n_440),
.Y(n_542)
);

CKINVDCx16_ASAP7_75t_R g544 ( 
.A(n_492),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_544),
.B(n_546),
.Y(n_566)
);

CKINVDCx20_ASAP7_75t_R g546 ( 
.A(n_500),
.Y(n_546)
);

XNOR2xp5_ASAP7_75t_L g548 ( 
.A(n_503),
.B(n_451),
.Y(n_548)
);

XNOR2xp5_ASAP7_75t_L g580 ( 
.A(n_548),
.B(n_471),
.Y(n_580)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_513),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_SL g550 ( 
.A1(n_498),
.A2(n_509),
.B1(n_497),
.B2(n_495),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_487),
.B(n_505),
.C(n_450),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_552),
.B(n_487),
.C(n_483),
.Y(n_553)
);

XNOR2xp5_ASAP7_75t_L g599 ( 
.A(n_553),
.B(n_581),
.Y(n_599)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_547),
.Y(n_554)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_554),
.Y(n_593)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_523),
.B(n_505),
.C(n_511),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g587 ( 
.A(n_555),
.B(n_557),
.C(n_558),
.Y(n_587)
);

XNOR2xp5_ASAP7_75t_SL g556 ( 
.A(n_535),
.B(n_511),
.Y(n_556)
);

XNOR2xp5_ASAP7_75t_SL g594 ( 
.A(n_556),
.B(n_570),
.Y(n_594)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_531),
.B(n_450),
.C(n_476),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_539),
.B(n_476),
.C(n_512),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_540),
.Y(n_559)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_559),
.Y(n_609)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_547),
.Y(n_561)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_561),
.Y(n_610)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_552),
.B(n_448),
.C(n_458),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g588 ( 
.A(n_563),
.B(n_567),
.C(n_571),
.Y(n_588)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_538),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_564),
.B(n_565),
.Y(n_598)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_521),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_548),
.B(n_458),
.C(n_479),
.Y(n_567)
);

OAI22xp5_ASAP7_75t_L g590 ( 
.A1(n_568),
.A2(n_577),
.B1(n_584),
.B2(n_572),
.Y(n_590)
);

OAI22xp5_ASAP7_75t_SL g569 ( 
.A1(n_525),
.A2(n_510),
.B1(n_475),
.B2(n_477),
.Y(n_569)
);

AOI22xp5_ASAP7_75t_SL g603 ( 
.A1(n_569),
.A2(n_583),
.B1(n_541),
.B2(n_543),
.Y(n_603)
);

XNOR2xp5_ASAP7_75t_SL g570 ( 
.A(n_528),
.B(n_466),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_517),
.B(n_458),
.C(n_506),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_517),
.B(n_458),
.C(n_475),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g596 ( 
.A(n_572),
.B(n_573),
.C(n_533),
.Y(n_596)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_528),
.B(n_442),
.C(n_456),
.Y(n_573)
);

XNOR2xp5_ASAP7_75t_SL g574 ( 
.A(n_550),
.B(n_442),
.Y(n_574)
);

XNOR2xp5_ASAP7_75t_SL g602 ( 
.A(n_574),
.B(n_579),
.Y(n_602)
);

XNOR2x1_ASAP7_75t_L g575 ( 
.A(n_532),
.B(n_443),
.Y(n_575)
);

XOR2xp5_ASAP7_75t_L g589 ( 
.A(n_575),
.B(n_580),
.Y(n_589)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_527),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_576),
.B(n_537),
.Y(n_591)
);

OAI22xp5_ASAP7_75t_L g577 ( 
.A1(n_522),
.A2(n_488),
.B1(n_501),
.B2(n_494),
.Y(n_577)
);

XNOR2xp5_ASAP7_75t_SL g579 ( 
.A(n_532),
.B(n_516),
.Y(n_579)
);

XNOR2xp5_ASAP7_75t_L g581 ( 
.A(n_542),
.B(n_489),
.Y(n_581)
);

OAI22xp5_ASAP7_75t_L g584 ( 
.A1(n_526),
.A2(n_485),
.B1(n_484),
.B2(n_481),
.Y(n_584)
);

OAI22xp5_ASAP7_75t_SL g585 ( 
.A1(n_582),
.A2(n_529),
.B1(n_532),
.B2(n_520),
.Y(n_585)
);

AOI22xp5_ASAP7_75t_L g614 ( 
.A1(n_585),
.A2(n_608),
.B1(n_581),
.B2(n_553),
.Y(n_614)
);

AOI21xp5_ASAP7_75t_L g586 ( 
.A1(n_575),
.A2(n_520),
.B(n_530),
.Y(n_586)
);

OAI22xp5_ASAP7_75t_L g611 ( 
.A1(n_586),
.A2(n_597),
.B1(n_604),
.B2(n_573),
.Y(n_611)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_590),
.Y(n_613)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_591),
.Y(n_615)
);

OAI21xp5_ASAP7_75t_SL g592 ( 
.A1(n_579),
.A2(n_530),
.B(n_518),
.Y(n_592)
);

MAJx2_ASAP7_75t_L g629 ( 
.A(n_592),
.B(n_596),
.C(n_445),
.Y(n_629)
);

INVxp67_ASAP7_75t_L g595 ( 
.A(n_566),
.Y(n_595)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_595),
.Y(n_618)
);

OAI22xp5_ASAP7_75t_L g597 ( 
.A1(n_578),
.A2(n_536),
.B1(n_527),
.B2(n_543),
.Y(n_597)
);

XNOR2xp5_ASAP7_75t_L g600 ( 
.A(n_557),
.B(n_530),
.Y(n_600)
);

XNOR2xp5_ASAP7_75t_L g617 ( 
.A(n_600),
.B(n_601),
.Y(n_617)
);

XNOR2xp5_ASAP7_75t_L g601 ( 
.A(n_558),
.B(n_530),
.Y(n_601)
);

OAI22xp5_ASAP7_75t_SL g625 ( 
.A1(n_603),
.A2(n_556),
.B1(n_423),
.B2(n_414),
.Y(n_625)
);

AOI21xp5_ASAP7_75t_L g604 ( 
.A1(n_571),
.A2(n_515),
.B(n_537),
.Y(n_604)
);

CKINVDCx20_ASAP7_75t_R g605 ( 
.A(n_569),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_605),
.B(n_607),
.Y(n_621)
);

XNOR2xp5_ASAP7_75t_L g606 ( 
.A(n_567),
.B(n_515),
.Y(n_606)
);

XNOR2xp5_ASAP7_75t_L g622 ( 
.A(n_606),
.B(n_563),
.Y(n_622)
);

MAJIxp5_ASAP7_75t_L g607 ( 
.A(n_560),
.B(n_467),
.C(n_536),
.Y(n_607)
);

OAI22xp5_ASAP7_75t_SL g608 ( 
.A1(n_574),
.A2(n_551),
.B1(n_545),
.B2(n_513),
.Y(n_608)
);

OR2x2_ASAP7_75t_L g641 ( 
.A(n_611),
.B(n_629),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_607),
.B(n_580),
.Y(n_612)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_612),
.Y(n_634)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_614),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_595),
.B(n_461),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_SL g645 ( 
.A(n_616),
.B(n_619),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_598),
.B(n_596),
.Y(n_619)
);

MAJIxp5_ASAP7_75t_L g620 ( 
.A(n_588),
.B(n_560),
.C(n_562),
.Y(n_620)
);

MAJIxp5_ASAP7_75t_L g633 ( 
.A(n_620),
.B(n_626),
.C(n_622),
.Y(n_633)
);

XNOR2xp5_ASAP7_75t_L g632 ( 
.A(n_622),
.B(n_625),
.Y(n_632)
);

AOI22xp5_ASAP7_75t_L g623 ( 
.A1(n_585),
.A2(n_570),
.B1(n_555),
.B2(n_562),
.Y(n_623)
);

OAI22xp5_ASAP7_75t_SL g646 ( 
.A1(n_623),
.A2(n_602),
.B1(n_589),
.B2(n_594),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_SL g624 ( 
.A(n_587),
.B(n_396),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_624),
.B(n_628),
.Y(n_637)
);

MAJIxp5_ASAP7_75t_L g626 ( 
.A(n_588),
.B(n_345),
.C(n_333),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_609),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_627),
.B(n_610),
.Y(n_640)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_608),
.Y(n_628)
);

XNOR2xp5_ASAP7_75t_L g630 ( 
.A(n_599),
.B(n_478),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_630),
.B(n_631),
.Y(n_639)
);

BUFx24_ASAP7_75t_SL g631 ( 
.A(n_604),
.Y(n_631)
);

XNOR2xp5_ASAP7_75t_L g650 ( 
.A(n_633),
.B(n_630),
.Y(n_650)
);

MAJIxp5_ASAP7_75t_L g635 ( 
.A(n_620),
.B(n_606),
.C(n_587),
.Y(n_635)
);

AOI21xp5_ASAP7_75t_L g655 ( 
.A1(n_635),
.A2(n_643),
.B(n_644),
.Y(n_655)
);

XOR2xp5_ASAP7_75t_L g638 ( 
.A(n_617),
.B(n_601),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_638),
.B(n_646),
.Y(n_659)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_640),
.Y(n_654)
);

AOI21xp5_ASAP7_75t_L g642 ( 
.A1(n_621),
.A2(n_592),
.B(n_586),
.Y(n_642)
);

OAI21xp5_ASAP7_75t_L g656 ( 
.A1(n_642),
.A2(n_641),
.B(n_649),
.Y(n_656)
);

OAI21xp5_ASAP7_75t_L g643 ( 
.A1(n_614),
.A2(n_603),
.B(n_593),
.Y(n_643)
);

MAJIxp5_ASAP7_75t_L g644 ( 
.A(n_617),
.B(n_599),
.C(n_600),
.Y(n_644)
);

MAJIxp5_ASAP7_75t_L g647 ( 
.A(n_612),
.B(n_589),
.C(n_602),
.Y(n_647)
);

AOI21xp5_ASAP7_75t_L g661 ( 
.A1(n_647),
.A2(n_635),
.B(n_643),
.Y(n_661)
);

OAI22xp5_ASAP7_75t_L g648 ( 
.A1(n_613),
.A2(n_594),
.B1(n_352),
.B2(n_359),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_648),
.B(n_629),
.Y(n_651)
);

OA21x2_ASAP7_75t_L g649 ( 
.A1(n_625),
.A2(n_359),
.B(n_345),
.Y(n_649)
);

AOI22xp5_ASAP7_75t_L g662 ( 
.A1(n_649),
.A2(n_642),
.B1(n_640),
.B2(n_637),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_650),
.B(n_652),
.Y(n_667)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_651),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_645),
.B(n_618),
.Y(n_652)
);

XOR2xp5_ASAP7_75t_L g653 ( 
.A(n_632),
.B(n_623),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_653),
.B(n_663),
.Y(n_668)
);

OR2x2_ASAP7_75t_L g671 ( 
.A(n_656),
.B(n_632),
.Y(n_671)
);

OAI22xp5_ASAP7_75t_SL g657 ( 
.A1(n_636),
.A2(n_615),
.B1(n_626),
.B2(n_341),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_657),
.B(n_658),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_SL g658 ( 
.A(n_639),
.B(n_333),
.Y(n_658)
);

OAI21xp5_ASAP7_75t_SL g660 ( 
.A1(n_634),
.A2(n_321),
.B(n_341),
.Y(n_660)
);

OAI21xp5_ASAP7_75t_SL g666 ( 
.A1(n_660),
.A2(n_661),
.B(n_641),
.Y(n_666)
);

AOI22xp5_ASAP7_75t_L g670 ( 
.A1(n_662),
.A2(n_656),
.B1(n_654),
.B2(n_649),
.Y(n_670)
);

BUFx24_ASAP7_75t_SL g663 ( 
.A(n_636),
.Y(n_663)
);

MAJIxp5_ASAP7_75t_L g664 ( 
.A(n_650),
.B(n_633),
.C(n_644),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_664),
.B(n_666),
.Y(n_674)
);

OAI21xp5_ASAP7_75t_SL g678 ( 
.A1(n_670),
.A2(n_671),
.B(n_646),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_655),
.B(n_638),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_672),
.B(n_659),
.Y(n_675)
);

MAJIxp5_ASAP7_75t_L g673 ( 
.A(n_664),
.B(n_659),
.C(n_653),
.Y(n_673)
);

XNOR2xp5_ASAP7_75t_L g681 ( 
.A(n_673),
.B(n_670),
.Y(n_681)
);

AOI21xp33_ASAP7_75t_L g680 ( 
.A1(n_675),
.A2(n_677),
.B(n_678),
.Y(n_680)
);

INVx6_ASAP7_75t_L g676 ( 
.A(n_667),
.Y(n_676)
);

AOI21xp5_ASAP7_75t_L g679 ( 
.A1(n_676),
.A2(n_665),
.B(n_669),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_668),
.B(n_662),
.Y(n_677)
);

OAI21xp5_ASAP7_75t_L g682 ( 
.A1(n_679),
.A2(n_674),
.B(n_678),
.Y(n_682)
);

AOI21xp5_ASAP7_75t_L g683 ( 
.A1(n_681),
.A2(n_671),
.B(n_647),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_682),
.Y(n_684)
);

MAJIxp5_ASAP7_75t_L g685 ( 
.A(n_684),
.B(n_683),
.C(n_680),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_685),
.B(n_363),
.Y(n_686)
);

AOI21xp5_ASAP7_75t_L g687 ( 
.A1(n_686),
.A2(n_321),
.B(n_363),
.Y(n_687)
);


endmodule