module real_aes_9855_n_266 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_266);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_266;
wire n_476;
wire n_887;
wire n_599;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1441;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_1382;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_619;
wire n_1095;
wire n_1284;
wire n_1250;
wire n_360;
wire n_1465;
wire n_859;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_411;
wire n_498;
wire n_1397;
wire n_765;
wire n_648;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_337;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_1392;
wire n_665;
wire n_991;
wire n_667;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_1014;
wire n_742;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1386;
wire n_406;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_985;
wire n_777;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_1179;
wire n_334;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_1462;
wire n_701;
wire n_809;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_689;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_1431;
wire n_721;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1162;
wire n_1463;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_285;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_1475;
wire n_977;
wire n_943;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_1470;
wire n_332;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1373;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_267;
wire n_1017;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1414;
wire n_1241;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_273;
wire n_1038;
wire n_276;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1191;
wire n_705;
wire n_1206;
wire n_1270;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1143;
wire n_929;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_1343;
wire n_1457;
wire n_719;
wire n_465;
wire n_1156;
wire n_988;
wire n_1466;
wire n_1396;
wire n_921;
wire n_1176;
wire n_640;
wire n_1151;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1420;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_372;
wire n_892;
wire n_578;
wire n_938;
wire n_327;
wire n_774;
wire n_559;
wire n_1049;
wire n_466;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_1100;
wire n_398;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_969;
wire n_1009;
wire n_1202;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_269;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_275;
wire n_536;
wire n_851;
wire n_470;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1436;
wire n_793;
wire n_1390;
wire n_272;
wire n_1412;
wire n_757;
wire n_803;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_1097;
wire n_703;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
INVx1_ASAP7_75t_L g557 ( .A(n_0), .Y(n_557) );
OAI22xp5_ASAP7_75t_L g603 ( .A1(n_0), .A2(n_164), .B1(n_281), .B2(n_299), .Y(n_603) );
AOI22xp33_ASAP7_75t_L g642 ( .A1(n_1), .A2(n_231), .B1(n_479), .B2(n_643), .Y(n_642) );
AOI22xp33_ASAP7_75t_L g662 ( .A1(n_1), .A2(n_231), .B1(n_321), .B2(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g753 ( .A(n_2), .Y(n_753) );
AOI22xp33_ASAP7_75t_L g765 ( .A1(n_2), .A2(n_141), .B1(n_412), .B2(n_766), .Y(n_765) );
INVx1_ASAP7_75t_L g1399 ( .A(n_3), .Y(n_1399) );
INVx1_ASAP7_75t_L g1218 ( .A(n_4), .Y(n_1218) );
AOI22xp33_ASAP7_75t_L g774 ( .A1(n_5), .A2(n_14), .B1(n_564), .B2(n_775), .Y(n_774) );
INVx1_ASAP7_75t_L g782 ( .A(n_5), .Y(n_782) );
INVx1_ASAP7_75t_L g863 ( .A(n_6), .Y(n_863) );
OAI22xp5_ASAP7_75t_L g923 ( .A1(n_7), .A2(n_173), .B1(n_529), .B2(n_533), .Y(n_923) );
AOI22xp33_ASAP7_75t_L g947 ( .A1(n_7), .A2(n_173), .B1(n_895), .B2(n_944), .Y(n_947) );
INVx1_ASAP7_75t_L g1057 ( .A(n_8), .Y(n_1057) );
INVx1_ASAP7_75t_L g1109 ( .A(n_9), .Y(n_1109) );
HB1xp67_ASAP7_75t_L g280 ( .A(n_10), .Y(n_280) );
INVx1_ASAP7_75t_L g433 ( .A(n_10), .Y(n_433) );
AND2x2_ASAP7_75t_L g1406 ( .A(n_10), .B(n_302), .Y(n_1406) );
NAND2xp5_ASAP7_75t_L g1420 ( .A(n_10), .B(n_199), .Y(n_1420) );
INVxp33_ASAP7_75t_L g1392 ( .A(n_11), .Y(n_1392) );
AOI21xp5_ASAP7_75t_L g1430 ( .A1(n_11), .A2(n_1028), .B(n_1431), .Y(n_1430) );
INVx1_ASAP7_75t_L g1396 ( .A(n_12), .Y(n_1396) );
OAI21xp33_ASAP7_75t_SL g686 ( .A1(n_13), .A2(n_544), .B(n_687), .Y(n_686) );
AOI22xp33_ASAP7_75t_L g721 ( .A1(n_13), .A2(n_124), .B1(n_722), .B2(n_724), .Y(n_721) );
INVx1_ASAP7_75t_L g783 ( .A(n_14), .Y(n_783) );
INVx1_ASAP7_75t_L g1401 ( .A(n_15), .Y(n_1401) );
OAI221xp5_ASAP7_75t_L g1413 ( .A1(n_15), .A2(n_264), .B1(n_1414), .B2(n_1421), .C(n_1423), .Y(n_1413) );
AOI22xp33_ASAP7_75t_L g934 ( .A1(n_16), .A2(n_207), .B1(n_412), .B2(n_663), .Y(n_934) );
AOI22xp33_ASAP7_75t_L g940 ( .A1(n_16), .A2(n_207), .B1(n_941), .B2(n_942), .Y(n_940) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_17), .A2(n_255), .B1(n_459), .B2(n_520), .Y(n_519) );
OAI22xp5_ASAP7_75t_L g528 ( .A1(n_17), .A2(n_255), .B1(n_529), .B2(n_533), .Y(n_528) );
INVx1_ASAP7_75t_L g691 ( .A(n_18), .Y(n_691) );
OAI222xp33_ASAP7_75t_L g699 ( .A1(n_18), .A2(n_29), .B1(n_253), .B2(n_327), .C1(n_496), .C2(n_669), .Y(n_699) );
AO22x2_ASAP7_75t_L g850 ( .A1(n_19), .A2(n_851), .B1(n_904), .B2(n_905), .Y(n_850) );
INVx1_ASAP7_75t_L g904 ( .A(n_19), .Y(n_904) );
AOI22xp33_ASAP7_75t_L g819 ( .A1(n_20), .A2(n_132), .B1(n_820), .B2(n_821), .Y(n_819) );
AOI22xp33_ASAP7_75t_L g836 ( .A1(n_20), .A2(n_132), .B1(n_837), .B2(n_839), .Y(n_836) );
CKINVDCx5p33_ASAP7_75t_R g747 ( .A(n_21), .Y(n_747) );
AOI22xp33_ASAP7_75t_SL g883 ( .A1(n_22), .A2(n_254), .B1(n_409), .B2(n_884), .Y(n_883) );
AOI22xp33_ASAP7_75t_L g891 ( .A1(n_22), .A2(n_254), .B1(n_376), .B2(n_738), .Y(n_891) );
INVx1_ASAP7_75t_L g751 ( .A(n_23), .Y(n_751) );
AOI22xp33_ASAP7_75t_L g762 ( .A1(n_23), .A2(n_263), .B1(n_763), .B2(n_764), .Y(n_762) );
AO221x2_ASAP7_75t_L g1189 ( .A1(n_24), .A2(n_58), .B1(n_1173), .B2(n_1182), .C(n_1190), .Y(n_1189) );
INVx1_ASAP7_75t_L g1206 ( .A(n_25), .Y(n_1206) );
INVxp67_ASAP7_75t_SL g814 ( .A(n_26), .Y(n_814) );
AOI22xp33_ASAP7_75t_L g844 ( .A1(n_26), .A2(n_204), .B1(n_770), .B2(n_845), .Y(n_844) );
INVxp33_ASAP7_75t_L g332 ( .A(n_27), .Y(n_332) );
AOI22xp33_ASAP7_75t_L g461 ( .A1(n_27), .A2(n_226), .B1(n_436), .B2(n_462), .Y(n_461) );
INVx2_ASAP7_75t_L g350 ( .A(n_28), .Y(n_350) );
AOI22xp33_ASAP7_75t_SL g737 ( .A1(n_29), .A2(n_171), .B1(n_731), .B2(n_738), .Y(n_737) );
AOI22xp33_ASAP7_75t_SL g1020 ( .A1(n_30), .A2(n_80), .B1(n_719), .B2(n_829), .Y(n_1020) );
AOI22xp33_ASAP7_75t_L g1033 ( .A1(n_30), .A2(n_80), .B1(n_736), .B2(n_740), .Y(n_1033) );
INVx1_ASAP7_75t_L g1191 ( .A(n_31), .Y(n_1191) );
CKINVDCx5p33_ASAP7_75t_R g547 ( .A(n_32), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g956 ( .A1(n_33), .A2(n_228), .B1(n_646), .B2(n_957), .Y(n_956) );
INVxp67_ASAP7_75t_SL g984 ( .A(n_33), .Y(n_984) );
INVxp67_ASAP7_75t_SL g1407 ( .A(n_34), .Y(n_1407) );
AOI22xp33_ASAP7_75t_L g1456 ( .A1(n_34), .A2(n_251), .B1(n_832), .B2(n_845), .Y(n_1456) );
AOI22xp33_ASAP7_75t_L g966 ( .A1(n_35), .A2(n_194), .B1(n_438), .B2(n_967), .Y(n_966) );
OAI211xp5_ASAP7_75t_SL g970 ( .A1(n_35), .A2(n_338), .B(n_971), .C(n_974), .Y(n_970) );
BUFx2_ASAP7_75t_L g343 ( .A(n_36), .Y(n_343) );
BUFx2_ASAP7_75t_L g396 ( .A(n_36), .Y(n_396) );
INVx1_ASAP7_75t_L g431 ( .A(n_36), .Y(n_431) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_37), .A2(n_49), .B1(n_562), .B2(n_565), .Y(n_561) );
OAI211xp5_ASAP7_75t_L g604 ( .A1(n_37), .A2(n_338), .B(n_605), .C(n_608), .Y(n_604) );
INVx1_ASAP7_75t_L g1251 ( .A(n_38), .Y(n_1251) );
AOI22xp33_ASAP7_75t_SL g657 ( .A1(n_39), .A2(n_110), .B1(n_459), .B2(n_658), .Y(n_657) );
INVxp67_ASAP7_75t_L g672 ( .A(n_39), .Y(n_672) );
INVx1_ASAP7_75t_L g693 ( .A(n_40), .Y(n_693) );
OAI22xp5_ASAP7_75t_L g698 ( .A1(n_40), .A2(n_171), .B1(n_281), .B2(n_299), .Y(n_698) );
INVxp33_ASAP7_75t_L g1394 ( .A(n_41), .Y(n_1394) );
AOI221xp5_ASAP7_75t_L g1428 ( .A1(n_41), .A2(n_97), .B1(n_722), .B2(n_933), .C(n_1429), .Y(n_1428) );
AOI22xp33_ASAP7_75t_L g954 ( .A1(n_42), .A2(n_179), .B1(n_412), .B2(n_648), .Y(n_954) );
AOI22xp33_ASAP7_75t_L g960 ( .A1(n_42), .A2(n_179), .B1(n_479), .B2(n_656), .Y(n_960) );
INVxp67_ASAP7_75t_SL g796 ( .A(n_43), .Y(n_796) );
OAI22xp5_ASAP7_75t_L g811 ( .A1(n_43), .A2(n_123), .B1(n_327), .B2(n_812), .Y(n_811) );
INVxp33_ASAP7_75t_SL g1000 ( .A(n_44), .Y(n_1000) );
AOI22xp33_ASAP7_75t_SL g1037 ( .A1(n_44), .A2(n_50), .B1(n_1038), .B2(n_1039), .Y(n_1037) );
INVx1_ASAP7_75t_L g1017 ( .A(n_45), .Y(n_1017) );
AOI22xp33_ASAP7_75t_L g1026 ( .A1(n_45), .A2(n_172), .B1(n_320), .B2(n_1027), .Y(n_1026) );
INVx1_ASAP7_75t_L g374 ( .A(n_46), .Y(n_374) );
AOI22xp33_ASAP7_75t_L g425 ( .A1(n_46), .A2(n_143), .B1(n_408), .B2(n_426), .Y(n_425) );
CKINVDCx16_ASAP7_75t_R g1203 ( .A(n_47), .Y(n_1203) );
INVx1_ASAP7_75t_L g1247 ( .A(n_48), .Y(n_1247) );
OAI22xp5_ASAP7_75t_L g611 ( .A1(n_49), .A2(n_106), .B1(n_529), .B2(n_533), .Y(n_611) );
INVxp33_ASAP7_75t_SL g1001 ( .A(n_50), .Y(n_1001) );
INVx1_ASAP7_75t_L g857 ( .A(n_51), .Y(n_857) );
INVx1_ASAP7_75t_L g1088 ( .A(n_52), .Y(n_1088) );
OAI211xp5_ASAP7_75t_L g1092 ( .A1(n_52), .A2(n_480), .B(n_544), .C(n_1093), .Y(n_1092) );
XNOR2xp5_ASAP7_75t_L g908 ( .A(n_53), .B(n_909), .Y(n_908) );
AOI22xp33_ASAP7_75t_L g407 ( .A1(n_54), .A2(n_145), .B1(n_408), .B2(n_412), .Y(n_407) );
AOI22xp33_ASAP7_75t_L g435 ( .A1(n_54), .A2(n_145), .B1(n_436), .B2(n_438), .Y(n_435) );
INVxp33_ASAP7_75t_SL g1008 ( .A(n_55), .Y(n_1008) );
AOI22xp33_ASAP7_75t_L g1036 ( .A1(n_55), .A2(n_56), .B1(n_754), .B2(n_837), .Y(n_1036) );
INVx1_ASAP7_75t_L g1003 ( .A(n_56), .Y(n_1003) );
AOI22xp33_ASAP7_75t_L g1124 ( .A1(n_57), .A2(n_62), .B1(n_1060), .B2(n_1125), .Y(n_1124) );
AOI22xp33_ASAP7_75t_L g1137 ( .A1(n_57), .A2(n_62), .B1(n_400), .B2(n_1138), .Y(n_1137) );
AOI22xp33_ASAP7_75t_L g655 ( .A1(n_59), .A2(n_233), .B1(n_438), .B2(n_656), .Y(n_655) );
INVxp33_ASAP7_75t_L g674 ( .A(n_59), .Y(n_674) );
AOI22xp33_ASAP7_75t_L g958 ( .A1(n_60), .A2(n_221), .B1(n_412), .B2(n_663), .Y(n_958) );
INVx1_ASAP7_75t_L g981 ( .A(n_60), .Y(n_981) );
OAI22xp5_ASAP7_75t_L g469 ( .A1(n_61), .A2(n_82), .B1(n_470), .B2(n_475), .Y(n_469) );
INVx1_ASAP7_75t_L g502 ( .A(n_61), .Y(n_502) );
INVx1_ASAP7_75t_L g1152 ( .A(n_63), .Y(n_1152) );
OAI22xp33_ASAP7_75t_L g484 ( .A1(n_64), .A2(n_244), .B1(n_485), .B2(n_486), .Y(n_484) );
AOI221xp5_ASAP7_75t_L g500 ( .A1(n_64), .A2(n_244), .B1(n_400), .B2(n_422), .C(n_501), .Y(n_500) );
INVxp33_ASAP7_75t_SL g1013 ( .A(n_65), .Y(n_1013) );
AOI22xp33_ASAP7_75t_L g1023 ( .A1(n_65), .A2(n_142), .B1(n_719), .B2(n_1024), .Y(n_1023) );
CKINVDCx16_ASAP7_75t_R g1165 ( .A(n_66), .Y(n_1165) );
INVx1_ASAP7_75t_L g600 ( .A(n_67), .Y(n_600) );
OAI211xp5_ASAP7_75t_SL g615 ( .A1(n_67), .A2(n_386), .B(n_616), .C(n_618), .Y(n_615) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_68), .A2(n_210), .B1(n_706), .B2(n_709), .Y(n_705) );
AOI22xp33_ASAP7_75t_L g728 ( .A1(n_68), .A2(n_222), .B1(n_729), .B2(n_731), .Y(n_728) );
AOI22xp33_ASAP7_75t_L g773 ( .A1(n_69), .A2(n_249), .B1(n_479), .B2(n_643), .Y(n_773) );
INVx1_ASAP7_75t_L g779 ( .A(n_69), .Y(n_779) );
OAI22xp5_ASAP7_75t_L g1044 ( .A1(n_70), .A2(n_1045), .B1(n_1095), .B2(n_1096), .Y(n_1044) );
INVx1_ASAP7_75t_L g1096 ( .A(n_70), .Y(n_1096) );
OAI22xp5_ASAP7_75t_L g1053 ( .A1(n_71), .A2(n_75), .B1(n_529), .B2(n_533), .Y(n_1053) );
AOI22xp33_ASAP7_75t_L g1066 ( .A1(n_71), .A2(n_75), .B1(n_658), .B2(n_895), .Y(n_1066) );
INVx1_ASAP7_75t_L g917 ( .A(n_72), .Y(n_917) );
INVx1_ASAP7_75t_L g920 ( .A(n_73), .Y(n_920) );
AOI22xp33_ASAP7_75t_L g936 ( .A1(n_73), .A2(n_128), .B1(n_722), .B2(n_763), .Y(n_936) );
AOI22xp33_ASAP7_75t_L g399 ( .A1(n_74), .A2(n_236), .B1(n_400), .B2(n_403), .Y(n_399) );
AOI22xp33_ASAP7_75t_L g440 ( .A1(n_74), .A2(n_236), .B1(n_441), .B2(n_444), .Y(n_440) );
INVx1_ASAP7_75t_L g1219 ( .A(n_76), .Y(n_1219) );
INVx1_ASAP7_75t_L g325 ( .A(n_77), .Y(n_325) );
CKINVDCx5p33_ASAP7_75t_R g609 ( .A(n_78), .Y(n_609) );
INVxp33_ASAP7_75t_SL g1115 ( .A(n_79), .Y(n_1115) );
AOI22xp33_ASAP7_75t_L g1140 ( .A1(n_79), .A2(n_243), .B1(n_321), .B2(n_491), .Y(n_1140) );
INVxp67_ASAP7_75t_SL g858 ( .A(n_81), .Y(n_858) );
AOI22xp33_ASAP7_75t_SL g886 ( .A1(n_81), .A2(n_202), .B1(n_490), .B2(n_887), .Y(n_886) );
INVx1_ASAP7_75t_L g527 ( .A(n_82), .Y(n_527) );
CKINVDCx16_ASAP7_75t_R g1171 ( .A(n_83), .Y(n_1171) );
AOI22xp5_ASAP7_75t_L g1187 ( .A1(n_84), .A2(n_139), .B1(n_1176), .B2(n_1179), .Y(n_1187) );
INVx1_ASAP7_75t_L g630 ( .A(n_85), .Y(n_630) );
OAI22xp5_ASAP7_75t_L g667 ( .A1(n_85), .A2(n_92), .B1(n_668), .B2(n_669), .Y(n_667) );
INVx1_ASAP7_75t_L g987 ( .A(n_86), .Y(n_987) );
INVx1_ASAP7_75t_L g394 ( .A(n_87), .Y(n_394) );
INVxp33_ASAP7_75t_SL g869 ( .A(n_88), .Y(n_869) );
AOI22xp33_ASAP7_75t_L g901 ( .A1(n_88), .A2(n_195), .B1(n_551), .B2(n_902), .Y(n_901) );
INVx1_ASAP7_75t_L g860 ( .A(n_89), .Y(n_860) );
AOI22xp33_ASAP7_75t_L g889 ( .A1(n_89), .A2(n_187), .B1(n_706), .B2(n_884), .Y(n_889) );
INVx1_ASAP7_75t_L g976 ( .A(n_90), .Y(n_976) );
AOI22xp33_ASAP7_75t_L g880 ( .A1(n_91), .A2(n_198), .B1(n_490), .B2(n_881), .Y(n_880) );
AOI22xp33_ASAP7_75t_L g892 ( .A1(n_91), .A2(n_198), .B1(n_893), .B2(n_896), .Y(n_892) );
INVx1_ASAP7_75t_L g632 ( .A(n_92), .Y(n_632) );
INVx1_ASAP7_75t_L g1058 ( .A(n_93), .Y(n_1058) );
AOI22xp33_ASAP7_75t_L g1021 ( .A1(n_94), .A2(n_104), .B1(n_320), .B2(n_409), .Y(n_1021) );
AOI22xp33_ASAP7_75t_L g1030 ( .A1(n_94), .A2(n_104), .B1(n_841), .B2(n_1031), .Y(n_1030) );
AOI22xp33_ASAP7_75t_L g1126 ( .A1(n_95), .A2(n_160), .B1(n_1127), .B2(n_1128), .Y(n_1126) );
AOI22xp33_ASAP7_75t_L g1133 ( .A1(n_95), .A2(n_160), .B1(n_1107), .B2(n_1134), .Y(n_1133) );
INVx1_ASAP7_75t_L g493 ( .A(n_96), .Y(n_493) );
INVxp67_ASAP7_75t_SL g1397 ( .A(n_97), .Y(n_1397) );
INVxp67_ASAP7_75t_SL g800 ( .A(n_98), .Y(n_800) );
AOI22xp33_ASAP7_75t_L g827 ( .A1(n_98), .A2(n_248), .B1(n_828), .B2(n_829), .Y(n_827) );
INVx1_ASAP7_75t_L g756 ( .A(n_99), .Y(n_756) );
OAI22xp33_ASAP7_75t_L g780 ( .A1(n_99), .A2(n_186), .B1(n_327), .B2(n_669), .Y(n_780) );
AOI22xp33_ASAP7_75t_L g965 ( .A1(n_100), .A2(n_147), .B1(n_559), .B2(n_564), .Y(n_965) );
OAI22xp5_ASAP7_75t_L g969 ( .A1(n_100), .A2(n_147), .B1(n_529), .B2(n_533), .Y(n_969) );
INVx1_ASAP7_75t_L g1086 ( .A(n_101), .Y(n_1086) );
OAI22xp5_ASAP7_75t_L g1091 ( .A1(n_101), .A2(n_151), .B1(n_470), .B2(n_485), .Y(n_1091) );
AOI22xp33_ASAP7_75t_L g1427 ( .A1(n_102), .A2(n_116), .B1(n_305), .B2(n_580), .Y(n_1427) );
AOI22xp33_ASAP7_75t_L g1448 ( .A1(n_102), .A2(n_116), .B1(n_832), .B2(n_1060), .Y(n_1448) );
CKINVDCx5p33_ASAP7_75t_R g610 ( .A(n_103), .Y(n_610) );
INVx1_ASAP7_75t_L g1205 ( .A(n_105), .Y(n_1205) );
INVx1_ASAP7_75t_L g560 ( .A(n_106), .Y(n_560) );
INVxp33_ASAP7_75t_SL g1103 ( .A(n_107), .Y(n_1103) );
AOI22xp33_ASAP7_75t_L g1130 ( .A1(n_107), .A2(n_242), .B1(n_1125), .B2(n_1131), .Y(n_1130) );
INVx1_ASAP7_75t_L g1004 ( .A(n_108), .Y(n_1004) );
AOI22xp33_ASAP7_75t_L g1059 ( .A1(n_109), .A2(n_153), .B1(n_770), .B2(n_1060), .Y(n_1059) );
INVxp67_ASAP7_75t_SL g1073 ( .A(n_109), .Y(n_1073) );
INVxp33_ASAP7_75t_L g671 ( .A(n_110), .Y(n_671) );
OAI22xp5_ASAP7_75t_L g695 ( .A1(n_111), .A2(n_130), .B1(n_470), .B2(n_485), .Y(n_695) );
AOI22xp33_ASAP7_75t_SL g718 ( .A1(n_111), .A2(n_130), .B1(n_409), .B2(n_719), .Y(n_718) );
AO221x2_ASAP7_75t_L g1216 ( .A1(n_112), .A2(n_178), .B1(n_1167), .B2(n_1173), .C(n_1217), .Y(n_1216) );
AOI22xp33_ASAP7_75t_L g759 ( .A1(n_113), .A2(n_230), .B1(n_424), .B2(n_646), .Y(n_759) );
AOI22xp33_ASAP7_75t_L g769 ( .A1(n_113), .A2(n_230), .B1(n_559), .B2(n_770), .Y(n_769) );
INVx1_ASAP7_75t_L g592 ( .A(n_114), .Y(n_592) );
OAI22xp5_ASAP7_75t_L g613 ( .A1(n_114), .A2(n_134), .B1(n_470), .B2(n_485), .Y(n_613) );
AO22x2_ASAP7_75t_L g620 ( .A1(n_115), .A2(n_621), .B1(n_677), .B2(n_678), .Y(n_620) );
INVx1_ASAP7_75t_L g677 ( .A(n_115), .Y(n_677) );
INVx1_ASAP7_75t_L g272 ( .A(n_117), .Y(n_272) );
XNOR2xp5_ASAP7_75t_L g537 ( .A(n_118), .B(n_538), .Y(n_537) );
AOI221xp5_ASAP7_75t_L g489 ( .A1(n_119), .A2(n_209), .B1(n_490), .B2(n_491), .C(n_492), .Y(n_489) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_119), .A2(n_209), .B1(n_459), .B2(n_460), .Y(n_515) );
INVx1_ASAP7_75t_L g483 ( .A(n_120), .Y(n_483) );
OAI211xp5_ASAP7_75t_L g1048 ( .A1(n_121), .A2(n_338), .B(n_1049), .C(n_1050), .Y(n_1048) );
INVx1_ASAP7_75t_L g1065 ( .A(n_121), .Y(n_1065) );
OAI22xp5_ASAP7_75t_L g977 ( .A1(n_122), .A2(n_194), .B1(n_281), .B2(n_299), .Y(n_977) );
OAI22xp33_ASAP7_75t_L g986 ( .A1(n_122), .A2(n_221), .B1(n_470), .B2(n_475), .Y(n_986) );
INVxp67_ASAP7_75t_SL g797 ( .A(n_123), .Y(n_797) );
INVxp67_ASAP7_75t_SL g694 ( .A(n_124), .Y(n_694) );
AOI22xp5_ASAP7_75t_L g1188 ( .A1(n_125), .A2(n_170), .B1(n_1173), .B2(n_1182), .Y(n_1188) );
INVx1_ASAP7_75t_L g634 ( .A(n_126), .Y(n_634) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_127), .A2(n_165), .B1(n_549), .B2(n_551), .Y(n_548) );
INVx1_ASAP7_75t_L g573 ( .A(n_127), .Y(n_573) );
INVxp67_ASAP7_75t_SL g919 ( .A(n_128), .Y(n_919) );
AOI22xp33_ASAP7_75t_L g823 ( .A1(n_129), .A2(n_158), .B1(n_712), .B2(n_824), .Y(n_823) );
AOI22xp33_ASAP7_75t_L g831 ( .A1(n_129), .A2(n_158), .B1(n_832), .B2(n_834), .Y(n_831) );
AOI22xp33_ASAP7_75t_L g641 ( .A1(n_131), .A2(n_137), .B1(n_443), .B2(n_460), .Y(n_641) );
AOI22xp33_ASAP7_75t_SL g661 ( .A1(n_131), .A2(n_137), .B1(n_424), .B2(n_646), .Y(n_661) );
INVx1_ASAP7_75t_L g294 ( .A(n_133), .Y(n_294) );
INVx1_ASAP7_75t_L g588 ( .A(n_134), .Y(n_588) );
CKINVDCx14_ASAP7_75t_R g466 ( .A(n_135), .Y(n_466) );
INVx1_ASAP7_75t_L g482 ( .A(n_136), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g711 ( .A1(n_138), .A2(n_222), .B1(n_712), .B2(n_714), .Y(n_711) );
AOI22xp33_ASAP7_75t_SL g733 ( .A1(n_138), .A2(n_210), .B1(n_734), .B2(n_736), .Y(n_733) );
INVxp33_ASAP7_75t_SL g624 ( .A(n_140), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_140), .A2(n_155), .B1(n_321), .B2(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g750 ( .A(n_141), .Y(n_750) );
INVxp67_ASAP7_75t_SL g1015 ( .A(n_142), .Y(n_1015) );
INVxp33_ASAP7_75t_L g346 ( .A(n_143), .Y(n_346) );
AOI22xp33_ASAP7_75t_L g952 ( .A1(n_144), .A2(n_149), .B1(n_646), .B2(n_953), .Y(n_952) );
AOI22xp33_ASAP7_75t_L g961 ( .A1(n_144), .A2(n_149), .B1(n_895), .B2(n_962), .Y(n_961) );
OAI22xp33_ASAP7_75t_L g921 ( .A1(n_146), .A2(n_189), .B1(n_470), .B2(n_475), .Y(n_921) );
AOI22xp33_ASAP7_75t_L g937 ( .A1(n_146), .A2(n_220), .B1(n_766), .B2(n_938), .Y(n_937) );
INVx1_ASAP7_75t_L g1005 ( .A(n_148), .Y(n_1005) );
AOI22xp5_ASAP7_75t_L g1468 ( .A1(n_150), .A2(n_1469), .B1(n_1470), .B2(n_1471), .Y(n_1468) );
CKINVDCx5p33_ASAP7_75t_R g1469 ( .A(n_150), .Y(n_1469) );
INVx1_ASAP7_75t_L g1079 ( .A(n_151), .Y(n_1079) );
INVxp67_ASAP7_75t_SL g358 ( .A(n_152), .Y(n_358) );
AOI22xp33_ASAP7_75t_L g420 ( .A1(n_152), .A2(n_203), .B1(n_421), .B2(n_422), .Y(n_420) );
INVxp67_ASAP7_75t_SL g1075 ( .A(n_153), .Y(n_1075) );
AOI22xp5_ASAP7_75t_L g1194 ( .A1(n_154), .A2(n_159), .B1(n_1176), .B2(n_1179), .Y(n_1194) );
INVxp67_ASAP7_75t_SL g627 ( .A(n_155), .Y(n_627) );
INVxp33_ASAP7_75t_SL g635 ( .A(n_156), .Y(n_635) );
AOI22xp33_ASAP7_75t_SL g645 ( .A1(n_156), .A2(n_174), .B1(n_424), .B2(n_646), .Y(n_645) );
AOI22xp33_ASAP7_75t_L g760 ( .A1(n_157), .A2(n_241), .B1(n_321), .B2(n_663), .Y(n_760) );
AOI22xp33_ASAP7_75t_L g768 ( .A1(n_157), .A2(n_241), .B1(n_479), .B2(n_643), .Y(n_768) );
INVx1_ASAP7_75t_L g303 ( .A(n_161), .Y(n_303) );
HB1xp67_ASAP7_75t_L g274 ( .A(n_162), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g1155 ( .A(n_162), .B(n_272), .Y(n_1155) );
AND3x2_ASAP7_75t_L g1170 ( .A(n_162), .B(n_272), .C(n_1158), .Y(n_1170) );
AOI22xp5_ASAP7_75t_L g1195 ( .A1(n_163), .A2(n_214), .B1(n_1167), .B2(n_1196), .Y(n_1195) );
OAI22xp5_ASAP7_75t_L g614 ( .A1(n_164), .A2(n_227), .B1(n_475), .B2(n_486), .Y(n_614) );
INVx1_ASAP7_75t_L g581 ( .A(n_165), .Y(n_581) );
INVxp33_ASAP7_75t_SL g802 ( .A(n_166), .Y(n_802) );
AOI22xp33_ASAP7_75t_L g826 ( .A1(n_166), .A2(n_237), .B1(n_320), .B2(n_820), .Y(n_826) );
INVx1_ASAP7_75t_L g916 ( .A(n_167), .Y(n_916) );
INVx2_ASAP7_75t_L g285 ( .A(n_168), .Y(n_285) );
AOI22xp5_ASAP7_75t_L g996 ( .A1(n_169), .A2(n_997), .B1(n_1040), .B2(n_1041), .Y(n_996) );
INVxp67_ASAP7_75t_L g1040 ( .A(n_169), .Y(n_1040) );
INVxp33_ASAP7_75t_SL g1012 ( .A(n_172), .Y(n_1012) );
INVxp33_ASAP7_75t_SL g625 ( .A(n_174), .Y(n_625) );
AOI22xp5_ASAP7_75t_L g1181 ( .A1(n_175), .A2(n_182), .B1(n_1173), .B2(n_1182), .Y(n_1181) );
INVx1_ASAP7_75t_L g1052 ( .A(n_176), .Y(n_1052) );
AOI22xp33_ASAP7_75t_L g932 ( .A1(n_177), .A2(n_201), .B1(n_595), .B2(n_933), .Y(n_932) );
AOI22xp33_ASAP7_75t_L g943 ( .A1(n_177), .A2(n_201), .B1(n_895), .B2(n_944), .Y(n_943) );
AOI21xp33_ASAP7_75t_L g1424 ( .A1(n_180), .A2(n_725), .B(n_1425), .Y(n_1424) );
INVxp67_ASAP7_75t_SL g1447 ( .A(n_180), .Y(n_1447) );
INVx1_ASAP7_75t_L g1158 ( .A(n_181), .Y(n_1158) );
INVxp67_ASAP7_75t_SL g309 ( .A(n_183), .Y(n_309) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_183), .A2(n_219), .B1(n_457), .B2(n_460), .Y(n_456) );
CKINVDCx16_ASAP7_75t_R g1202 ( .A(n_184), .Y(n_1202) );
OAI211xp5_ASAP7_75t_L g924 ( .A1(n_185), .A2(n_338), .B(n_925), .C(n_926), .Y(n_924) );
AOI22xp33_ASAP7_75t_L g946 ( .A1(n_185), .A2(n_261), .B1(n_643), .B2(n_942), .Y(n_946) );
INVx1_ASAP7_75t_L g755 ( .A(n_186), .Y(n_755) );
INVxp33_ASAP7_75t_SL g854 ( .A(n_187), .Y(n_854) );
INVx1_ASAP7_75t_L g1009 ( .A(n_188), .Y(n_1009) );
OAI22xp5_ASAP7_75t_L g929 ( .A1(n_189), .A2(n_261), .B1(n_281), .B2(n_299), .Y(n_929) );
INVx1_ASAP7_75t_L g1249 ( .A(n_190), .Y(n_1249) );
INVxp33_ASAP7_75t_SL g702 ( .A(n_191), .Y(n_702) );
AOI22xp33_ASAP7_75t_L g739 ( .A1(n_191), .A2(n_245), .B1(n_736), .B2(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g1437 ( .A(n_192), .Y(n_1437) );
INVxp67_ASAP7_75t_SL g808 ( .A(n_193), .Y(n_808) );
AOI22xp33_ASAP7_75t_L g840 ( .A1(n_193), .A2(n_232), .B1(n_628), .B2(n_841), .Y(n_840) );
INVxp33_ASAP7_75t_SL g870 ( .A(n_195), .Y(n_870) );
INVx1_ASAP7_75t_L g517 ( .A(n_196), .Y(n_517) );
OAI22xp5_ASAP7_75t_L g1047 ( .A1(n_197), .A2(n_262), .B1(n_281), .B2(n_299), .Y(n_1047) );
INVx1_ASAP7_75t_L g1063 ( .A(n_197), .Y(n_1063) );
INVx1_ASAP7_75t_L g287 ( .A(n_199), .Y(n_287) );
INVx2_ASAP7_75t_L g302 ( .A(n_199), .Y(n_302) );
OAI211xp5_ASAP7_75t_L g476 ( .A1(n_200), .A2(n_477), .B(n_480), .C(n_481), .Y(n_476) );
INVx1_ASAP7_75t_L g505 ( .A(n_200), .Y(n_505) );
INVxp33_ASAP7_75t_SL g855 ( .A(n_202), .Y(n_855) );
INVxp67_ASAP7_75t_SL g368 ( .A(n_203), .Y(n_368) );
INVxp33_ASAP7_75t_SL g815 ( .A(n_204), .Y(n_815) );
AO22x2_ASAP7_75t_L g791 ( .A1(n_205), .A2(n_792), .B1(n_847), .B2(n_848), .Y(n_791) );
CKINVDCx14_ASAP7_75t_R g847 ( .A(n_205), .Y(n_847) );
INVxp67_ASAP7_75t_SL g1121 ( .A(n_206), .Y(n_1121) );
AOI22xp33_ASAP7_75t_L g1139 ( .A1(n_206), .A2(n_246), .B1(n_400), .B2(n_1134), .Y(n_1139) );
AOI22xp5_ASAP7_75t_L g1175 ( .A1(n_208), .A2(n_235), .B1(n_1176), .B2(n_1179), .Y(n_1175) );
XNOR2xp5_ASAP7_75t_L g1388 ( .A(n_208), .B(n_1389), .Y(n_1388) );
AOI22xp33_ASAP7_75t_L g1463 ( .A1(n_208), .A2(n_1464), .B1(n_1467), .B2(n_1472), .Y(n_1463) );
XNOR2xp5_ASAP7_75t_L g743 ( .A(n_211), .B(n_744), .Y(n_743) );
CKINVDCx20_ASAP7_75t_R g311 ( .A(n_212), .Y(n_311) );
INVx1_ASAP7_75t_L g495 ( .A(n_213), .Y(n_495) );
INVx1_ASAP7_75t_L g1435 ( .A(n_215), .Y(n_1435) );
INVx1_ASAP7_75t_L g1112 ( .A(n_216), .Y(n_1112) );
CKINVDCx5p33_ASAP7_75t_R g542 ( .A(n_217), .Y(n_542) );
INVx1_ASAP7_75t_L g1106 ( .A(n_218), .Y(n_1106) );
AOI22xp33_ASAP7_75t_L g1129 ( .A1(n_218), .A2(n_239), .B1(n_375), .B2(n_1060), .Y(n_1129) );
INVxp67_ASAP7_75t_SL g337 ( .A(n_219), .Y(n_337) );
INVx1_ASAP7_75t_L g913 ( .A(n_220), .Y(n_913) );
INVx1_ASAP7_75t_L g799 ( .A(n_223), .Y(n_799) );
INVx1_ASAP7_75t_L g1051 ( .A(n_224), .Y(n_1051) );
AO22x2_ASAP7_75t_L g1098 ( .A1(n_225), .A2(n_1099), .B1(n_1100), .B2(n_1142), .Y(n_1098) );
INVx1_ASAP7_75t_L g1099 ( .A(n_225), .Y(n_1099) );
INVxp67_ASAP7_75t_SL g319 ( .A(n_226), .Y(n_319) );
INVx1_ASAP7_75t_L g597 ( .A(n_227), .Y(n_597) );
INVx1_ASAP7_75t_L g985 ( .A(n_228), .Y(n_985) );
INVx1_ASAP7_75t_L g1159 ( .A(n_229), .Y(n_1159) );
NAND2xp5_ASAP7_75t_L g1163 ( .A(n_229), .B(n_1157), .Y(n_1163) );
INVxp33_ASAP7_75t_SL g806 ( .A(n_232), .Y(n_806) );
INVxp67_ASAP7_75t_SL g666 ( .A(n_233), .Y(n_666) );
INVx1_ASAP7_75t_L g864 ( .A(n_234), .Y(n_864) );
INVx1_ASAP7_75t_L g795 ( .A(n_237), .Y(n_795) );
INVx1_ASAP7_75t_L g975 ( .A(n_238), .Y(n_975) );
INVxp67_ASAP7_75t_SL g1104 ( .A(n_239), .Y(n_1104) );
CKINVDCx5p33_ASAP7_75t_R g1426 ( .A(n_240), .Y(n_1426) );
INVxp33_ASAP7_75t_SL g1111 ( .A(n_242), .Y(n_1111) );
INVx1_ASAP7_75t_L g1117 ( .A(n_243), .Y(n_1117) );
INVxp33_ASAP7_75t_L g701 ( .A(n_245), .Y(n_701) );
INVxp33_ASAP7_75t_SL g1119 ( .A(n_246), .Y(n_1119) );
INVx2_ASAP7_75t_L g284 ( .A(n_247), .Y(n_284) );
INVxp67_ASAP7_75t_SL g803 ( .A(n_248), .Y(n_803) );
INVx1_ASAP7_75t_L g785 ( .A(n_249), .Y(n_785) );
INVxp33_ASAP7_75t_SL g877 ( .A(n_250), .Y(n_877) );
AOI22xp33_ASAP7_75t_L g898 ( .A1(n_250), .A2(n_265), .B1(n_754), .B2(n_899), .Y(n_898) );
INVxp67_ASAP7_75t_SL g1404 ( .A(n_251), .Y(n_1404) );
XOR2xp5_ASAP7_75t_L g681 ( .A(n_252), .B(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g688 ( .A(n_253), .Y(n_688) );
BUFx3_ASAP7_75t_L g355 ( .A(n_256), .Y(n_355) );
INVx1_ASAP7_75t_L g372 ( .A(n_256), .Y(n_372) );
BUFx3_ASAP7_75t_L g357 ( .A(n_257), .Y(n_357) );
INVx1_ASAP7_75t_L g363 ( .A(n_257), .Y(n_363) );
INVx1_ASAP7_75t_L g1081 ( .A(n_258), .Y(n_1081) );
OAI22xp33_ASAP7_75t_L g1094 ( .A1(n_258), .A2(n_262), .B1(n_475), .B2(n_486), .Y(n_1094) );
INVx1_ASAP7_75t_L g518 ( .A(n_259), .Y(n_518) );
INVx1_ASAP7_75t_L g1108 ( .A(n_260), .Y(n_1108) );
INVx1_ASAP7_75t_L g748 ( .A(n_263), .Y(n_748) );
INVx1_ASAP7_75t_L g1400 ( .A(n_264), .Y(n_1400) );
INVx1_ASAP7_75t_L g872 ( .A(n_265), .Y(n_872) );
AOI21xp5_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_288), .B(n_1144), .Y(n_266) );
INVx2_ASAP7_75t_SL g267 ( .A(n_268), .Y(n_267) );
INVx1_ASAP7_75t_SL g268 ( .A(n_269), .Y(n_268) );
AND2x4_ASAP7_75t_L g269 ( .A(n_270), .B(n_275), .Y(n_269) );
AND2x4_ASAP7_75t_L g1462 ( .A(n_270), .B(n_276), .Y(n_1462) );
NOR2xp33_ASAP7_75t_SL g270 ( .A(n_271), .B(n_273), .Y(n_270) );
INVx1_ASAP7_75t_SL g1466 ( .A(n_271), .Y(n_1466) );
NAND2xp5_ASAP7_75t_L g1475 ( .A(n_271), .B(n_273), .Y(n_1475) );
HB1xp67_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g1465 ( .A(n_273), .B(n_1466), .Y(n_1465) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g276 ( .A(n_277), .B(n_281), .Y(n_276) );
INVxp67_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
OR2x6_ASAP7_75t_L g342 ( .A(n_278), .B(n_343), .Y(n_342) );
OR2x2_ASAP7_75t_L g676 ( .A(n_278), .B(n_343), .Y(n_676) );
HB1xp67_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g418 ( .A(n_279), .B(n_287), .Y(n_418) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
OR2x2_ASAP7_75t_L g571 ( .A(n_280), .B(n_301), .Y(n_571) );
INVx8_ASAP7_75t_L g331 ( .A(n_281), .Y(n_331) );
OR2x6_ASAP7_75t_L g281 ( .A(n_282), .B(n_286), .Y(n_281) );
OR2x6_ASAP7_75t_L g299 ( .A(n_282), .B(n_300), .Y(n_299) );
HB1xp67_ASAP7_75t_L g494 ( .A(n_282), .Y(n_494) );
INVx2_ASAP7_75t_SL g504 ( .A(n_282), .Y(n_504) );
INVx2_ASAP7_75t_SL g584 ( .A(n_282), .Y(n_584) );
BUFx6f_ASAP7_75t_L g1070 ( .A(n_282), .Y(n_1070) );
INVx1_ASAP7_75t_L g1085 ( .A(n_282), .Y(n_1085) );
OAI21xp33_ASAP7_75t_L g1425 ( .A1(n_282), .A2(n_418), .B(n_1426), .Y(n_1425) );
BUFx6f_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
INVx2_ASAP7_75t_L g306 ( .A(n_284), .Y(n_306) );
INVx1_ASAP7_75t_L g315 ( .A(n_284), .Y(n_315) );
INVx1_ASAP7_75t_L g323 ( .A(n_284), .Y(n_323) );
AND2x4_ASAP7_75t_L g336 ( .A(n_284), .B(n_324), .Y(n_336) );
AND2x2_ASAP7_75t_L g411 ( .A(n_284), .B(n_285), .Y(n_411) );
INVx1_ASAP7_75t_L g308 ( .A(n_285), .Y(n_308) );
INVx2_ASAP7_75t_L g324 ( .A(n_285), .Y(n_324) );
INVx1_ASAP7_75t_L g329 ( .A(n_285), .Y(n_329) );
INVx1_ASAP7_75t_L g498 ( .A(n_285), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_285), .B(n_306), .Y(n_532) );
AND2x4_ASAP7_75t_L g328 ( .A(n_286), .B(n_329), .Y(n_328) );
INVx2_ASAP7_75t_SL g286 ( .A(n_287), .Y(n_286) );
OR2x2_ASAP7_75t_L g669 ( .A(n_287), .B(n_314), .Y(n_669) );
OR2x2_ASAP7_75t_L g812 ( .A(n_287), .B(n_314), .Y(n_812) );
OAI22xp33_ASAP7_75t_L g288 ( .A1(n_289), .A2(n_990), .B1(n_991), .B2(n_1143), .Y(n_288) );
INVx1_ASAP7_75t_L g1143 ( .A(n_289), .Y(n_1143) );
XNOR2xp5_ASAP7_75t_L g289 ( .A(n_290), .B(n_789), .Y(n_289) );
XNOR2xp5_ASAP7_75t_L g290 ( .A(n_291), .B(n_535), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
XNOR2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_465), .Y(n_292) );
XNOR2xp5_ASAP7_75t_L g293 ( .A(n_294), .B(n_295), .Y(n_293) );
OAI22xp5_ASAP7_75t_L g1190 ( .A1(n_294), .A2(n_1154), .B1(n_1162), .B2(n_1191), .Y(n_1190) );
AOI221xp5_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_341), .B1(n_344), .B2(n_390), .C(n_397), .Y(n_295) );
NAND4xp25_ASAP7_75t_L g296 ( .A(n_297), .B(n_310), .C(n_330), .D(n_338), .Y(n_296) );
AOI22xp33_ASAP7_75t_SL g297 ( .A1(n_298), .A2(n_303), .B1(n_304), .B2(n_309), .Y(n_297) );
AOI22xp33_ASAP7_75t_L g526 ( .A1(n_298), .A2(n_331), .B1(n_517), .B2(n_527), .Y(n_526) );
AOI22xp33_ASAP7_75t_SL g784 ( .A1(n_298), .A2(n_331), .B1(n_747), .B2(n_785), .Y(n_784) );
AOI22xp33_ASAP7_75t_L g1007 ( .A1(n_298), .A2(n_331), .B1(n_1008), .B2(n_1009), .Y(n_1007) );
AOI22xp33_ASAP7_75t_L g1110 ( .A1(n_298), .A2(n_331), .B1(n_1111), .B2(n_1112), .Y(n_1110) );
INVx4_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx5_ASAP7_75t_L g675 ( .A(n_299), .Y(n_675) );
AND2x4_ASAP7_75t_L g304 ( .A(n_300), .B(n_305), .Y(n_304) );
AND2x4_ASAP7_75t_L g333 ( .A(n_300), .B(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g530 ( .A(n_300), .Y(n_530) );
AND2x4_ASAP7_75t_L g534 ( .A(n_300), .B(n_334), .Y(n_534) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g318 ( .A(n_302), .Y(n_318) );
AOI22xp33_ASAP7_75t_L g364 ( .A1(n_303), .A2(n_365), .B1(n_368), .B2(n_369), .Y(n_364) );
AOI22xp33_ASAP7_75t_SL g670 ( .A1(n_304), .A2(n_333), .B1(n_671), .B2(n_672), .Y(n_670) );
AOI22xp33_ASAP7_75t_L g700 ( .A1(n_304), .A2(n_333), .B1(n_701), .B2(n_702), .Y(n_700) );
AOI22xp33_ASAP7_75t_SL g781 ( .A1(n_304), .A2(n_333), .B1(n_782), .B2(n_783), .Y(n_781) );
AOI22xp5_ASAP7_75t_L g813 ( .A1(n_304), .A2(n_534), .B1(n_814), .B2(n_815), .Y(n_813) );
AOI22xp33_ASAP7_75t_L g868 ( .A1(n_304), .A2(n_333), .B1(n_869), .B2(n_870), .Y(n_868) );
AOI22xp33_ASAP7_75t_L g999 ( .A1(n_304), .A2(n_534), .B1(n_1000), .B2(n_1001), .Y(n_999) );
AOI22xp33_ASAP7_75t_L g1102 ( .A1(n_304), .A2(n_534), .B1(n_1103), .B2(n_1104), .Y(n_1102) );
BUFx6f_ASAP7_75t_L g402 ( .A(n_305), .Y(n_402) );
BUFx2_ASAP7_75t_L g421 ( .A(n_305), .Y(n_421) );
BUFx2_ASAP7_75t_L g490 ( .A(n_305), .Y(n_490) );
BUFx6f_ASAP7_75t_L g646 ( .A(n_305), .Y(n_646) );
INVx1_ASAP7_75t_L g713 ( .A(n_305), .Y(n_713) );
INVx1_ASAP7_75t_L g720 ( .A(n_305), .Y(n_720) );
BUFx6f_ASAP7_75t_L g763 ( .A(n_305), .Y(n_763) );
AND2x2_ASAP7_75t_L g1405 ( .A(n_305), .B(n_1406), .Y(n_1405) );
AND2x4_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
INVx1_ASAP7_75t_L g1422 ( .A(n_306), .Y(n_1422) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
AOI222xp33_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_312), .B1(n_319), .B2(n_320), .C1(n_325), .C2(n_326), .Y(n_310) );
AOI222xp33_ASAP7_75t_L g373 ( .A1(n_311), .A2(n_325), .B1(n_374), .B2(n_375), .C1(n_379), .C2(n_384), .Y(n_373) );
AOI222xp33_ASAP7_75t_L g523 ( .A1(n_312), .A2(n_328), .B1(n_482), .B2(n_483), .C1(n_518), .C2(n_524), .Y(n_523) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_312), .A2(n_328), .B1(n_609), .B2(n_610), .Y(n_608) );
AOI222xp33_ASAP7_75t_L g871 ( .A1(n_312), .A2(n_326), .B1(n_863), .B2(n_864), .C1(n_872), .C2(n_873), .Y(n_871) );
AOI22xp33_ASAP7_75t_L g926 ( .A1(n_312), .A2(n_916), .B1(n_917), .B2(n_927), .Y(n_926) );
AOI22xp33_ASAP7_75t_L g974 ( .A1(n_312), .A2(n_328), .B1(n_975), .B2(n_976), .Y(n_974) );
AOI22xp33_ASAP7_75t_L g1050 ( .A1(n_312), .A2(n_927), .B1(n_1051), .B2(n_1052), .Y(n_1050) );
AOI222xp33_ASAP7_75t_L g1105 ( .A1(n_312), .A2(n_328), .B1(n_1106), .B2(n_1107), .C1(n_1108), .C2(n_1109), .Y(n_1105) );
AND2x4_ASAP7_75t_L g312 ( .A(n_313), .B(n_316), .Y(n_312) );
AND2x4_ASAP7_75t_L g1006 ( .A(n_313), .B(n_316), .Y(n_1006) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g497 ( .A(n_315), .B(n_498), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_315), .B(n_498), .Y(n_607) );
INVxp67_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g340 ( .A(n_317), .Y(n_340) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
NAND2x1p5_ASAP7_75t_L g432 ( .A(n_318), .B(n_433), .Y(n_432) );
AOI211xp5_ASAP7_75t_L g665 ( .A1(n_320), .A2(n_339), .B(n_666), .C(n_667), .Y(n_665) );
AOI211xp5_ASAP7_75t_L g778 ( .A1(n_320), .A2(n_339), .B(n_779), .C(n_780), .Y(n_778) );
BUFx6f_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx2_ASAP7_75t_SL g427 ( .A(n_321), .Y(n_427) );
BUFx6f_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
AND2x4_ASAP7_75t_L g339 ( .A(n_322), .B(n_340), .Y(n_339) );
BUFx3_ASAP7_75t_L g413 ( .A(n_322), .Y(n_413) );
BUFx3_ASAP7_75t_L g525 ( .A(n_322), .Y(n_525) );
BUFx6f_ASAP7_75t_L g725 ( .A(n_322), .Y(n_725) );
INVx1_ASAP7_75t_L g810 ( .A(n_322), .Y(n_810) );
BUFx2_ASAP7_75t_L g875 ( .A(n_322), .Y(n_875) );
AND2x4_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx2_ASAP7_75t_L g668 ( .A(n_328), .Y(n_668) );
INVx2_ASAP7_75t_L g928 ( .A(n_328), .Y(n_928) );
AOI222xp33_ASAP7_75t_L g1002 ( .A1(n_328), .A2(n_725), .B1(n_1003), .B2(n_1004), .C1(n_1005), .C2(n_1006), .Y(n_1002) );
INVx1_ASAP7_75t_L g1416 ( .A(n_329), .Y(n_1416) );
AOI22xp33_ASAP7_75t_SL g330 ( .A1(n_331), .A2(n_332), .B1(n_333), .B2(n_337), .Y(n_330) );
AOI22xp33_ASAP7_75t_SL g673 ( .A1(n_331), .A2(n_634), .B1(n_674), .B2(n_675), .Y(n_673) );
AOI22xp5_ASAP7_75t_L g805 ( .A1(n_331), .A2(n_675), .B1(n_799), .B2(n_806), .Y(n_805) );
AOI22xp33_ASAP7_75t_L g876 ( .A1(n_331), .A2(n_675), .B1(n_857), .B2(n_877), .Y(n_876) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx3_ASAP7_75t_L g406 ( .A(n_336), .Y(n_406) );
BUFx6f_ASAP7_75t_L g424 ( .A(n_336), .Y(n_424) );
INVx1_ASAP7_75t_L g717 ( .A(n_336), .Y(n_717) );
NAND3xp33_ASAP7_75t_L g522 ( .A(n_338), .B(n_523), .C(n_526), .Y(n_522) );
NAND4xp25_ASAP7_75t_SL g867 ( .A(n_338), .B(n_868), .C(n_871), .D(n_876), .Y(n_867) );
NAND4xp25_ASAP7_75t_L g998 ( .A(n_338), .B(n_999), .C(n_1002), .D(n_1007), .Y(n_998) );
NAND4xp25_ASAP7_75t_L g1101 ( .A(n_338), .B(n_1102), .C(n_1105), .D(n_1110), .Y(n_1101) );
CKINVDCx11_ASAP7_75t_R g338 ( .A(n_339), .Y(n_338) );
NOR3xp33_ASAP7_75t_L g697 ( .A(n_339), .B(n_698), .C(n_699), .Y(n_697) );
AOI211xp5_ASAP7_75t_L g807 ( .A1(n_339), .A2(n_808), .B(n_809), .C(n_811), .Y(n_807) );
OAI21xp5_ASAP7_75t_L g521 ( .A1(n_341), .A2(n_522), .B(n_528), .Y(n_521) );
OAI31xp33_ASAP7_75t_SL g602 ( .A1(n_341), .A2(n_603), .A3(n_604), .B(n_611), .Y(n_602) );
AOI221x1_ASAP7_75t_L g851 ( .A1(n_341), .A2(n_852), .B1(n_866), .B2(n_867), .C(n_878), .Y(n_851) );
OAI31xp33_ASAP7_75t_L g922 ( .A1(n_341), .A2(n_923), .A3(n_924), .B(n_929), .Y(n_922) );
OAI31xp33_ASAP7_75t_SL g968 ( .A1(n_341), .A2(n_969), .A3(n_970), .B(n_977), .Y(n_968) );
AOI221xp5_ASAP7_75t_L g997 ( .A1(n_341), .A2(n_392), .B1(n_998), .B2(n_1010), .C(n_1018), .Y(n_997) );
OAI31xp33_ASAP7_75t_L g1046 ( .A1(n_341), .A2(n_1047), .A3(n_1048), .B(n_1053), .Y(n_1046) );
AOI221x1_ASAP7_75t_L g1100 ( .A1(n_341), .A2(n_392), .B1(n_1101), .B2(n_1113), .C(n_1122), .Y(n_1100) );
CKINVDCx16_ASAP7_75t_R g341 ( .A(n_342), .Y(n_341) );
AOI31xp33_ASAP7_75t_L g777 ( .A1(n_342), .A2(n_778), .A3(n_781), .B(n_784), .Y(n_777) );
AND2x4_ASAP7_75t_L g453 ( .A(n_343), .B(n_454), .Y(n_453) );
AND2x4_ASAP7_75t_L g654 ( .A(n_343), .B(n_454), .Y(n_654) );
NAND4xp25_ASAP7_75t_L g344 ( .A(n_345), .B(n_364), .C(n_373), .D(n_386), .Y(n_344) );
AOI22xp33_ASAP7_75t_L g345 ( .A1(n_346), .A2(n_347), .B1(n_358), .B2(n_359), .Y(n_345) );
AOI22xp33_ASAP7_75t_L g623 ( .A1(n_347), .A2(n_359), .B1(n_624), .B2(n_625), .Y(n_623) );
AOI22xp5_ASAP7_75t_L g749 ( .A1(n_347), .A2(n_359), .B1(n_750), .B2(n_751), .Y(n_749) );
AOI22xp33_ASAP7_75t_L g801 ( .A1(n_347), .A2(n_359), .B1(n_802), .B2(n_803), .Y(n_801) );
AOI22xp33_ASAP7_75t_L g853 ( .A1(n_347), .A2(n_359), .B1(n_854), .B2(n_855), .Y(n_853) );
AOI22xp33_ASAP7_75t_L g1011 ( .A1(n_347), .A2(n_359), .B1(n_1012), .B2(n_1013), .Y(n_1011) );
HB1xp67_ASAP7_75t_L g1120 ( .A(n_347), .Y(n_1120) );
AND2x4_ASAP7_75t_L g347 ( .A(n_348), .B(n_351), .Y(n_347) );
AND2x6_ASAP7_75t_L g369 ( .A(n_348), .B(n_370), .Y(n_369) );
AND2x4_ASAP7_75t_L g1393 ( .A(n_348), .B(n_351), .Y(n_1393) );
INVx1_ASAP7_75t_SL g348 ( .A(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g689 ( .A(n_349), .B(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g361 ( .A(n_350), .Y(n_361) );
HB1xp67_ASAP7_75t_L g367 ( .A(n_350), .Y(n_367) );
AND2x2_ASAP7_75t_L g449 ( .A(n_350), .B(n_394), .Y(n_449) );
INVx2_ASAP7_75t_L g455 ( .A(n_350), .Y(n_455) );
INVx2_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx2_ASAP7_75t_L g437 ( .A(n_352), .Y(n_437) );
BUFx6f_ASAP7_75t_L g735 ( .A(n_352), .Y(n_735) );
INVx2_ASAP7_75t_L g838 ( .A(n_352), .Y(n_838) );
INVx2_ASAP7_75t_SL g843 ( .A(n_352), .Y(n_843) );
HB1xp67_ASAP7_75t_L g900 ( .A(n_352), .Y(n_900) );
INVx1_ASAP7_75t_L g967 ( .A(n_352), .Y(n_967) );
INVx6_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
AND2x4_ASAP7_75t_L g365 ( .A(n_353), .B(n_366), .Y(n_365) );
INVx2_ASAP7_75t_L g644 ( .A(n_353), .Y(n_644) );
BUFx2_ASAP7_75t_L g941 ( .A(n_353), .Y(n_941) );
AND2x4_ASAP7_75t_L g353 ( .A(n_354), .B(n_356), .Y(n_353) );
INVx1_ASAP7_75t_L g385 ( .A(n_354), .Y(n_385) );
INVx2_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
AND2x4_ASAP7_75t_L g362 ( .A(n_355), .B(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g378 ( .A(n_355), .B(n_357), .Y(n_378) );
INVx1_ASAP7_75t_L g383 ( .A(n_356), .Y(n_383) );
INVx2_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AND2x4_ASAP7_75t_L g371 ( .A(n_357), .B(n_372), .Y(n_371) );
CKINVDCx6p67_ASAP7_75t_R g485 ( .A(n_359), .Y(n_485) );
AOI22xp5_ASAP7_75t_L g918 ( .A1(n_359), .A2(n_369), .B1(n_919), .B2(n_920), .Y(n_918) );
AOI22xp5_ASAP7_75t_L g983 ( .A1(n_359), .A2(n_369), .B1(n_984), .B2(n_985), .Y(n_983) );
AOI22xp33_ASAP7_75t_L g1118 ( .A1(n_359), .A2(n_1119), .B1(n_1120), .B2(n_1121), .Y(n_1118) );
AOI22xp33_ASAP7_75t_L g1391 ( .A1(n_359), .A2(n_1392), .B1(n_1393), .B2(n_1394), .Y(n_1391) );
AND2x6_ASAP7_75t_L g359 ( .A(n_360), .B(n_362), .Y(n_359) );
INVx1_ASAP7_75t_L g388 ( .A(n_360), .Y(n_388) );
INVx1_ASAP7_75t_L g471 ( .A(n_360), .Y(n_471) );
AND2x2_ASAP7_75t_L g478 ( .A(n_360), .B(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
AND2x6_ASAP7_75t_L g384 ( .A(n_361), .B(n_385), .Y(n_384) );
BUFx6f_ASAP7_75t_L g443 ( .A(n_362), .Y(n_443) );
BUFx3_ASAP7_75t_L g459 ( .A(n_362), .Y(n_459) );
BUFx6f_ASAP7_75t_L g564 ( .A(n_362), .Y(n_564) );
BUFx2_ASAP7_75t_L g740 ( .A(n_362), .Y(n_740) );
INVx2_ASAP7_75t_SL g771 ( .A(n_362), .Y(n_771) );
BUFx6f_ASAP7_75t_L g833 ( .A(n_362), .Y(n_833) );
BUFx6f_ASAP7_75t_L g895 ( .A(n_362), .Y(n_895) );
HB1xp67_ASAP7_75t_L g902 ( .A(n_362), .Y(n_902) );
INVx1_ASAP7_75t_L g474 ( .A(n_363), .Y(n_474) );
INVx4_ASAP7_75t_L g475 ( .A(n_365), .Y(n_475) );
AOI22xp33_ASAP7_75t_L g633 ( .A1(n_365), .A2(n_369), .B1(n_634), .B2(n_635), .Y(n_633) );
AOI22xp33_ASAP7_75t_L g692 ( .A1(n_365), .A2(n_369), .B1(n_693), .B2(n_694), .Y(n_692) );
AOI22xp5_ASAP7_75t_L g746 ( .A1(n_365), .A2(n_369), .B1(n_747), .B2(n_748), .Y(n_746) );
AOI22xp33_ASAP7_75t_L g798 ( .A1(n_365), .A2(n_369), .B1(n_799), .B2(n_800), .Y(n_798) );
AOI22xp33_ASAP7_75t_L g856 ( .A1(n_365), .A2(n_369), .B1(n_857), .B2(n_858), .Y(n_856) );
AOI22xp33_ASAP7_75t_L g1014 ( .A1(n_365), .A2(n_369), .B1(n_1009), .B2(n_1015), .Y(n_1014) );
AOI22xp33_ASAP7_75t_L g1114 ( .A1(n_365), .A2(n_369), .B1(n_1112), .B2(n_1115), .Y(n_1114) );
AOI22xp33_ASAP7_75t_L g1395 ( .A1(n_365), .A2(n_369), .B1(n_1396), .B2(n_1397), .Y(n_1395) );
AND2x4_ASAP7_75t_L g380 ( .A(n_366), .B(n_381), .Y(n_380) );
AND2x2_ASAP7_75t_SL g631 ( .A(n_366), .B(n_381), .Y(n_631) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx4_ASAP7_75t_L g486 ( .A(n_369), .Y(n_486) );
BUFx6f_ASAP7_75t_L g460 ( .A(n_370), .Y(n_460) );
INVx2_ASAP7_75t_L g552 ( .A(n_370), .Y(n_552) );
BUFx6f_ASAP7_75t_L g559 ( .A(n_370), .Y(n_559) );
INVx1_ASAP7_75t_L g776 ( .A(n_370), .Y(n_776) );
INVx1_ASAP7_75t_L g835 ( .A(n_370), .Y(n_835) );
INVx1_ASAP7_75t_L g846 ( .A(n_370), .Y(n_846) );
BUFx6f_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g445 ( .A(n_371), .Y(n_445) );
BUFx6f_ASAP7_75t_L g520 ( .A(n_371), .Y(n_520) );
INVx2_ASAP7_75t_L g660 ( .A(n_371), .Y(n_660) );
INVx1_ASAP7_75t_L g963 ( .A(n_371), .Y(n_963) );
INVx1_ASAP7_75t_L g473 ( .A(n_372), .Y(n_473) );
AOI222xp33_ASAP7_75t_L g1116 ( .A1(n_375), .A2(n_379), .B1(n_384), .B2(n_1108), .C1(n_1109), .C2(n_1117), .Y(n_1116) );
BUFx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
BUFx4f_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
BUFx6f_ASAP7_75t_L g464 ( .A(n_377), .Y(n_464) );
INVx1_ASAP7_75t_L g629 ( .A(n_377), .Y(n_629) );
INVx2_ASAP7_75t_SL g732 ( .A(n_377), .Y(n_732) );
BUFx3_ASAP7_75t_L g754 ( .A(n_377), .Y(n_754) );
INVx1_ASAP7_75t_L g915 ( .A(n_377), .Y(n_915) );
BUFx6f_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
BUFx6f_ASAP7_75t_L g389 ( .A(n_378), .Y(n_389) );
AOI222xp33_ASAP7_75t_L g859 ( .A1(n_379), .A2(n_384), .B1(n_860), .B2(n_861), .C1(n_863), .C2(n_864), .Y(n_859) );
BUFx4f_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AOI22xp33_ASAP7_75t_L g481 ( .A1(n_380), .A2(n_384), .B1(n_482), .B2(n_483), .Y(n_481) );
AOI22xp33_ASAP7_75t_L g618 ( .A1(n_380), .A2(n_384), .B1(n_609), .B2(n_610), .Y(n_618) );
AOI222xp33_ASAP7_75t_L g794 ( .A1(n_380), .A2(n_384), .B1(n_565), .B2(n_795), .C1(n_796), .C2(n_797), .Y(n_794) );
AOI22xp33_ASAP7_75t_L g1093 ( .A1(n_380), .A2(n_384), .B1(n_1051), .B2(n_1052), .Y(n_1093) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g690 ( .A(n_382), .Y(n_690) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
AOI222xp33_ASAP7_75t_L g626 ( .A1(n_384), .A2(n_627), .B1(n_628), .B2(n_630), .C1(n_631), .C2(n_632), .Y(n_626) );
AOI22xp5_ASAP7_75t_L g687 ( .A1(n_384), .A2(n_688), .B1(n_689), .B2(n_691), .Y(n_687) );
AOI222xp33_ASAP7_75t_L g752 ( .A1(n_384), .A2(n_631), .B1(n_753), .B2(n_754), .C1(n_755), .C2(n_756), .Y(n_752) );
AOI222xp33_ASAP7_75t_L g912 ( .A1(n_384), .A2(n_631), .B1(n_913), .B2(n_914), .C1(n_916), .C2(n_917), .Y(n_912) );
AOI222xp33_ASAP7_75t_L g980 ( .A1(n_384), .A2(n_689), .B1(n_975), .B2(n_976), .C1(n_981), .C2(n_982), .Y(n_980) );
AOI222xp33_ASAP7_75t_L g1016 ( .A1(n_384), .A2(n_438), .B1(n_631), .B2(n_1004), .C1(n_1005), .C2(n_1017), .Y(n_1016) );
AOI222xp33_ASAP7_75t_L g1398 ( .A1(n_384), .A2(n_631), .B1(n_754), .B2(n_1399), .C1(n_1400), .C2(n_1401), .Y(n_1398) );
NAND4xp25_ASAP7_75t_L g745 ( .A(n_386), .B(n_746), .C(n_749), .D(n_752), .Y(n_745) );
BUFx2_ASAP7_75t_L g865 ( .A(n_386), .Y(n_865) );
NAND4xp25_ASAP7_75t_L g1390 ( .A(n_386), .B(n_1391), .C(n_1395), .D(n_1398), .Y(n_1390) );
INVx5_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
CKINVDCx8_ASAP7_75t_R g480 ( .A(n_387), .Y(n_480) );
NOR2xp33_ASAP7_75t_SL g685 ( .A(n_387), .B(n_686), .Y(n_685) );
AND2x4_ASAP7_75t_L g387 ( .A(n_388), .B(n_389), .Y(n_387) );
INVx2_ASAP7_75t_L g439 ( .A(n_389), .Y(n_439) );
BUFx6f_ASAP7_75t_L g479 ( .A(n_389), .Y(n_479) );
INVx1_ASAP7_75t_L g566 ( .A(n_389), .Y(n_566) );
BUFx6f_ASAP7_75t_L g1032 ( .A(n_389), .Y(n_1032) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
OAI31xp33_ASAP7_75t_SL g612 ( .A1(n_392), .A2(n_613), .A3(n_614), .B(n_615), .Y(n_612) );
OAI21xp5_ASAP7_75t_L g683 ( .A1(n_392), .A2(n_684), .B(n_695), .Y(n_683) );
AOI211x1_ASAP7_75t_SL g792 ( .A1(n_392), .A2(n_793), .B(n_804), .C(n_816), .Y(n_792) );
BUFx6f_ASAP7_75t_L g866 ( .A(n_392), .Y(n_866) );
AND2x4_ASAP7_75t_L g392 ( .A(n_393), .B(n_395), .Y(n_392) );
AND2x4_ASAP7_75t_L g487 ( .A(n_393), .B(n_395), .Y(n_487) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
AND2x4_ASAP7_75t_L g454 ( .A(n_394), .B(n_455), .Y(n_454) );
BUFx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx2_ASAP7_75t_L g417 ( .A(n_396), .Y(n_417) );
OR2x6_ASAP7_75t_L g570 ( .A(n_396), .B(n_571), .Y(n_570) );
NAND4xp25_ASAP7_75t_L g397 ( .A(n_398), .B(n_419), .C(n_434), .D(n_450), .Y(n_397) );
NAND3xp33_ASAP7_75t_L g398 ( .A(n_399), .B(n_407), .C(n_414), .Y(n_398) );
INVx3_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx2_ASAP7_75t_SL g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
BUFx3_ASAP7_75t_L g1138 ( .A(n_405), .Y(n_1138) );
INVx3_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx3_ASAP7_75t_L g580 ( .A(n_406), .Y(n_580) );
BUFx6f_ASAP7_75t_L g723 ( .A(n_406), .Y(n_723) );
BUFx3_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx2_ASAP7_75t_SL g708 ( .A(n_410), .Y(n_708) );
INVx2_ASAP7_75t_SL g1028 ( .A(n_410), .Y(n_1028) );
INVx3_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
BUFx6f_ASAP7_75t_L g650 ( .A(n_411), .Y(n_650) );
BUFx6f_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g710 ( .A(n_413), .Y(n_710) );
AND2x4_ASAP7_75t_L g1436 ( .A(n_413), .B(n_1409), .Y(n_1436) );
NAND3xp33_ASAP7_75t_L g879 ( .A(n_414), .B(n_880), .C(n_883), .Y(n_879) );
AOI33xp33_ASAP7_75t_L g1132 ( .A1(n_414), .A2(n_1133), .A3(n_1137), .B1(n_1139), .B2(n_1140), .B3(n_1141), .Y(n_1132) );
INVx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
BUFx3_ASAP7_75t_L g499 ( .A(n_416), .Y(n_499) );
AOI33xp33_ASAP7_75t_L g653 ( .A1(n_416), .A2(n_654), .A3(n_655), .B1(n_657), .B2(n_661), .B3(n_662), .Y(n_653) );
NAND3xp33_ASAP7_75t_L g758 ( .A(n_416), .B(n_759), .C(n_760), .Y(n_758) );
NAND3xp33_ASAP7_75t_L g931 ( .A(n_416), .B(n_932), .C(n_934), .Y(n_931) );
NAND3xp33_ASAP7_75t_L g951 ( .A(n_416), .B(n_952), .C(n_954), .Y(n_951) );
NAND3xp33_ASAP7_75t_L g1019 ( .A(n_416), .B(n_1020), .C(n_1021), .Y(n_1019) );
AND2x4_ASAP7_75t_L g416 ( .A(n_417), .B(n_418), .Y(n_416) );
OR2x6_ASAP7_75t_L g447 ( .A(n_417), .B(n_448), .Y(n_447) );
OR2x2_ASAP7_75t_L g508 ( .A(n_417), .B(n_448), .Y(n_508) );
OR2x2_ASAP7_75t_L g639 ( .A(n_417), .B(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_L g651 ( .A(n_417), .B(n_652), .Y(n_651) );
AND2x4_ASAP7_75t_L g704 ( .A(n_417), .B(n_418), .Y(n_704) );
BUFx2_ASAP7_75t_L g1444 ( .A(n_417), .Y(n_1444) );
NAND3xp33_ASAP7_75t_L g419 ( .A(n_420), .B(n_425), .C(n_428), .Y(n_419) );
INVxp67_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx2_ASAP7_75t_SL g423 ( .A(n_424), .Y(n_423) );
BUFx3_ASAP7_75t_L g491 ( .A(n_424), .Y(n_491) );
INVx2_ASAP7_75t_SL g882 ( .A(n_424), .Y(n_882) );
INVx4_ASAP7_75t_L g888 ( .A(n_424), .Y(n_888) );
INVx2_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
CKINVDCx8_ASAP7_75t_R g601 ( .A(n_428), .Y(n_601) );
AOI33xp33_ASAP7_75t_L g817 ( .A1(n_428), .A2(n_818), .A3(n_819), .B1(n_823), .B2(n_826), .B3(n_827), .Y(n_817) );
NAND3xp33_ASAP7_75t_L g885 ( .A(n_428), .B(n_886), .C(n_889), .Y(n_885) );
NAND3xp33_ASAP7_75t_L g935 ( .A(n_428), .B(n_936), .C(n_937), .Y(n_935) );
NAND3xp33_ASAP7_75t_L g1022 ( .A(n_428), .B(n_1023), .C(n_1026), .Y(n_1022) );
INVx5_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx6_ASAP7_75t_L g506 ( .A(n_429), .Y(n_506) );
OR2x6_ASAP7_75t_L g429 ( .A(n_430), .B(n_432), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g652 ( .A(n_432), .Y(n_652) );
NAND3xp33_ASAP7_75t_L g434 ( .A(n_435), .B(n_440), .C(n_446), .Y(n_434) );
BUFx3_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g862 ( .A(n_438), .Y(n_862) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx3_ASAP7_75t_L g839 ( .A(n_439), .Y(n_839) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx2_ASAP7_75t_SL g550 ( .A(n_443), .Y(n_550) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g736 ( .A(n_445), .Y(n_736) );
NAND3xp33_ASAP7_75t_L g890 ( .A(n_446), .B(n_891), .C(n_892), .Y(n_890) );
CKINVDCx5p33_ASAP7_75t_R g446 ( .A(n_447), .Y(n_446) );
OAI22xp5_ASAP7_75t_L g540 ( .A1(n_447), .A2(n_452), .B1(n_541), .B2(n_553), .Y(n_540) );
INVx2_ASAP7_75t_L g727 ( .A(n_447), .Y(n_727) );
CKINVDCx5p33_ASAP7_75t_R g1034 ( .A(n_447), .Y(n_1034) );
OAI22xp5_ASAP7_75t_L g1055 ( .A1(n_447), .A2(n_1056), .B1(n_1062), .B2(n_1067), .Y(n_1055) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g640 ( .A(n_449), .Y(n_640) );
NAND3xp33_ASAP7_75t_L g450 ( .A(n_451), .B(n_456), .C(n_461), .Y(n_450) );
AOI33xp33_ASAP7_75t_L g1123 ( .A1(n_451), .A2(n_727), .A3(n_1124), .B1(n_1126), .B2(n_1129), .B3(n_1130), .Y(n_1123) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
OAI22xp5_ASAP7_75t_SL g507 ( .A1(n_452), .A2(n_508), .B1(n_509), .B2(n_516), .Y(n_507) );
INVx4_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
BUFx4f_ASAP7_75t_L g741 ( .A(n_453), .Y(n_741) );
BUFx4f_ASAP7_75t_L g903 ( .A(n_453), .Y(n_903) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx2_ASAP7_75t_SL g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
HB1xp67_ASAP7_75t_L g1128 ( .A(n_464), .Y(n_1128) );
XNOR2xp5_ASAP7_75t_L g465 ( .A(n_466), .B(n_467), .Y(n_465) );
NAND3x1_ASAP7_75t_SL g467 ( .A(n_468), .B(n_488), .C(n_521), .Y(n_467) );
OAI31xp33_ASAP7_75t_L g468 ( .A1(n_469), .A2(n_476), .A3(n_484), .B(n_487), .Y(n_468) );
OR2x2_ASAP7_75t_L g470 ( .A(n_471), .B(n_472), .Y(n_470) );
INVx2_ASAP7_75t_L g511 ( .A(n_472), .Y(n_511) );
BUFx2_ASAP7_75t_L g543 ( .A(n_472), .Y(n_543) );
INVx1_ASAP7_75t_L g556 ( .A(n_472), .Y(n_556) );
OR2x2_ASAP7_75t_L g472 ( .A(n_473), .B(n_474), .Y(n_472) );
AND2x2_ASAP7_75t_L g514 ( .A(n_473), .B(n_474), .Y(n_514) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
NAND4xp25_ASAP7_75t_L g622 ( .A(n_480), .B(n_623), .C(n_626), .D(n_633), .Y(n_622) );
NAND4xp25_ASAP7_75t_SL g793 ( .A(n_480), .B(n_794), .C(n_798), .D(n_801), .Y(n_793) );
NAND3xp33_ASAP7_75t_SL g911 ( .A(n_480), .B(n_912), .C(n_918), .Y(n_911) );
NAND3xp33_ASAP7_75t_SL g979 ( .A(n_480), .B(n_980), .C(n_983), .Y(n_979) );
NAND4xp25_ASAP7_75t_SL g1010 ( .A(n_480), .B(n_1011), .C(n_1014), .D(n_1016), .Y(n_1010) );
AOI211x1_ASAP7_75t_L g621 ( .A1(n_487), .A2(n_622), .B(n_636), .C(n_664), .Y(n_621) );
AOI211xp5_ASAP7_75t_L g744 ( .A1(n_487), .A2(n_745), .B(n_757), .C(n_777), .Y(n_744) );
OAI21xp5_ASAP7_75t_L g910 ( .A1(n_487), .A2(n_911), .B(n_921), .Y(n_910) );
OAI21xp5_ASAP7_75t_SL g978 ( .A1(n_487), .A2(n_979), .B(n_986), .Y(n_978) );
OAI31xp33_ASAP7_75t_SL g1090 ( .A1(n_487), .A2(n_1091), .A3(n_1092), .B(n_1094), .Y(n_1090) );
AOI221xp5_ASAP7_75t_L g488 ( .A1(n_489), .A2(n_499), .B1(n_500), .B2(n_506), .C(n_507), .Y(n_488) );
OAI22xp33_ASAP7_75t_L g492 ( .A1(n_493), .A2(n_494), .B1(n_495), .B2(n_496), .Y(n_492) );
OAI221xp5_ASAP7_75t_L g509 ( .A1(n_493), .A2(n_495), .B1(n_510), .B2(n_512), .C(n_515), .Y(n_509) );
OAI22xp33_ASAP7_75t_SL g501 ( .A1(n_496), .A2(n_502), .B1(n_503), .B2(n_505), .Y(n_501) );
INVx1_ASAP7_75t_L g586 ( .A(n_496), .Y(n_586) );
BUFx2_ASAP7_75t_L g1049 ( .A(n_496), .Y(n_1049) );
OAI21xp5_ASAP7_75t_SL g1429 ( .A1(n_496), .A2(n_1399), .B(n_1430), .Y(n_1429) );
INVx3_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
BUFx2_ASAP7_75t_L g599 ( .A(n_497), .Y(n_599) );
INVx2_ASAP7_75t_L g973 ( .A(n_497), .Y(n_973) );
INVx2_ASAP7_75t_L g1087 ( .A(n_497), .Y(n_1087) );
INVx3_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
AOI33xp33_ASAP7_75t_L g703 ( .A1(n_506), .A2(n_704), .A3(n_705), .B1(n_711), .B2(n_718), .B3(n_721), .Y(n_703) );
NAND3xp33_ASAP7_75t_L g955 ( .A(n_506), .B(n_956), .C(n_958), .Y(n_955) );
INVx1_ASAP7_75t_L g1089 ( .A(n_506), .Y(n_1089) );
OAI221xp5_ASAP7_75t_L g516 ( .A1(n_510), .A2(n_512), .B1(n_517), .B2(n_518), .C(n_519), .Y(n_516) );
OAI221xp5_ASAP7_75t_L g1056 ( .A1(n_510), .A2(n_616), .B1(n_1057), .B2(n_1058), .C(n_1059), .Y(n_1056) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
HB1xp67_ASAP7_75t_L g1452 ( .A(n_511), .Y(n_1452) );
BUFx3_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g617 ( .A(n_513), .Y(n_617) );
OAI221xp5_ASAP7_75t_SL g1446 ( .A1(n_513), .A2(n_555), .B1(n_1426), .B2(n_1447), .C(n_1448), .Y(n_1446) );
INVx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g546 ( .A(n_514), .Y(n_546) );
BUFx2_ASAP7_75t_L g1455 ( .A(n_514), .Y(n_1455) );
BUFx6f_ASAP7_75t_L g944 ( .A(n_520), .Y(n_944) );
BUFx3_ASAP7_75t_L g1039 ( .A(n_520), .Y(n_1039) );
BUFx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
OR2x2_ASAP7_75t_L g529 ( .A(n_530), .B(n_531), .Y(n_529) );
BUFx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g576 ( .A(n_532), .Y(n_576) );
INVx1_ASAP7_75t_L g591 ( .A(n_532), .Y(n_591) );
INVx5_ASAP7_75t_SL g533 ( .A(n_534), .Y(n_533) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_536), .A2(n_680), .B1(n_787), .B2(n_788), .Y(n_535) );
INVx1_ASAP7_75t_L g787 ( .A(n_536), .Y(n_787) );
AOI22xp5_ASAP7_75t_L g536 ( .A1(n_537), .A2(n_619), .B1(n_620), .B2(n_679), .Y(n_536) );
INVx1_ASAP7_75t_L g679 ( .A(n_537), .Y(n_679) );
NAND3xp33_ASAP7_75t_L g538 ( .A(n_539), .B(n_602), .C(n_612), .Y(n_538) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_540), .B(n_567), .Y(n_539) );
OAI221xp5_ASAP7_75t_L g541 ( .A1(n_542), .A2(n_543), .B1(n_544), .B2(n_547), .C(n_548), .Y(n_541) );
OAI22xp33_ASAP7_75t_L g582 ( .A1(n_542), .A2(n_547), .B1(n_583), .B2(n_585), .Y(n_582) );
OAI221xp5_ASAP7_75t_L g1062 ( .A1(n_543), .A2(n_1063), .B1(n_1064), .B2(n_1065), .C(n_1066), .Y(n_1062) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
BUFx2_ASAP7_75t_L g1064 ( .A(n_546), .Y(n_1064) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g896 ( .A(n_552), .Y(n_896) );
OAI221xp5_ASAP7_75t_L g553 ( .A1(n_554), .A2(n_557), .B1(n_558), .B2(n_560), .C(n_561), .Y(n_553) );
BUFx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx2_ASAP7_75t_L g730 ( .A(n_564), .Y(n_730) );
BUFx2_ASAP7_75t_L g1125 ( .A(n_564), .Y(n_1125) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
OAI33xp33_ASAP7_75t_L g567 ( .A1(n_568), .A2(n_572), .A3(n_582), .B1(n_587), .B2(n_593), .B3(n_601), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
OAI33xp33_ASAP7_75t_L g1068 ( .A1(n_570), .A2(n_1069), .A3(n_1072), .B1(n_1078), .B2(n_1083), .B3(n_1089), .Y(n_1068) );
OAI22xp5_ASAP7_75t_L g572 ( .A1(n_573), .A2(n_574), .B1(n_577), .B2(n_581), .Y(n_572) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx2_ASAP7_75t_SL g1074 ( .A(n_575), .Y(n_1074) );
INVx2_ASAP7_75t_L g1080 ( .A(n_575), .Y(n_1080) );
BUFx3_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx2_ASAP7_75t_L g596 ( .A(n_580), .Y(n_596) );
INVx2_ASAP7_75t_L g825 ( .A(n_580), .Y(n_825) );
OAI22xp33_ASAP7_75t_L g587 ( .A1(n_583), .A2(n_588), .B1(n_589), .B2(n_592), .Y(n_587) );
INVx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
HB1xp67_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
OAI22xp33_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_597), .B1(n_598), .B2(n_600), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx2_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVx2_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g925 ( .A(n_599), .Y(n_925) );
INVx1_ASAP7_75t_L g1071 ( .A(n_599), .Y(n_1071) );
INVx1_ASAP7_75t_L g1141 ( .A(n_601), .Y(n_1141) );
BUFx3_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
BUFx6f_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx2_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g678 ( .A(n_621), .Y(n_678) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_637), .B(n_653), .Y(n_636) );
AOI33xp33_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_641), .A3(n_642), .B1(n_645), .B2(n_647), .B3(n_651), .Y(n_637) );
NAND3xp33_ASAP7_75t_L g767 ( .A(n_638), .B(n_768), .C(n_769), .Y(n_767) );
NAND3xp33_ASAP7_75t_L g939 ( .A(n_638), .B(n_940), .C(n_943), .Y(n_939) );
NAND3xp33_ASAP7_75t_L g959 ( .A(n_638), .B(n_960), .C(n_961), .Y(n_959) );
INVx3_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx2_ASAP7_75t_SL g656 ( .A(n_644), .Y(n_656) );
INVx2_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx2_ASAP7_75t_SL g663 ( .A(n_649), .Y(n_663) );
INVx3_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
BUFx2_ASAP7_75t_L g766 ( .A(n_650), .Y(n_766) );
BUFx6f_ASAP7_75t_L g1136 ( .A(n_650), .Y(n_1136) );
AND2x4_ASAP7_75t_L g1438 ( .A(n_650), .B(n_1406), .Y(n_1438) );
NAND3xp33_ASAP7_75t_L g761 ( .A(n_651), .B(n_762), .C(n_765), .Y(n_761) );
INVx1_ASAP7_75t_L g1431 ( .A(n_652), .Y(n_1431) );
NAND3xp33_ASAP7_75t_L g772 ( .A(n_654), .B(n_773), .C(n_774), .Y(n_772) );
AOI33xp33_ASAP7_75t_L g830 ( .A1(n_654), .A2(n_727), .A3(n_831), .B1(n_836), .B2(n_840), .B3(n_844), .Y(n_830) );
NAND3xp33_ASAP7_75t_L g945 ( .A(n_654), .B(n_946), .C(n_947), .Y(n_945) );
NAND3xp33_ASAP7_75t_L g964 ( .A(n_654), .B(n_965), .C(n_966), .Y(n_964) );
BUFx2_ASAP7_75t_L g1131 ( .A(n_656), .Y(n_1131) );
BUFx2_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx2_ASAP7_75t_L g1061 ( .A(n_659), .Y(n_1061) );
INVx2_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
AOI31xp33_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_670), .A3(n_673), .B(n_676), .Y(n_664) );
AO21x1_ASAP7_75t_SL g696 ( .A1(n_676), .A2(n_697), .B(n_700), .Y(n_696) );
AOI31xp33_ASAP7_75t_L g804 ( .A1(n_676), .A2(n_805), .A3(n_807), .B(n_813), .Y(n_804) );
INVx1_ASAP7_75t_L g788 ( .A(n_680), .Y(n_788) );
AO22x2_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_742), .B1(n_743), .B2(n_786), .Y(n_680) );
INVx1_ASAP7_75t_L g786 ( .A(n_681), .Y(n_786) );
NAND4xp25_ASAP7_75t_L g682 ( .A(n_683), .B(n_696), .C(n_703), .D(n_726), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_685), .B(n_692), .Y(n_684) );
BUFx2_ASAP7_75t_L g818 ( .A(n_704), .Y(n_818) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
BUFx2_ASAP7_75t_L g820 ( .A(n_708), .Y(n_820) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx2_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g1025 ( .A(n_716), .Y(n_1025) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx2_ASAP7_75t_L g1411 ( .A(n_717), .Y(n_1411) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g828 ( .A(n_720), .Y(n_828) );
INVx1_ASAP7_75t_L g933 ( .A(n_720), .Y(n_933) );
INVx1_ASAP7_75t_L g1082 ( .A(n_722), .Y(n_1082) );
INVx2_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx2_ASAP7_75t_SL g764 ( .A(n_723), .Y(n_764) );
INVx2_ASAP7_75t_L g953 ( .A(n_723), .Y(n_953) );
INVx2_ASAP7_75t_L g957 ( .A(n_723), .Y(n_957) );
INVx3_ASAP7_75t_L g1077 ( .A(n_723), .Y(n_1077) );
BUFx2_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx2_ASAP7_75t_SL g822 ( .A(n_725), .Y(n_822) );
AOI33xp33_ASAP7_75t_L g726 ( .A1(n_727), .A2(n_728), .A3(n_733), .B1(n_737), .B2(n_739), .B3(n_741), .Y(n_726) );
INVx1_ASAP7_75t_L g1449 ( .A(n_727), .Y(n_1449) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g942 ( .A(n_732), .Y(n_942) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx4_ASAP7_75t_L g738 ( .A(n_735), .Y(n_738) );
CKINVDCx5p33_ASAP7_75t_R g1067 ( .A(n_741), .Y(n_1067) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
NAND4xp25_ASAP7_75t_L g757 ( .A(n_758), .B(n_761), .C(n_767), .D(n_772), .Y(n_757) );
INVx2_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVx1_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
AO22x1_ASAP7_75t_L g789 ( .A1(n_790), .A2(n_907), .B1(n_988), .B2(n_989), .Y(n_789) );
INVx1_ASAP7_75t_L g988 ( .A(n_790), .Y(n_988) );
AOI22xp5_ASAP7_75t_L g790 ( .A1(n_791), .A2(n_849), .B1(n_850), .B2(n_906), .Y(n_790) );
INVx1_ASAP7_75t_L g906 ( .A(n_791), .Y(n_906) );
INVx1_ASAP7_75t_L g848 ( .A(n_792), .Y(n_848) );
INVx2_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g816 ( .A(n_817), .B(n_830), .Y(n_816) );
INVx2_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
INVx2_ASAP7_75t_L g938 ( .A(n_822), .Y(n_938) );
INVx2_ASAP7_75t_SL g824 ( .A(n_825), .Y(n_824) );
INVx2_ASAP7_75t_L g829 ( .A(n_825), .Y(n_829) );
BUFx4f_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
INVx1_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
HB1xp67_ASAP7_75t_L g1127 ( .A(n_837), .Y(n_1127) );
BUFx6f_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
INVx2_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
INVx1_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
INVx1_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
INVx1_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
INVx1_ASAP7_75t_L g905 ( .A(n_851), .Y(n_905) );
NAND4xp25_ASAP7_75t_L g852 ( .A(n_853), .B(n_856), .C(n_859), .D(n_865), .Y(n_852) );
INVx1_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
NAND4xp25_ASAP7_75t_SL g1113 ( .A(n_865), .B(n_1114), .C(n_1116), .D(n_1118), .Y(n_1113) );
AOI221x1_ASAP7_75t_L g1389 ( .A1(n_866), .A2(n_1390), .B1(n_1402), .B2(n_1442), .C(n_1445), .Y(n_1389) );
INVx1_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
INVx1_ASAP7_75t_L g884 ( .A(n_874), .Y(n_884) );
INVx1_ASAP7_75t_L g1107 ( .A(n_874), .Y(n_1107) );
INVx1_ASAP7_75t_L g874 ( .A(n_875), .Y(n_874) );
NAND4xp25_ASAP7_75t_L g878 ( .A(n_879), .B(n_885), .C(n_890), .D(n_897), .Y(n_878) );
INVx1_ASAP7_75t_L g881 ( .A(n_882), .Y(n_881) );
INVx2_ASAP7_75t_L g887 ( .A(n_888), .Y(n_887) );
INVx2_ASAP7_75t_SL g893 ( .A(n_894), .Y(n_893) );
INVx2_ASAP7_75t_L g894 ( .A(n_895), .Y(n_894) );
BUFx3_ASAP7_75t_L g1038 ( .A(n_895), .Y(n_1038) );
NAND3xp33_ASAP7_75t_L g897 ( .A(n_898), .B(n_901), .C(n_903), .Y(n_897) );
INVx1_ASAP7_75t_L g899 ( .A(n_900), .Y(n_899) );
NAND3xp33_ASAP7_75t_L g1035 ( .A(n_903), .B(n_1036), .C(n_1037), .Y(n_1035) );
OAI22xp5_ASAP7_75t_L g1250 ( .A1(n_904), .A2(n_1251), .B1(n_1252), .B2(n_1253), .Y(n_1250) );
INVx2_ASAP7_75t_L g989 ( .A(n_907), .Y(n_989) );
XOR2x2_ASAP7_75t_L g907 ( .A(n_908), .B(n_948), .Y(n_907) );
NAND3x1_ASAP7_75t_L g909 ( .A(n_910), .B(n_922), .C(n_930), .Y(n_909) );
INVx1_ASAP7_75t_L g914 ( .A(n_915), .Y(n_914) );
INVx1_ASAP7_75t_L g982 ( .A(n_915), .Y(n_982) );
INVx1_ASAP7_75t_L g927 ( .A(n_928), .Y(n_927) );
AND4x1_ASAP7_75t_L g930 ( .A(n_931), .B(n_935), .C(n_939), .D(n_945), .Y(n_930) );
XOR2xp5_ASAP7_75t_L g948 ( .A(n_949), .B(n_987), .Y(n_948) );
NAND3xp33_ASAP7_75t_L g949 ( .A(n_950), .B(n_968), .C(n_978), .Y(n_949) );
AND4x1_ASAP7_75t_L g950 ( .A(n_951), .B(n_955), .C(n_959), .D(n_964), .Y(n_950) );
INVx2_ASAP7_75t_L g962 ( .A(n_963), .Y(n_962) );
INVx1_ASAP7_75t_L g971 ( .A(n_972), .Y(n_971) );
INVx1_ASAP7_75t_L g972 ( .A(n_973), .Y(n_972) );
OR2x6_ASAP7_75t_L g1433 ( .A(n_973), .B(n_1418), .Y(n_1433) );
INVx1_ASAP7_75t_L g990 ( .A(n_991), .Y(n_990) );
OAI22xp5_ASAP7_75t_L g991 ( .A1(n_992), .A2(n_993), .B1(n_1097), .B2(n_1098), .Y(n_991) );
INVx1_ASAP7_75t_L g992 ( .A(n_993), .Y(n_992) );
AOI22xp5_ASAP7_75t_L g993 ( .A1(n_994), .A2(n_995), .B1(n_1042), .B2(n_1043), .Y(n_993) );
INVx1_ASAP7_75t_L g994 ( .A(n_995), .Y(n_994) );
HB1xp67_ASAP7_75t_L g995 ( .A(n_996), .Y(n_995) );
INVx1_ASAP7_75t_L g1041 ( .A(n_997), .Y(n_1041) );
NAND4xp25_ASAP7_75t_SL g1018 ( .A(n_1019), .B(n_1022), .C(n_1029), .D(n_1035), .Y(n_1018) );
INVx1_ASAP7_75t_L g1024 ( .A(n_1025), .Y(n_1024) );
BUFx2_ASAP7_75t_L g1027 ( .A(n_1028), .Y(n_1027) );
NAND2xp5_ASAP7_75t_L g1440 ( .A(n_1028), .B(n_1441), .Y(n_1440) );
NAND3xp33_ASAP7_75t_L g1029 ( .A(n_1030), .B(n_1033), .C(n_1034), .Y(n_1029) );
BUFx6f_ASAP7_75t_L g1031 ( .A(n_1032), .Y(n_1031) );
INVx1_ASAP7_75t_L g1042 ( .A(n_1043), .Y(n_1042) );
HB1xp67_ASAP7_75t_L g1043 ( .A(n_1044), .Y(n_1043) );
INVx1_ASAP7_75t_L g1095 ( .A(n_1045), .Y(n_1095) );
NAND3xp33_ASAP7_75t_L g1045 ( .A(n_1046), .B(n_1054), .C(n_1090), .Y(n_1045) );
NOR2xp33_ASAP7_75t_L g1054 ( .A(n_1055), .B(n_1068), .Y(n_1054) );
OAI22xp33_ASAP7_75t_L g1069 ( .A1(n_1057), .A2(n_1058), .B1(n_1070), .B2(n_1071), .Y(n_1069) );
INVx2_ASAP7_75t_SL g1060 ( .A(n_1061), .Y(n_1060) );
OAI22xp5_ASAP7_75t_L g1445 ( .A1(n_1067), .A2(n_1446), .B1(n_1449), .B2(n_1450), .Y(n_1445) );
OAI22xp5_ASAP7_75t_L g1072 ( .A1(n_1073), .A2(n_1074), .B1(n_1075), .B2(n_1076), .Y(n_1072) );
INVx1_ASAP7_75t_L g1076 ( .A(n_1077), .Y(n_1076) );
OAI22xp5_ASAP7_75t_SL g1078 ( .A1(n_1079), .A2(n_1080), .B1(n_1081), .B2(n_1082), .Y(n_1078) );
OAI22xp33_ASAP7_75t_L g1083 ( .A1(n_1084), .A2(n_1086), .B1(n_1087), .B2(n_1088), .Y(n_1083) );
INVx2_ASAP7_75t_L g1084 ( .A(n_1085), .Y(n_1084) );
INVx2_ASAP7_75t_SL g1097 ( .A(n_1098), .Y(n_1097) );
OAI22xp33_ASAP7_75t_L g1151 ( .A1(n_1099), .A2(n_1152), .B1(n_1153), .B2(n_1160), .Y(n_1151) );
INVx1_ASAP7_75t_L g1142 ( .A(n_1100), .Y(n_1142) );
NAND2xp5_ASAP7_75t_L g1122 ( .A(n_1123), .B(n_1132), .Y(n_1122) );
INVx1_ASAP7_75t_L g1134 ( .A(n_1135), .Y(n_1134) );
INVx1_ASAP7_75t_L g1135 ( .A(n_1136), .Y(n_1135) );
OAI221xp5_ASAP7_75t_SL g1144 ( .A1(n_1145), .A2(n_1383), .B1(n_1386), .B2(n_1457), .C(n_1463), .Y(n_1144) );
AND5x1_ASAP7_75t_L g1145 ( .A(n_1146), .B(n_1293), .C(n_1331), .D(n_1343), .E(n_1366), .Y(n_1145) );
A2O1A1Ixp33_ASAP7_75t_L g1146 ( .A1(n_1147), .A2(n_1149), .B(n_1236), .C(n_1269), .Y(n_1146) );
OAI211xp5_ASAP7_75t_L g1147 ( .A1(n_1148), .A2(n_1183), .B(n_1223), .C(n_1225), .Y(n_1147) );
OR2x2_ASAP7_75t_L g1148 ( .A(n_1149), .B(n_1174), .Y(n_1148) );
INVx1_ASAP7_75t_L g1234 ( .A(n_1149), .Y(n_1234) );
INVx3_ASAP7_75t_L g1255 ( .A(n_1149), .Y(n_1255) );
AND2x2_ASAP7_75t_L g1265 ( .A(n_1149), .B(n_1215), .Y(n_1265) );
AND2x2_ASAP7_75t_L g1267 ( .A(n_1149), .B(n_1268), .Y(n_1267) );
AND2x2_ASAP7_75t_L g1323 ( .A(n_1149), .B(n_1279), .Y(n_1323) );
AND2x2_ASAP7_75t_L g1325 ( .A(n_1149), .B(n_1174), .Y(n_1325) );
INVx3_ASAP7_75t_L g1149 ( .A(n_1150), .Y(n_1149) );
AND2x2_ASAP7_75t_L g1235 ( .A(n_1150), .B(n_1174), .Y(n_1235) );
OR2x2_ASAP7_75t_L g1257 ( .A(n_1150), .B(n_1258), .Y(n_1257) );
OR2x2_ASAP7_75t_L g1150 ( .A(n_1151), .B(n_1164), .Y(n_1150) );
OAI22xp5_ASAP7_75t_L g1204 ( .A1(n_1153), .A2(n_1162), .B1(n_1205), .B2(n_1206), .Y(n_1204) );
OAI22xp33_ASAP7_75t_L g1217 ( .A1(n_1153), .A2(n_1162), .B1(n_1218), .B2(n_1219), .Y(n_1217) );
BUFx3_ASAP7_75t_L g1252 ( .A(n_1153), .Y(n_1252) );
BUFx6f_ASAP7_75t_L g1153 ( .A(n_1154), .Y(n_1153) );
OR2x2_ASAP7_75t_L g1154 ( .A(n_1155), .B(n_1156), .Y(n_1154) );
OR2x2_ASAP7_75t_L g1162 ( .A(n_1155), .B(n_1163), .Y(n_1162) );
INVx1_ASAP7_75t_L g1178 ( .A(n_1155), .Y(n_1178) );
INVx1_ASAP7_75t_L g1177 ( .A(n_1156), .Y(n_1177) );
NAND2xp5_ASAP7_75t_L g1156 ( .A(n_1157), .B(n_1159), .Y(n_1156) );
INVx1_ASAP7_75t_L g1157 ( .A(n_1158), .Y(n_1157) );
INVx1_ASAP7_75t_L g1169 ( .A(n_1159), .Y(n_1169) );
HB1xp67_ASAP7_75t_L g1253 ( .A(n_1160), .Y(n_1253) );
INVx1_ASAP7_75t_L g1160 ( .A(n_1161), .Y(n_1160) );
INVx1_ASAP7_75t_L g1161 ( .A(n_1162), .Y(n_1161) );
INVx1_ASAP7_75t_L g1180 ( .A(n_1163), .Y(n_1180) );
OAI22xp5_ASAP7_75t_L g1164 ( .A1(n_1165), .A2(n_1166), .B1(n_1171), .B2(n_1172), .Y(n_1164) );
INVx1_ASAP7_75t_L g1166 ( .A(n_1167), .Y(n_1166) );
INVx1_ASAP7_75t_L g1248 ( .A(n_1167), .Y(n_1248) );
AND2x4_ASAP7_75t_L g1167 ( .A(n_1168), .B(n_1170), .Y(n_1167) );
AND2x2_ASAP7_75t_L g1182 ( .A(n_1168), .B(n_1170), .Y(n_1182) );
INVx1_ASAP7_75t_L g1168 ( .A(n_1169), .Y(n_1168) );
AND2x4_ASAP7_75t_L g1173 ( .A(n_1169), .B(n_1170), .Y(n_1173) );
OAI22xp5_ASAP7_75t_L g1200 ( .A1(n_1172), .A2(n_1201), .B1(n_1202), .B2(n_1203), .Y(n_1200) );
INVx1_ASAP7_75t_SL g1172 ( .A(n_1173), .Y(n_1172) );
INVx2_ASAP7_75t_L g1197 ( .A(n_1173), .Y(n_1197) );
AND2x2_ASAP7_75t_L g1231 ( .A(n_1174), .B(n_1215), .Y(n_1231) );
OR2x2_ASAP7_75t_L g1242 ( .A(n_1174), .B(n_1215), .Y(n_1242) );
OR2x2_ASAP7_75t_L g1258 ( .A(n_1174), .B(n_1216), .Y(n_1258) );
INVx2_ASAP7_75t_L g1268 ( .A(n_1174), .Y(n_1268) );
AND2x2_ASAP7_75t_L g1279 ( .A(n_1174), .B(n_1216), .Y(n_1279) );
OAI211xp5_ASAP7_75t_L g1307 ( .A1(n_1174), .A2(n_1308), .B(n_1310), .C(n_1313), .Y(n_1307) );
OAI221xp5_ASAP7_75t_L g1333 ( .A1(n_1174), .A2(n_1223), .B1(n_1334), .B2(n_1336), .C(n_1337), .Y(n_1333) );
OAI211xp5_ASAP7_75t_L g1345 ( .A1(n_1174), .A2(n_1346), .B(n_1348), .C(n_1354), .Y(n_1345) );
AND2x4_ASAP7_75t_L g1174 ( .A(n_1175), .B(n_1181), .Y(n_1174) );
AND2x4_ASAP7_75t_L g1176 ( .A(n_1177), .B(n_1178), .Y(n_1176) );
AND2x4_ASAP7_75t_L g1179 ( .A(n_1178), .B(n_1180), .Y(n_1179) );
HB1xp67_ASAP7_75t_L g1474 ( .A(n_1180), .Y(n_1474) );
INVx1_ASAP7_75t_L g1201 ( .A(n_1182), .Y(n_1201) );
AOI211xp5_ASAP7_75t_L g1183 ( .A1(n_1184), .A2(n_1192), .B(n_1207), .C(n_1210), .Y(n_1183) );
AOI21xp33_ASAP7_75t_L g1287 ( .A1(n_1184), .A2(n_1288), .B(n_1290), .Y(n_1287) );
AOI21xp5_ASAP7_75t_L g1341 ( .A1(n_1184), .A2(n_1290), .B(n_1327), .Y(n_1341) );
INVx1_ASAP7_75t_L g1184 ( .A(n_1185), .Y(n_1184) );
AND2x2_ASAP7_75t_L g1240 ( .A(n_1185), .B(n_1208), .Y(n_1240) );
AND2x2_ASAP7_75t_L g1283 ( .A(n_1185), .B(n_1198), .Y(n_1283) );
NAND2xp5_ASAP7_75t_L g1295 ( .A(n_1185), .B(n_1192), .Y(n_1295) );
NAND2xp5_ASAP7_75t_L g1305 ( .A(n_1185), .B(n_1193), .Y(n_1305) );
AND2x2_ASAP7_75t_L g1185 ( .A(n_1186), .B(n_1189), .Y(n_1185) );
OR2x2_ASAP7_75t_L g1209 ( .A(n_1186), .B(n_1189), .Y(n_1209) );
AND2x2_ASAP7_75t_L g1221 ( .A(n_1186), .B(n_1222), .Y(n_1221) );
NOR2xp33_ASAP7_75t_L g1229 ( .A(n_1186), .B(n_1230), .Y(n_1229) );
INVx1_ASAP7_75t_L g1263 ( .A(n_1186), .Y(n_1263) );
AND2x2_ASAP7_75t_L g1340 ( .A(n_1186), .B(n_1199), .Y(n_1340) );
AND2x2_ASAP7_75t_L g1186 ( .A(n_1187), .B(n_1188), .Y(n_1186) );
INVx1_ASAP7_75t_L g1222 ( .A(n_1189), .Y(n_1222) );
AND2x2_ASAP7_75t_L g1262 ( .A(n_1189), .B(n_1263), .Y(n_1262) );
AND2x2_ASAP7_75t_L g1278 ( .A(n_1189), .B(n_1198), .Y(n_1278) );
NOR2xp33_ASAP7_75t_L g1289 ( .A(n_1189), .B(n_1198), .Y(n_1289) );
AND2x2_ASAP7_75t_L g1319 ( .A(n_1189), .B(n_1192), .Y(n_1319) );
NAND2xp5_ASAP7_75t_L g1261 ( .A(n_1192), .B(n_1262), .Y(n_1261) );
NAND2xp5_ASAP7_75t_L g1299 ( .A(n_1192), .B(n_1300), .Y(n_1299) );
AND2x2_ASAP7_75t_L g1192 ( .A(n_1193), .B(n_1198), .Y(n_1192) );
INVx4_ASAP7_75t_L g1208 ( .A(n_1193), .Y(n_1208) );
INVx2_ASAP7_75t_L g1212 ( .A(n_1193), .Y(n_1212) );
OR2x2_ASAP7_75t_L g1223 ( .A(n_1193), .B(n_1224), .Y(n_1223) );
OR2x2_ASAP7_75t_L g1276 ( .A(n_1193), .B(n_1209), .Y(n_1276) );
OR2x2_ASAP7_75t_L g1330 ( .A(n_1193), .B(n_1213), .Y(n_1330) );
NAND2xp5_ASAP7_75t_L g1346 ( .A(n_1193), .B(n_1347), .Y(n_1346) );
NOR2xp33_ASAP7_75t_L g1357 ( .A(n_1193), .B(n_1198), .Y(n_1357) );
AND2x6_ASAP7_75t_L g1193 ( .A(n_1194), .B(n_1195), .Y(n_1193) );
INVx2_ASAP7_75t_L g1196 ( .A(n_1197), .Y(n_1196) );
OAI22xp5_ASAP7_75t_L g1246 ( .A1(n_1197), .A2(n_1247), .B1(n_1248), .B2(n_1249), .Y(n_1246) );
OR2x2_ASAP7_75t_L g1228 ( .A(n_1198), .B(n_1222), .Y(n_1228) );
AND2x2_ASAP7_75t_L g1260 ( .A(n_1198), .B(n_1222), .Y(n_1260) );
NOR2xp33_ASAP7_75t_L g1304 ( .A(n_1198), .B(n_1305), .Y(n_1304) );
AND2x2_ASAP7_75t_L g1306 ( .A(n_1198), .B(n_1262), .Y(n_1306) );
AND2x2_ASAP7_75t_L g1335 ( .A(n_1198), .B(n_1240), .Y(n_1335) );
CKINVDCx6p67_ASAP7_75t_R g1198 ( .A(n_1199), .Y(n_1198) );
OR2x2_ASAP7_75t_L g1224 ( .A(n_1199), .B(n_1209), .Y(n_1224) );
NAND2xp5_ASAP7_75t_L g1239 ( .A(n_1199), .B(n_1240), .Y(n_1239) );
OR2x2_ASAP7_75t_L g1286 ( .A(n_1199), .B(n_1263), .Y(n_1286) );
AND2x2_ASAP7_75t_L g1309 ( .A(n_1199), .B(n_1262), .Y(n_1309) );
AND2x2_ASAP7_75t_L g1328 ( .A(n_1199), .B(n_1300), .Y(n_1328) );
AND2x2_ASAP7_75t_L g1347 ( .A(n_1199), .B(n_1221), .Y(n_1347) );
AND2x2_ASAP7_75t_L g1365 ( .A(n_1199), .B(n_1263), .Y(n_1365) );
OR2x6_ASAP7_75t_SL g1199 ( .A(n_1200), .B(n_1204), .Y(n_1199) );
NOR2xp33_ASAP7_75t_L g1207 ( .A(n_1208), .B(n_1209), .Y(n_1207) );
NAND2xp5_ASAP7_75t_L g1230 ( .A(n_1208), .B(n_1231), .Y(n_1230) );
INVx1_ASAP7_75t_L g1292 ( .A(n_1208), .Y(n_1292) );
AND2x2_ASAP7_75t_L g1314 ( .A(n_1208), .B(n_1315), .Y(n_1314) );
AND2x2_ASAP7_75t_L g1371 ( .A(n_1208), .B(n_1365), .Y(n_1371) );
INVx1_ASAP7_75t_L g1300 ( .A(n_1209), .Y(n_1300) );
NOR2xp33_ASAP7_75t_L g1210 ( .A(n_1211), .B(n_1220), .Y(n_1210) );
INVx1_ASAP7_75t_L g1312 ( .A(n_1211), .Y(n_1312) );
NAND2xp5_ASAP7_75t_L g1211 ( .A(n_1212), .B(n_1213), .Y(n_1211) );
INVx2_ASAP7_75t_L g1227 ( .A(n_1212), .Y(n_1227) );
AND2x2_ASAP7_75t_L g1277 ( .A(n_1212), .B(n_1278), .Y(n_1277) );
AND2x2_ASAP7_75t_L g1284 ( .A(n_1212), .B(n_1285), .Y(n_1284) );
NAND2xp5_ASAP7_75t_L g1308 ( .A(n_1212), .B(n_1309), .Y(n_1308) );
OAI21xp33_ASAP7_75t_L g1326 ( .A1(n_1212), .A2(n_1288), .B(n_1327), .Y(n_1326) );
NAND2xp5_ASAP7_75t_L g1339 ( .A(n_1212), .B(n_1340), .Y(n_1339) );
NOR2xp33_ASAP7_75t_L g1351 ( .A(n_1212), .B(n_1268), .Y(n_1351) );
INVx1_ASAP7_75t_L g1213 ( .A(n_1214), .Y(n_1213) );
INVx1_ASAP7_75t_L g1233 ( .A(n_1214), .Y(n_1233) );
O2A1O1Ixp33_ASAP7_75t_L g1282 ( .A1(n_1214), .A2(n_1283), .B(n_1284), .C(n_1287), .Y(n_1282) );
NOR2xp33_ASAP7_75t_L g1363 ( .A(n_1214), .B(n_1364), .Y(n_1363) );
INVx2_ASAP7_75t_SL g1214 ( .A(n_1215), .Y(n_1214) );
INVx2_ASAP7_75t_SL g1215 ( .A(n_1216), .Y(n_1215) );
HB1xp67_ASAP7_75t_L g1298 ( .A(n_1216), .Y(n_1298) );
NOR2xp33_ASAP7_75t_L g1321 ( .A(n_1220), .B(n_1322), .Y(n_1321) );
NOR3xp33_ASAP7_75t_L g1329 ( .A(n_1220), .B(n_1255), .C(n_1330), .Y(n_1329) );
INVx1_ASAP7_75t_L g1220 ( .A(n_1221), .Y(n_1220) );
OAI222xp33_ASAP7_75t_L g1256 ( .A1(n_1224), .A2(n_1257), .B1(n_1259), .B2(n_1261), .C1(n_1264), .C2(n_1266), .Y(n_1256) );
NOR2xp33_ASAP7_75t_L g1342 ( .A(n_1224), .B(n_1257), .Y(n_1342) );
OAI22xp5_ASAP7_75t_L g1225 ( .A1(n_1226), .A2(n_1229), .B1(n_1232), .B2(n_1235), .Y(n_1225) );
NOR2x1_ASAP7_75t_L g1226 ( .A(n_1227), .B(n_1228), .Y(n_1226) );
NAND2xp5_ASAP7_75t_L g1364 ( .A(n_1227), .B(n_1365), .Y(n_1364) );
NOR2x1_ASAP7_75t_R g1377 ( .A(n_1227), .B(n_1378), .Y(n_1377) );
OR2x2_ASAP7_75t_L g1382 ( .A(n_1227), .B(n_1242), .Y(n_1382) );
AOI221xp5_ASAP7_75t_L g1274 ( .A1(n_1231), .A2(n_1275), .B1(n_1277), .B2(n_1279), .C(n_1280), .Y(n_1274) );
AND2x2_ASAP7_75t_L g1280 ( .A(n_1231), .B(n_1281), .Y(n_1280) );
A2O1A1Ixp33_ASAP7_75t_L g1337 ( .A1(n_1231), .A2(n_1245), .B(n_1338), .C(n_1341), .Y(n_1337) );
AND2x2_ASAP7_75t_L g1232 ( .A(n_1233), .B(n_1234), .Y(n_1232) );
O2A1O1Ixp33_ASAP7_75t_SL g1293 ( .A1(n_1234), .A2(n_1294), .B(n_1307), .C(n_1316), .Y(n_1293) );
INVxp67_ASAP7_75t_SL g1236 ( .A(n_1237), .Y(n_1236) );
OAI211xp5_ASAP7_75t_L g1269 ( .A1(n_1237), .A2(n_1270), .B(n_1274), .C(n_1282), .Y(n_1269) );
AOI21xp5_ASAP7_75t_L g1237 ( .A1(n_1238), .A2(n_1254), .B(n_1256), .Y(n_1237) );
OAI21xp5_ASAP7_75t_SL g1238 ( .A1(n_1239), .A2(n_1241), .B(n_1243), .Y(n_1238) );
OAI21xp5_ASAP7_75t_SL g1301 ( .A1(n_1241), .A2(n_1302), .B(n_1306), .Y(n_1301) );
OAI21xp33_ASAP7_75t_SL g1317 ( .A1(n_1241), .A2(n_1318), .B(n_1319), .Y(n_1317) );
INVx2_ASAP7_75t_L g1241 ( .A(n_1242), .Y(n_1241) );
NOR2xp33_ASAP7_75t_L g1352 ( .A(n_1242), .B(n_1353), .Y(n_1352) );
CKINVDCx14_ASAP7_75t_R g1243 ( .A(n_1244), .Y(n_1243) );
INVx1_ASAP7_75t_L g1244 ( .A(n_1245), .Y(n_1244) );
NAND2xp5_ASAP7_75t_L g1254 ( .A(n_1245), .B(n_1255), .Y(n_1254) );
CKINVDCx5p33_ASAP7_75t_R g1272 ( .A(n_1245), .Y(n_1272) );
AOI31xp33_ASAP7_75t_L g1316 ( .A1(n_1245), .A2(n_1317), .A3(n_1320), .B(n_1324), .Y(n_1316) );
OR2x6_ASAP7_75t_SL g1245 ( .A(n_1246), .B(n_1250), .Y(n_1245) );
BUFx2_ASAP7_75t_SL g1385 ( .A(n_1253), .Y(n_1385) );
INVx1_ASAP7_75t_L g1344 ( .A(n_1254), .Y(n_1344) );
INVx1_ASAP7_75t_SL g1273 ( .A(n_1255), .Y(n_1273) );
INVx1_ASAP7_75t_L g1332 ( .A(n_1257), .Y(n_1332) );
INVx1_ASAP7_75t_L g1315 ( .A(n_1258), .Y(n_1315) );
INVx1_ASAP7_75t_L g1259 ( .A(n_1260), .Y(n_1259) );
NAND2xp5_ASAP7_75t_L g1313 ( .A(n_1260), .B(n_1314), .Y(n_1313) );
INVx1_ASAP7_75t_L g1281 ( .A(n_1261), .Y(n_1281) );
INVx1_ASAP7_75t_L g1378 ( .A(n_1262), .Y(n_1378) );
INVx1_ASAP7_75t_L g1264 ( .A(n_1265), .Y(n_1264) );
AOI221xp5_ASAP7_75t_L g1324 ( .A1(n_1265), .A2(n_1284), .B1(n_1325), .B2(n_1326), .C(n_1329), .Y(n_1324) );
INVx1_ASAP7_75t_L g1266 ( .A(n_1267), .Y(n_1266) );
AOI21xp5_ASAP7_75t_L g1320 ( .A1(n_1267), .A2(n_1283), .B(n_1321), .Y(n_1320) );
NOR2xp33_ASAP7_75t_L g1336 ( .A(n_1267), .B(n_1298), .Y(n_1336) );
A2O1A1Ixp33_ASAP7_75t_L g1294 ( .A1(n_1268), .A2(n_1295), .B(n_1296), .C(n_1301), .Y(n_1294) );
NAND2xp5_ASAP7_75t_L g1362 ( .A(n_1268), .B(n_1272), .Y(n_1362) );
INVx1_ASAP7_75t_L g1270 ( .A(n_1271), .Y(n_1270) );
NAND2xp5_ASAP7_75t_L g1271 ( .A(n_1272), .B(n_1273), .Y(n_1271) );
OAI21xp33_ASAP7_75t_L g1369 ( .A1(n_1272), .A2(n_1298), .B(n_1370), .Y(n_1369) );
AOI21xp5_ASAP7_75t_L g1376 ( .A1(n_1272), .A2(n_1315), .B(n_1377), .Y(n_1376) );
INVx1_ASAP7_75t_L g1275 ( .A(n_1276), .Y(n_1275) );
INVx1_ASAP7_75t_L g1373 ( .A(n_1277), .Y(n_1373) );
AND2x2_ASAP7_75t_L g1291 ( .A(n_1279), .B(n_1292), .Y(n_1291) );
INVx1_ASAP7_75t_L g1375 ( .A(n_1279), .Y(n_1375) );
INVx1_ASAP7_75t_L g1374 ( .A(n_1284), .Y(n_1374) );
NOR2xp33_ASAP7_75t_L g1350 ( .A(n_1285), .B(n_1309), .Y(n_1350) );
INVx1_ASAP7_75t_L g1285 ( .A(n_1286), .Y(n_1285) );
INVx1_ASAP7_75t_L g1288 ( .A(n_1289), .Y(n_1288) );
INVx1_ASAP7_75t_L g1290 ( .A(n_1291), .Y(n_1290) );
AND2x2_ASAP7_75t_L g1359 ( .A(n_1295), .B(n_1360), .Y(n_1359) );
INVx1_ASAP7_75t_L g1367 ( .A(n_1296), .Y(n_1367) );
OR2x2_ASAP7_75t_L g1296 ( .A(n_1297), .B(n_1299), .Y(n_1296) );
OAI21xp33_ASAP7_75t_L g1354 ( .A1(n_1297), .A2(n_1355), .B(n_1358), .Y(n_1354) );
INVx1_ASAP7_75t_L g1297 ( .A(n_1298), .Y(n_1297) );
INVx1_ASAP7_75t_L g1360 ( .A(n_1298), .Y(n_1360) );
NAND2xp5_ASAP7_75t_L g1356 ( .A(n_1300), .B(n_1357), .Y(n_1356) );
NAND2xp5_ASAP7_75t_L g1380 ( .A(n_1300), .B(n_1381), .Y(n_1380) );
AOI211xp5_ASAP7_75t_L g1331 ( .A1(n_1302), .A2(n_1332), .B(n_1333), .C(n_1342), .Y(n_1331) );
INVx1_ASAP7_75t_L g1302 ( .A(n_1303), .Y(n_1302) );
INVx1_ASAP7_75t_L g1303 ( .A(n_1304), .Y(n_1303) );
INVx1_ASAP7_75t_L g1318 ( .A(n_1308), .Y(n_1318) );
AND2x2_ASAP7_75t_L g1311 ( .A(n_1309), .B(n_1312), .Y(n_1311) );
INVxp67_ASAP7_75t_L g1310 ( .A(n_1311), .Y(n_1310) );
INVx1_ASAP7_75t_L g1322 ( .A(n_1323), .Y(n_1322) );
INVx1_ASAP7_75t_L g1327 ( .A(n_1328), .Y(n_1327) );
INVx1_ASAP7_75t_L g1334 ( .A(n_1335), .Y(n_1334) );
INVx1_ASAP7_75t_L g1338 ( .A(n_1339), .Y(n_1338) );
AOI22xp5_ASAP7_75t_L g1343 ( .A1(n_1344), .A2(n_1345), .B1(n_1361), .B2(n_1363), .Y(n_1343) );
INVx1_ASAP7_75t_L g1368 ( .A(n_1346), .Y(n_1368) );
INVx1_ASAP7_75t_L g1353 ( .A(n_1347), .Y(n_1353) );
AOI21xp5_ASAP7_75t_L g1348 ( .A1(n_1349), .A2(n_1351), .B(n_1352), .Y(n_1348) );
INVx1_ASAP7_75t_L g1349 ( .A(n_1350), .Y(n_1349) );
INVx1_ASAP7_75t_L g1355 ( .A(n_1356), .Y(n_1355) );
INVxp67_ASAP7_75t_SL g1358 ( .A(n_1359), .Y(n_1358) );
INVx1_ASAP7_75t_L g1361 ( .A(n_1362), .Y(n_1361) );
OAI321xp33_ASAP7_75t_L g1366 ( .A1(n_1362), .A2(n_1367), .A3(n_1368), .B1(n_1369), .B2(n_1372), .C(n_1379), .Y(n_1366) );
INVxp33_ASAP7_75t_L g1370 ( .A(n_1371), .Y(n_1370) );
A2O1A1Ixp33_ASAP7_75t_L g1372 ( .A1(n_1373), .A2(n_1374), .B(n_1375), .C(n_1376), .Y(n_1372) );
INVx1_ASAP7_75t_L g1379 ( .A(n_1380), .Y(n_1379) );
INVx1_ASAP7_75t_L g1381 ( .A(n_1382), .Y(n_1381) );
CKINVDCx5p33_ASAP7_75t_R g1383 ( .A(n_1384), .Y(n_1383) );
INVx1_ASAP7_75t_SL g1384 ( .A(n_1385), .Y(n_1384) );
INVx1_ASAP7_75t_L g1386 ( .A(n_1387), .Y(n_1386) );
INVx1_ASAP7_75t_L g1387 ( .A(n_1388), .Y(n_1387) );
HB1xp67_ASAP7_75t_L g1470 ( .A(n_1389), .Y(n_1470) );
AOI222xp33_ASAP7_75t_L g1434 ( .A1(n_1396), .A2(n_1435), .B1(n_1436), .B2(n_1437), .C1(n_1438), .C2(n_1439), .Y(n_1434) );
NAND3xp33_ASAP7_75t_L g1402 ( .A(n_1403), .B(n_1412), .C(n_1434), .Y(n_1402) );
AOI22xp5_ASAP7_75t_L g1403 ( .A1(n_1404), .A2(n_1405), .B1(n_1407), .B2(n_1408), .Y(n_1403) );
INVx2_ASAP7_75t_L g1410 ( .A(n_1406), .Y(n_1410) );
AND2x4_ASAP7_75t_L g1408 ( .A(n_1409), .B(n_1411), .Y(n_1408) );
INVx1_ASAP7_75t_L g1409 ( .A(n_1410), .Y(n_1409) );
NOR3xp33_ASAP7_75t_L g1412 ( .A(n_1413), .B(n_1428), .C(n_1432), .Y(n_1412) );
NAND2x1p5_ASAP7_75t_L g1414 ( .A(n_1415), .B(n_1417), .Y(n_1414) );
INVx2_ASAP7_75t_L g1415 ( .A(n_1416), .Y(n_1415) );
INVx1_ASAP7_75t_L g1417 ( .A(n_1418), .Y(n_1417) );
OR2x6_ASAP7_75t_L g1421 ( .A(n_1418), .B(n_1422), .Y(n_1421) );
INVx1_ASAP7_75t_L g1441 ( .A(n_1418), .Y(n_1441) );
INVx2_ASAP7_75t_L g1418 ( .A(n_1419), .Y(n_1418) );
INVx1_ASAP7_75t_L g1419 ( .A(n_1420), .Y(n_1419) );
NAND2xp5_ASAP7_75t_L g1423 ( .A(n_1424), .B(n_1427), .Y(n_1423) );
INVx2_ASAP7_75t_L g1432 ( .A(n_1433), .Y(n_1432) );
OAI221xp5_ASAP7_75t_SL g1450 ( .A1(n_1435), .A2(n_1437), .B1(n_1451), .B2(n_1453), .C(n_1456), .Y(n_1450) );
INVx1_ASAP7_75t_L g1439 ( .A(n_1440), .Y(n_1439) );
INVx2_ASAP7_75t_L g1442 ( .A(n_1443), .Y(n_1442) );
CKINVDCx8_ASAP7_75t_R g1443 ( .A(n_1444), .Y(n_1443) );
INVx1_ASAP7_75t_L g1451 ( .A(n_1452), .Y(n_1451) );
HB1xp67_ASAP7_75t_L g1453 ( .A(n_1454), .Y(n_1453) );
INVx2_ASAP7_75t_SL g1454 ( .A(n_1455), .Y(n_1454) );
INVx1_ASAP7_75t_SL g1457 ( .A(n_1458), .Y(n_1457) );
INVx1_ASAP7_75t_L g1458 ( .A(n_1459), .Y(n_1458) );
INVx1_ASAP7_75t_L g1459 ( .A(n_1460), .Y(n_1459) );
INVx1_ASAP7_75t_L g1460 ( .A(n_1461), .Y(n_1460) );
INVx1_ASAP7_75t_L g1461 ( .A(n_1462), .Y(n_1461) );
BUFx2_ASAP7_75t_L g1464 ( .A(n_1465), .Y(n_1464) );
OAI21xp5_ASAP7_75t_L g1473 ( .A1(n_1466), .A2(n_1474), .B(n_1475), .Y(n_1473) );
INVxp33_ASAP7_75t_L g1467 ( .A(n_1468), .Y(n_1467) );
INVx1_ASAP7_75t_L g1471 ( .A(n_1470), .Y(n_1471) );
HB1xp67_ASAP7_75t_L g1472 ( .A(n_1473), .Y(n_1472) );
endmodule