module fake_jpeg_20544_n_290 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_290);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_290;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_228;
wire n_178;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_22),
.B(n_8),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_41),
.B(n_22),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_20),
.B(n_0),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_43),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_20),
.B(n_0),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_24),
.A2(n_36),
.B1(n_23),
.B2(n_26),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_47),
.A2(n_26),
.B1(n_21),
.B2(n_32),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_46),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_51),
.B(n_56),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_45),
.A2(n_24),
.B1(n_36),
.B2(n_23),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_52),
.A2(n_54),
.B1(n_57),
.B2(n_60),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_45),
.A2(n_24),
.B1(n_36),
.B2(n_23),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_46),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_41),
.A2(n_21),
.B1(n_34),
.B2(n_19),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_45),
.A2(n_21),
.B1(n_34),
.B2(n_19),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_20),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_71),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_63),
.A2(n_75),
.B1(n_31),
.B2(n_35),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_32),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_65),
.B(n_66),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_39),
.B(n_22),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_43),
.B(n_33),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_43),
.B(n_17),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_73),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_39),
.B(n_29),
.Y(n_74)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_40),
.A2(n_28),
.B1(n_17),
.B2(n_29),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_44),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_76),
.B(n_63),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_49),
.A2(n_40),
.B1(n_44),
.B2(n_47),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_81),
.A2(n_89),
.B1(n_102),
.B2(n_103),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_83),
.B(n_53),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_76),
.A2(n_40),
.B1(n_47),
.B2(n_38),
.Y(n_89)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_91),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_49),
.B(n_33),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_92),
.B(n_95),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_50),
.A2(n_38),
.B1(n_28),
.B2(n_31),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_93),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_71),
.B(n_22),
.Y(n_95)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_59),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_96),
.B(n_98),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_61),
.B(n_22),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_101),
.Y(n_127)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_50),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_69),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_99),
.Y(n_116)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_64),
.Y(n_100)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_100),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_67),
.B(n_22),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_68),
.A2(n_38),
.B1(n_35),
.B2(n_27),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_68),
.B(n_30),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_104),
.B(n_105),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_66),
.B(n_30),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_70),
.A2(n_31),
.B1(n_35),
.B2(n_27),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_106),
.A2(n_107),
.B1(n_112),
.B2(n_51),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_70),
.A2(n_35),
.B1(n_27),
.B2(n_25),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_55),
.Y(n_108)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_108),
.Y(n_126)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_69),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_109),
.B(n_110),
.Y(n_124)
);

INVx13_ASAP7_75t_L g110 ( 
.A(n_62),
.Y(n_110)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_69),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_58),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_66),
.A2(n_30),
.B1(n_18),
.B2(n_25),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_117),
.A2(n_121),
.B1(n_81),
.B2(n_112),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_77),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_118),
.B(n_120),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_91),
.Y(n_120)
);

O2A1O1Ixp33_ASAP7_75t_L g121 ( 
.A1(n_83),
.A2(n_56),
.B(n_72),
.C(n_55),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_122),
.B(n_132),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_94),
.B(n_53),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_123),
.A2(n_108),
.B(n_79),
.Y(n_152)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_100),
.Y(n_128)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_128),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_88),
.A2(n_72),
.B1(n_25),
.B2(n_27),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_130),
.A2(n_82),
.B1(n_48),
.B2(n_87),
.Y(n_162)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_104),
.Y(n_131)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_131),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_78),
.B(n_53),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_78),
.B(n_58),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_133),
.B(n_138),
.Y(n_153)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_80),
.Y(n_134)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_134),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_135),
.Y(n_146)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_80),
.Y(n_137)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_137),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_92),
.B(n_58),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_97),
.B(n_10),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_139),
.B(n_90),
.Y(n_156)
);

A2O1A1Ixp33_ASAP7_75t_L g140 ( 
.A1(n_85),
.A2(n_25),
.B(n_48),
.C(n_30),
.Y(n_140)
);

OAI31xp33_ASAP7_75t_SL g159 ( 
.A1(n_140),
.A2(n_48),
.A3(n_59),
.B(n_110),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_116),
.Y(n_142)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_142),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_143),
.A2(n_147),
.B1(n_157),
.B2(n_164),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_118),
.B(n_90),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_144),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_119),
.B(n_95),
.C(n_105),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_145),
.B(n_139),
.C(n_129),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_117),
.A2(n_85),
.B1(n_101),
.B2(n_79),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_122),
.B(n_48),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_149),
.A2(n_165),
.B(n_140),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_125),
.A2(n_84),
.B1(n_96),
.B2(n_86),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_150),
.A2(n_162),
.B1(n_166),
.B2(n_114),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_152),
.B(n_156),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_136),
.A2(n_98),
.B1(n_86),
.B2(n_99),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_127),
.B(n_13),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_158),
.B(n_168),
.Y(n_185)
);

O2A1O1Ixp33_ASAP7_75t_L g180 ( 
.A1(n_159),
.A2(n_167),
.B(n_114),
.C(n_115),
.Y(n_180)
);

OA22x2_ASAP7_75t_L g160 ( 
.A1(n_131),
.A2(n_109),
.B1(n_84),
.B2(n_111),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_160),
.B(n_161),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_123),
.A2(n_9),
.B1(n_16),
.B2(n_15),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_133),
.B(n_138),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_163),
.B(n_170),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_136),
.A2(n_8),
.B1(n_15),
.B2(n_14),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_140),
.A2(n_0),
.B(n_1),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_132),
.A2(n_82),
.B1(n_87),
.B2(n_3),
.Y(n_166)
);

A2O1A1Ixp33_ASAP7_75t_SL g167 ( 
.A1(n_120),
.A2(n_82),
.B(n_2),
.C(n_3),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_127),
.B(n_6),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_124),
.B(n_6),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_171),
.A2(n_175),
.B1(n_189),
.B2(n_196),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_172),
.B(n_184),
.C(n_192),
.Y(n_204)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_155),
.Y(n_174)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_174),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_164),
.A2(n_129),
.B1(n_115),
.B2(n_128),
.Y(n_175)
);

INVx13_ASAP7_75t_L g176 ( 
.A(n_142),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_176),
.B(n_183),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_177),
.A2(n_180),
.B(n_165),
.Y(n_209)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_155),
.Y(n_181)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_181),
.Y(n_206)
);

AND2x6_ASAP7_75t_L g183 ( 
.A(n_147),
.B(n_121),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_145),
.B(n_119),
.C(n_123),
.Y(n_184)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_169),
.Y(n_186)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_186),
.Y(n_211)
);

CKINVDCx12_ASAP7_75t_R g187 ( 
.A(n_146),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_187),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_143),
.A2(n_121),
.B1(n_113),
.B2(n_134),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_169),
.Y(n_190)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_190),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_148),
.B(n_137),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_191),
.B(n_194),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_153),
.B(n_126),
.C(n_113),
.Y(n_192)
);

OR2x2_ASAP7_75t_L g194 ( 
.A(n_151),
.B(n_124),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_141),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_195),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_157),
.A2(n_126),
.B1(n_135),
.B2(n_116),
.Y(n_196)
);

INVx13_ASAP7_75t_L g197 ( 
.A(n_167),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_197),
.B(n_160),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_174),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_202),
.B(n_207),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_182),
.B(n_153),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_203),
.B(n_215),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_181),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_209),
.A2(n_1),
.B(n_2),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_191),
.B(n_148),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_210),
.B(n_212),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_183),
.A2(n_154),
.B1(n_159),
.B2(n_141),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_213),
.A2(n_179),
.B1(n_166),
.B2(n_149),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_188),
.B(n_160),
.Y(n_214)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_214),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_184),
.B(n_152),
.C(n_156),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_194),
.B(n_160),
.Y(n_216)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_216),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_193),
.A2(n_180),
.B1(n_196),
.B2(n_179),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_217),
.A2(n_177),
.B1(n_193),
.B2(n_192),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_186),
.Y(n_218)
);

AOI21xp33_ASAP7_75t_L g226 ( 
.A1(n_218),
.A2(n_195),
.B(n_154),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_190),
.Y(n_220)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_220),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_222),
.A2(n_231),
.B1(n_234),
.B2(n_219),
.Y(n_245)
);

AO22x1_ASAP7_75t_L g223 ( 
.A1(n_199),
.A2(n_197),
.B1(n_179),
.B2(n_167),
.Y(n_223)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_223),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_224),
.A2(n_225),
.B1(n_227),
.B2(n_210),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_199),
.B(n_185),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_226),
.A2(n_238),
.B(n_209),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_203),
.B(n_185),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_215),
.B(n_182),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_228),
.B(n_204),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_213),
.A2(n_149),
.B1(n_178),
.B2(n_173),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_230),
.A2(n_206),
.B1(n_200),
.B2(n_220),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_217),
.A2(n_178),
.B1(n_172),
.B2(n_161),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_201),
.A2(n_173),
.B1(n_167),
.B2(n_176),
.Y(n_234)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_205),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_236),
.B(n_207),
.Y(n_241)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_239),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_241),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_235),
.A2(n_208),
.B1(n_201),
.B2(n_218),
.Y(n_242)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_242),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_221),
.A2(n_202),
.B(n_205),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_243),
.B(n_247),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_244),
.B(n_245),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_246),
.B(n_250),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_221),
.A2(n_219),
.B(n_211),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_229),
.B(n_211),
.Y(n_248)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_248),
.Y(n_259)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_237),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_249),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_229),
.B(n_206),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_251),
.B(n_252),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_228),
.B(n_204),
.Y(n_252)
);

A2O1A1Ixp33_ASAP7_75t_SL g260 ( 
.A1(n_242),
.A2(n_224),
.B(n_230),
.C(n_223),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_260),
.A2(n_240),
.B1(n_245),
.B2(n_232),
.Y(n_265)
);

BUFx24_ASAP7_75t_SL g262 ( 
.A(n_246),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_262),
.B(n_198),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_264),
.B(n_268),
.Y(n_275)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_265),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_259),
.B(n_251),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_266),
.B(n_267),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_261),
.B(n_252),
.C(n_233),
.Y(n_267)
);

OAI322xp33_ASAP7_75t_L g268 ( 
.A1(n_254),
.A2(n_239),
.A3(n_260),
.B1(n_231),
.B2(n_258),
.C1(n_233),
.C2(n_240),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_263),
.B(n_248),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_269),
.B(n_270),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_257),
.B(n_236),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_253),
.B(n_247),
.C(n_243),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_271),
.B(n_250),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_271),
.A2(n_241),
.B(n_255),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_276),
.B(n_277),
.Y(n_278)
);

AOI322xp5_ASAP7_75t_L g279 ( 
.A1(n_277),
.A2(n_272),
.A3(n_249),
.B1(n_275),
.B2(n_200),
.C1(n_260),
.C2(n_274),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_279),
.A2(n_280),
.B1(n_281),
.B2(n_223),
.Y(n_283)
);

AOI322xp5_ASAP7_75t_L g280 ( 
.A1(n_273),
.A2(n_265),
.A3(n_270),
.B1(n_256),
.B2(n_198),
.C1(n_222),
.C2(n_234),
.Y(n_280)
);

OAI21x1_ASAP7_75t_L g281 ( 
.A1(n_273),
.A2(n_238),
.B(n_267),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_278),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_282),
.A2(n_7),
.B(n_10),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_283),
.B(n_284),
.C(n_5),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_278),
.B(n_116),
.Y(n_284)
);

AOI321xp33_ASAP7_75t_SL g287 ( 
.A1(n_285),
.A2(n_286),
.A3(n_5),
.B1(n_10),
.B2(n_9),
.C(n_4),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_287),
.A2(n_4),
.B1(n_8),
.B2(n_9),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_288),
.B(n_12),
.C(n_2),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_289),
.B(n_1),
.Y(n_290)
);


endmodule