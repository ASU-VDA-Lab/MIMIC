module fake_netlist_5_529_n_1623 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1623);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1623;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_155;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_156;
wire n_1078;
wire n_775;
wire n_219;
wire n_157;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_675;
wire n_888;
wire n_1167;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_887;
wire n_154;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1293;
wire n_965;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_284;
wire n_1128;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_254;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_433;
wire n_368;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1534;
wire n_560;
wire n_1354;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_233;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_562;
wire n_1436;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_153;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_833;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1419;
wire n_338;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_253;
wire n_1116;
wire n_1212;
wire n_1541;
wire n_172;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1514;
wire n_1335;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_768;
wire n_1475;
wire n_1302;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_685;
wire n_598;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_462;
wire n_1193;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1245;
wire n_846;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1540;
wire n_229;
wire n_437;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_45),
.Y(n_153)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_50),
.Y(n_154)
);

BUFx5_ASAP7_75t_L g155 ( 
.A(n_86),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_2),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_17),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_43),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_143),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_126),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_74),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_52),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_110),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_29),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_136),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_51),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_43),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_7),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_139),
.Y(n_169)
);

INVx2_ASAP7_75t_SL g170 ( 
.A(n_12),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_140),
.Y(n_171)
);

INVx2_ASAP7_75t_SL g172 ( 
.A(n_36),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_56),
.Y(n_173)
);

INVx2_ASAP7_75t_SL g174 ( 
.A(n_70),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_87),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_117),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_48),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_76),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_98),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_39),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_6),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_85),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_92),
.Y(n_183)
);

BUFx5_ASAP7_75t_L g184 ( 
.A(n_63),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_93),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_46),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_45),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_40),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_19),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_23),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_23),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_90),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_7),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_148),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_147),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_65),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_78),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_3),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_18),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_68),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_35),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_53),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_12),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_122),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_62),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_120),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_88),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_75),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_26),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_19),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_2),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_102),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_72),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_100),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_13),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_118),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_97),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_14),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_3),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_79),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_115),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_1),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_14),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_33),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_35),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_135),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_108),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_113),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_61),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_54),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_64),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_125),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_142),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_77),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_121),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_8),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_39),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_131),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_18),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_21),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_38),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_116),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_80),
.Y(n_243)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_99),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_11),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_144),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_55),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_58),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_89),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_47),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_30),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_109),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_25),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_6),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_5),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_73),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_29),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_152),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_101),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_27),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_81),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_5),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_49),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_51),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_137),
.Y(n_265)
);

BUFx8_ASAP7_75t_SL g266 ( 
.A(n_130),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_42),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_42),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_123),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_71),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_37),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_59),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_151),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_138),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_40),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_60),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_38),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_119),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_49),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_16),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_34),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_150),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_44),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_28),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_0),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_141),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_82),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_67),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_105),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_145),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g291 ( 
.A(n_32),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_33),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_114),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_28),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_4),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_83),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_95),
.Y(n_297)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_36),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_9),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_127),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_20),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_298),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_271),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_178),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_298),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_291),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_298),
.Y(n_307)
);

NOR2xp67_ASAP7_75t_L g308 ( 
.A(n_170),
.B(n_0),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_167),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_156),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_167),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_186),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_187),
.Y(n_313)
);

NOR2xp67_ASAP7_75t_L g314 ( 
.A(n_170),
.B(n_1),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_182),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_177),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_183),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_214),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_297),
.B(n_4),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_256),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_199),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_190),
.Y(n_322)
);

INVxp33_ASAP7_75t_SL g323 ( 
.A(n_157),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_191),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_174),
.B(n_8),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_266),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_238),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_177),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_174),
.B(n_9),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_203),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_224),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_209),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_224),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_279),
.Y(n_334)
);

HB1xp67_ASAP7_75t_L g335 ( 
.A(n_157),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_279),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_242),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_210),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_164),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_166),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_168),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_188),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_193),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_218),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_185),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_222),
.Y(n_346)
);

CKINVDCx16_ASAP7_75t_R g347 ( 
.A(n_153),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_192),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_223),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_176),
.B(n_10),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_194),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_225),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_198),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_211),
.Y(n_354)
);

INVxp67_ASAP7_75t_SL g355 ( 
.A(n_244),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_236),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_219),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_239),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_245),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_237),
.Y(n_360)
);

OR2x2_ASAP7_75t_L g361 ( 
.A(n_250),
.B(n_10),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_254),
.Y(n_362)
);

INVxp33_ASAP7_75t_SL g363 ( 
.A(n_162),
.Y(n_363)
);

BUFx6f_ASAP7_75t_SL g364 ( 
.A(n_244),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_240),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_275),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_199),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_241),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_155),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_253),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_251),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_255),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_305),
.B(n_176),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_337),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_321),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_337),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_308),
.B(n_172),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_307),
.B(n_197),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_321),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_367),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_367),
.Y(n_381)
);

NAND3xp33_ASAP7_75t_L g382 ( 
.A(n_329),
.B(n_172),
.C(n_253),
.Y(n_382)
);

AND2x4_ASAP7_75t_L g383 ( 
.A(n_302),
.B(n_197),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_370),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_370),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_337),
.Y(n_386)
);

AND2x2_ASAP7_75t_SL g387 ( 
.A(n_350),
.B(n_269),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_337),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_337),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_355),
.B(n_159),
.Y(n_390)
);

NAND2xp33_ASAP7_75t_L g391 ( 
.A(n_325),
.B(n_267),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_319),
.B(n_195),
.Y(n_392)
);

CKINVDCx8_ASAP7_75t_R g393 ( 
.A(n_347),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_369),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_302),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_369),
.Y(n_396)
);

AND2x4_ASAP7_75t_L g397 ( 
.A(n_309),
.B(n_269),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_339),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_340),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_341),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_342),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_343),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_353),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_354),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_357),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_311),
.B(n_267),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_358),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_359),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_335),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_362),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_316),
.B(n_159),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_366),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_328),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_331),
.Y(n_414)
);

INVx3_ASAP7_75t_L g415 ( 
.A(n_361),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_361),
.A2(n_180),
.B1(n_294),
.B2(n_215),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_333),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_334),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_336),
.B(n_160),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_310),
.Y(n_420)
);

CKINVDCx6p67_ASAP7_75t_R g421 ( 
.A(n_326),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_314),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_364),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_364),
.Y(n_424)
);

BUFx3_ASAP7_75t_L g425 ( 
.A(n_345),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_364),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_306),
.B(n_165),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_312),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_312),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_313),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_313),
.Y(n_431)
);

INVx1_ASAP7_75t_SL g432 ( 
.A(n_322),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_322),
.B(n_169),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_324),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_324),
.B(n_160),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_330),
.Y(n_436)
);

HB1xp67_ASAP7_75t_L g437 ( 
.A(n_330),
.Y(n_437)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_394),
.Y(n_438)
);

BUFx10_ASAP7_75t_L g439 ( 
.A(n_392),
.Y(n_439)
);

INVx1_ASAP7_75t_SL g440 ( 
.A(n_432),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_415),
.B(n_332),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_394),
.Y(n_442)
);

AOI22xp33_ASAP7_75t_L g443 ( 
.A1(n_387),
.A2(n_363),
.B1(n_323),
.B2(n_277),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_394),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_417),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_417),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_374),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_394),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_394),
.Y(n_449)
);

NAND3xp33_ASAP7_75t_L g450 ( 
.A(n_392),
.B(n_338),
.C(n_332),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_417),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_435),
.B(n_348),
.Y(n_452)
);

INVx3_ASAP7_75t_L g453 ( 
.A(n_394),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_417),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_394),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_415),
.B(n_338),
.Y(n_456)
);

INVx3_ASAP7_75t_L g457 ( 
.A(n_394),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_396),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_435),
.B(n_351),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_428),
.B(n_430),
.Y(n_460)
);

AND2x2_ASAP7_75t_SL g461 ( 
.A(n_387),
.B(n_242),
.Y(n_461)
);

OR2x2_ASAP7_75t_L g462 ( 
.A(n_415),
.B(n_303),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_396),
.Y(n_463)
);

NAND2xp33_ASAP7_75t_L g464 ( 
.A(n_436),
.B(n_344),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_395),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g466 ( 
.A(n_415),
.B(n_344),
.Y(n_466)
);

BUFx3_ASAP7_75t_L g467 ( 
.A(n_413),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_415),
.B(n_346),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_396),
.Y(n_469)
);

HB1xp67_ASAP7_75t_L g470 ( 
.A(n_409),
.Y(n_470)
);

INVx2_ASAP7_75t_SL g471 ( 
.A(n_433),
.Y(n_471)
);

BUFx2_ASAP7_75t_L g472 ( 
.A(n_409),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_396),
.Y(n_473)
);

BUFx4f_ASAP7_75t_L g474 ( 
.A(n_387),
.Y(n_474)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_390),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_395),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_396),
.Y(n_477)
);

NOR2x1p5_ASAP7_75t_L g478 ( 
.A(n_423),
.B(n_162),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_396),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_416),
.A2(n_201),
.B1(n_189),
.B2(n_158),
.Y(n_480)
);

INVx3_ASAP7_75t_L g481 ( 
.A(n_396),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_396),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_373),
.B(n_346),
.Y(n_483)
);

INVxp67_ASAP7_75t_L g484 ( 
.A(n_437),
.Y(n_484)
);

BUFx3_ASAP7_75t_L g485 ( 
.A(n_413),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_374),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_436),
.B(n_349),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_414),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_374),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_390),
.B(n_349),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_398),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_422),
.B(n_352),
.Y(n_492)
);

NOR2x1p5_ASAP7_75t_L g493 ( 
.A(n_423),
.B(n_181),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_374),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_428),
.B(n_352),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_436),
.B(n_356),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_422),
.B(n_356),
.Y(n_497)
);

INVx5_ASAP7_75t_L g498 ( 
.A(n_374),
.Y(n_498)
);

BUFx2_ASAP7_75t_L g499 ( 
.A(n_437),
.Y(n_499)
);

BUFx6f_ASAP7_75t_L g500 ( 
.A(n_374),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_398),
.Y(n_501)
);

BUFx2_ASAP7_75t_L g502 ( 
.A(n_429),
.Y(n_502)
);

NAND3xp33_ASAP7_75t_L g503 ( 
.A(n_391),
.B(n_365),
.C(n_360),
.Y(n_503)
);

BUFx10_ASAP7_75t_L g504 ( 
.A(n_436),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_436),
.B(n_360),
.Y(n_505)
);

OR2x6_ASAP7_75t_L g506 ( 
.A(n_429),
.B(n_436),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_L g507 ( 
.A1(n_429),
.A2(n_327),
.B1(n_371),
.B2(n_368),
.Y(n_507)
);

AOI22xp33_ASAP7_75t_L g508 ( 
.A1(n_391),
.A2(n_382),
.B1(n_427),
.B2(n_397),
.Y(n_508)
);

OAI21xp33_ASAP7_75t_SL g509 ( 
.A1(n_377),
.A2(n_154),
.B(n_196),
.Y(n_509)
);

AOI22xp33_ASAP7_75t_L g510 ( 
.A1(n_382),
.A2(n_242),
.B1(n_248),
.B2(n_289),
.Y(n_510)
);

INVx2_ASAP7_75t_SL g511 ( 
.A(n_433),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_433),
.B(n_365),
.Y(n_512)
);

BUFx3_ASAP7_75t_L g513 ( 
.A(n_418),
.Y(n_513)
);

BUFx6f_ASAP7_75t_SL g514 ( 
.A(n_430),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_436),
.B(n_368),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_376),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_376),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_376),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_376),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_373),
.B(n_371),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_373),
.B(n_372),
.Y(n_521)
);

BUFx3_ASAP7_75t_L g522 ( 
.A(n_418),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_378),
.B(n_372),
.Y(n_523)
);

INVx4_ASAP7_75t_L g524 ( 
.A(n_374),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_388),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_398),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_378),
.B(n_270),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_398),
.Y(n_528)
);

AND2x6_ASAP7_75t_L g529 ( 
.A(n_424),
.B(n_242),
.Y(n_529)
);

AOI22xp33_ASAP7_75t_L g530 ( 
.A1(n_427),
.A2(n_397),
.B1(n_383),
.B2(n_377),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_374),
.Y(n_531)
);

OR2x2_ASAP7_75t_L g532 ( 
.A(n_416),
.B(n_257),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_429),
.B(n_411),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_386),
.Y(n_534)
);

AND2x4_ASAP7_75t_L g535 ( 
.A(n_397),
.B(n_212),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_431),
.B(n_320),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_386),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_388),
.Y(n_538)
);

AND2x6_ASAP7_75t_L g539 ( 
.A(n_424),
.B(n_242),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_401),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_401),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_431),
.B(n_318),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_388),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_401),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_411),
.B(n_200),
.Y(n_545)
);

BUFx6f_ASAP7_75t_SL g546 ( 
.A(n_434),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_402),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_402),
.Y(n_548)
);

INVx3_ASAP7_75t_L g549 ( 
.A(n_386),
.Y(n_549)
);

AOI22xp5_ASAP7_75t_L g550 ( 
.A1(n_434),
.A2(n_181),
.B1(n_281),
.B2(n_283),
.Y(n_550)
);

BUFx3_ASAP7_75t_L g551 ( 
.A(n_399),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_386),
.Y(n_552)
);

AOI21x1_ASAP7_75t_L g553 ( 
.A1(n_383),
.A2(n_233),
.B(n_261),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_419),
.B(n_202),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_386),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_386),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_386),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_386),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_419),
.B(n_204),
.Y(n_559)
);

INVx3_ASAP7_75t_L g560 ( 
.A(n_389),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_397),
.B(n_205),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_389),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_436),
.B(n_317),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_421),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_397),
.B(n_206),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_389),
.Y(n_566)
);

NOR2x1p5_ASAP7_75t_L g567 ( 
.A(n_426),
.B(n_264),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_389),
.Y(n_568)
);

INVxp67_ASAP7_75t_SL g569 ( 
.A(n_389),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_389),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_389),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_432),
.B(n_315),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_402),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_402),
.Y(n_574)
);

INVx4_ASAP7_75t_L g575 ( 
.A(n_389),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_404),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_404),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_404),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_404),
.Y(n_579)
);

NOR3xp33_ASAP7_75t_L g580 ( 
.A(n_507),
.B(n_450),
.C(n_503),
.Y(n_580)
);

INVxp67_ASAP7_75t_L g581 ( 
.A(n_472),
.Y(n_581)
);

INVx8_ASAP7_75t_L g582 ( 
.A(n_514),
.Y(n_582)
);

AOI22xp5_ASAP7_75t_L g583 ( 
.A1(n_471),
.A2(n_304),
.B1(n_427),
.B2(n_426),
.Y(n_583)
);

OR2x2_ASAP7_75t_L g584 ( 
.A(n_462),
.B(n_425),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_533),
.B(n_404),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_475),
.B(n_420),
.Y(n_586)
);

AOI22xp33_ASAP7_75t_L g587 ( 
.A1(n_461),
.A2(n_383),
.B1(n_406),
.B2(n_289),
.Y(n_587)
);

HB1xp67_ASAP7_75t_L g588 ( 
.A(n_502),
.Y(n_588)
);

INVxp67_ASAP7_75t_L g589 ( 
.A(n_472),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_461),
.B(n_404),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_474),
.B(n_461),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_502),
.B(n_404),
.Y(n_592)
);

BUFx6f_ASAP7_75t_L g593 ( 
.A(n_551),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_441),
.B(n_404),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_441),
.B(n_456),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_551),
.Y(n_596)
);

AOI22xp5_ASAP7_75t_L g597 ( 
.A1(n_471),
.A2(n_258),
.B1(n_259),
.B2(n_213),
.Y(n_597)
);

NAND3xp33_ASAP7_75t_L g598 ( 
.A(n_443),
.B(n_420),
.C(n_399),
.Y(n_598)
);

AOI21xp5_ASAP7_75t_L g599 ( 
.A1(n_569),
.A2(n_383),
.B(n_405),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_456),
.B(n_466),
.Y(n_600)
);

BUFx6f_ASAP7_75t_SL g601 ( 
.A(n_439),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_474),
.B(n_248),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_474),
.B(n_248),
.Y(n_603)
);

NAND2x1p5_ASAP7_75t_L g604 ( 
.A(n_474),
.B(n_216),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_466),
.B(n_383),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_488),
.Y(n_606)
);

O2A1O1Ixp5_ASAP7_75t_L g607 ( 
.A1(n_468),
.A2(n_274),
.B(n_276),
.C(n_287),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_440),
.B(n_425),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_511),
.B(n_248),
.Y(n_609)
);

NOR3xp33_ASAP7_75t_SL g610 ( 
.A(n_509),
.B(n_299),
.C(n_280),
.Y(n_610)
);

INVx2_ASAP7_75t_SL g611 ( 
.A(n_462),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_511),
.B(n_248),
.Y(n_612)
);

INVx4_ASAP7_75t_L g613 ( 
.A(n_551),
.Y(n_613)
);

AOI22xp33_ASAP7_75t_L g614 ( 
.A1(n_510),
.A2(n_506),
.B1(n_439),
.B2(n_476),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_460),
.B(n_400),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_439),
.B(n_393),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_504),
.B(n_289),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_490),
.B(n_226),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_545),
.B(n_249),
.Y(n_619)
);

INVx2_ASAP7_75t_SL g620 ( 
.A(n_483),
.Y(n_620)
);

OAI22xp5_ASAP7_75t_L g621 ( 
.A1(n_506),
.A2(n_288),
.B1(n_300),
.B2(n_171),
.Y(n_621)
);

NOR2xp67_ASAP7_75t_L g622 ( 
.A(n_484),
.B(n_425),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_554),
.B(n_406),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_559),
.B(n_406),
.Y(n_624)
);

INVx2_ASAP7_75t_SL g625 ( 
.A(n_483),
.Y(n_625)
);

NAND2x1_ASAP7_75t_L g626 ( 
.A(n_506),
.B(n_289),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_465),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_530),
.B(n_405),
.Y(n_628)
);

AOI22xp33_ASAP7_75t_L g629 ( 
.A1(n_506),
.A2(n_439),
.B1(n_476),
.B2(n_465),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_470),
.B(n_425),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_508),
.B(n_405),
.Y(n_631)
);

INVx2_ASAP7_75t_SL g632 ( 
.A(n_499),
.Y(n_632)
);

AO22x2_ASAP7_75t_L g633 ( 
.A1(n_532),
.A2(n_407),
.B1(n_410),
.B2(n_403),
.Y(n_633)
);

INVxp67_ASAP7_75t_SL g634 ( 
.A(n_438),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_492),
.B(n_400),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_467),
.B(n_408),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_485),
.B(n_408),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_485),
.Y(n_638)
);

AOI22xp33_ASAP7_75t_L g639 ( 
.A1(n_506),
.A2(n_289),
.B1(n_184),
.B2(n_155),
.Y(n_639)
);

AOI22xp5_ASAP7_75t_L g640 ( 
.A1(n_452),
.A2(n_221),
.B1(n_232),
.B2(n_234),
.Y(n_640)
);

CKINVDCx11_ASAP7_75t_R g641 ( 
.A(n_499),
.Y(n_641)
);

AOI21xp5_ASAP7_75t_L g642 ( 
.A1(n_561),
.A2(n_408),
.B(n_412),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_485),
.B(n_375),
.Y(n_643)
);

INVx3_ASAP7_75t_L g644 ( 
.A(n_513),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_513),
.B(n_375),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_504),
.B(n_155),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_445),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_513),
.Y(n_648)
);

HB1xp67_ASAP7_75t_L g649 ( 
.A(n_520),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_522),
.B(n_379),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_504),
.B(n_155),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_522),
.B(n_527),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_495),
.B(n_393),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_512),
.B(n_393),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_497),
.B(n_161),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_521),
.B(n_161),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_522),
.B(n_379),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_504),
.B(n_155),
.Y(n_658)
);

AND2x4_ASAP7_75t_L g659 ( 
.A(n_535),
.B(n_380),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_535),
.B(n_380),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_445),
.Y(n_661)
);

INVx8_ASAP7_75t_L g662 ( 
.A(n_514),
.Y(n_662)
);

AOI22xp5_ASAP7_75t_L g663 ( 
.A1(n_459),
.A2(n_207),
.B1(n_208),
.B2(n_217),
.Y(n_663)
);

BUFx3_ASAP7_75t_L g664 ( 
.A(n_535),
.Y(n_664)
);

AND2x4_ASAP7_75t_L g665 ( 
.A(n_535),
.B(n_381),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_523),
.B(n_155),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_565),
.B(n_381),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_438),
.B(n_384),
.Y(n_668)
);

AOI22xp5_ASAP7_75t_L g669 ( 
.A1(n_464),
.A2(n_220),
.B1(n_227),
.B2(n_228),
.Y(n_669)
);

NAND3xp33_ASAP7_75t_L g670 ( 
.A(n_480),
.B(n_260),
.C(n_262),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_446),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_487),
.B(n_155),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_438),
.B(n_385),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_453),
.B(n_385),
.Y(n_674)
);

NOR2xp67_ASAP7_75t_L g675 ( 
.A(n_563),
.B(n_230),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_453),
.B(n_231),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_446),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_453),
.B(n_235),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_453),
.B(n_243),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_496),
.B(n_155),
.Y(n_680)
);

CKINVDCx11_ASAP7_75t_R g681 ( 
.A(n_564),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_505),
.B(n_163),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_515),
.B(n_184),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_457),
.B(n_246),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_457),
.B(n_247),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_572),
.B(n_421),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_457),
.B(n_252),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_451),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_514),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_509),
.B(n_163),
.Y(n_690)
);

BUFx5_ASAP7_75t_L g691 ( 
.A(n_576),
.Y(n_691)
);

INVxp33_ASAP7_75t_L g692 ( 
.A(n_532),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_454),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_457),
.B(n_171),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_550),
.B(n_173),
.Y(n_695)
);

AND2x6_ASAP7_75t_SL g696 ( 
.A(n_536),
.B(n_264),
.Y(n_696)
);

INVx4_ASAP7_75t_L g697 ( 
.A(n_447),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_481),
.B(n_173),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_491),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_542),
.B(n_421),
.Y(n_700)
);

NOR2xp67_ASAP7_75t_L g701 ( 
.A(n_550),
.B(n_175),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_481),
.B(n_175),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_481),
.B(n_179),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_444),
.B(n_184),
.Y(n_704)
);

NAND2xp33_ASAP7_75t_L g705 ( 
.A(n_529),
.B(n_184),
.Y(n_705)
);

HB1xp67_ASAP7_75t_L g706 ( 
.A(n_478),
.Y(n_706)
);

NOR2xp67_ASAP7_75t_L g707 ( 
.A(n_480),
.B(n_179),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_501),
.Y(n_708)
);

O2A1O1Ixp33_ASAP7_75t_L g709 ( 
.A1(n_501),
.A2(n_282),
.B(n_272),
.C(n_296),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_526),
.Y(n_710)
);

A2O1A1Ixp33_ASAP7_75t_L g711 ( 
.A1(n_526),
.A2(n_282),
.B(n_229),
.C(n_296),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_444),
.B(n_184),
.Y(n_712)
);

BUFx10_ASAP7_75t_L g713 ( 
.A(n_478),
.Y(n_713)
);

AND2x4_ASAP7_75t_L g714 ( 
.A(n_493),
.B(n_229),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_528),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_444),
.B(n_184),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_514),
.B(n_265),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_463),
.B(n_272),
.Y(n_718)
);

AOI21xp5_ASAP7_75t_L g719 ( 
.A1(n_442),
.A2(n_273),
.B(n_286),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_463),
.B(n_184),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_481),
.B(n_265),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_546),
.B(n_273),
.Y(n_722)
);

NAND2x1p5_ASAP7_75t_L g723 ( 
.A(n_493),
.B(n_103),
.Y(n_723)
);

NOR2xp67_ASAP7_75t_L g724 ( 
.A(n_540),
.B(n_278),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_463),
.B(n_184),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_469),
.B(n_278),
.Y(n_726)
);

AND2x6_ASAP7_75t_SL g727 ( 
.A(n_546),
.B(n_268),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_540),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_541),
.Y(n_729)
);

BUFx6f_ASAP7_75t_L g730 ( 
.A(n_447),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_541),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_SL g732 ( 
.A(n_546),
.B(n_286),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_544),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_442),
.B(n_290),
.Y(n_734)
);

BUFx6f_ASAP7_75t_L g735 ( 
.A(n_447),
.Y(n_735)
);

AOI21xp5_ASAP7_75t_L g736 ( 
.A1(n_594),
.A2(n_524),
.B(n_575),
.Y(n_736)
);

BUFx2_ASAP7_75t_L g737 ( 
.A(n_608),
.Y(n_737)
);

AOI21xp5_ASAP7_75t_L g738 ( 
.A1(n_585),
.A2(n_524),
.B(n_575),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_649),
.B(n_546),
.Y(n_739)
);

AOI21xp5_ASAP7_75t_L g740 ( 
.A1(n_605),
.A2(n_524),
.B(n_575),
.Y(n_740)
);

NAND2x1p5_ASAP7_75t_L g741 ( 
.A(n_613),
.B(n_644),
.Y(n_741)
);

O2A1O1Ixp33_ASAP7_75t_L g742 ( 
.A1(n_595),
.A2(n_574),
.B(n_548),
.C(n_544),
.Y(n_742)
);

INVxp67_ASAP7_75t_L g743 ( 
.A(n_586),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_600),
.B(n_448),
.Y(n_744)
);

BUFx2_ASAP7_75t_L g745 ( 
.A(n_632),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_629),
.B(n_448),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_649),
.B(n_547),
.Y(n_747)
);

O2A1O1Ixp5_ASAP7_75t_L g748 ( 
.A1(n_602),
.A2(n_603),
.B(n_666),
.C(n_672),
.Y(n_748)
);

OAI21xp5_ASAP7_75t_L g749 ( 
.A1(n_590),
.A2(n_458),
.B(n_449),
.Y(n_749)
);

AOI21xp5_ASAP7_75t_L g750 ( 
.A1(n_592),
.A2(n_524),
.B(n_575),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_629),
.B(n_449),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_627),
.Y(n_752)
);

AOI21xp5_ASAP7_75t_L g753 ( 
.A1(n_628),
.A2(n_455),
.B(n_458),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_588),
.B(n_547),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_615),
.B(n_455),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_580),
.B(n_473),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_588),
.B(n_548),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_692),
.B(n_573),
.Y(n_758)
);

AOI21xp5_ASAP7_75t_L g759 ( 
.A1(n_697),
.A2(n_473),
.B(n_477),
.Y(n_759)
);

AOI21xp5_ASAP7_75t_L g760 ( 
.A1(n_697),
.A2(n_482),
.B(n_479),
.Y(n_760)
);

O2A1O1Ixp33_ASAP7_75t_L g761 ( 
.A1(n_631),
.A2(n_573),
.B(n_574),
.C(n_567),
.Y(n_761)
);

AOI21xp5_ASAP7_75t_L g762 ( 
.A1(n_652),
.A2(n_482),
.B(n_479),
.Y(n_762)
);

NOR2x1p5_ASAP7_75t_L g763 ( 
.A(n_689),
.B(n_268),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_586),
.B(n_567),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_593),
.B(n_477),
.Y(n_765)
);

AOI21x1_ASAP7_75t_L g766 ( 
.A1(n_646),
.A2(n_579),
.B(n_576),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_593),
.B(n_469),
.Y(n_767)
);

AOI21xp5_ASAP7_75t_L g768 ( 
.A1(n_644),
.A2(n_469),
.B(n_500),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_615),
.B(n_549),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_653),
.B(n_280),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_623),
.B(n_549),
.Y(n_771)
);

AND2x2_ASAP7_75t_L g772 ( 
.A(n_620),
.B(n_281),
.Y(n_772)
);

OAI21xp5_ASAP7_75t_L g773 ( 
.A1(n_602),
.A2(n_553),
.B(n_579),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_624),
.B(n_549),
.Y(n_774)
);

NOR2xp67_ASAP7_75t_L g775 ( 
.A(n_581),
.B(n_577),
.Y(n_775)
);

AOI21xp5_ASAP7_75t_L g776 ( 
.A1(n_603),
.A2(n_678),
.B(n_676),
.Y(n_776)
);

AOI21xp5_ASAP7_75t_L g777 ( 
.A1(n_679),
.A2(n_537),
.B(n_447),
.Y(n_777)
);

INVx2_ASAP7_75t_SL g778 ( 
.A(n_630),
.Y(n_778)
);

AOI22xp5_ASAP7_75t_L g779 ( 
.A1(n_591),
.A2(n_529),
.B1(n_539),
.B2(n_578),
.Y(n_779)
);

A2O1A1Ixp33_ASAP7_75t_L g780 ( 
.A1(n_695),
.A2(n_283),
.B(n_284),
.C(n_299),
.Y(n_780)
);

AOI22x1_ASAP7_75t_L g781 ( 
.A1(n_634),
.A2(n_531),
.B1(n_486),
.B2(n_571),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_688),
.Y(n_782)
);

BUFx2_ASAP7_75t_SL g783 ( 
.A(n_622),
.Y(n_783)
);

O2A1O1Ixp5_ASAP7_75t_L g784 ( 
.A1(n_666),
.A2(n_553),
.B(n_578),
.C(n_577),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_596),
.Y(n_785)
);

BUFx6f_ASAP7_75t_L g786 ( 
.A(n_730),
.Y(n_786)
);

AOI21xp5_ASAP7_75t_L g787 ( 
.A1(n_684),
.A2(n_500),
.B(n_537),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_625),
.B(n_549),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_635),
.B(n_560),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_593),
.B(n_486),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_693),
.Y(n_791)
);

BUFx4f_ASAP7_75t_SL g792 ( 
.A(n_616),
.Y(n_792)
);

AOI21xp5_ASAP7_75t_L g793 ( 
.A1(n_685),
.A2(n_500),
.B(n_537),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_635),
.B(n_560),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_606),
.Y(n_795)
);

OAI21xp5_ASAP7_75t_L g796 ( 
.A1(n_591),
.A2(n_571),
.B(n_570),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_611),
.B(n_560),
.Y(n_797)
);

AOI21xp5_ASAP7_75t_L g798 ( 
.A1(n_687),
.A2(n_500),
.B(n_537),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_618),
.B(n_655),
.Y(n_799)
);

AOI21xp5_ASAP7_75t_L g800 ( 
.A1(n_730),
.A2(n_500),
.B(n_537),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_655),
.B(n_486),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_589),
.B(n_263),
.Y(n_802)
);

AOI21xp5_ASAP7_75t_L g803 ( 
.A1(n_730),
.A2(n_500),
.B(n_537),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_667),
.B(n_489),
.Y(n_804)
);

AOI33xp33_ASAP7_75t_L g805 ( 
.A1(n_583),
.A2(n_714),
.A3(n_639),
.B1(n_587),
.B2(n_614),
.B3(n_686),
.Y(n_805)
);

AOI21xp5_ASAP7_75t_L g806 ( 
.A1(n_730),
.A2(n_447),
.B(n_570),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_735),
.A2(n_447),
.B(n_570),
.Y(n_807)
);

CKINVDCx16_ASAP7_75t_R g808 ( 
.A(n_700),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_638),
.B(n_494),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_695),
.B(n_301),
.Y(n_810)
);

AOI21xp5_ASAP7_75t_L g811 ( 
.A1(n_735),
.A2(n_571),
.B(n_568),
.Y(n_811)
);

NAND3xp33_ASAP7_75t_L g812 ( 
.A(n_682),
.B(n_290),
.C(n_293),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_648),
.B(n_494),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_614),
.B(n_494),
.Y(n_814)
);

BUFx3_ASAP7_75t_L g815 ( 
.A(n_582),
.Y(n_815)
);

OAI21xp5_ASAP7_75t_L g816 ( 
.A1(n_660),
.A2(n_651),
.B(n_646),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_691),
.B(n_531),
.Y(n_817)
);

NOR2xp67_ASAP7_75t_L g818 ( 
.A(n_717),
.B(n_516),
.Y(n_818)
);

AOI21xp5_ASAP7_75t_L g819 ( 
.A1(n_735),
.A2(n_568),
.B(n_566),
.Y(n_819)
);

BUFx3_ASAP7_75t_L g820 ( 
.A(n_582),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_584),
.B(n_284),
.Y(n_821)
);

OAI22xp5_ASAP7_75t_L g822 ( 
.A1(n_604),
.A2(n_517),
.B1(n_518),
.B2(n_519),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_L g823 ( 
.A(n_654),
.B(n_285),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_619),
.B(n_643),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_735),
.A2(n_568),
.B(n_566),
.Y(n_825)
);

AOI21xp5_ASAP7_75t_L g826 ( 
.A1(n_617),
.A2(n_566),
.B(n_562),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_617),
.A2(n_562),
.B(n_558),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_645),
.B(n_562),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_650),
.B(n_558),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_657),
.B(n_558),
.Y(n_830)
);

OAI21xp5_ASAP7_75t_L g831 ( 
.A1(n_651),
.A2(n_557),
.B(n_556),
.Y(n_831)
);

AOI22xp5_ASAP7_75t_L g832 ( 
.A1(n_682),
.A2(n_529),
.B1(n_539),
.B2(n_555),
.Y(n_832)
);

NOR2xp33_ASAP7_75t_L g833 ( 
.A(n_670),
.B(n_285),
.Y(n_833)
);

INVx3_ASAP7_75t_L g834 ( 
.A(n_664),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_701),
.B(n_292),
.Y(n_835)
);

BUFx2_ASAP7_75t_L g836 ( 
.A(n_633),
.Y(n_836)
);

BUFx4f_ASAP7_75t_L g837 ( 
.A(n_582),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_659),
.B(n_665),
.Y(n_838)
);

OAI21xp5_ASAP7_75t_L g839 ( 
.A1(n_658),
.A2(n_557),
.B(n_556),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_665),
.B(n_556),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_587),
.B(n_555),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_708),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_636),
.A2(n_552),
.B(n_531),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_707),
.B(n_292),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_675),
.B(n_552),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_637),
.B(n_534),
.Y(n_846)
);

INVx11_ASAP7_75t_L g847 ( 
.A(n_641),
.Y(n_847)
);

NAND2xp33_ASAP7_75t_L g848 ( 
.A(n_662),
.B(n_539),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_656),
.B(n_295),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_642),
.B(n_534),
.Y(n_850)
);

OAI21xp5_ASAP7_75t_L g851 ( 
.A1(n_599),
.A2(n_543),
.B(n_525),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_691),
.B(n_543),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_668),
.A2(n_674),
.B(n_673),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_691),
.B(n_538),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_722),
.B(n_295),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_647),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_694),
.A2(n_698),
.B(n_721),
.Y(n_857)
);

BUFx6f_ASAP7_75t_L g858 ( 
.A(n_662),
.Y(n_858)
);

BUFx6f_ASAP7_75t_L g859 ( 
.A(n_662),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_691),
.B(n_539),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_702),
.A2(n_498),
.B(n_293),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_703),
.A2(n_498),
.B(n_529),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_691),
.B(n_529),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_691),
.B(n_529),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_661),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_626),
.A2(n_498),
.B(n_539),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_598),
.B(n_11),
.Y(n_867)
);

O2A1O1Ixp5_ASAP7_75t_L g868 ( 
.A1(n_680),
.A2(n_539),
.B(n_57),
.C(n_66),
.Y(n_868)
);

AND2x4_ASAP7_75t_L g869 ( 
.A(n_706),
.B(n_539),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_734),
.A2(n_498),
.B(n_149),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_671),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_604),
.B(n_498),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_680),
.A2(n_146),
.B(n_134),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_731),
.Y(n_874)
);

OAI21xp5_ASAP7_75t_L g875 ( 
.A1(n_609),
.A2(n_133),
.B(n_132),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_733),
.B(n_13),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_690),
.B(n_15),
.Y(n_877)
);

OAI21xp5_ASAP7_75t_L g878 ( 
.A1(n_609),
.A2(n_129),
.B(n_128),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_690),
.B(n_15),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_677),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_706),
.B(n_16),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_732),
.B(n_124),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_SL g883 ( 
.A(n_639),
.B(n_112),
.Y(n_883)
);

O2A1O1Ixp5_ASAP7_75t_L g884 ( 
.A1(n_683),
.A2(n_111),
.B(n_107),
.C(n_106),
.Y(n_884)
);

O2A1O1Ixp33_ASAP7_75t_L g885 ( 
.A1(n_711),
.A2(n_17),
.B(n_20),
.C(n_21),
.Y(n_885)
);

OAI21xp33_ASAP7_75t_L g886 ( 
.A1(n_640),
.A2(n_22),
.B(n_24),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_683),
.A2(n_612),
.B(n_726),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_612),
.A2(n_104),
.B(n_96),
.Y(n_888)
);

O2A1O1Ixp33_ASAP7_75t_L g889 ( 
.A1(n_726),
.A2(n_22),
.B(n_24),
.C(n_25),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_699),
.B(n_94),
.Y(n_890)
);

NOR3xp33_ASAP7_75t_L g891 ( 
.A(n_722),
.B(n_27),
.C(n_30),
.Y(n_891)
);

AOI21xp33_ASAP7_75t_L g892 ( 
.A1(n_663),
.A2(n_31),
.B(n_34),
.Y(n_892)
);

OAI21xp5_ASAP7_75t_L g893 ( 
.A1(n_710),
.A2(n_91),
.B(n_84),
.Y(n_893)
);

OAI321xp33_ASAP7_75t_L g894 ( 
.A1(n_723),
.A2(n_31),
.A3(n_37),
.B1(n_41),
.B2(n_44),
.C(n_46),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_715),
.B(n_729),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_728),
.B(n_41),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_718),
.A2(n_69),
.B(n_48),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_714),
.B(n_47),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_724),
.B(n_50),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_633),
.B(n_52),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_704),
.A2(n_725),
.B(n_712),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_782),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_776),
.A2(n_774),
.B(n_771),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_857),
.A2(n_845),
.B(n_824),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_736),
.A2(n_621),
.B(n_725),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_SL g906 ( 
.A(n_764),
.B(n_597),
.Y(n_906)
);

AOI22xp5_ASAP7_75t_L g907 ( 
.A1(n_810),
.A2(n_633),
.B1(n_601),
.B2(n_669),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_782),
.Y(n_908)
);

OAI22xp5_ASAP7_75t_L g909 ( 
.A1(n_799),
.A2(n_601),
.B1(n_723),
.B2(n_610),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_755),
.B(n_610),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_747),
.B(n_712),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_847),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_743),
.B(n_739),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_740),
.A2(n_720),
.B(n_704),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_770),
.B(n_713),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_804),
.A2(n_750),
.B(n_738),
.Y(n_916)
);

A2O1A1Ixp33_ASAP7_75t_L g917 ( 
.A1(n_810),
.A2(n_709),
.B(n_607),
.C(n_720),
.Y(n_917)
);

OAI22xp5_ASAP7_75t_L g918 ( 
.A1(n_841),
.A2(n_789),
.B1(n_794),
.B2(n_769),
.Y(n_918)
);

NOR3xp33_ASAP7_75t_SL g919 ( 
.A(n_780),
.B(n_696),
.C(n_716),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_L g920 ( 
.A(n_737),
.B(n_713),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_L g921 ( 
.A(n_808),
.B(n_681),
.Y(n_921)
);

O2A1O1Ixp33_ASAP7_75t_L g922 ( 
.A1(n_877),
.A2(n_716),
.B(n_719),
.C(n_705),
.Y(n_922)
);

BUFx6f_ASAP7_75t_L g923 ( 
.A(n_858),
.Y(n_923)
);

NOR3xp33_ASAP7_75t_L g924 ( 
.A(n_833),
.B(n_727),
.C(n_849),
.Y(n_924)
);

NAND2x1p5_ASAP7_75t_L g925 ( 
.A(n_858),
.B(n_859),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_747),
.B(n_805),
.Y(n_926)
);

HB1xp67_ASAP7_75t_L g927 ( 
.A(n_745),
.Y(n_927)
);

BUFx2_ASAP7_75t_L g928 ( 
.A(n_836),
.Y(n_928)
);

BUFx6f_ASAP7_75t_L g929 ( 
.A(n_858),
.Y(n_929)
);

INVx4_ASAP7_75t_L g930 ( 
.A(n_858),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_R g931 ( 
.A(n_837),
.B(n_859),
.Y(n_931)
);

OAI22xp5_ASAP7_75t_L g932 ( 
.A1(n_838),
.A2(n_739),
.B1(n_801),
.B2(n_791),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_778),
.B(n_855),
.Y(n_933)
);

AOI22xp33_ASAP7_75t_L g934 ( 
.A1(n_879),
.A2(n_867),
.B1(n_833),
.B2(n_886),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_SL g935 ( 
.A(n_834),
.B(n_805),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_834),
.B(n_758),
.Y(n_936)
);

A2O1A1Ixp33_ASAP7_75t_SL g937 ( 
.A1(n_758),
.A2(n_761),
.B(n_867),
.C(n_849),
.Y(n_937)
);

INVx1_ASAP7_75t_SL g938 ( 
.A(n_772),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_L g939 ( 
.A(n_792),
.B(n_821),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_791),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_792),
.Y(n_941)
);

CKINVDCx14_ASAP7_75t_R g942 ( 
.A(n_835),
.Y(n_942)
);

NOR2xp67_ASAP7_75t_SL g943 ( 
.A(n_859),
.B(n_894),
.Y(n_943)
);

AND2x4_ASAP7_75t_L g944 ( 
.A(n_815),
.B(n_820),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_856),
.Y(n_945)
);

A2O1A1Ixp33_ASAP7_75t_SL g946 ( 
.A1(n_823),
.A2(n_821),
.B(n_881),
.C(n_893),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_752),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_853),
.A2(n_872),
.B(n_816),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_754),
.B(n_757),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_872),
.A2(n_887),
.B(n_787),
.Y(n_950)
);

OAI22xp5_ASAP7_75t_L g951 ( 
.A1(n_814),
.A2(n_883),
.B1(n_741),
.B2(n_842),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_R g952 ( 
.A(n_837),
.B(n_859),
.Y(n_952)
);

OAI22xp5_ASAP7_75t_L g953 ( 
.A1(n_814),
.A2(n_883),
.B1(n_741),
.B2(n_874),
.Y(n_953)
);

INVxp67_ASAP7_75t_L g954 ( 
.A(n_881),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_777),
.A2(n_793),
.B(n_798),
.Y(n_955)
);

INVx6_ASAP7_75t_L g956 ( 
.A(n_815),
.Y(n_956)
);

OAI21xp33_ASAP7_75t_L g957 ( 
.A1(n_823),
.A2(n_802),
.B(n_780),
.Y(n_957)
);

AOI22xp33_ASAP7_75t_SL g958 ( 
.A1(n_844),
.A2(n_898),
.B1(n_802),
.B2(n_783),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_817),
.A2(n_749),
.B(n_829),
.Y(n_959)
);

OAI21xp5_ASAP7_75t_L g960 ( 
.A1(n_748),
.A2(n_746),
.B(n_751),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_865),
.Y(n_961)
);

AO32x2_ASAP7_75t_L g962 ( 
.A1(n_822),
.A2(n_756),
.A3(n_746),
.B1(n_751),
.B2(n_773),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_754),
.B(n_757),
.Y(n_963)
);

OR2x6_ASAP7_75t_L g964 ( 
.A(n_820),
.B(n_869),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_817),
.A2(n_828),
.B(n_830),
.Y(n_965)
);

BUFx2_ASAP7_75t_L g966 ( 
.A(n_900),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_860),
.A2(n_863),
.B(n_864),
.Y(n_967)
);

A2O1A1Ixp33_ASAP7_75t_L g968 ( 
.A1(n_812),
.A2(n_892),
.B(n_901),
.C(n_756),
.Y(n_968)
);

O2A1O1Ixp33_ASAP7_75t_L g969 ( 
.A1(n_891),
.A2(n_876),
.B(n_889),
.C(n_882),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_800),
.A2(n_803),
.B(n_846),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_768),
.A2(n_854),
.B(n_852),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_763),
.B(n_775),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_788),
.B(n_880),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_852),
.A2(n_854),
.B(n_850),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_788),
.B(n_785),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_744),
.A2(n_767),
.B(n_840),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_895),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_882),
.Y(n_978)
);

OAI21xp5_ASAP7_75t_L g979 ( 
.A1(n_753),
.A2(n_796),
.B(n_762),
.Y(n_979)
);

O2A1O1Ixp33_ASAP7_75t_L g980 ( 
.A1(n_899),
.A2(n_896),
.B(n_885),
.C(n_744),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_SL g981 ( 
.A(n_869),
.B(n_818),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_797),
.B(n_795),
.Y(n_982)
);

INVx1_ASAP7_75t_SL g983 ( 
.A(n_871),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_767),
.A2(n_790),
.B(n_765),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_809),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_790),
.A2(n_765),
.B(n_807),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_L g987 ( 
.A(n_813),
.B(n_766),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_806),
.A2(n_851),
.B(n_759),
.Y(n_988)
);

OAI22xp5_ASAP7_75t_L g989 ( 
.A1(n_786),
.A2(n_781),
.B1(n_779),
.B2(n_832),
.Y(n_989)
);

INVx3_ASAP7_75t_L g990 ( 
.A(n_786),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_786),
.B(n_742),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_843),
.B(n_831),
.Y(n_992)
);

OAI22xp5_ASAP7_75t_L g993 ( 
.A1(n_839),
.A2(n_875),
.B1(n_878),
.B2(n_890),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_760),
.A2(n_811),
.B(n_819),
.Y(n_994)
);

BUFx8_ASAP7_75t_SL g995 ( 
.A(n_884),
.Y(n_995)
);

AND2x4_ASAP7_75t_L g996 ( 
.A(n_890),
.B(n_827),
.Y(n_996)
);

INVx4_ASAP7_75t_L g997 ( 
.A(n_848),
.Y(n_997)
);

OAI22xp5_ASAP7_75t_L g998 ( 
.A1(n_826),
.A2(n_825),
.B1(n_861),
.B2(n_897),
.Y(n_998)
);

A2O1A1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_784),
.A2(n_873),
.B(n_868),
.C(n_870),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_862),
.A2(n_888),
.B(n_866),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_L g1001 ( 
.A(n_810),
.B(n_440),
.Y(n_1001)
);

NAND3xp33_ASAP7_75t_L g1002 ( 
.A(n_810),
.B(n_392),
.C(n_695),
.Y(n_1002)
);

BUFx12f_ASAP7_75t_L g1003 ( 
.A(n_745),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_776),
.A2(n_506),
.B(n_474),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_810),
.B(n_440),
.Y(n_1005)
);

NOR2xp67_ASAP7_75t_L g1006 ( 
.A(n_812),
.B(n_581),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_782),
.Y(n_1007)
);

AO21x1_ASAP7_75t_L g1008 ( 
.A1(n_877),
.A2(n_879),
.B(n_603),
.Y(n_1008)
);

A2O1A1Ixp33_ASAP7_75t_SL g1009 ( 
.A1(n_810),
.A2(n_460),
.B(n_563),
.C(n_452),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_810),
.B(n_440),
.Y(n_1010)
);

A2O1A1Ixp33_ASAP7_75t_L g1011 ( 
.A1(n_810),
.A2(n_474),
.B(n_799),
.C(n_805),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_799),
.B(n_595),
.Y(n_1012)
);

O2A1O1Ixp33_ASAP7_75t_L g1013 ( 
.A1(n_810),
.A2(n_879),
.B(n_877),
.C(n_780),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_776),
.A2(n_506),
.B(n_474),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_776),
.A2(n_506),
.B(n_474),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_799),
.B(n_595),
.Y(n_1016)
);

BUFx2_ASAP7_75t_L g1017 ( 
.A(n_745),
.Y(n_1017)
);

O2A1O1Ixp33_ASAP7_75t_L g1018 ( 
.A1(n_810),
.A2(n_879),
.B(n_877),
.C(n_780),
.Y(n_1018)
);

CKINVDCx16_ASAP7_75t_R g1019 ( 
.A(n_808),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_776),
.A2(n_506),
.B(n_474),
.Y(n_1020)
);

NOR2xp33_ASAP7_75t_R g1021 ( 
.A(n_808),
.B(n_304),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_776),
.A2(n_506),
.B(n_474),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_L g1023 ( 
.A(n_810),
.B(n_440),
.Y(n_1023)
);

AOI22xp5_ASAP7_75t_L g1024 ( 
.A1(n_810),
.A2(n_764),
.B1(n_459),
.B2(n_452),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_764),
.B(n_440),
.Y(n_1025)
);

INVxp67_ASAP7_75t_L g1026 ( 
.A(n_745),
.Y(n_1026)
);

INVxp67_ASAP7_75t_L g1027 ( 
.A(n_745),
.Y(n_1027)
);

AND3x2_ASAP7_75t_L g1028 ( 
.A(n_810),
.B(n_732),
.C(n_695),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_SL g1029 ( 
.A(n_764),
.B(n_440),
.Y(n_1029)
);

HB1xp67_ASAP7_75t_L g1030 ( 
.A(n_745),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_947),
.Y(n_1031)
);

OAI21x1_ASAP7_75t_L g1032 ( 
.A1(n_986),
.A2(n_970),
.B(n_950),
.Y(n_1032)
);

NOR2xp33_ASAP7_75t_L g1033 ( 
.A(n_1002),
.B(n_1001),
.Y(n_1033)
);

AOI21x1_ASAP7_75t_L g1034 ( 
.A1(n_1004),
.A2(n_1015),
.B(n_1014),
.Y(n_1034)
);

NOR2xp33_ASAP7_75t_L g1035 ( 
.A(n_1005),
.B(n_1010),
.Y(n_1035)
);

OAI22x1_ASAP7_75t_L g1036 ( 
.A1(n_1024),
.A2(n_1023),
.B1(n_978),
.B2(n_907),
.Y(n_1036)
);

AOI22xp5_ASAP7_75t_L g1037 ( 
.A1(n_924),
.A2(n_939),
.B1(n_957),
.B2(n_1028),
.Y(n_1037)
);

OR2x2_ASAP7_75t_L g1038 ( 
.A(n_938),
.B(n_1019),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_904),
.A2(n_903),
.B(n_1022),
.Y(n_1039)
);

OAI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_1011),
.A2(n_968),
.B(n_1013),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_SL g1041 ( 
.A(n_958),
.B(n_933),
.Y(n_1041)
);

AND2x2_ASAP7_75t_L g1042 ( 
.A(n_966),
.B(n_954),
.Y(n_1042)
);

NAND2x1p5_ASAP7_75t_L g1043 ( 
.A(n_930),
.B(n_923),
.Y(n_1043)
);

AO31x2_ASAP7_75t_L g1044 ( 
.A1(n_1008),
.A2(n_993),
.A3(n_918),
.B(n_989),
.Y(n_1044)
);

OAI21x1_ASAP7_75t_L g1045 ( 
.A1(n_988),
.A2(n_955),
.B(n_1000),
.Y(n_1045)
);

OAI21x1_ASAP7_75t_L g1046 ( 
.A1(n_971),
.A2(n_994),
.B(n_984),
.Y(n_1046)
);

OAI21x1_ASAP7_75t_L g1047 ( 
.A1(n_916),
.A2(n_976),
.B(n_974),
.Y(n_1047)
);

BUFx3_ASAP7_75t_L g1048 ( 
.A(n_1003),
.Y(n_1048)
);

OAI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_1018),
.A2(n_934),
.B(n_960),
.Y(n_1049)
);

CKINVDCx11_ASAP7_75t_R g1050 ( 
.A(n_1017),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_1012),
.B(n_1016),
.Y(n_1051)
);

A2O1A1Ixp33_ASAP7_75t_L g1052 ( 
.A1(n_946),
.A2(n_969),
.B(n_1009),
.C(n_937),
.Y(n_1052)
);

O2A1O1Ixp33_ASAP7_75t_L g1053 ( 
.A1(n_906),
.A2(n_913),
.B(n_1025),
.C(n_1029),
.Y(n_1053)
);

OAI21x1_ASAP7_75t_L g1054 ( 
.A1(n_967),
.A2(n_1020),
.B(n_914),
.Y(n_1054)
);

OR2x2_ASAP7_75t_L g1055 ( 
.A(n_1030),
.B(n_1026),
.Y(n_1055)
);

A2O1A1Ixp33_ASAP7_75t_L g1056 ( 
.A1(n_980),
.A2(n_917),
.B(n_910),
.C(n_926),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_SL g1057 ( 
.A(n_949),
.B(n_963),
.Y(n_1057)
);

INVxp67_ASAP7_75t_SL g1058 ( 
.A(n_1027),
.Y(n_1058)
);

OAI22xp5_ASAP7_75t_L g1059 ( 
.A1(n_949),
.A2(n_963),
.B1(n_926),
.B2(n_911),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_948),
.A2(n_959),
.B(n_992),
.Y(n_1060)
);

AO31x2_ASAP7_75t_L g1061 ( 
.A1(n_999),
.A2(n_951),
.A3(n_953),
.B(n_998),
.Y(n_1061)
);

AO21x1_ASAP7_75t_L g1062 ( 
.A1(n_932),
.A2(n_991),
.B(n_910),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_908),
.Y(n_1063)
);

A2O1A1Ixp33_ASAP7_75t_L g1064 ( 
.A1(n_977),
.A2(n_919),
.B(n_922),
.C(n_909),
.Y(n_1064)
);

OR2x2_ASAP7_75t_L g1065 ( 
.A(n_928),
.B(n_983),
.Y(n_1065)
);

O2A1O1Ixp33_ASAP7_75t_SL g1066 ( 
.A1(n_935),
.A2(n_911),
.B(n_991),
.C(n_981),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_992),
.A2(n_965),
.B(n_979),
.Y(n_1067)
);

OAI22x1_ASAP7_75t_L g1068 ( 
.A1(n_941),
.A2(n_936),
.B1(n_920),
.B2(n_1007),
.Y(n_1068)
);

A2O1A1Ixp33_ASAP7_75t_L g1069 ( 
.A1(n_1006),
.A2(n_982),
.B(n_905),
.C(n_943),
.Y(n_1069)
);

NOR2xp67_ASAP7_75t_L g1070 ( 
.A(n_915),
.B(n_912),
.Y(n_1070)
);

INVxp67_ASAP7_75t_L g1071 ( 
.A(n_921),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_940),
.Y(n_1072)
);

AND2x2_ASAP7_75t_L g1073 ( 
.A(n_942),
.B(n_972),
.Y(n_1073)
);

A2O1A1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_987),
.A2(n_996),
.B(n_975),
.C(n_973),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_996),
.A2(n_997),
.B(n_985),
.Y(n_1075)
);

INVx1_ASAP7_75t_SL g1076 ( 
.A(n_1021),
.Y(n_1076)
);

OAI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_964),
.A2(n_997),
.B1(n_945),
.B2(n_961),
.Y(n_1077)
);

OR2x2_ASAP7_75t_L g1078 ( 
.A(n_964),
.B(n_944),
.Y(n_1078)
);

INVx2_ASAP7_75t_SL g1079 ( 
.A(n_956),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_990),
.B(n_995),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_L g1081 ( 
.A(n_956),
.B(n_964),
.Y(n_1081)
);

CKINVDCx6p67_ASAP7_75t_R g1082 ( 
.A(n_944),
.Y(n_1082)
);

AO31x2_ASAP7_75t_L g1083 ( 
.A1(n_962),
.A2(n_930),
.A3(n_925),
.B(n_929),
.Y(n_1083)
);

OAI21x1_ASAP7_75t_L g1084 ( 
.A1(n_962),
.A2(n_931),
.B(n_952),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_962),
.Y(n_1085)
);

A2O1A1Ixp33_ASAP7_75t_L g1086 ( 
.A1(n_923),
.A2(n_1002),
.B(n_957),
.C(n_810),
.Y(n_1086)
);

A2O1A1Ixp33_ASAP7_75t_L g1087 ( 
.A1(n_923),
.A2(n_1002),
.B(n_957),
.C(n_810),
.Y(n_1087)
);

OAI21x1_ASAP7_75t_L g1088 ( 
.A1(n_929),
.A2(n_986),
.B(n_970),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_929),
.B(n_956),
.Y(n_1089)
);

OAI21x1_ASAP7_75t_L g1090 ( 
.A1(n_986),
.A2(n_970),
.B(n_950),
.Y(n_1090)
);

OAI21x1_ASAP7_75t_L g1091 ( 
.A1(n_986),
.A2(n_970),
.B(n_950),
.Y(n_1091)
);

AOI221xp5_ASAP7_75t_SL g1092 ( 
.A1(n_934),
.A2(n_957),
.B1(n_886),
.B2(n_780),
.C(n_810),
.Y(n_1092)
);

BUFx3_ASAP7_75t_L g1093 ( 
.A(n_1003),
.Y(n_1093)
);

AND2x2_ASAP7_75t_L g1094 ( 
.A(n_1001),
.B(n_770),
.Y(n_1094)
);

OAI21x1_ASAP7_75t_L g1095 ( 
.A1(n_986),
.A2(n_970),
.B(n_950),
.Y(n_1095)
);

AOI22xp5_ASAP7_75t_L g1096 ( 
.A1(n_1002),
.A2(n_1005),
.B1(n_1010),
.B2(n_1001),
.Y(n_1096)
);

INVx4_ASAP7_75t_L g1097 ( 
.A(n_923),
.Y(n_1097)
);

BUFx8_ASAP7_75t_L g1098 ( 
.A(n_1017),
.Y(n_1098)
);

AO31x2_ASAP7_75t_L g1099 ( 
.A1(n_1008),
.A2(n_993),
.A3(n_918),
.B(n_989),
.Y(n_1099)
);

OAI21x1_ASAP7_75t_L g1100 ( 
.A1(n_986),
.A2(n_970),
.B(n_950),
.Y(n_1100)
);

OR2x2_ASAP7_75t_L g1101 ( 
.A(n_938),
.B(n_440),
.Y(n_1101)
);

NAND2x1p5_ASAP7_75t_L g1102 ( 
.A(n_930),
.B(n_858),
.Y(n_1102)
);

OAI21xp33_ASAP7_75t_L g1103 ( 
.A1(n_1002),
.A2(n_810),
.B(n_1001),
.Y(n_1103)
);

AND2x2_ASAP7_75t_L g1104 ( 
.A(n_1001),
.B(n_770),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_904),
.A2(n_903),
.B(n_1004),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_SL g1106 ( 
.A(n_1001),
.B(n_1005),
.Y(n_1106)
);

CKINVDCx11_ASAP7_75t_R g1107 ( 
.A(n_1003),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_902),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_904),
.A2(n_903),
.B(n_1004),
.Y(n_1109)
);

OAI22xp5_ASAP7_75t_L g1110 ( 
.A1(n_1002),
.A2(n_934),
.B1(n_963),
.B2(n_949),
.Y(n_1110)
);

A2O1A1Ixp33_ASAP7_75t_L g1111 ( 
.A1(n_1002),
.A2(n_957),
.B(n_810),
.C(n_1013),
.Y(n_1111)
);

NOR2xp33_ASAP7_75t_L g1112 ( 
.A(n_1002),
.B(n_1001),
.Y(n_1112)
);

AOI22xp5_ASAP7_75t_L g1113 ( 
.A1(n_1002),
.A2(n_1005),
.B1(n_1010),
.B2(n_1001),
.Y(n_1113)
);

A2O1A1Ixp33_ASAP7_75t_L g1114 ( 
.A1(n_1002),
.A2(n_957),
.B(n_810),
.C(n_1013),
.Y(n_1114)
);

AOI221x1_ASAP7_75t_L g1115 ( 
.A1(n_1002),
.A2(n_957),
.B1(n_810),
.B2(n_924),
.C(n_879),
.Y(n_1115)
);

OAI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_1002),
.A2(n_1011),
.B(n_968),
.Y(n_1116)
);

O2A1O1Ixp33_ASAP7_75t_L g1117 ( 
.A1(n_1002),
.A2(n_810),
.B(n_946),
.C(n_1001),
.Y(n_1117)
);

INVxp67_ASAP7_75t_L g1118 ( 
.A(n_927),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_904),
.A2(n_916),
.B(n_955),
.Y(n_1119)
);

AO32x2_ASAP7_75t_L g1120 ( 
.A1(n_918),
.A2(n_932),
.A3(n_993),
.B1(n_953),
.B2(n_951),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_947),
.Y(n_1121)
);

BUFx2_ASAP7_75t_SL g1122 ( 
.A(n_944),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_904),
.A2(n_916),
.B(n_955),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_947),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_904),
.A2(n_903),
.B(n_1004),
.Y(n_1125)
);

OAI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_1002),
.A2(n_1011),
.B(n_968),
.Y(n_1126)
);

AND2x2_ASAP7_75t_L g1127 ( 
.A(n_1001),
.B(n_770),
.Y(n_1127)
);

INVxp67_ASAP7_75t_L g1128 ( 
.A(n_927),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_904),
.A2(n_903),
.B(n_1004),
.Y(n_1129)
);

INVx2_ASAP7_75t_SL g1130 ( 
.A(n_1003),
.Y(n_1130)
);

OAI21x1_ASAP7_75t_L g1131 ( 
.A1(n_986),
.A2(n_970),
.B(n_950),
.Y(n_1131)
);

OAI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_1002),
.A2(n_1011),
.B(n_968),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_904),
.A2(n_903),
.B(n_1004),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_SL g1134 ( 
.A1(n_1011),
.A2(n_591),
.B(n_883),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_904),
.A2(n_903),
.B(n_1004),
.Y(n_1135)
);

HB1xp67_ASAP7_75t_L g1136 ( 
.A(n_1017),
.Y(n_1136)
);

O2A1O1Ixp33_ASAP7_75t_L g1137 ( 
.A1(n_1002),
.A2(n_810),
.B(n_946),
.C(n_1001),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_947),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_904),
.A2(n_903),
.B(n_1004),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_904),
.A2(n_903),
.B(n_1004),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_947),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_904),
.A2(n_916),
.B(n_955),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_902),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_947),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_904),
.A2(n_903),
.B(n_1004),
.Y(n_1145)
);

AOI221x1_ASAP7_75t_L g1146 ( 
.A1(n_1002),
.A2(n_957),
.B1(n_810),
.B2(n_924),
.C(n_879),
.Y(n_1146)
);

CKINVDCx11_ASAP7_75t_R g1147 ( 
.A(n_1003),
.Y(n_1147)
);

BUFx12f_ASAP7_75t_L g1148 ( 
.A(n_912),
.Y(n_1148)
);

OR2x2_ASAP7_75t_L g1149 ( 
.A(n_938),
.B(n_440),
.Y(n_1149)
);

AO31x2_ASAP7_75t_L g1150 ( 
.A1(n_1008),
.A2(n_993),
.A3(n_918),
.B(n_989),
.Y(n_1150)
);

O2A1O1Ixp33_ASAP7_75t_L g1151 ( 
.A1(n_1002),
.A2(n_810),
.B(n_946),
.C(n_1001),
.Y(n_1151)
);

INVx3_ASAP7_75t_L g1152 ( 
.A(n_930),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1012),
.B(n_1016),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_904),
.A2(n_916),
.B(n_955),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_947),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1012),
.B(n_1016),
.Y(n_1156)
);

OAI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_1002),
.A2(n_1011),
.B(n_968),
.Y(n_1157)
);

OAI21x1_ASAP7_75t_L g1158 ( 
.A1(n_986),
.A2(n_970),
.B(n_950),
.Y(n_1158)
);

BUFx6f_ASAP7_75t_L g1159 ( 
.A(n_923),
.Y(n_1159)
);

AOI22xp33_ASAP7_75t_L g1160 ( 
.A1(n_1103),
.A2(n_1035),
.B1(n_1112),
.B2(n_1033),
.Y(n_1160)
);

INVx6_ASAP7_75t_L g1161 ( 
.A(n_1098),
.Y(n_1161)
);

BUFx3_ASAP7_75t_L g1162 ( 
.A(n_1098),
.Y(n_1162)
);

AOI22xp33_ASAP7_75t_SL g1163 ( 
.A1(n_1110),
.A2(n_1049),
.B1(n_1040),
.B2(n_1104),
.Y(n_1163)
);

BUFx4f_ASAP7_75t_SL g1164 ( 
.A(n_1148),
.Y(n_1164)
);

OAI22xp33_ASAP7_75t_L g1165 ( 
.A1(n_1096),
.A2(n_1113),
.B1(n_1051),
.B2(n_1156),
.Y(n_1165)
);

BUFx10_ASAP7_75t_L g1166 ( 
.A(n_1079),
.Y(n_1166)
);

OAI22xp33_ASAP7_75t_L g1167 ( 
.A1(n_1051),
.A2(n_1153),
.B1(n_1156),
.B2(n_1106),
.Y(n_1167)
);

OAI22xp5_ASAP7_75t_L g1168 ( 
.A1(n_1153),
.A2(n_1037),
.B1(n_1111),
.B2(n_1114),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1031),
.Y(n_1169)
);

BUFx12f_ASAP7_75t_L g1170 ( 
.A(n_1107),
.Y(n_1170)
);

AOI22xp33_ASAP7_75t_L g1171 ( 
.A1(n_1110),
.A2(n_1036),
.B1(n_1049),
.B2(n_1041),
.Y(n_1171)
);

INVx8_ASAP7_75t_L g1172 ( 
.A(n_1159),
.Y(n_1172)
);

BUFx2_ASAP7_75t_L g1173 ( 
.A(n_1136),
.Y(n_1173)
);

INVx6_ASAP7_75t_L g1174 ( 
.A(n_1097),
.Y(n_1174)
);

BUFx12f_ASAP7_75t_L g1175 ( 
.A(n_1147),
.Y(n_1175)
);

BUFx12f_ASAP7_75t_L g1176 ( 
.A(n_1050),
.Y(n_1176)
);

AOI22xp33_ASAP7_75t_L g1177 ( 
.A1(n_1116),
.A2(n_1132),
.B1(n_1157),
.B2(n_1126),
.Y(n_1177)
);

CKINVDCx11_ASAP7_75t_R g1178 ( 
.A(n_1076),
.Y(n_1178)
);

CKINVDCx20_ASAP7_75t_R g1179 ( 
.A(n_1082),
.Y(n_1179)
);

AOI22xp33_ASAP7_75t_L g1180 ( 
.A1(n_1116),
.A2(n_1126),
.B1(n_1157),
.B2(n_1132),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_1076),
.Y(n_1181)
);

INVx1_ASAP7_75t_SL g1182 ( 
.A(n_1101),
.Y(n_1182)
);

OAI22xp5_ASAP7_75t_L g1183 ( 
.A1(n_1080),
.A2(n_1149),
.B1(n_1094),
.B2(n_1127),
.Y(n_1183)
);

OAI21xp5_ASAP7_75t_SL g1184 ( 
.A1(n_1117),
.A2(n_1151),
.B(n_1137),
.Y(n_1184)
);

BUFx12f_ASAP7_75t_L g1185 ( 
.A(n_1130),
.Y(n_1185)
);

AOI22xp33_ASAP7_75t_L g1186 ( 
.A1(n_1040),
.A2(n_1059),
.B1(n_1057),
.B2(n_1062),
.Y(n_1186)
);

AOI22xp33_ASAP7_75t_L g1187 ( 
.A1(n_1059),
.A2(n_1042),
.B1(n_1068),
.B2(n_1092),
.Y(n_1187)
);

OAI22xp5_ASAP7_75t_L g1188 ( 
.A1(n_1080),
.A2(n_1087),
.B1(n_1086),
.B2(n_1065),
.Y(n_1188)
);

AOI22xp33_ASAP7_75t_L g1189 ( 
.A1(n_1092),
.A2(n_1121),
.B1(n_1155),
.B2(n_1141),
.Y(n_1189)
);

BUFx12f_ASAP7_75t_L g1190 ( 
.A(n_1038),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1124),
.Y(n_1191)
);

BUFx2_ASAP7_75t_L g1192 ( 
.A(n_1058),
.Y(n_1192)
);

INVx6_ASAP7_75t_L g1193 ( 
.A(n_1097),
.Y(n_1193)
);

AOI22xp33_ASAP7_75t_L g1194 ( 
.A1(n_1138),
.A2(n_1144),
.B1(n_1072),
.B2(n_1063),
.Y(n_1194)
);

BUFx2_ASAP7_75t_L g1195 ( 
.A(n_1118),
.Y(n_1195)
);

BUFx12f_ASAP7_75t_L g1196 ( 
.A(n_1055),
.Y(n_1196)
);

CKINVDCx6p67_ASAP7_75t_R g1197 ( 
.A(n_1048),
.Y(n_1197)
);

AOI22xp33_ASAP7_75t_L g1198 ( 
.A1(n_1071),
.A2(n_1108),
.B1(n_1143),
.B2(n_1077),
.Y(n_1198)
);

AOI22xp33_ASAP7_75t_L g1199 ( 
.A1(n_1077),
.A2(n_1075),
.B1(n_1115),
.B2(n_1146),
.Y(n_1199)
);

OAI22xp5_ASAP7_75t_L g1200 ( 
.A1(n_1064),
.A2(n_1070),
.B1(n_1074),
.B2(n_1128),
.Y(n_1200)
);

AND2x2_ASAP7_75t_L g1201 ( 
.A(n_1073),
.B(n_1078),
.Y(n_1201)
);

BUFx2_ASAP7_75t_SL g1202 ( 
.A(n_1093),
.Y(n_1202)
);

BUFx4f_ASAP7_75t_SL g1203 ( 
.A(n_1159),
.Y(n_1203)
);

AOI22xp5_ASAP7_75t_L g1204 ( 
.A1(n_1081),
.A2(n_1122),
.B1(n_1069),
.B2(n_1066),
.Y(n_1204)
);

BUFx6f_ASAP7_75t_L g1205 ( 
.A(n_1043),
.Y(n_1205)
);

OR2x2_ASAP7_75t_L g1206 ( 
.A(n_1089),
.B(n_1056),
.Y(n_1206)
);

INVx8_ASAP7_75t_L g1207 ( 
.A(n_1152),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1083),
.Y(n_1208)
);

INVx3_ASAP7_75t_SL g1209 ( 
.A(n_1053),
.Y(n_1209)
);

CKINVDCx6p67_ASAP7_75t_R g1210 ( 
.A(n_1102),
.Y(n_1210)
);

INVxp67_ASAP7_75t_L g1211 ( 
.A(n_1084),
.Y(n_1211)
);

CKINVDCx11_ASAP7_75t_R g1212 ( 
.A(n_1085),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1075),
.Y(n_1213)
);

AOI21xp33_ASAP7_75t_L g1214 ( 
.A1(n_1052),
.A2(n_1067),
.B(n_1046),
.Y(n_1214)
);

HB1xp67_ASAP7_75t_L g1215 ( 
.A(n_1061),
.Y(n_1215)
);

BUFx4f_ASAP7_75t_SL g1216 ( 
.A(n_1134),
.Y(n_1216)
);

INVx4_ASAP7_75t_L g1217 ( 
.A(n_1088),
.Y(n_1217)
);

AOI22xp33_ASAP7_75t_L g1218 ( 
.A1(n_1060),
.A2(n_1139),
.B1(n_1109),
.B2(n_1039),
.Y(n_1218)
);

INVx3_ASAP7_75t_L g1219 ( 
.A(n_1034),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1044),
.Y(n_1220)
);

AOI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_1105),
.A2(n_1135),
.B1(n_1145),
.B2(n_1125),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_1129),
.Y(n_1222)
);

AOI22xp5_ASAP7_75t_L g1223 ( 
.A1(n_1133),
.A2(n_1140),
.B1(n_1054),
.B2(n_1142),
.Y(n_1223)
);

OAI22xp5_ASAP7_75t_L g1224 ( 
.A1(n_1119),
.A2(n_1154),
.B1(n_1123),
.B2(n_1142),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1099),
.Y(n_1225)
);

OAI22xp33_ASAP7_75t_L g1226 ( 
.A1(n_1120),
.A2(n_1150),
.B1(n_1154),
.B2(n_1123),
.Y(n_1226)
);

OAI22xp33_ASAP7_75t_SL g1227 ( 
.A1(n_1120),
.A2(n_1119),
.B1(n_1061),
.B2(n_1047),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1061),
.B(n_1045),
.Y(n_1228)
);

BUFx10_ASAP7_75t_L g1229 ( 
.A(n_1120),
.Y(n_1229)
);

OAI22xp5_ASAP7_75t_L g1230 ( 
.A1(n_1032),
.A2(n_1090),
.B1(n_1091),
.B2(n_1095),
.Y(n_1230)
);

INVxp67_ASAP7_75t_SL g1231 ( 
.A(n_1100),
.Y(n_1231)
);

AOI22xp33_ASAP7_75t_L g1232 ( 
.A1(n_1131),
.A2(n_1002),
.B1(n_1103),
.B2(n_1035),
.Y(n_1232)
);

BUFx4_ASAP7_75t_SL g1233 ( 
.A(n_1158),
.Y(n_1233)
);

OAI22xp5_ASAP7_75t_L g1234 ( 
.A1(n_1035),
.A2(n_1002),
.B1(n_1005),
.B2(n_1001),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1031),
.Y(n_1235)
);

AOI22xp33_ASAP7_75t_L g1236 ( 
.A1(n_1103),
.A2(n_1002),
.B1(n_1035),
.B2(n_1033),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1031),
.Y(n_1237)
);

BUFx2_ASAP7_75t_L g1238 ( 
.A(n_1098),
.Y(n_1238)
);

INVx6_ASAP7_75t_L g1239 ( 
.A(n_1098),
.Y(n_1239)
);

BUFx4_ASAP7_75t_SL g1240 ( 
.A(n_1048),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1031),
.Y(n_1241)
);

OAI22xp33_ASAP7_75t_L g1242 ( 
.A1(n_1096),
.A2(n_1002),
.B1(n_1113),
.B2(n_1035),
.Y(n_1242)
);

BUFx2_ASAP7_75t_SL g1243 ( 
.A(n_1070),
.Y(n_1243)
);

AOI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_1035),
.A2(n_1002),
.B1(n_1005),
.B2(n_1001),
.Y(n_1244)
);

OAI22xp5_ASAP7_75t_L g1245 ( 
.A1(n_1035),
.A2(n_1002),
.B1(n_1005),
.B2(n_1001),
.Y(n_1245)
);

INVx4_ASAP7_75t_L g1246 ( 
.A(n_1159),
.Y(n_1246)
);

AOI22xp33_ASAP7_75t_L g1247 ( 
.A1(n_1103),
.A2(n_1002),
.B1(n_1035),
.B2(n_1033),
.Y(n_1247)
);

BUFx2_ASAP7_75t_L g1248 ( 
.A(n_1098),
.Y(n_1248)
);

INVx3_ASAP7_75t_L g1249 ( 
.A(n_1097),
.Y(n_1249)
);

BUFx8_ASAP7_75t_L g1250 ( 
.A(n_1148),
.Y(n_1250)
);

AOI22xp33_ASAP7_75t_L g1251 ( 
.A1(n_1103),
.A2(n_1002),
.B1(n_1035),
.B2(n_1033),
.Y(n_1251)
);

INVx6_ASAP7_75t_L g1252 ( 
.A(n_1098),
.Y(n_1252)
);

INVx6_ASAP7_75t_L g1253 ( 
.A(n_1098),
.Y(n_1253)
);

BUFx2_ASAP7_75t_SL g1254 ( 
.A(n_1070),
.Y(n_1254)
);

OAI22xp5_ASAP7_75t_L g1255 ( 
.A1(n_1035),
.A2(n_1002),
.B1(n_1005),
.B2(n_1001),
.Y(n_1255)
);

AOI22xp33_ASAP7_75t_SL g1256 ( 
.A1(n_1035),
.A2(n_1002),
.B1(n_810),
.B2(n_1033),
.Y(n_1256)
);

INVx3_ASAP7_75t_L g1257 ( 
.A(n_1097),
.Y(n_1257)
);

AOI22xp33_ASAP7_75t_L g1258 ( 
.A1(n_1103),
.A2(n_1002),
.B1(n_1035),
.B2(n_1033),
.Y(n_1258)
);

AOI22xp33_ASAP7_75t_L g1259 ( 
.A1(n_1103),
.A2(n_1002),
.B1(n_1035),
.B2(n_1033),
.Y(n_1259)
);

INVx6_ASAP7_75t_L g1260 ( 
.A(n_1098),
.Y(n_1260)
);

BUFx3_ASAP7_75t_L g1261 ( 
.A(n_1098),
.Y(n_1261)
);

OAI22xp5_ASAP7_75t_L g1262 ( 
.A1(n_1035),
.A2(n_1002),
.B1(n_1005),
.B2(n_1001),
.Y(n_1262)
);

AND2x2_ASAP7_75t_L g1263 ( 
.A(n_1163),
.B(n_1177),
.Y(n_1263)
);

AND2x4_ASAP7_75t_L g1264 ( 
.A(n_1213),
.B(n_1211),
.Y(n_1264)
);

OAI21x1_ASAP7_75t_L g1265 ( 
.A1(n_1230),
.A2(n_1224),
.B(n_1219),
.Y(n_1265)
);

AO21x2_ASAP7_75t_L g1266 ( 
.A1(n_1214),
.A2(n_1221),
.B(n_1223),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1208),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1220),
.Y(n_1268)
);

INVxp67_ASAP7_75t_L g1269 ( 
.A(n_1173),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1225),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1215),
.Y(n_1271)
);

OA21x2_ASAP7_75t_L g1272 ( 
.A1(n_1218),
.A2(n_1199),
.B(n_1186),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1215),
.Y(n_1273)
);

OR2x2_ASAP7_75t_L g1274 ( 
.A(n_1184),
.B(n_1211),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1229),
.Y(n_1275)
);

HB1xp67_ASAP7_75t_L g1276 ( 
.A(n_1192),
.Y(n_1276)
);

NAND2x1p5_ASAP7_75t_L g1277 ( 
.A(n_1204),
.B(n_1217),
.Y(n_1277)
);

AO22x1_ASAP7_75t_L g1278 ( 
.A1(n_1209),
.A2(n_1262),
.B1(n_1245),
.B2(n_1255),
.Y(n_1278)
);

INVx2_ASAP7_75t_SL g1279 ( 
.A(n_1233),
.Y(n_1279)
);

BUFx2_ASAP7_75t_L g1280 ( 
.A(n_1222),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1165),
.B(n_1177),
.Y(n_1281)
);

AOI21x1_ASAP7_75t_L g1282 ( 
.A1(n_1228),
.A2(n_1168),
.B(n_1200),
.Y(n_1282)
);

BUFx12f_ASAP7_75t_L g1283 ( 
.A(n_1178),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1169),
.Y(n_1284)
);

OAI21x1_ASAP7_75t_L g1285 ( 
.A1(n_1218),
.A2(n_1231),
.B(n_1199),
.Y(n_1285)
);

INVx1_ASAP7_75t_SL g1286 ( 
.A(n_1209),
.Y(n_1286)
);

HB1xp67_ASAP7_75t_L g1287 ( 
.A(n_1206),
.Y(n_1287)
);

INVx4_ASAP7_75t_L g1288 ( 
.A(n_1216),
.Y(n_1288)
);

AOI22xp5_ASAP7_75t_L g1289 ( 
.A1(n_1256),
.A2(n_1242),
.B1(n_1234),
.B2(n_1244),
.Y(n_1289)
);

OR2x2_ASAP7_75t_L g1290 ( 
.A(n_1180),
.B(n_1187),
.Y(n_1290)
);

INVx3_ASAP7_75t_L g1291 ( 
.A(n_1216),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_1191),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_1235),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1237),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1241),
.Y(n_1295)
);

INVx2_ASAP7_75t_L g1296 ( 
.A(n_1231),
.Y(n_1296)
);

OA21x2_ASAP7_75t_L g1297 ( 
.A1(n_1186),
.A2(n_1180),
.B(n_1171),
.Y(n_1297)
);

INVx4_ASAP7_75t_L g1298 ( 
.A(n_1205),
.Y(n_1298)
);

BUFx2_ASAP7_75t_SL g1299 ( 
.A(n_1179),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_1178),
.Y(n_1300)
);

O2A1O1Ixp33_ASAP7_75t_SL g1301 ( 
.A1(n_1242),
.A2(n_1165),
.B(n_1167),
.C(n_1188),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1227),
.Y(n_1302)
);

AND2x2_ASAP7_75t_L g1303 ( 
.A(n_1163),
.B(n_1171),
.Y(n_1303)
);

HB1xp67_ASAP7_75t_L g1304 ( 
.A(n_1182),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1187),
.B(n_1232),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1226),
.Y(n_1306)
);

INVx1_ASAP7_75t_SL g1307 ( 
.A(n_1195),
.Y(n_1307)
);

OAI21x1_ASAP7_75t_L g1308 ( 
.A1(n_1189),
.A2(n_1194),
.B(n_1198),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1226),
.Y(n_1309)
);

AOI22xp33_ASAP7_75t_L g1310 ( 
.A1(n_1256),
.A2(n_1160),
.B1(n_1247),
.B2(n_1236),
.Y(n_1310)
);

OR2x6_ASAP7_75t_L g1311 ( 
.A(n_1243),
.B(n_1254),
.Y(n_1311)
);

OR2x2_ASAP7_75t_L g1312 ( 
.A(n_1183),
.B(n_1167),
.Y(n_1312)
);

OAI21x1_ASAP7_75t_L g1313 ( 
.A1(n_1189),
.A2(n_1194),
.B(n_1198),
.Y(n_1313)
);

BUFx3_ASAP7_75t_L g1314 ( 
.A(n_1196),
.Y(n_1314)
);

BUFx10_ASAP7_75t_L g1315 ( 
.A(n_1161),
.Y(n_1315)
);

INVx2_ASAP7_75t_SL g1316 ( 
.A(n_1207),
.Y(n_1316)
);

HB1xp67_ASAP7_75t_L g1317 ( 
.A(n_1201),
.Y(n_1317)
);

INVx2_ASAP7_75t_L g1318 ( 
.A(n_1212),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1212),
.Y(n_1319)
);

INVx2_ASAP7_75t_SL g1320 ( 
.A(n_1207),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1236),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1247),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1251),
.Y(n_1323)
);

AOI221xp5_ASAP7_75t_L g1324 ( 
.A1(n_1160),
.A2(n_1259),
.B1(n_1258),
.B2(n_1251),
.C(n_1181),
.Y(n_1324)
);

BUFx4f_ASAP7_75t_SL g1325 ( 
.A(n_1170),
.Y(n_1325)
);

OA21x2_ASAP7_75t_L g1326 ( 
.A1(n_1285),
.A2(n_1265),
.B(n_1302),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1317),
.B(n_1190),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1284),
.Y(n_1328)
);

OAI21xp5_ASAP7_75t_L g1329 ( 
.A1(n_1289),
.A2(n_1259),
.B(n_1258),
.Y(n_1329)
);

OR2x2_ASAP7_75t_L g1330 ( 
.A(n_1287),
.B(n_1238),
.Y(n_1330)
);

NOR2x1_ASAP7_75t_SL g1331 ( 
.A(n_1279),
.B(n_1176),
.Y(n_1331)
);

NOR2xp33_ASAP7_75t_L g1332 ( 
.A(n_1280),
.B(n_1286),
.Y(n_1332)
);

NAND2xp33_ASAP7_75t_SL g1333 ( 
.A(n_1280),
.B(n_1179),
.Y(n_1333)
);

AOI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1301),
.A2(n_1172),
.B(n_1257),
.Y(n_1334)
);

OR2x2_ASAP7_75t_L g1335 ( 
.A(n_1276),
.B(n_1248),
.Y(n_1335)
);

OAI21xp5_ASAP7_75t_L g1336 ( 
.A1(n_1289),
.A2(n_1257),
.B(n_1249),
.Y(n_1336)
);

NOR2xp33_ASAP7_75t_L g1337 ( 
.A(n_1286),
.B(n_1164),
.Y(n_1337)
);

OAI21xp5_ASAP7_75t_L g1338 ( 
.A1(n_1310),
.A2(n_1281),
.B(n_1324),
.Y(n_1338)
);

A2O1A1Ixp33_ASAP7_75t_L g1339 ( 
.A1(n_1324),
.A2(n_1261),
.B(n_1162),
.C(n_1202),
.Y(n_1339)
);

OA21x2_ASAP7_75t_L g1340 ( 
.A1(n_1285),
.A2(n_1210),
.B(n_1203),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1274),
.B(n_1166),
.Y(n_1341)
);

O2A1O1Ixp33_ASAP7_75t_L g1342 ( 
.A1(n_1281),
.A2(n_1261),
.B(n_1162),
.C(n_1240),
.Y(n_1342)
);

AOI22xp5_ASAP7_75t_L g1343 ( 
.A1(n_1278),
.A2(n_1161),
.B1(n_1253),
.B2(n_1252),
.Y(n_1343)
);

NAND3xp33_ASAP7_75t_L g1344 ( 
.A(n_1278),
.B(n_1321),
.C(n_1323),
.Y(n_1344)
);

OA21x2_ASAP7_75t_L g1345 ( 
.A1(n_1285),
.A2(n_1203),
.B(n_1172),
.Y(n_1345)
);

OR2x2_ASAP7_75t_L g1346 ( 
.A(n_1274),
.B(n_1197),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1318),
.B(n_1246),
.Y(n_1347)
);

OAI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_1322),
.A2(n_1240),
.B(n_1193),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1318),
.B(n_1161),
.Y(n_1349)
);

NAND3xp33_ASAP7_75t_L g1350 ( 
.A(n_1323),
.B(n_1250),
.C(n_1260),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1318),
.B(n_1239),
.Y(n_1351)
);

OA21x2_ASAP7_75t_L g1352 ( 
.A1(n_1265),
.A2(n_1193),
.B(n_1174),
.Y(n_1352)
);

A2O1A1Ixp33_ASAP7_75t_L g1353 ( 
.A1(n_1303),
.A2(n_1239),
.B(n_1253),
.C(n_1252),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1319),
.B(n_1239),
.Y(n_1354)
);

AOI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1266),
.A2(n_1174),
.B(n_1260),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1319),
.B(n_1260),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1319),
.B(n_1252),
.Y(n_1357)
);

AOI21xp5_ASAP7_75t_L g1358 ( 
.A1(n_1266),
.A2(n_1174),
.B(n_1164),
.Y(n_1358)
);

O2A1O1Ixp33_ASAP7_75t_L g1359 ( 
.A1(n_1303),
.A2(n_1185),
.B(n_1250),
.C(n_1175),
.Y(n_1359)
);

A2O1A1Ixp33_ASAP7_75t_L g1360 ( 
.A1(n_1263),
.A2(n_1312),
.B(n_1308),
.C(n_1313),
.Y(n_1360)
);

AO32x2_ASAP7_75t_L g1361 ( 
.A1(n_1298),
.A2(n_1320),
.A3(n_1288),
.B1(n_1302),
.B2(n_1316),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1292),
.B(n_1293),
.Y(n_1362)
);

AO32x2_ASAP7_75t_L g1363 ( 
.A1(n_1298),
.A2(n_1320),
.A3(n_1288),
.B1(n_1316),
.B2(n_1309),
.Y(n_1363)
);

NOR2x1_ASAP7_75t_SL g1364 ( 
.A(n_1311),
.B(n_1282),
.Y(n_1364)
);

A2O1A1Ixp33_ASAP7_75t_L g1365 ( 
.A1(n_1308),
.A2(n_1313),
.B(n_1290),
.C(n_1305),
.Y(n_1365)
);

OA21x2_ASAP7_75t_L g1366 ( 
.A1(n_1306),
.A2(n_1309),
.B(n_1282),
.Y(n_1366)
);

CKINVDCx20_ASAP7_75t_R g1367 ( 
.A(n_1325),
.Y(n_1367)
);

AOI211xp5_ASAP7_75t_L g1368 ( 
.A1(n_1305),
.A2(n_1307),
.B(n_1304),
.C(n_1269),
.Y(n_1368)
);

NOR2xp33_ASAP7_75t_L g1369 ( 
.A(n_1300),
.B(n_1307),
.Y(n_1369)
);

OAI21xp5_ASAP7_75t_L g1370 ( 
.A1(n_1297),
.A2(n_1272),
.B(n_1277),
.Y(n_1370)
);

NOR2xp33_ASAP7_75t_L g1371 ( 
.A(n_1283),
.B(n_1299),
.Y(n_1371)
);

NOR2xp33_ASAP7_75t_L g1372 ( 
.A(n_1283),
.B(n_1299),
.Y(n_1372)
);

AO32x2_ASAP7_75t_L g1373 ( 
.A1(n_1298),
.A2(n_1320),
.A3(n_1306),
.B1(n_1271),
.B2(n_1273),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1370),
.B(n_1266),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1362),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1328),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1373),
.B(n_1264),
.Y(n_1377)
);

NOR2xp33_ASAP7_75t_L g1378 ( 
.A(n_1329),
.B(n_1311),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1362),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1365),
.B(n_1264),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1373),
.B(n_1264),
.Y(n_1381)
);

OAI22xp5_ASAP7_75t_L g1382 ( 
.A1(n_1329),
.A2(n_1297),
.B1(n_1272),
.B2(n_1291),
.Y(n_1382)
);

INVxp67_ASAP7_75t_SL g1383 ( 
.A(n_1366),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1326),
.B(n_1296),
.Y(n_1384)
);

OR2x2_ASAP7_75t_L g1385 ( 
.A(n_1326),
.B(n_1296),
.Y(n_1385)
);

OR2x2_ASAP7_75t_L g1386 ( 
.A(n_1366),
.B(n_1267),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1345),
.B(n_1268),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1360),
.B(n_1294),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1363),
.B(n_1270),
.Y(n_1389)
);

AOI221xp5_ASAP7_75t_L g1390 ( 
.A1(n_1338),
.A2(n_1344),
.B1(n_1339),
.B2(n_1368),
.C(n_1342),
.Y(n_1390)
);

INVx3_ASAP7_75t_L g1391 ( 
.A(n_1352),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1368),
.B(n_1294),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1361),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_1363),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1344),
.B(n_1295),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1361),
.Y(n_1396)
);

NOR2x1p5_ASAP7_75t_L g1397 ( 
.A(n_1350),
.B(n_1291),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1394),
.B(n_1340),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1376),
.Y(n_1399)
);

BUFx3_ASAP7_75t_L g1400 ( 
.A(n_1389),
.Y(n_1400)
);

BUFx3_ASAP7_75t_L g1401 ( 
.A(n_1389),
.Y(n_1401)
);

INVx2_ASAP7_75t_L g1402 ( 
.A(n_1385),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1376),
.Y(n_1403)
);

OAI31xp33_ASAP7_75t_SL g1404 ( 
.A1(n_1390),
.A2(n_1338),
.A3(n_1350),
.B(n_1336),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1394),
.B(n_1377),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1375),
.B(n_1379),
.Y(n_1406)
);

NOR2xp33_ASAP7_75t_L g1407 ( 
.A(n_1378),
.B(n_1346),
.Y(n_1407)
);

INVx5_ASAP7_75t_L g1408 ( 
.A(n_1391),
.Y(n_1408)
);

OAI221xp5_ASAP7_75t_SL g1409 ( 
.A1(n_1390),
.A2(n_1342),
.B1(n_1343),
.B2(n_1359),
.C(n_1358),
.Y(n_1409)
);

BUFx3_ASAP7_75t_L g1410 ( 
.A(n_1389),
.Y(n_1410)
);

AOI22xp33_ASAP7_75t_SL g1411 ( 
.A1(n_1378),
.A2(n_1297),
.B1(n_1272),
.B2(n_1332),
.Y(n_1411)
);

INVx2_ASAP7_75t_SL g1412 ( 
.A(n_1384),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1394),
.B(n_1364),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1375),
.B(n_1358),
.Y(n_1414)
);

OAI21xp5_ASAP7_75t_L g1415 ( 
.A1(n_1382),
.A2(n_1297),
.B(n_1355),
.Y(n_1415)
);

NOR2xp33_ASAP7_75t_L g1416 ( 
.A(n_1392),
.B(n_1341),
.Y(n_1416)
);

AND2x2_ASAP7_75t_SL g1417 ( 
.A(n_1380),
.B(n_1272),
.Y(n_1417)
);

OAI211xp5_ASAP7_75t_L g1418 ( 
.A1(n_1382),
.A2(n_1333),
.B(n_1336),
.C(n_1353),
.Y(n_1418)
);

INVxp67_ASAP7_75t_L g1419 ( 
.A(n_1383),
.Y(n_1419)
);

AOI22xp33_ASAP7_75t_L g1420 ( 
.A1(n_1397),
.A2(n_1395),
.B1(n_1388),
.B2(n_1283),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1387),
.Y(n_1421)
);

INVxp67_ASAP7_75t_SL g1422 ( 
.A(n_1386),
.Y(n_1422)
);

OR2x2_ASAP7_75t_L g1423 ( 
.A(n_1393),
.B(n_1275),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1400),
.B(n_1381),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_1412),
.Y(n_1425)
);

NOR2x1p5_ASAP7_75t_L g1426 ( 
.A(n_1400),
.B(n_1380),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1419),
.B(n_1395),
.Y(n_1427)
);

INVx1_ASAP7_75t_SL g1428 ( 
.A(n_1414),
.Y(n_1428)
);

INVx3_ASAP7_75t_L g1429 ( 
.A(n_1408),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1412),
.Y(n_1430)
);

AND2x2_ASAP7_75t_SL g1431 ( 
.A(n_1417),
.B(n_1388),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1412),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1419),
.B(n_1375),
.Y(n_1433)
);

OR2x2_ASAP7_75t_L g1434 ( 
.A(n_1400),
.B(n_1393),
.Y(n_1434)
);

OR2x2_ASAP7_75t_L g1435 ( 
.A(n_1400),
.B(n_1393),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1399),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1399),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1399),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1403),
.Y(n_1439)
);

INVxp33_ASAP7_75t_L g1440 ( 
.A(n_1407),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1400),
.B(n_1381),
.Y(n_1441)
);

HB1xp67_ASAP7_75t_L g1442 ( 
.A(n_1419),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1401),
.B(n_1381),
.Y(n_1443)
);

NOR2xp33_ASAP7_75t_L g1444 ( 
.A(n_1407),
.B(n_1330),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1401),
.B(n_1396),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1401),
.B(n_1396),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1403),
.Y(n_1447)
);

AND2x4_ASAP7_75t_L g1448 ( 
.A(n_1408),
.B(n_1391),
.Y(n_1448)
);

OR2x2_ASAP7_75t_L g1449 ( 
.A(n_1401),
.B(n_1396),
.Y(n_1449)
);

OR2x2_ASAP7_75t_L g1450 ( 
.A(n_1401),
.B(n_1410),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1406),
.B(n_1414),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1410),
.B(n_1374),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1410),
.B(n_1374),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1406),
.B(n_1414),
.Y(n_1454)
);

OAI21xp5_ASAP7_75t_L g1455 ( 
.A1(n_1418),
.A2(n_1392),
.B(n_1374),
.Y(n_1455)
);

NOR2x1_ASAP7_75t_L g1456 ( 
.A(n_1418),
.B(n_1397),
.Y(n_1456)
);

HB1xp67_ASAP7_75t_L g1457 ( 
.A(n_1442),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1442),
.Y(n_1458)
);

NOR2x1p5_ASAP7_75t_SL g1459 ( 
.A(n_1450),
.B(n_1402),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1450),
.Y(n_1460)
);

OAI21xp33_ASAP7_75t_L g1461 ( 
.A1(n_1455),
.A2(n_1404),
.B(n_1417),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1426),
.B(n_1410),
.Y(n_1462)
);

NOR2x1p5_ASAP7_75t_SL g1463 ( 
.A(n_1450),
.B(n_1402),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1436),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1436),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1437),
.Y(n_1466)
);

OR2x2_ASAP7_75t_L g1467 ( 
.A(n_1428),
.B(n_1423),
.Y(n_1467)
);

AOI32xp33_ASAP7_75t_SL g1468 ( 
.A1(n_1427),
.A2(n_1416),
.A3(n_1422),
.B1(n_1371),
.B2(n_1372),
.Y(n_1468)
);

OR2x2_ASAP7_75t_L g1469 ( 
.A(n_1428),
.B(n_1423),
.Y(n_1469)
);

AND2x4_ASAP7_75t_L g1470 ( 
.A(n_1424),
.B(n_1410),
.Y(n_1470)
);

HB1xp67_ASAP7_75t_L g1471 ( 
.A(n_1434),
.Y(n_1471)
);

INVxp67_ASAP7_75t_SL g1472 ( 
.A(n_1456),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1426),
.B(n_1405),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1440),
.B(n_1416),
.Y(n_1474)
);

NAND2xp33_ASAP7_75t_L g1475 ( 
.A(n_1456),
.B(n_1397),
.Y(n_1475)
);

OR2x2_ASAP7_75t_L g1476 ( 
.A(n_1451),
.B(n_1423),
.Y(n_1476)
);

OR2x2_ASAP7_75t_L g1477 ( 
.A(n_1451),
.B(n_1423),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1438),
.Y(n_1478)
);

OAI32xp33_ASAP7_75t_L g1479 ( 
.A1(n_1455),
.A2(n_1415),
.A3(n_1420),
.B1(n_1413),
.B2(n_1398),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1424),
.B(n_1405),
.Y(n_1480)
);

OR2x2_ASAP7_75t_L g1481 ( 
.A(n_1454),
.B(n_1421),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1439),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1440),
.B(n_1404),
.Y(n_1483)
);

NAND2x1p5_ASAP7_75t_L g1484 ( 
.A(n_1429),
.B(n_1431),
.Y(n_1484)
);

NOR2xp33_ASAP7_75t_L g1485 ( 
.A(n_1444),
.B(n_1409),
.Y(n_1485)
);

BUFx2_ASAP7_75t_L g1486 ( 
.A(n_1424),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1447),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1444),
.B(n_1404),
.Y(n_1488)
);

NOR2xp67_ASAP7_75t_L g1489 ( 
.A(n_1429),
.B(n_1408),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1434),
.Y(n_1490)
);

INVx1_ASAP7_75t_SL g1491 ( 
.A(n_1431),
.Y(n_1491)
);

HB1xp67_ASAP7_75t_L g1492 ( 
.A(n_1434),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1431),
.B(n_1417),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1435),
.Y(n_1494)
);

OR2x2_ASAP7_75t_L g1495 ( 
.A(n_1460),
.B(n_1454),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_SL g1496 ( 
.A(n_1461),
.B(n_1431),
.Y(n_1496)
);

INVx3_ASAP7_75t_SL g1497 ( 
.A(n_1470),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1472),
.B(n_1427),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1462),
.B(n_1441),
.Y(n_1499)
);

OR2x2_ASAP7_75t_L g1500 ( 
.A(n_1460),
.B(n_1435),
.Y(n_1500)
);

NAND2x1p5_ASAP7_75t_L g1501 ( 
.A(n_1489),
.B(n_1417),
.Y(n_1501)
);

OAI31xp33_ASAP7_75t_L g1502 ( 
.A1(n_1485),
.A2(n_1409),
.A3(n_1418),
.B(n_1420),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1488),
.B(n_1445),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1462),
.B(n_1441),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1457),
.Y(n_1505)
);

OR2x2_ASAP7_75t_L g1506 ( 
.A(n_1494),
.B(n_1490),
.Y(n_1506)
);

OAI21xp5_ASAP7_75t_L g1507 ( 
.A1(n_1485),
.A2(n_1409),
.B(n_1417),
.Y(n_1507)
);

AND3x2_ASAP7_75t_L g1508 ( 
.A(n_1483),
.B(n_1337),
.C(n_1369),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1486),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1471),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1473),
.B(n_1441),
.Y(n_1511)
);

NAND4xp75_ASAP7_75t_L g1512 ( 
.A(n_1459),
.B(n_1415),
.C(n_1348),
.D(n_1453),
.Y(n_1512)
);

NOR2xp67_ASAP7_75t_L g1513 ( 
.A(n_1470),
.B(n_1492),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1473),
.B(n_1470),
.Y(n_1514)
);

AND2x4_ASAP7_75t_SL g1515 ( 
.A(n_1480),
.B(n_1315),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1484),
.B(n_1443),
.Y(n_1516)
);

INVxp67_ASAP7_75t_SL g1517 ( 
.A(n_1475),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1458),
.B(n_1445),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1464),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1484),
.B(n_1443),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1467),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1480),
.B(n_1443),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1491),
.B(n_1452),
.Y(n_1523)
);

NAND2x1_ASAP7_75t_L g1524 ( 
.A(n_1493),
.B(n_1452),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1475),
.B(n_1452),
.Y(n_1525)
);

HB1xp67_ASAP7_75t_L g1526 ( 
.A(n_1465),
.Y(n_1526)
);

INVx1_ASAP7_75t_SL g1527 ( 
.A(n_1474),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1476),
.B(n_1453),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1466),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1526),
.Y(n_1530)
);

OAI22xp5_ASAP7_75t_L g1531 ( 
.A1(n_1507),
.A2(n_1411),
.B1(n_1468),
.B2(n_1415),
.Y(n_1531)
);

OA22x2_ASAP7_75t_L g1532 ( 
.A1(n_1508),
.A2(n_1453),
.B1(n_1446),
.B2(n_1445),
.Y(n_1532)
);

A2O1A1Ixp33_ASAP7_75t_L g1533 ( 
.A1(n_1502),
.A2(n_1479),
.B(n_1463),
.C(n_1411),
.Y(n_1533)
);

AOI221xp5_ASAP7_75t_L g1534 ( 
.A1(n_1507),
.A2(n_1411),
.B1(n_1422),
.B2(n_1467),
.C(n_1469),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1514),
.B(n_1497),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1527),
.B(n_1413),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1526),
.Y(n_1537)
);

INVx2_ASAP7_75t_SL g1538 ( 
.A(n_1497),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1527),
.B(n_1413),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1519),
.Y(n_1540)
);

NAND2x1_ASAP7_75t_L g1541 ( 
.A(n_1513),
.B(n_1446),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1514),
.B(n_1446),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1519),
.Y(n_1543)
);

AOI21xp33_ASAP7_75t_SL g1544 ( 
.A1(n_1502),
.A2(n_1469),
.B(n_1351),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1529),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1529),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1510),
.Y(n_1547)
);

OAI32xp33_ASAP7_75t_L g1548 ( 
.A1(n_1496),
.A2(n_1449),
.A3(n_1435),
.B1(n_1477),
.B2(n_1476),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1510),
.Y(n_1549)
);

HB1xp67_ASAP7_75t_L g1550 ( 
.A(n_1513),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1517),
.B(n_1413),
.Y(n_1551)
);

OR2x2_ASAP7_75t_L g1552 ( 
.A(n_1503),
.B(n_1449),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1505),
.Y(n_1553)
);

OAI21xp5_ASAP7_75t_SL g1554 ( 
.A1(n_1508),
.A2(n_1348),
.B(n_1349),
.Y(n_1554)
);

OR2x2_ASAP7_75t_L g1555 ( 
.A(n_1538),
.B(n_1503),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1538),
.B(n_1517),
.Y(n_1556)
);

OAI221xp5_ASAP7_75t_L g1557 ( 
.A1(n_1533),
.A2(n_1524),
.B1(n_1497),
.B2(n_1498),
.C(n_1525),
.Y(n_1557)
);

INVx1_ASAP7_75t_SL g1558 ( 
.A(n_1535),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1544),
.B(n_1505),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1550),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1541),
.Y(n_1561)
);

NAND2x1_ASAP7_75t_L g1562 ( 
.A(n_1530),
.B(n_1525),
.Y(n_1562)
);

AOI21xp5_ASAP7_75t_L g1563 ( 
.A1(n_1533),
.A2(n_1498),
.B(n_1524),
.Y(n_1563)
);

O2A1O1Ixp33_ASAP7_75t_L g1564 ( 
.A1(n_1531),
.A2(n_1509),
.B(n_1518),
.C(n_1521),
.Y(n_1564)
);

INVxp67_ASAP7_75t_L g1565 ( 
.A(n_1550),
.Y(n_1565)
);

AND2x4_ASAP7_75t_L g1566 ( 
.A(n_1537),
.B(n_1509),
.Y(n_1566)
);

AOI21xp5_ASAP7_75t_L g1567 ( 
.A1(n_1554),
.A2(n_1509),
.B(n_1521),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1540),
.Y(n_1568)
);

INVx1_ASAP7_75t_SL g1569 ( 
.A(n_1547),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_1542),
.Y(n_1570)
);

OR2x2_ASAP7_75t_L g1571 ( 
.A(n_1552),
.B(n_1518),
.Y(n_1571)
);

OAI21xp33_ASAP7_75t_L g1572 ( 
.A1(n_1534),
.A2(n_1532),
.B(n_1551),
.Y(n_1572)
);

NOR4xp25_ASAP7_75t_L g1573 ( 
.A(n_1553),
.B(n_1521),
.C(n_1506),
.D(n_1523),
.Y(n_1573)
);

OR2x2_ASAP7_75t_L g1574 ( 
.A(n_1559),
.B(n_1549),
.Y(n_1574)
);

AOI21xp5_ASAP7_75t_L g1575 ( 
.A1(n_1564),
.A2(n_1534),
.B(n_1532),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1558),
.B(n_1499),
.Y(n_1576)
);

AOI22xp5_ASAP7_75t_L g1577 ( 
.A1(n_1557),
.A2(n_1512),
.B1(n_1523),
.B2(n_1520),
.Y(n_1577)
);

AOI21xp33_ASAP7_75t_SL g1578 ( 
.A1(n_1573),
.A2(n_1548),
.B(n_1501),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1560),
.Y(n_1579)
);

INVx1_ASAP7_75t_SL g1580 ( 
.A(n_1569),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1566),
.B(n_1543),
.Y(n_1581)
);

AOI221xp5_ASAP7_75t_L g1582 ( 
.A1(n_1573),
.A2(n_1546),
.B1(n_1545),
.B2(n_1539),
.C(n_1536),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1570),
.B(n_1561),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1566),
.B(n_1499),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1565),
.B(n_1504),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1576),
.B(n_1556),
.Y(n_1586)
);

NOR3xp33_ASAP7_75t_L g1587 ( 
.A(n_1585),
.B(n_1572),
.C(n_1555),
.Y(n_1587)
);

OAI21xp33_ASAP7_75t_L g1588 ( 
.A1(n_1575),
.A2(n_1563),
.B(n_1562),
.Y(n_1588)
);

NAND5xp2_ASAP7_75t_L g1589 ( 
.A(n_1577),
.B(n_1567),
.C(n_1568),
.D(n_1501),
.E(n_1520),
.Y(n_1589)
);

NAND4xp25_ASAP7_75t_L g1590 ( 
.A(n_1583),
.B(n_1569),
.C(n_1571),
.D(n_1516),
.Y(n_1590)
);

AOI221xp5_ASAP7_75t_L g1591 ( 
.A1(n_1578),
.A2(n_1516),
.B1(n_1506),
.B2(n_1504),
.C(n_1511),
.Y(n_1591)
);

INVx5_ASAP7_75t_L g1592 ( 
.A(n_1580),
.Y(n_1592)
);

NOR4xp25_ASAP7_75t_L g1593 ( 
.A(n_1580),
.B(n_1500),
.C(n_1495),
.D(n_1511),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1581),
.Y(n_1594)
);

OAI211xp5_ASAP7_75t_L g1595 ( 
.A1(n_1588),
.A2(n_1582),
.B(n_1574),
.C(n_1579),
.Y(n_1595)
);

NOR3xp33_ASAP7_75t_L g1596 ( 
.A(n_1586),
.B(n_1584),
.C(n_1512),
.Y(n_1596)
);

AOI221xp5_ASAP7_75t_L g1597 ( 
.A1(n_1593),
.A2(n_1500),
.B1(n_1528),
.B2(n_1501),
.C(n_1522),
.Y(n_1597)
);

AOI211xp5_ASAP7_75t_L g1598 ( 
.A1(n_1589),
.A2(n_1495),
.B(n_1528),
.C(n_1522),
.Y(n_1598)
);

AOI221xp5_ASAP7_75t_L g1599 ( 
.A1(n_1587),
.A2(n_1515),
.B1(n_1422),
.B2(n_1429),
.C(n_1482),
.Y(n_1599)
);

NOR4xp25_ASAP7_75t_L g1600 ( 
.A(n_1595),
.B(n_1594),
.C(n_1590),
.D(n_1592),
.Y(n_1600)
);

AOI222xp33_ASAP7_75t_L g1601 ( 
.A1(n_1597),
.A2(n_1591),
.B1(n_1592),
.B2(n_1463),
.C1(n_1515),
.C2(n_1398),
.Y(n_1601)
);

OAI211xp5_ASAP7_75t_SL g1602 ( 
.A1(n_1596),
.A2(n_1335),
.B(n_1429),
.C(n_1449),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1598),
.B(n_1515),
.Y(n_1603)
);

AOI211xp5_ASAP7_75t_L g1604 ( 
.A1(n_1599),
.A2(n_1354),
.B(n_1356),
.C(n_1357),
.Y(n_1604)
);

OAI221xp5_ASAP7_75t_L g1605 ( 
.A1(n_1595),
.A2(n_1429),
.B1(n_1314),
.B2(n_1477),
.C(n_1481),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1603),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1605),
.Y(n_1607)
);

AOI22xp5_ASAP7_75t_L g1608 ( 
.A1(n_1601),
.A2(n_1367),
.B1(n_1314),
.B2(n_1448),
.Y(n_1608)
);

OAI22xp33_ASAP7_75t_L g1609 ( 
.A1(n_1600),
.A2(n_1430),
.B1(n_1425),
.B2(n_1481),
.Y(n_1609)
);

INVx2_ASAP7_75t_SL g1610 ( 
.A(n_1602),
.Y(n_1610)
);

OAI22xp33_ASAP7_75t_L g1611 ( 
.A1(n_1608),
.A2(n_1430),
.B1(n_1425),
.B2(n_1432),
.Y(n_1611)
);

OAI211xp5_ASAP7_75t_L g1612 ( 
.A1(n_1606),
.A2(n_1604),
.B(n_1314),
.C(n_1408),
.Y(n_1612)
);

INVxp67_ASAP7_75t_L g1613 ( 
.A(n_1607),
.Y(n_1613)
);

AOI22xp33_ASAP7_75t_L g1614 ( 
.A1(n_1613),
.A2(n_1610),
.B1(n_1609),
.B2(n_1448),
.Y(n_1614)
);

AO22x2_ASAP7_75t_L g1615 ( 
.A1(n_1614),
.A2(n_1612),
.B1(n_1611),
.B2(n_1487),
.Y(n_1615)
);

AOI22xp5_ASAP7_75t_L g1616 ( 
.A1(n_1615),
.A2(n_1448),
.B1(n_1315),
.B2(n_1478),
.Y(n_1616)
);

INVxp67_ASAP7_75t_L g1617 ( 
.A(n_1616),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1617),
.Y(n_1618)
);

NAND2x1p5_ASAP7_75t_L g1619 ( 
.A(n_1618),
.B(n_1327),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1619),
.B(n_1331),
.Y(n_1620)
);

HB1xp67_ASAP7_75t_L g1621 ( 
.A(n_1620),
.Y(n_1621)
);

AOI221xp5_ASAP7_75t_L g1622 ( 
.A1(n_1621),
.A2(n_1448),
.B1(n_1433),
.B2(n_1425),
.C(n_1430),
.Y(n_1622)
);

AOI211xp5_ASAP7_75t_L g1623 ( 
.A1(n_1622),
.A2(n_1347),
.B(n_1398),
.C(n_1334),
.Y(n_1623)
);


endmodule