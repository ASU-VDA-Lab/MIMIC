module real_aes_6917_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_363;
wire n_182;
wire n_754;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_434;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_756;
wire n_598;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_420;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_314;
wire n_252;
wire n_283;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g108 ( .A(n_0), .Y(n_108) );
INVx1_ASAP7_75t_L g509 ( .A(n_1), .Y(n_509) );
INVx1_ASAP7_75t_L g266 ( .A(n_2), .Y(n_266) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_3), .A2(n_38), .B1(n_185), .B2(n_537), .Y(n_536) );
AOI21xp33_ASAP7_75t_L g173 ( .A1(n_4), .A2(n_174), .B(n_175), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_5), .B(n_172), .Y(n_486) );
AND2x6_ASAP7_75t_L g147 ( .A(n_6), .B(n_148), .Y(n_147) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_7), .A2(n_242), .B(n_243), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_8), .B(n_114), .Y(n_113) );
NOR2xp33_ASAP7_75t_L g450 ( .A(n_8), .B(n_39), .Y(n_450) );
INVx1_ASAP7_75t_L g182 ( .A(n_9), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_10), .B(n_234), .Y(n_233) );
INVx1_ASAP7_75t_L g144 ( .A(n_11), .Y(n_144) );
INVx1_ASAP7_75t_L g505 ( .A(n_12), .Y(n_505) );
INVx1_ASAP7_75t_L g248 ( .A(n_13), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_14), .B(n_150), .Y(n_543) );
AOI222xp33_ASAP7_75t_SL g454 ( .A1(n_15), .A2(n_455), .B1(n_456), .B2(n_465), .C1(n_752), .C2(n_753), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_16), .B(n_140), .Y(n_514) );
XNOR2xp5_ASAP7_75t_L g122 ( .A(n_17), .B(n_123), .Y(n_122) );
AO32x2_ASAP7_75t_L g534 ( .A1(n_17), .A2(n_139), .A3(n_172), .B1(n_497), .B2(n_535), .Y(n_534) );
NAND2xp5_ASAP7_75t_SL g546 ( .A(n_18), .B(n_185), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_19), .B(n_193), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_20), .B(n_140), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_21), .A2(n_50), .B1(n_185), .B2(n_537), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_22), .B(n_174), .Y(n_202) );
AOI22xp33_ASAP7_75t_SL g557 ( .A1(n_23), .A2(n_77), .B1(n_150), .B2(n_185), .Y(n_557) );
NAND2xp5_ASAP7_75t_SL g529 ( .A(n_24), .B(n_185), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_25), .B(n_170), .Y(n_196) );
OAI22xp5_ASAP7_75t_SL g456 ( .A1(n_26), .A2(n_457), .B1(n_458), .B2(n_464), .Y(n_456) );
INVx1_ASAP7_75t_L g464 ( .A(n_26), .Y(n_464) );
A2O1A1Ixp33_ASAP7_75t_L g245 ( .A1(n_27), .A2(n_246), .B(n_247), .C(n_249), .Y(n_245) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_28), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_29), .B(n_187), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_30), .B(n_180), .Y(n_267) );
INVx1_ASAP7_75t_L g158 ( .A(n_31), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_32), .B(n_187), .Y(n_531) );
INVx2_ASAP7_75t_L g152 ( .A(n_33), .Y(n_152) );
NAND2xp5_ASAP7_75t_SL g491 ( .A(n_34), .B(n_185), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_35), .B(n_187), .Y(n_548) );
AOI22xp5_ASAP7_75t_L g127 ( .A1(n_36), .A2(n_42), .B1(n_128), .B2(n_129), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_36), .Y(n_129) );
A2O1A1Ixp33_ASAP7_75t_L g203 ( .A1(n_37), .A2(n_147), .B(n_159), .C(n_204), .Y(n_203) );
INVx1_ASAP7_75t_L g114 ( .A(n_39), .Y(n_114) );
INVx1_ASAP7_75t_L g156 ( .A(n_40), .Y(n_156) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_41), .B(n_180), .Y(n_219) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_42), .Y(n_128) );
NAND2xp5_ASAP7_75t_SL g479 ( .A(n_43), .B(n_185), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_44), .A2(n_88), .B1(n_210), .B2(n_537), .Y(n_556) );
NAND2xp5_ASAP7_75t_SL g482 ( .A(n_45), .B(n_185), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_46), .B(n_185), .Y(n_506) );
CKINVDCx16_ASAP7_75t_R g162 ( .A(n_47), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_48), .B(n_484), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_49), .B(n_174), .Y(n_236) );
AOI22xp33_ASAP7_75t_SL g518 ( .A1(n_51), .A2(n_60), .B1(n_150), .B2(n_185), .Y(n_518) );
AOI22xp5_ASAP7_75t_L g149 ( .A1(n_52), .A2(n_150), .B1(n_153), .B2(n_159), .Y(n_149) );
CKINVDCx20_ASAP7_75t_R g213 ( .A(n_53), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g496 ( .A(n_54), .B(n_185), .Y(n_496) );
CKINVDCx16_ASAP7_75t_R g263 ( .A(n_55), .Y(n_263) );
NAND2xp5_ASAP7_75t_SL g542 ( .A(n_56), .B(n_185), .Y(n_542) );
A2O1A1Ixp33_ASAP7_75t_L g178 ( .A1(n_57), .A2(n_179), .B(n_181), .C(n_184), .Y(n_178) );
CKINVDCx20_ASAP7_75t_R g223 ( .A(n_58), .Y(n_223) );
INVx1_ASAP7_75t_L g176 ( .A(n_59), .Y(n_176) );
INVx1_ASAP7_75t_L g148 ( .A(n_61), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_62), .B(n_185), .Y(n_510) );
INVx1_ASAP7_75t_L g143 ( .A(n_63), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_64), .Y(n_120) );
AO32x2_ASAP7_75t_L g554 ( .A1(n_65), .A2(n_172), .A3(n_228), .B1(n_497), .B2(n_555), .Y(n_554) );
INVx1_ASAP7_75t_L g494 ( .A(n_66), .Y(n_494) );
OAI22xp5_ASAP7_75t_SL g125 ( .A1(n_67), .A2(n_126), .B1(n_127), .B2(n_130), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_67), .Y(n_130) );
INVx1_ASAP7_75t_L g526 ( .A(n_68), .Y(n_526) );
A2O1A1Ixp33_ASAP7_75t_SL g192 ( .A1(n_69), .A2(n_184), .B(n_193), .C(n_194), .Y(n_192) );
INVxp67_ASAP7_75t_L g195 ( .A(n_70), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_71), .B(n_150), .Y(n_527) );
INVx1_ASAP7_75t_L g112 ( .A(n_72), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g167 ( .A(n_73), .Y(n_167) );
INVx1_ASAP7_75t_L g216 ( .A(n_74), .Y(n_216) );
OAI22xp5_ASAP7_75t_L g461 ( .A1(n_75), .A2(n_102), .B1(n_462), .B2(n_463), .Y(n_461) );
CKINVDCx20_ASAP7_75t_R g462 ( .A(n_75), .Y(n_462) );
NAND2xp5_ASAP7_75t_SL g451 ( .A(n_76), .B(n_452), .Y(n_451) );
AOI22xp5_ASAP7_75t_L g104 ( .A1(n_78), .A2(n_105), .B1(n_115), .B2(n_757), .Y(n_104) );
A2O1A1Ixp33_ASAP7_75t_L g217 ( .A1(n_79), .A2(n_147), .B(n_159), .C(n_218), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_80), .B(n_537), .Y(n_547) );
NAND2xp5_ASAP7_75t_SL g530 ( .A(n_81), .B(n_150), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_82), .B(n_206), .Y(n_205) );
INVx2_ASAP7_75t_L g141 ( .A(n_83), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_84), .B(n_193), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_85), .B(n_150), .Y(n_480) );
A2O1A1Ixp33_ASAP7_75t_L g264 ( .A1(n_86), .A2(n_147), .B(n_159), .C(n_265), .Y(n_264) );
INVx2_ASAP7_75t_L g109 ( .A(n_87), .Y(n_109) );
OR2x2_ASAP7_75t_L g447 ( .A(n_87), .B(n_448), .Y(n_447) );
OR2x2_ASAP7_75t_L g468 ( .A(n_87), .B(n_449), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_89), .A2(n_103), .B1(n_150), .B2(n_151), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_90), .B(n_187), .Y(n_186) );
CKINVDCx20_ASAP7_75t_R g270 ( .A(n_91), .Y(n_270) );
A2O1A1Ixp33_ASAP7_75t_L g230 ( .A1(n_92), .A2(n_147), .B(n_159), .C(n_231), .Y(n_230) );
CKINVDCx20_ASAP7_75t_R g238 ( .A(n_93), .Y(n_238) );
INVx1_ASAP7_75t_L g191 ( .A(n_94), .Y(n_191) );
CKINVDCx16_ASAP7_75t_R g244 ( .A(n_95), .Y(n_244) );
NAND2xp5_ASAP7_75t_SL g232 ( .A(n_96), .B(n_206), .Y(n_232) );
AOI22xp5_ASAP7_75t_L g458 ( .A1(n_97), .A2(n_459), .B1(n_460), .B2(n_461), .Y(n_458) );
CKINVDCx20_ASAP7_75t_R g459 ( .A(n_97), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_98), .B(n_150), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_99), .B(n_172), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_100), .B(n_112), .Y(n_111) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_101), .A2(n_174), .B(n_190), .Y(n_189) );
CKINVDCx16_ASAP7_75t_R g463 ( .A(n_102), .Y(n_463) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g758 ( .A(n_106), .Y(n_758) );
OR2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_113), .Y(n_106) );
NAND3xp33_ASAP7_75t_SL g107 ( .A(n_108), .B(n_109), .C(n_110), .Y(n_107) );
AND2x2_ASAP7_75t_L g449 ( .A(n_108), .B(n_450), .Y(n_449) );
OR2x2_ASAP7_75t_L g751 ( .A(n_109), .B(n_449), .Y(n_751) );
NOR2x2_ASAP7_75t_L g752 ( .A(n_109), .B(n_448), .Y(n_752) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
OA21x2_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_121), .B(n_453), .Y(n_115) );
INVx1_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
INVx1_ASAP7_75t_SL g117 ( .A(n_118), .Y(n_117) );
BUFx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_L g756 ( .A(n_120), .Y(n_756) );
OAI21x1_ASAP7_75t_SL g121 ( .A1(n_122), .A2(n_444), .B(n_451), .Y(n_121) );
OAI22xp5_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_125), .B1(n_131), .B2(n_132), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_125), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_127), .Y(n_126) );
OAI22xp5_ASAP7_75t_SL g465 ( .A1(n_131), .A2(n_466), .B1(n_469), .B2(n_749), .Y(n_465) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
OAI22xp5_ASAP7_75t_SL g753 ( .A1(n_132), .A2(n_466), .B1(n_754), .B2(n_755), .Y(n_753) );
AND3x1_ASAP7_75t_L g132 ( .A(n_133), .B(n_369), .C(n_418), .Y(n_132) );
NOR3xp33_ASAP7_75t_SL g133 ( .A(n_134), .B(n_276), .C(n_314), .Y(n_133) );
OAI222xp33_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_197), .B1(n_251), .B2(n_257), .C1(n_271), .C2(n_274), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_136), .B(n_168), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_136), .B(n_344), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_136), .B(n_319), .Y(n_410) );
BUFx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
OR2x2_ASAP7_75t_L g287 ( .A(n_137), .B(n_188), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_137), .B(n_169), .Y(n_295) );
AND2x2_ASAP7_75t_L g330 ( .A(n_137), .B(n_307), .Y(n_330) );
OR2x2_ASAP7_75t_L g354 ( .A(n_137), .B(n_169), .Y(n_354) );
OR2x2_ASAP7_75t_L g362 ( .A(n_137), .B(n_261), .Y(n_362) );
AND2x2_ASAP7_75t_L g365 ( .A(n_137), .B(n_188), .Y(n_365) );
INVx3_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
OR2x2_ASAP7_75t_L g259 ( .A(n_138), .B(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g273 ( .A(n_138), .B(n_188), .Y(n_273) );
AND2x2_ASAP7_75t_L g323 ( .A(n_138), .B(n_261), .Y(n_323) );
AND2x2_ASAP7_75t_L g336 ( .A(n_138), .B(n_169), .Y(n_336) );
NOR2xp33_ASAP7_75t_L g443 ( .A(n_138), .B(n_422), .Y(n_443) );
AO21x2_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_145), .B(n_166), .Y(n_138) );
NOR2xp33_ASAP7_75t_L g166 ( .A(n_139), .B(n_167), .Y(n_166) );
INVx2_ASAP7_75t_L g211 ( .A(n_139), .Y(n_211) );
AO21x2_ASAP7_75t_L g261 ( .A1(n_139), .A2(n_262), .B(n_269), .Y(n_261) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_140), .Y(n_172) );
AND2x2_ASAP7_75t_L g140 ( .A(n_141), .B(n_142), .Y(n_140) );
AND2x2_ASAP7_75t_SL g187 ( .A(n_141), .B(n_142), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_143), .B(n_144), .Y(n_142) );
OAI22xp33_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_149), .B1(n_162), .B2(n_163), .Y(n_145) );
O2A1O1Ixp33_ASAP7_75t_L g175 ( .A1(n_146), .A2(n_176), .B(n_177), .C(n_178), .Y(n_175) );
O2A1O1Ixp33_ASAP7_75t_L g190 ( .A1(n_146), .A2(n_177), .B(n_191), .C(n_192), .Y(n_190) );
O2A1O1Ixp33_ASAP7_75t_L g243 ( .A1(n_146), .A2(n_177), .B(n_244), .C(n_245), .Y(n_243) );
INVx4_ASAP7_75t_SL g146 ( .A(n_147), .Y(n_146) );
NAND2x1p5_ASAP7_75t_L g163 ( .A(n_147), .B(n_164), .Y(n_163) );
AND2x4_ASAP7_75t_L g174 ( .A(n_147), .B(n_164), .Y(n_174) );
OAI21xp5_ASAP7_75t_L g477 ( .A1(n_147), .A2(n_478), .B(n_481), .Y(n_477) );
BUFx3_ASAP7_75t_L g497 ( .A(n_147), .Y(n_497) );
OAI21xp5_ASAP7_75t_L g503 ( .A1(n_147), .A2(n_504), .B(n_508), .Y(n_503) );
OAI21xp5_ASAP7_75t_L g524 ( .A1(n_147), .A2(n_525), .B(n_528), .Y(n_524) );
OAI21xp5_ASAP7_75t_L g540 ( .A1(n_147), .A2(n_541), .B(n_545), .Y(n_540) );
INVx2_ASAP7_75t_L g268 ( .A(n_150), .Y(n_268) );
INVx3_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g160 ( .A(n_152), .Y(n_160) );
INVx1_ASAP7_75t_L g165 ( .A(n_152), .Y(n_165) );
OAI22xp5_ASAP7_75t_SL g153 ( .A1(n_154), .A2(n_156), .B1(n_157), .B2(n_158), .Y(n_153) );
INVx2_ASAP7_75t_L g157 ( .A(n_154), .Y(n_157) );
INVx4_ASAP7_75t_L g246 ( .A(n_154), .Y(n_246) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx1_ASAP7_75t_L g161 ( .A(n_155), .Y(n_161) );
AND2x2_ASAP7_75t_L g164 ( .A(n_155), .B(n_165), .Y(n_164) );
BUFx6f_ASAP7_75t_L g180 ( .A(n_155), .Y(n_180) );
INVx3_ASAP7_75t_L g183 ( .A(n_155), .Y(n_183) );
INVx1_ASAP7_75t_L g193 ( .A(n_155), .Y(n_193) );
INVx5_ASAP7_75t_L g177 ( .A(n_159), .Y(n_177) );
AND2x6_ASAP7_75t_L g159 ( .A(n_160), .B(n_161), .Y(n_159) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_160), .Y(n_185) );
BUFx3_ASAP7_75t_L g210 ( .A(n_160), .Y(n_210) );
INVx1_ASAP7_75t_L g537 ( .A(n_160), .Y(n_537) );
OAI21xp5_ASAP7_75t_L g215 ( .A1(n_163), .A2(n_216), .B(n_217), .Y(n_215) );
OAI21xp5_ASAP7_75t_L g262 ( .A1(n_163), .A2(n_263), .B(n_264), .Y(n_262) );
INVx1_ASAP7_75t_L g484 ( .A(n_165), .Y(n_484) );
O2A1O1Ixp33_ASAP7_75t_L g361 ( .A1(n_168), .A2(n_362), .B(n_363), .C(n_366), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_168), .B(n_391), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_168), .B(n_306), .Y(n_428) );
AND2x2_ASAP7_75t_L g168 ( .A(n_169), .B(n_188), .Y(n_168) );
AND2x2_ASAP7_75t_SL g272 ( .A(n_169), .B(n_273), .Y(n_272) );
INVx2_ASAP7_75t_L g286 ( .A(n_169), .Y(n_286) );
AND2x2_ASAP7_75t_L g313 ( .A(n_169), .B(n_307), .Y(n_313) );
INVx1_ASAP7_75t_SL g321 ( .A(n_169), .Y(n_321) );
AND2x2_ASAP7_75t_L g344 ( .A(n_169), .B(n_345), .Y(n_344) );
BUFx2_ASAP7_75t_L g422 ( .A(n_169), .Y(n_422) );
OA21x2_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_173), .B(n_186), .Y(n_169) );
INVx3_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
NOR2xp33_ASAP7_75t_SL g212 ( .A(n_171), .B(n_213), .Y(n_212) );
NAND3xp33_ASAP7_75t_L g515 ( .A(n_171), .B(n_497), .C(n_516), .Y(n_515) );
AO21x1_ASAP7_75t_L g560 ( .A1(n_171), .A2(n_516), .B(n_561), .Y(n_560) );
INVx4_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
OA21x2_ASAP7_75t_L g188 ( .A1(n_172), .A2(n_189), .B(n_196), .Y(n_188) );
OA21x2_ASAP7_75t_L g476 ( .A1(n_172), .A2(n_477), .B(n_486), .Y(n_476) );
BUFx2_ASAP7_75t_L g242 ( .A(n_174), .Y(n_242) );
O2A1O1Ixp5_ASAP7_75t_L g493 ( .A1(n_179), .A2(n_494), .B(n_495), .C(n_496), .Y(n_493) );
AOI21xp5_ASAP7_75t_L g545 ( .A1(n_179), .A2(n_546), .B(n_547), .Y(n_545) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx4_ASAP7_75t_L g234 ( .A(n_180), .Y(n_234) );
OAI22xp5_ASAP7_75t_L g516 ( .A1(n_180), .A2(n_485), .B1(n_517), .B2(n_518), .Y(n_516) );
OAI22xp5_ASAP7_75t_L g535 ( .A1(n_180), .A2(n_485), .B1(n_536), .B2(n_538), .Y(n_535) );
OAI22xp5_ASAP7_75t_SL g555 ( .A1(n_180), .A2(n_183), .B1(n_556), .B2(n_557), .Y(n_555) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_182), .B(n_183), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_183), .B(n_195), .Y(n_194) );
INVx5_ASAP7_75t_L g206 ( .A(n_183), .Y(n_206) );
O2A1O1Ixp5_ASAP7_75t_SL g525 ( .A1(n_184), .A2(n_206), .B(n_526), .C(n_527), .Y(n_525) );
INVx3_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
HB1xp67_ASAP7_75t_L g235 ( .A(n_185), .Y(n_235) );
INVx1_ASAP7_75t_L g224 ( .A(n_187), .Y(n_224) );
INVx2_ASAP7_75t_L g228 ( .A(n_187), .Y(n_228) );
OA21x2_ASAP7_75t_L g240 ( .A1(n_187), .A2(n_241), .B(n_250), .Y(n_240) );
OA21x2_ASAP7_75t_L g523 ( .A1(n_187), .A2(n_524), .B(n_531), .Y(n_523) );
OA21x2_ASAP7_75t_L g539 ( .A1(n_187), .A2(n_540), .B(n_548), .Y(n_539) );
BUFx2_ASAP7_75t_L g258 ( .A(n_188), .Y(n_258) );
INVx1_ASAP7_75t_L g320 ( .A(n_188), .Y(n_320) );
INVx3_ASAP7_75t_L g345 ( .A(n_188), .Y(n_345) );
INVx1_ASAP7_75t_L g544 ( .A(n_193), .Y(n_544) );
NAND2xp5_ASAP7_75t_SL g278 ( .A(n_197), .B(n_279), .Y(n_278) );
OR2x2_ASAP7_75t_L g197 ( .A(n_198), .B(n_225), .Y(n_197) );
INVx1_ASAP7_75t_L g341 ( .A(n_198), .Y(n_341) );
OAI32xp33_ASAP7_75t_L g347 ( .A1(n_198), .A2(n_286), .A3(n_348), .B1(n_349), .B2(n_350), .Y(n_347) );
OAI22xp5_ASAP7_75t_L g351 ( .A1(n_198), .A2(n_352), .B1(n_355), .B2(n_360), .Y(n_351) );
INVx4_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
AND2x2_ASAP7_75t_L g289 ( .A(n_199), .B(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g367 ( .A(n_199), .B(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g437 ( .A(n_199), .B(n_383), .Y(n_437) );
AND2x2_ASAP7_75t_L g199 ( .A(n_200), .B(n_214), .Y(n_199) );
AND2x2_ASAP7_75t_L g252 ( .A(n_200), .B(n_253), .Y(n_252) );
INVx2_ASAP7_75t_L g282 ( .A(n_200), .Y(n_282) );
INVx1_ASAP7_75t_L g301 ( .A(n_200), .Y(n_301) );
OR2x2_ASAP7_75t_L g309 ( .A(n_200), .B(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g316 ( .A(n_200), .B(n_290), .Y(n_316) );
NOR2xp33_ASAP7_75t_L g324 ( .A(n_200), .B(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g337 ( .A(n_200), .B(n_255), .Y(n_337) );
INVx3_ASAP7_75t_L g359 ( .A(n_200), .Y(n_359) );
AND2x2_ASAP7_75t_L g384 ( .A(n_200), .B(n_256), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g432 ( .A(n_200), .B(n_349), .Y(n_432) );
OR2x6_ASAP7_75t_L g200 ( .A(n_201), .B(n_212), .Y(n_200) );
AOI21xp5_ASAP7_75t_SL g201 ( .A1(n_202), .A2(n_203), .B(n_211), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_207), .B(n_208), .Y(n_204) );
O2A1O1Ixp33_ASAP7_75t_L g265 ( .A1(n_206), .A2(n_266), .B(n_267), .C(n_268), .Y(n_265) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_206), .A2(n_479), .B(n_480), .Y(n_478) );
INVx2_ASAP7_75t_L g485 ( .A(n_206), .Y(n_485) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_206), .A2(n_491), .B(n_492), .Y(n_490) );
AOI21xp5_ASAP7_75t_L g218 ( .A1(n_208), .A2(n_219), .B(n_220), .Y(n_218) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
INVx1_ASAP7_75t_L g249 ( .A(n_210), .Y(n_249) );
INVx1_ASAP7_75t_L g221 ( .A(n_211), .Y(n_221) );
OA21x2_ASAP7_75t_L g488 ( .A1(n_211), .A2(n_489), .B(n_498), .Y(n_488) );
OA21x2_ASAP7_75t_L g502 ( .A1(n_211), .A2(n_503), .B(n_511), .Y(n_502) );
INVx2_ASAP7_75t_L g256 ( .A(n_214), .Y(n_256) );
AND2x2_ASAP7_75t_L g388 ( .A(n_214), .B(n_226), .Y(n_388) );
AO21x2_ASAP7_75t_L g214 ( .A1(n_215), .A2(n_221), .B(n_222), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_223), .B(n_224), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g237 ( .A(n_224), .B(n_238), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g269 ( .A(n_224), .B(n_270), .Y(n_269) );
INVx2_ASAP7_75t_L g430 ( .A(n_225), .Y(n_430) );
OR2x2_ASAP7_75t_L g225 ( .A(n_226), .B(n_239), .Y(n_225) );
INVx1_ASAP7_75t_L g275 ( .A(n_226), .Y(n_275) );
AND2x2_ASAP7_75t_L g302 ( .A(n_226), .B(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_226), .B(n_256), .Y(n_310) );
AND2x2_ASAP7_75t_L g368 ( .A(n_226), .B(n_291), .Y(n_368) );
INVx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVx1_ASAP7_75t_L g254 ( .A(n_227), .Y(n_254) );
AND2x2_ASAP7_75t_L g281 ( .A(n_227), .B(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g290 ( .A(n_227), .B(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_227), .B(n_256), .Y(n_356) );
AO21x2_ASAP7_75t_L g227 ( .A1(n_228), .A2(n_229), .B(n_237), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_230), .B(n_236), .Y(n_229) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_233), .B(n_235), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_239), .B(n_284), .Y(n_283) );
INVx2_ASAP7_75t_L g303 ( .A(n_239), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_239), .B(n_256), .Y(n_349) );
AND2x2_ASAP7_75t_L g358 ( .A(n_239), .B(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g383 ( .A(n_239), .Y(n_383) );
INVx2_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_L g255 ( .A(n_240), .B(n_256), .Y(n_255) );
INVx1_ASAP7_75t_L g291 ( .A(n_240), .Y(n_291) );
NOR2xp33_ASAP7_75t_L g247 ( .A(n_246), .B(n_248), .Y(n_247) );
INVx1_ASAP7_75t_L g507 ( .A(n_246), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_246), .A2(n_529), .B(n_530), .Y(n_528) );
OAI22xp5_ASAP7_75t_L g419 ( .A1(n_251), .A2(n_261), .B1(n_420), .B2(n_423), .Y(n_419) );
INVx1_ASAP7_75t_SL g251 ( .A(n_252), .Y(n_251) );
OAI21xp5_ASAP7_75t_SL g442 ( .A1(n_253), .A2(n_364), .B(n_443), .Y(n_442) );
AND2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g376 ( .A(n_254), .B(n_359), .Y(n_376) );
INVx1_ASAP7_75t_L g401 ( .A(n_254), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_255), .B(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g328 ( .A(n_255), .B(n_281), .Y(n_328) );
INVx2_ASAP7_75t_L g284 ( .A(n_256), .Y(n_284) );
INVx1_ASAP7_75t_L g334 ( .A(n_256), .Y(n_334) );
OAI221xp5_ASAP7_75t_L g425 ( .A1(n_257), .A2(n_409), .B1(n_426), .B2(n_429), .C(n_431), .Y(n_425) );
OR2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
INVx1_ASAP7_75t_L g296 ( .A(n_258), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_258), .B(n_307), .Y(n_348) );
NOR2xp33_ASAP7_75t_L g317 ( .A(n_259), .B(n_318), .Y(n_317) );
OR2x2_ASAP7_75t_L g350 ( .A(n_259), .B(n_296), .Y(n_350) );
INVx3_ASAP7_75t_SL g391 ( .A(n_259), .Y(n_391) );
AND2x2_ASAP7_75t_L g335 ( .A(n_260), .B(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g364 ( .A(n_260), .B(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_260), .B(n_273), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_260), .B(n_319), .Y(n_405) );
INVx3_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVx3_ASAP7_75t_L g307 ( .A(n_261), .Y(n_307) );
OAI322xp33_ASAP7_75t_L g402 ( .A1(n_261), .A2(n_333), .A3(n_355), .B1(n_403), .B2(n_405), .C1(n_406), .C2(n_407), .Y(n_402) );
O2A1O1Ixp33_ASAP7_75t_L g504 ( .A1(n_268), .A2(n_505), .B(n_506), .C(n_507), .Y(n_504) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AOI21xp33_ASAP7_75t_L g426 ( .A1(n_272), .A2(n_275), .B(n_427), .Y(n_426) );
NOR2xp33_ASAP7_75t_SL g352 ( .A(n_273), .B(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g374 ( .A(n_273), .B(n_286), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_273), .B(n_313), .Y(n_389) );
INVxp67_ASAP7_75t_L g340 ( .A(n_275), .Y(n_340) );
AOI211xp5_ASAP7_75t_L g346 ( .A1(n_275), .A2(n_347), .B(n_351), .C(n_361), .Y(n_346) );
OAI221xp5_ASAP7_75t_SL g276 ( .A1(n_277), .A2(n_285), .B1(n_288), .B2(n_292), .C(n_297), .Y(n_276) );
INVxp67_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
OR2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_283), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g300 ( .A(n_284), .B(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g417 ( .A(n_284), .Y(n_417) );
OAI221xp5_ASAP7_75t_L g433 ( .A1(n_285), .A2(n_434), .B1(n_439), .B2(n_440), .C(n_442), .Y(n_433) );
OR2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_286), .B(n_330), .Y(n_329) );
INVx1_ASAP7_75t_SL g333 ( .A(n_286), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_286), .B(n_364), .Y(n_371) );
AND2x2_ASAP7_75t_L g413 ( .A(n_286), .B(n_391), .Y(n_413) );
NOR2xp33_ASAP7_75t_L g311 ( .A(n_287), .B(n_312), .Y(n_311) );
OAI22xp33_ASAP7_75t_L g408 ( .A1(n_287), .A2(n_299), .B1(n_409), .B2(n_410), .Y(n_408) );
OR2x2_ASAP7_75t_L g439 ( .A(n_287), .B(n_307), .Y(n_439) );
CKINVDCx16_ASAP7_75t_R g288 ( .A(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g416 ( .A(n_290), .Y(n_416) );
AND2x2_ASAP7_75t_L g441 ( .A(n_290), .B(n_384), .Y(n_441) );
INVxp67_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
NOR2xp33_ASAP7_75t_SL g293 ( .A(n_294), .B(n_296), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
OR2x2_ASAP7_75t_L g305 ( .A(n_295), .B(n_306), .Y(n_305) );
AOI22xp5_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_304), .B1(n_308), .B2(n_311), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_300), .B(n_302), .Y(n_299) );
INVx1_ASAP7_75t_L g372 ( .A(n_300), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_300), .B(n_340), .Y(n_407) );
AOI322xp5_ASAP7_75t_L g331 ( .A1(n_302), .A2(n_332), .A3(n_334), .B1(n_335), .B2(n_337), .C1(n_338), .C2(n_342), .Y(n_331) );
INVxp67_ASAP7_75t_L g325 ( .A(n_303), .Y(n_325) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
OAI22xp5_ASAP7_75t_L g326 ( .A1(n_305), .A2(n_310), .B1(n_327), .B2(n_329), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_306), .B(n_319), .Y(n_406) );
INVx1_ASAP7_75t_SL g306 ( .A(n_307), .Y(n_306) );
NOR2xp33_ASAP7_75t_L g415 ( .A(n_307), .B(n_345), .Y(n_415) );
NOR2xp33_ASAP7_75t_L g421 ( .A(n_307), .B(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
OR2x2_ASAP7_75t_L g403 ( .A(n_309), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_SL g312 ( .A(n_313), .Y(n_312) );
NAND3xp33_ASAP7_75t_SL g314 ( .A(n_315), .B(n_331), .C(n_346), .Y(n_314) );
AOI221xp5_ASAP7_75t_L g315 ( .A1(n_316), .A2(n_317), .B1(n_322), .B2(n_324), .C(n_326), .Y(n_315) );
AND2x2_ASAP7_75t_L g322 ( .A(n_318), .B(n_323), .Y(n_322) );
INVx3_ASAP7_75t_SL g318 ( .A(n_319), .Y(n_318) );
AND2x4_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
AND2x2_ASAP7_75t_L g332 ( .A(n_323), .B(n_333), .Y(n_332) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_325), .Y(n_404) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_330), .B(n_344), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_333), .B(n_391), .Y(n_397) );
NOR2xp33_ASAP7_75t_L g393 ( .A(n_334), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_SL g409 ( .A(n_337), .Y(n_409) );
AND2x2_ASAP7_75t_L g424 ( .A(n_337), .B(n_401), .Y(n_424) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
AOI211xp5_ASAP7_75t_L g418 ( .A1(n_348), .A2(n_419), .B(n_425), .C(n_433), .Y(n_418) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
OR2x2_ASAP7_75t_L g355 ( .A(n_356), .B(n_357), .Y(n_355) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g387 ( .A(n_358), .B(n_388), .Y(n_387) );
NAND2x1_ASAP7_75t_SL g429 ( .A(n_359), .B(n_430), .Y(n_429) );
CKINVDCx16_ASAP7_75t_R g399 ( .A(n_362), .Y(n_399) );
INVx1_ASAP7_75t_SL g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g394 ( .A(n_368), .Y(n_394) );
AND2x2_ASAP7_75t_L g398 ( .A(n_368), .B(n_384), .Y(n_398) );
NOR5xp2_ASAP7_75t_L g369 ( .A(n_370), .B(n_385), .C(n_402), .D(n_408), .E(n_411), .Y(n_369) );
OAI221xp5_ASAP7_75t_L g370 ( .A1(n_371), .A2(n_372), .B1(n_373), .B2(n_375), .C(n_377), .Y(n_370) );
INVx2_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_374), .B(n_432), .Y(n_431) );
INVxp67_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_378), .B(n_380), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_382), .B(n_384), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
AND2x2_ASAP7_75t_L g400 ( .A(n_384), .B(n_401), .Y(n_400) );
OAI221xp5_ASAP7_75t_SL g385 ( .A1(n_386), .A2(n_389), .B1(n_390), .B2(n_392), .C(n_395), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
AOI22xp33_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_398), .B1(n_399), .B2(n_400), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g438 ( .A(n_398), .Y(n_438) );
AOI211xp5_ASAP7_75t_SL g411 ( .A1(n_412), .A2(n_414), .B(n_416), .C(n_417), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVxp67_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_436), .B(n_438), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
CKINVDCx14_ASAP7_75t_R g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_SL g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_SL g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g452 ( .A(n_447), .Y(n_452) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
NAND3xp33_ASAP7_75t_L g453 ( .A(n_451), .B(n_454), .C(n_756), .Y(n_453) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
CKINVDCx14_ASAP7_75t_R g460 ( .A(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g754 ( .A(n_469), .Y(n_754) );
NAND2x1p5_ASAP7_75t_L g469 ( .A(n_470), .B(n_673), .Y(n_469) );
AND2x2_ASAP7_75t_SL g470 ( .A(n_471), .B(n_631), .Y(n_470) );
NOR4xp25_ASAP7_75t_L g471 ( .A(n_472), .B(n_571), .C(n_607), .D(n_621), .Y(n_471) );
OAI221xp5_ASAP7_75t_SL g472 ( .A1(n_473), .A2(n_519), .B1(n_549), .B2(n_558), .C(n_562), .Y(n_472) );
NAND2xp5_ASAP7_75t_SL g705 ( .A(n_473), .B(n_706), .Y(n_705) );
OR2x2_ASAP7_75t_L g473 ( .A(n_474), .B(n_499), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_476), .B(n_487), .Y(n_475) );
AND2x2_ASAP7_75t_L g568 ( .A(n_476), .B(n_488), .Y(n_568) );
INVx3_ASAP7_75t_L g576 ( .A(n_476), .Y(n_576) );
AND2x2_ASAP7_75t_L g630 ( .A(n_476), .B(n_502), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_476), .B(n_501), .Y(n_666) );
AND2x2_ASAP7_75t_L g724 ( .A(n_476), .B(n_586), .Y(n_724) );
AOI21xp5_ASAP7_75t_L g481 ( .A1(n_482), .A2(n_483), .B(n_485), .Y(n_481) );
INVx2_ASAP7_75t_L g495 ( .A(n_484), .Y(n_495) );
O2A1O1Ixp33_ASAP7_75t_L g508 ( .A1(n_485), .A2(n_495), .B(n_509), .C(n_510), .Y(n_508) );
AND2x2_ASAP7_75t_L g559 ( .A(n_487), .B(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g573 ( .A(n_487), .B(n_502), .Y(n_573) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_488), .B(n_502), .Y(n_588) );
AND2x2_ASAP7_75t_L g600 ( .A(n_488), .B(n_576), .Y(n_600) );
OR2x2_ASAP7_75t_L g602 ( .A(n_488), .B(n_560), .Y(n_602) );
AND2x2_ASAP7_75t_L g637 ( .A(n_488), .B(n_560), .Y(n_637) );
HB1xp67_ASAP7_75t_L g682 ( .A(n_488), .Y(n_682) );
INVx1_ASAP7_75t_L g690 ( .A(n_488), .Y(n_690) );
OAI21xp5_ASAP7_75t_L g489 ( .A1(n_490), .A2(n_493), .B(n_497), .Y(n_489) );
OAI221xp5_ASAP7_75t_L g607 ( .A1(n_499), .A2(n_608), .B1(n_612), .B2(n_616), .C(n_617), .Y(n_607) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
AND2x2_ASAP7_75t_L g567 ( .A(n_500), .B(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g500 ( .A(n_501), .B(n_512), .Y(n_500) );
INVx2_ASAP7_75t_L g566 ( .A(n_501), .Y(n_566) );
AND2x2_ASAP7_75t_L g619 ( .A(n_501), .B(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g638 ( .A(n_501), .B(n_576), .Y(n_638) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
AND2x2_ASAP7_75t_L g701 ( .A(n_502), .B(n_576), .Y(n_701) );
AND2x2_ASAP7_75t_L g623 ( .A(n_512), .B(n_568), .Y(n_623) );
OAI322xp33_ASAP7_75t_L g691 ( .A1(n_512), .A2(n_647), .A3(n_692), .B1(n_694), .B2(n_697), .C1(n_699), .C2(n_703), .Y(n_691) );
INVx3_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
NOR2x1_ASAP7_75t_L g574 ( .A(n_513), .B(n_575), .Y(n_574) );
INVx2_ASAP7_75t_L g587 ( .A(n_513), .Y(n_587) );
AND2x2_ASAP7_75t_L g696 ( .A(n_513), .B(n_576), .Y(n_696) );
AND2x2_ASAP7_75t_L g728 ( .A(n_513), .B(n_600), .Y(n_728) );
OR2x2_ASAP7_75t_L g731 ( .A(n_513), .B(n_732), .Y(n_731) );
AND2x4_ASAP7_75t_L g513 ( .A(n_514), .B(n_515), .Y(n_513) );
INVx1_ASAP7_75t_L g561 ( .A(n_514), .Y(n_561) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_532), .Y(n_520) );
INVx1_ASAP7_75t_L g744 ( .A(n_521), .Y(n_744) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
OR2x2_ASAP7_75t_L g551 ( .A(n_522), .B(n_539), .Y(n_551) );
INVx2_ASAP7_75t_L g584 ( .A(n_522), .Y(n_584) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx2_ASAP7_75t_L g606 ( .A(n_523), .Y(n_606) );
HB1xp67_ASAP7_75t_L g614 ( .A(n_523), .Y(n_614) );
OR2x2_ASAP7_75t_L g738 ( .A(n_523), .B(n_739), .Y(n_738) );
AND2x2_ASAP7_75t_L g563 ( .A(n_532), .B(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g603 ( .A(n_532), .B(n_604), .Y(n_603) );
AND2x2_ASAP7_75t_L g655 ( .A(n_532), .B(n_656), .Y(n_655) );
AND2x2_ASAP7_75t_L g532 ( .A(n_533), .B(n_539), .Y(n_532) );
AND2x2_ASAP7_75t_L g552 ( .A(n_533), .B(n_553), .Y(n_552) );
NOR2xp67_ASAP7_75t_L g610 ( .A(n_533), .B(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g664 ( .A(n_533), .B(n_554), .Y(n_664) );
OR2x2_ASAP7_75t_L g672 ( .A(n_533), .B(n_606), .Y(n_672) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
BUFx2_ASAP7_75t_L g581 ( .A(n_534), .Y(n_581) );
AND2x2_ASAP7_75t_L g591 ( .A(n_534), .B(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g615 ( .A(n_534), .B(n_539), .Y(n_615) );
AND2x2_ASAP7_75t_L g679 ( .A(n_534), .B(n_554), .Y(n_679) );
NOR2xp33_ASAP7_75t_L g569 ( .A(n_539), .B(n_570), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_539), .B(n_584), .Y(n_583) );
INVx2_ASAP7_75t_L g592 ( .A(n_539), .Y(n_592) );
INVx1_ASAP7_75t_L g597 ( .A(n_539), .Y(n_597) );
AND2x2_ASAP7_75t_L g609 ( .A(n_539), .B(n_610), .Y(n_609) );
HB1xp67_ASAP7_75t_L g687 ( .A(n_539), .Y(n_687) );
INVx1_ASAP7_75t_L g739 ( .A(n_539), .Y(n_739) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_542), .A2(n_543), .B(n_544), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_550), .B(n_552), .Y(n_549) );
AND2x2_ASAP7_75t_L g716 ( .A(n_550), .B(n_625), .Y(n_716) );
INVx2_ASAP7_75t_SL g550 ( .A(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g643 ( .A(n_552), .B(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g742 ( .A(n_552), .B(n_677), .Y(n_742) );
INVx1_ASAP7_75t_L g564 ( .A(n_553), .Y(n_564) );
AND2x2_ASAP7_75t_L g590 ( .A(n_553), .B(n_584), .Y(n_590) );
BUFx2_ASAP7_75t_L g649 ( .A(n_553), .Y(n_649) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
BUFx6f_ASAP7_75t_L g570 ( .A(n_554), .Y(n_570) );
INVx1_ASAP7_75t_L g580 ( .A(n_554), .Y(n_580) );
NOR2xp67_ASAP7_75t_L g718 ( .A(n_558), .B(n_565), .Y(n_718) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
AOI32xp33_ASAP7_75t_L g562 ( .A1(n_559), .A2(n_563), .A3(n_565), .B1(n_567), .B2(n_569), .Y(n_562) );
AND2x2_ASAP7_75t_L g702 ( .A(n_559), .B(n_575), .Y(n_702) );
AND2x2_ASAP7_75t_L g740 ( .A(n_559), .B(n_638), .Y(n_740) );
INVx1_ASAP7_75t_L g620 ( .A(n_560), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_564), .B(n_626), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_565), .B(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_565), .B(n_568), .Y(n_616) );
NAND2xp5_ASAP7_75t_SL g719 ( .A(n_565), .B(n_637), .Y(n_719) );
OR2x2_ASAP7_75t_L g733 ( .A(n_565), .B(n_602), .Y(n_733) );
INVx3_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g660 ( .A(n_566), .B(n_568), .Y(n_660) );
OR2x2_ASAP7_75t_L g669 ( .A(n_566), .B(n_656), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_568), .B(n_619), .Y(n_641) );
INVx2_ASAP7_75t_L g656 ( .A(n_570), .Y(n_656) );
OR2x2_ASAP7_75t_L g671 ( .A(n_570), .B(n_672), .Y(n_671) );
AND2x2_ASAP7_75t_L g686 ( .A(n_570), .B(n_687), .Y(n_686) );
A2O1A1Ixp33_ASAP7_75t_L g743 ( .A1(n_570), .A2(n_663), .B(n_744), .C(n_745), .Y(n_743) );
OAI321xp33_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_577), .A3(n_582), .B1(n_585), .B2(n_589), .C(n_593), .Y(n_571) );
INVx1_ASAP7_75t_L g684 ( .A(n_572), .Y(n_684) );
NAND2x1p5_ASAP7_75t_L g572 ( .A(n_573), .B(n_574), .Y(n_572) );
AND2x2_ASAP7_75t_L g695 ( .A(n_573), .B(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g647 ( .A(n_575), .Y(n_647) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_576), .B(n_690), .Y(n_707) );
OAI221xp5_ASAP7_75t_L g714 ( .A1(n_577), .A2(n_715), .B1(n_717), .B2(n_719), .C(n_720), .Y(n_714) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_581), .Y(n_578) );
AND2x2_ASAP7_75t_L g652 ( .A(n_579), .B(n_626), .Y(n_652) );
HB1xp67_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_580), .B(n_606), .Y(n_605) );
INVx2_ASAP7_75t_L g625 ( .A(n_581), .Y(n_625) );
A2O1A1Ixp33_ASAP7_75t_L g667 ( .A1(n_582), .A2(n_623), .B(n_668), .C(n_670), .Y(n_667) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g634 ( .A(n_584), .B(n_591), .Y(n_634) );
BUFx2_ASAP7_75t_L g644 ( .A(n_584), .Y(n_644) );
INVx1_ASAP7_75t_L g659 ( .A(n_584), .Y(n_659) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
NOR2xp33_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
OR2x2_ASAP7_75t_L g665 ( .A(n_587), .B(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g748 ( .A(n_587), .Y(n_748) );
INVx1_ASAP7_75t_L g741 ( .A(n_588), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
AND2x2_ASAP7_75t_L g594 ( .A(n_590), .B(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g698 ( .A(n_590), .B(n_615), .Y(n_698) );
INVx1_ASAP7_75t_L g627 ( .A(n_591), .Y(n_627) );
AOI22xp5_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_598), .B1(n_601), .B2(n_603), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_595), .B(n_711), .Y(n_710) );
INVxp67_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
AND2x4_ASAP7_75t_L g663 ( .A(n_596), .B(n_664), .Y(n_663) );
BUFx3_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_SL g626 ( .A(n_597), .B(n_606), .Y(n_626) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g618 ( .A(n_600), .B(n_619), .Y(n_618) );
INVx1_ASAP7_75t_SL g601 ( .A(n_602), .Y(n_601) );
OR2x2_ASAP7_75t_L g628 ( .A(n_602), .B(n_629), .Y(n_628) );
INVx1_ASAP7_75t_SL g604 ( .A(n_605), .Y(n_604) );
OAI221xp5_ASAP7_75t_L g722 ( .A1(n_605), .A2(n_723), .B1(n_725), .B2(n_726), .C(n_727), .Y(n_722) );
INVx1_ASAP7_75t_L g611 ( .A(n_606), .Y(n_611) );
HB1xp67_ASAP7_75t_L g677 ( .A(n_606), .Y(n_677) );
INVx1_ASAP7_75t_SL g608 ( .A(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_609), .B(n_728), .Y(n_727) );
OAI21xp5_ASAP7_75t_L g617 ( .A1(n_610), .A2(n_615), .B(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_613), .B(n_623), .Y(n_720) );
AND2x2_ASAP7_75t_L g613 ( .A(n_614), .B(n_615), .Y(n_613) );
INVx1_ASAP7_75t_L g689 ( .A(n_614), .Y(n_689) );
AND2x2_ASAP7_75t_L g648 ( .A(n_615), .B(n_649), .Y(n_648) );
INVx2_ASAP7_75t_L g737 ( .A(n_615), .Y(n_737) );
INVx1_ASAP7_75t_L g653 ( .A(n_618), .Y(n_653) );
INVx1_ASAP7_75t_L g708 ( .A(n_619), .Y(n_708) );
OAI22xp5_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_624), .B1(n_627), .B2(n_628), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_625), .B(n_626), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_625), .B(n_659), .Y(n_658) );
INVx2_ASAP7_75t_L g693 ( .A(n_626), .Y(n_693) );
NAND2xp5_ASAP7_75t_SL g730 ( .A(n_626), .B(n_664), .Y(n_730) );
OR2x2_ASAP7_75t_L g703 ( .A(n_627), .B(n_656), .Y(n_703) );
INVx1_ASAP7_75t_L g642 ( .A(n_628), .Y(n_642) );
INVx1_ASAP7_75t_SL g629 ( .A(n_630), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_630), .B(n_681), .Y(n_680) );
NOR3xp33_ASAP7_75t_L g631 ( .A(n_632), .B(n_650), .C(n_661), .Y(n_631) );
OAI211xp5_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_635), .B(n_639), .C(n_645), .Y(n_632) );
INVxp67_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
AOI221xp5_ASAP7_75t_L g704 ( .A1(n_634), .A2(n_705), .B1(n_709), .B2(n_712), .C(n_714), .Y(n_704) );
INVx1_ASAP7_75t_SL g635 ( .A(n_636), .Y(n_635) );
AND2x2_ASAP7_75t_L g636 ( .A(n_637), .B(n_638), .Y(n_636) );
AND2x2_ASAP7_75t_L g646 ( .A(n_637), .B(n_647), .Y(n_646) );
AND2x2_ASAP7_75t_L g700 ( .A(n_637), .B(n_701), .Y(n_700) );
OAI211xp5_ASAP7_75t_L g685 ( .A1(n_638), .A2(n_686), .B(n_688), .C(n_690), .Y(n_685) );
INVx2_ASAP7_75t_L g732 ( .A(n_638), .Y(n_732) );
OAI21xp5_ASAP7_75t_SL g639 ( .A1(n_640), .A2(n_642), .B(n_643), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
AND2x2_ASAP7_75t_L g711 ( .A(n_644), .B(n_664), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_646), .B(n_648), .Y(n_645) );
OAI21xp5_ASAP7_75t_SL g650 ( .A1(n_651), .A2(n_653), .B(n_654), .Y(n_650) );
INVxp67_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
OAI21xp5_ASAP7_75t_SL g654 ( .A1(n_655), .A2(n_657), .B(n_660), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_655), .B(n_684), .Y(n_683) );
INVxp67_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_660), .B(n_747), .Y(n_746) );
OAI21xp33_ASAP7_75t_L g661 ( .A1(n_662), .A2(n_665), .B(n_667), .Y(n_661) );
INVx1_ASAP7_75t_SL g662 ( .A(n_663), .Y(n_662) );
AND2x2_ASAP7_75t_L g688 ( .A(n_664), .B(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
AND4x1_ASAP7_75t_L g673 ( .A(n_674), .B(n_704), .C(n_721), .D(n_743), .Y(n_673) );
NOR2xp33_ASAP7_75t_L g674 ( .A(n_675), .B(n_691), .Y(n_674) );
OAI211xp5_ASAP7_75t_SL g675 ( .A1(n_676), .A2(n_680), .B(n_683), .C(n_685), .Y(n_675) );
OR2x2_ASAP7_75t_L g676 ( .A(n_677), .B(n_678), .Y(n_676) );
INVx1_ASAP7_75t_SL g678 ( .A(n_679), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_679), .B(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
NOR2xp33_ASAP7_75t_L g712 ( .A(n_690), .B(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
NOR2xp33_ASAP7_75t_L g699 ( .A(n_700), .B(n_702), .Y(n_699) );
INVx1_ASAP7_75t_L g725 ( .A(n_700), .Y(n_725) );
INVx2_ASAP7_75t_SL g713 ( .A(n_701), .Y(n_713) );
OR2x2_ASAP7_75t_L g706 ( .A(n_707), .B(n_708), .Y(n_706) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g726 ( .A(n_711), .Y(n_726) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
NOR2xp33_ASAP7_75t_SL g721 ( .A(n_722), .B(n_729), .Y(n_721) );
INVx1_ASAP7_75t_SL g723 ( .A(n_724), .Y(n_723) );
OAI221xp5_ASAP7_75t_SL g729 ( .A1(n_730), .A2(n_731), .B1(n_733), .B2(n_734), .C(n_735), .Y(n_729) );
AOI22xp5_ASAP7_75t_L g735 ( .A1(n_736), .A2(n_740), .B1(n_741), .B2(n_742), .Y(n_735) );
NAND2xp5_ASAP7_75t_SL g736 ( .A(n_737), .B(n_738), .Y(n_736) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx2_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx2_ASAP7_75t_L g755 ( .A(n_750), .Y(n_755) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx1_ASAP7_75t_SL g757 ( .A(n_758), .Y(n_757) );
endmodule