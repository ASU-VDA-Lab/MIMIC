module real_aes_1733_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_635;
wire n_792;
wire n_386;
wire n_503;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_555;
wire n_364;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_537;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_527;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_789;
wire n_268;
wire n_544;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_809;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_797;
wire n_668;
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_0), .B(n_153), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_1), .A2(n_147), .B(n_195), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g120 ( .A(n_2), .B(n_121), .Y(n_120) );
NAND2xp5_ASAP7_75t_SL g239 ( .A(n_3), .B(n_164), .Y(n_239) );
INVx1_ASAP7_75t_L g152 ( .A(n_4), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_5), .B(n_164), .Y(n_203) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_6), .B(n_216), .Y(n_507) );
INVx1_ASAP7_75t_L g550 ( .A(n_7), .Y(n_550) );
CKINVDCx16_ASAP7_75t_R g121 ( .A(n_8), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g564 ( .A(n_9), .Y(n_564) );
NAND2xp33_ASAP7_75t_L g215 ( .A(n_10), .B(n_162), .Y(n_215) );
INVx2_ASAP7_75t_L g144 ( .A(n_11), .Y(n_144) );
AOI221x1_ASAP7_75t_L g146 ( .A1(n_12), .A2(n_24), .B1(n_147), .B2(n_153), .C(n_160), .Y(n_146) );
CKINVDCx16_ASAP7_75t_R g114 ( .A(n_13), .Y(n_114) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_14), .B(n_153), .Y(n_211) );
AO21x2_ASAP7_75t_L g208 ( .A1(n_15), .A2(n_209), .B(n_210), .Y(n_208) );
INVx1_ASAP7_75t_L g516 ( .A(n_16), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_17), .B(n_142), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_18), .B(n_164), .Y(n_223) );
AO21x1_ASAP7_75t_L g234 ( .A1(n_19), .A2(n_153), .B(n_235), .Y(n_234) );
INVx1_ASAP7_75t_L g118 ( .A(n_20), .Y(n_118) );
INVx1_ASAP7_75t_L g514 ( .A(n_21), .Y(n_514) );
INVx1_ASAP7_75t_SL g500 ( .A(n_22), .Y(n_500) );
NAND2xp5_ASAP7_75t_SL g478 ( .A(n_23), .B(n_154), .Y(n_478) );
NAND2x1_ASAP7_75t_L g172 ( .A(n_25), .B(n_164), .Y(n_172) );
AOI33xp33_ASAP7_75t_L g531 ( .A1(n_26), .A2(n_55), .A3(n_466), .B1(n_475), .B2(n_532), .B3(n_533), .Y(n_531) );
NAND2x1_ASAP7_75t_L g202 ( .A(n_27), .B(n_162), .Y(n_202) );
INVx1_ASAP7_75t_L g558 ( .A(n_28), .Y(n_558) );
OR2x2_ASAP7_75t_L g145 ( .A(n_29), .B(n_90), .Y(n_145) );
OA21x2_ASAP7_75t_L g178 ( .A1(n_29), .A2(n_90), .B(n_144), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_30), .B(n_491), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_31), .B(n_162), .Y(n_197) );
AOI22xp5_ASAP7_75t_L g793 ( .A1(n_32), .A2(n_33), .B1(n_794), .B2(n_795), .Y(n_793) );
CKINVDCx20_ASAP7_75t_R g794 ( .A(n_32), .Y(n_794) );
INVx1_ASAP7_75t_L g795 ( .A(n_33), .Y(n_795) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_34), .B(n_164), .Y(n_214) );
OAI22xp5_ASAP7_75t_SL g130 ( .A1(n_35), .A2(n_36), .B1(n_131), .B2(n_132), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g132 ( .A(n_35), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_36), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_37), .B(n_162), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g182 ( .A1(n_38), .A2(n_147), .B(n_183), .Y(n_182) );
AND2x2_ASAP7_75t_L g148 ( .A(n_39), .B(n_149), .Y(n_148) );
AND2x2_ASAP7_75t_L g159 ( .A(n_39), .B(n_152), .Y(n_159) );
INVx1_ASAP7_75t_L g474 ( .A(n_39), .Y(n_474) );
OR2x6_ASAP7_75t_L g116 ( .A(n_40), .B(n_117), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g560 ( .A(n_41), .Y(n_560) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_42), .B(n_153), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_43), .B(n_491), .Y(n_538) );
AOI221xp5_ASAP7_75t_L g103 ( .A1(n_44), .A2(n_104), .B1(n_122), .B2(n_446), .C(n_449), .Y(n_103) );
OAI22xp5_ASAP7_75t_SL g126 ( .A1(n_44), .A2(n_88), .B1(n_127), .B2(n_128), .Y(n_126) );
INVxp67_ASAP7_75t_L g127 ( .A(n_44), .Y(n_127) );
AOI22xp5_ASAP7_75t_L g462 ( .A1(n_44), .A2(n_177), .B1(n_216), .B2(n_463), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_45), .B(n_480), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_46), .B(n_154), .Y(n_501) );
CKINVDCx20_ASAP7_75t_R g227 ( .A(n_47), .Y(n_227) );
CKINVDCx20_ASAP7_75t_R g807 ( .A(n_48), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_49), .B(n_162), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g552 ( .A(n_50), .B(n_209), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_51), .B(n_154), .Y(n_551) );
AOI21xp5_ASAP7_75t_L g200 ( .A1(n_52), .A2(n_147), .B(n_201), .Y(n_200) );
CKINVDCx5p33_ASAP7_75t_R g470 ( .A(n_53), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_54), .B(n_162), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_56), .B(n_154), .Y(n_542) );
INVx1_ASAP7_75t_L g151 ( .A(n_57), .Y(n_151) );
INVx1_ASAP7_75t_L g156 ( .A(n_57), .Y(n_156) );
AND2x2_ASAP7_75t_L g543 ( .A(n_58), .B(n_142), .Y(n_543) );
AOI221xp5_ASAP7_75t_L g548 ( .A1(n_59), .A2(n_77), .B1(n_472), .B2(n_491), .C(n_549), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_60), .B(n_491), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_61), .B(n_164), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_62), .B(n_177), .Y(n_566) );
AOI21xp5_ASAP7_75t_SL g486 ( .A1(n_63), .A2(n_472), .B(n_487), .Y(n_486) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_64), .A2(n_147), .B(n_171), .Y(n_170) );
INVx1_ASAP7_75t_L g510 ( .A(n_65), .Y(n_510) );
AO21x1_ASAP7_75t_L g236 ( .A1(n_66), .A2(n_147), .B(n_237), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_67), .B(n_153), .Y(n_193) );
INVx1_ASAP7_75t_L g541 ( .A(n_68), .Y(n_541) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_69), .B(n_153), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g539 ( .A1(n_70), .A2(n_472), .B(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g187 ( .A(n_71), .B(n_143), .Y(n_187) );
INVx1_ASAP7_75t_L g149 ( .A(n_72), .Y(n_149) );
INVx1_ASAP7_75t_L g158 ( .A(n_72), .Y(n_158) );
AND2x2_ASAP7_75t_L g206 ( .A(n_73), .B(n_176), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_74), .B(n_491), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_75), .B(n_442), .Y(n_441) );
AOI22xp5_ASAP7_75t_L g788 ( .A1(n_76), .A2(n_789), .B1(n_790), .B2(n_791), .Y(n_788) );
CKINVDCx20_ASAP7_75t_R g789 ( .A(n_76), .Y(n_789) );
AND2x2_ASAP7_75t_L g502 ( .A(n_78), .B(n_176), .Y(n_502) );
INVx1_ASAP7_75t_L g511 ( .A(n_79), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_80), .A2(n_472), .B(n_499), .Y(n_498) );
OAI22xp5_ASAP7_75t_SL g791 ( .A1(n_81), .A2(n_792), .B1(n_793), .B2(n_796), .Y(n_791) );
CKINVDCx20_ASAP7_75t_R g796 ( .A(n_81), .Y(n_796) );
A2O1A1Ixp33_ASAP7_75t_L g471 ( .A1(n_82), .A2(n_472), .B(n_477), .C(n_482), .Y(n_471) );
INVx1_ASAP7_75t_L g119 ( .A(n_83), .Y(n_119) );
AND2x2_ASAP7_75t_L g191 ( .A(n_84), .B(n_176), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_85), .B(n_153), .Y(n_225) );
AND2x2_ASAP7_75t_SL g484 ( .A(n_86), .B(n_176), .Y(n_484) );
AOI22xp5_ASAP7_75t_L g528 ( .A1(n_87), .A2(n_472), .B1(n_529), .B2(n_530), .Y(n_528) );
INVx1_ASAP7_75t_L g128 ( .A(n_88), .Y(n_128) );
AND2x2_ASAP7_75t_L g235 ( .A(n_89), .B(n_216), .Y(n_235) );
AND2x2_ASAP7_75t_L g179 ( .A(n_91), .B(n_176), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_92), .B(n_162), .Y(n_224) );
INVx1_ASAP7_75t_L g488 ( .A(n_93), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_94), .B(n_164), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_95), .B(n_162), .Y(n_161) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_96), .A2(n_147), .B(n_222), .Y(n_221) );
AND2x2_ASAP7_75t_L g535 ( .A(n_97), .B(n_176), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_98), .B(n_164), .Y(n_196) );
A2O1A1Ixp33_ASAP7_75t_L g555 ( .A1(n_99), .A2(n_556), .B(n_557), .C(n_559), .Y(n_555) );
BUFx2_ASAP7_75t_SL g110 ( .A(n_100), .Y(n_110) );
BUFx2_ASAP7_75t_L g448 ( .A(n_100), .Y(n_448) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_101), .A2(n_147), .B(n_213), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_102), .B(n_154), .Y(n_489) );
INVx1_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
AOI21xp5_ASAP7_75t_L g107 ( .A1(n_108), .A2(n_111), .B(n_120), .Y(n_107) );
CKINVDCx11_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
CKINVDCx8_ASAP7_75t_R g109 ( .A(n_110), .Y(n_109) );
INVx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
BUFx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
BUFx2_ASAP7_75t_L g124 ( .A(n_113), .Y(n_124) );
BUFx3_ASAP7_75t_L g445 ( .A(n_113), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_114), .B(n_115), .Y(n_113) );
OR2x6_ASAP7_75t_SL g784 ( .A(n_114), .B(n_115), .Y(n_784) );
AND2x6_ASAP7_75t_SL g787 ( .A(n_114), .B(n_116), .Y(n_787) );
OR2x2_ASAP7_75t_L g808 ( .A(n_114), .B(n_116), .Y(n_808) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_116), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g117 ( .A(n_118), .B(n_119), .Y(n_117) );
OR2x2_ASAP7_75t_SL g447 ( .A(n_120), .B(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g814 ( .A(n_120), .Y(n_814) );
OAI21x1_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_125), .B(n_441), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
AND2x2_ASAP7_75t_L g811 ( .A(n_124), .B(n_812), .Y(n_811) );
AOI22xp33_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_129), .B1(n_439), .B2(n_440), .Y(n_125) );
INVx1_ASAP7_75t_L g439 ( .A(n_126), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_129), .Y(n_440) );
XOR2x1_ASAP7_75t_L g129 ( .A(n_130), .B(n_133), .Y(n_129) );
INVx3_ASAP7_75t_L g785 ( .A(n_133), .Y(n_785) );
OAI22xp5_ASAP7_75t_SL g799 ( .A1(n_133), .A2(n_800), .B1(n_802), .B2(n_803), .Y(n_799) );
AND2x4_ASAP7_75t_L g133 ( .A(n_134), .B(n_351), .Y(n_133) );
AND4x1_ASAP7_75t_L g134 ( .A(n_135), .B(n_263), .C(n_290), .D(n_325), .Y(n_134) );
AOI221xp5_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_188), .B1(n_228), .B2(n_243), .C(n_247), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_138), .B(n_167), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_138), .B(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
OR2x2_ASAP7_75t_L g304 ( .A(n_139), .B(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g359 ( .A(n_139), .B(n_314), .Y(n_359) );
BUFx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
AND2x2_ASAP7_75t_L g262 ( .A(n_140), .B(n_180), .Y(n_262) );
AND2x4_ASAP7_75t_L g298 ( .A(n_140), .B(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g312 ( .A(n_140), .B(n_313), .Y(n_312) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx2_ASAP7_75t_L g229 ( .A(n_141), .Y(n_229) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_141), .Y(n_401) );
OA21x2_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_146), .B(n_166), .Y(n_141) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_142), .A2(n_193), .B(n_194), .Y(n_192) );
CKINVDCx5p33_ASAP7_75t_R g205 ( .A(n_142), .Y(n_205) );
OA21x2_ASAP7_75t_L g275 ( .A1(n_142), .A2(n_146), .B(n_166), .Y(n_275) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
AND2x2_ASAP7_75t_SL g143 ( .A(n_144), .B(n_145), .Y(n_143) );
AND2x4_ASAP7_75t_L g216 ( .A(n_144), .B(n_145), .Y(n_216) );
AND2x6_ASAP7_75t_L g147 ( .A(n_148), .B(n_150), .Y(n_147) );
BUFx3_ASAP7_75t_L g469 ( .A(n_148), .Y(n_469) );
AND2x6_ASAP7_75t_L g162 ( .A(n_149), .B(n_155), .Y(n_162) );
INVx2_ASAP7_75t_L g476 ( .A(n_149), .Y(n_476) );
AND2x4_ASAP7_75t_L g472 ( .A(n_150), .B(n_473), .Y(n_472) );
AND2x2_ASAP7_75t_L g150 ( .A(n_151), .B(n_152), .Y(n_150) );
AND2x4_ASAP7_75t_L g164 ( .A(n_151), .B(n_157), .Y(n_164) );
INVx2_ASAP7_75t_L g466 ( .A(n_151), .Y(n_466) );
HB1xp67_ASAP7_75t_L g467 ( .A(n_152), .Y(n_467) );
AND2x4_ASAP7_75t_L g153 ( .A(n_154), .B(n_159), .Y(n_153) );
INVx1_ASAP7_75t_L g512 ( .A(n_154), .Y(n_512) );
AND2x4_ASAP7_75t_L g154 ( .A(n_155), .B(n_157), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx5_ASAP7_75t_L g165 ( .A(n_159), .Y(n_165) );
HB1xp67_ASAP7_75t_L g559 ( .A(n_159), .Y(n_559) );
AOI21xp5_ASAP7_75t_L g160 ( .A1(n_161), .A2(n_163), .B(n_165), .Y(n_160) );
INVxp67_ASAP7_75t_L g515 ( .A(n_162), .Y(n_515) );
INVxp67_ASAP7_75t_L g517 ( .A(n_164), .Y(n_517) );
AOI21xp5_ASAP7_75t_L g171 ( .A1(n_165), .A2(n_172), .B(n_173), .Y(n_171) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_165), .A2(n_184), .B(n_185), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g195 ( .A1(n_165), .A2(n_196), .B(n_197), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_165), .A2(n_202), .B(n_203), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_165), .A2(n_214), .B(n_215), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_165), .A2(n_223), .B(n_224), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_165), .A2(n_238), .B(n_239), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_165), .A2(n_478), .B(n_479), .Y(n_477) );
O2A1O1Ixp33_ASAP7_75t_L g487 ( .A1(n_165), .A2(n_481), .B(n_488), .C(n_489), .Y(n_487) );
O2A1O1Ixp33_ASAP7_75t_SL g499 ( .A1(n_165), .A2(n_481), .B(n_500), .C(n_501), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g518 ( .A(n_165), .B(n_216), .Y(n_518) );
INVx1_ASAP7_75t_L g529 ( .A(n_165), .Y(n_529) );
O2A1O1Ixp33_ASAP7_75t_L g540 ( .A1(n_165), .A2(n_481), .B(n_541), .C(n_542), .Y(n_540) );
O2A1O1Ixp33_ASAP7_75t_SL g549 ( .A1(n_165), .A2(n_481), .B(n_550), .C(n_551), .Y(n_549) );
A2O1A1Ixp33_ASAP7_75t_SL g256 ( .A1(n_167), .A2(n_229), .B(n_257), .C(n_261), .Y(n_256) );
AND2x2_ASAP7_75t_L g277 ( .A(n_167), .B(n_278), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_167), .B(n_229), .Y(n_417) );
AND2x2_ASAP7_75t_L g167 ( .A(n_168), .B(n_180), .Y(n_167) );
INVx2_ASAP7_75t_L g297 ( .A(n_168), .Y(n_297) );
BUFx3_ASAP7_75t_L g313 ( .A(n_168), .Y(n_313) );
INVxp67_ASAP7_75t_L g317 ( .A(n_168), .Y(n_317) );
AO21x2_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_175), .B(n_179), .Y(n_168) );
AO21x2_ASAP7_75t_L g267 ( .A1(n_169), .A2(n_175), .B(n_179), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_170), .B(n_174), .Y(n_169) );
AO21x2_ASAP7_75t_L g180 ( .A1(n_175), .A2(n_181), .B(n_187), .Y(n_180) );
AO21x2_ASAP7_75t_L g242 ( .A1(n_175), .A2(n_181), .B(n_187), .Y(n_242) );
AO21x2_ASAP7_75t_L g536 ( .A1(n_175), .A2(n_537), .B(n_543), .Y(n_536) );
OAI22xp5_ASAP7_75t_L g554 ( .A1(n_175), .A2(n_176), .B1(n_555), .B2(n_560), .Y(n_554) );
AO21x2_ASAP7_75t_L g573 ( .A1(n_175), .A2(n_537), .B(n_543), .Y(n_573) );
INVx3_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx4_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_177), .B(n_563), .Y(n_562) );
INVx3_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
BUFx4f_ASAP7_75t_L g209 ( .A(n_178), .Y(n_209) );
INVx2_ASAP7_75t_L g296 ( .A(n_180), .Y(n_296) );
AND2x2_ASAP7_75t_L g302 ( .A(n_180), .B(n_275), .Y(n_302) );
AND2x2_ASAP7_75t_L g328 ( .A(n_180), .B(n_297), .Y(n_328) );
NAND2xp5_ASAP7_75t_SL g181 ( .A(n_182), .B(n_186), .Y(n_181) );
AOI211xp5_ASAP7_75t_L g325 ( .A1(n_188), .A2(n_326), .B(n_329), .C(n_339), .Y(n_325) );
AND2x2_ASAP7_75t_SL g188 ( .A(n_189), .B(n_207), .Y(n_188) );
OAI321xp33_ASAP7_75t_L g300 ( .A1(n_189), .A2(n_248), .A3(n_301), .B1(n_303), .B2(n_304), .C(n_306), .Y(n_300) );
AND2x2_ASAP7_75t_L g421 ( .A(n_189), .B(n_396), .Y(n_421) );
INVx1_ASAP7_75t_L g424 ( .A(n_189), .Y(n_424) );
AND2x2_ASAP7_75t_L g189 ( .A(n_190), .B(n_198), .Y(n_189) );
INVx5_ASAP7_75t_L g246 ( .A(n_190), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_190), .B(n_260), .Y(n_259) );
NOR2x1_ASAP7_75t_SL g291 ( .A(n_190), .B(n_292), .Y(n_291) );
BUFx2_ASAP7_75t_L g336 ( .A(n_190), .Y(n_336) );
AND2x2_ASAP7_75t_L g438 ( .A(n_190), .B(n_208), .Y(n_438) );
OR2x6_ASAP7_75t_L g190 ( .A(n_191), .B(n_192), .Y(n_190) );
AND2x2_ASAP7_75t_L g245 ( .A(n_198), .B(n_246), .Y(n_245) );
HB1xp67_ASAP7_75t_L g255 ( .A(n_198), .Y(n_255) );
INVx4_ASAP7_75t_L g260 ( .A(n_198), .Y(n_260) );
AO21x2_ASAP7_75t_L g198 ( .A1(n_199), .A2(n_205), .B(n_206), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_200), .B(n_204), .Y(n_199) );
AO21x2_ASAP7_75t_L g495 ( .A1(n_205), .A2(n_496), .B(n_502), .Y(n_495) );
INVx1_ASAP7_75t_L g303 ( .A(n_207), .Y(n_303) );
A2O1A1Ixp33_ASAP7_75t_R g406 ( .A1(n_207), .A2(n_245), .B(n_277), .C(n_407), .Y(n_406) );
AND2x2_ASAP7_75t_L g426 ( .A(n_207), .B(n_251), .Y(n_426) );
AND2x2_ASAP7_75t_L g207 ( .A(n_208), .B(n_217), .Y(n_207) );
INVx1_ASAP7_75t_L g244 ( .A(n_208), .Y(n_244) );
INVx2_ASAP7_75t_L g250 ( .A(n_208), .Y(n_250) );
OR2x2_ASAP7_75t_L g269 ( .A(n_208), .B(n_260), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_208), .B(n_292), .Y(n_338) );
BUFx3_ASAP7_75t_L g345 ( .A(n_208), .Y(n_345) );
INVx2_ASAP7_75t_SL g482 ( .A(n_209), .Y(n_482) );
OA21x2_ASAP7_75t_L g547 ( .A1(n_209), .A2(n_548), .B(n_552), .Y(n_547) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_212), .B(n_216), .Y(n_210) );
INVx1_ASAP7_75t_SL g219 ( .A(n_216), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_216), .B(n_241), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_216), .A2(n_486), .B(n_490), .Y(n_485) );
INVx1_ASAP7_75t_L g308 ( .A(n_217), .Y(n_308) );
HB1xp67_ASAP7_75t_L g321 ( .A(n_217), .Y(n_321) );
INVx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVx1_ASAP7_75t_L g254 ( .A(n_218), .Y(n_254) );
INVx1_ASAP7_75t_L g363 ( .A(n_218), .Y(n_363) );
AO21x2_ASAP7_75t_L g218 ( .A1(n_219), .A2(n_220), .B(n_226), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_219), .B(n_227), .Y(n_226) );
AO21x2_ASAP7_75t_L g292 ( .A1(n_219), .A2(n_220), .B(n_226), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_221), .B(n_225), .Y(n_220) );
AND2x2_ASAP7_75t_L g264 ( .A(n_228), .B(n_265), .Y(n_264) );
OAI31xp33_ASAP7_75t_L g415 ( .A1(n_228), .A2(n_416), .A3(n_418), .B(n_421), .Y(n_415) );
INVx1_ASAP7_75t_SL g433 ( .A(n_228), .Y(n_433) );
AND2x4_ASAP7_75t_L g228 ( .A(n_229), .B(n_230), .Y(n_228) );
AOI21xp33_ASAP7_75t_L g247 ( .A1(n_229), .A2(n_248), .B(n_256), .Y(n_247) );
NAND2x1_ASAP7_75t_L g327 ( .A(n_229), .B(n_328), .Y(n_327) );
INVx1_ASAP7_75t_SL g356 ( .A(n_229), .Y(n_356) );
INVx2_ASAP7_75t_L g305 ( .A(n_230), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_230), .B(n_288), .Y(n_385) );
NOR2xp33_ASAP7_75t_L g397 ( .A(n_230), .B(n_287), .Y(n_397) );
NOR2xp33_ASAP7_75t_SL g405 ( .A(n_230), .B(n_356), .Y(n_405) );
AND2x4_ASAP7_75t_L g230 ( .A(n_231), .B(n_242), .Y(n_230) );
AND2x2_ASAP7_75t_SL g274 ( .A(n_231), .B(n_275), .Y(n_274) );
OR2x2_ASAP7_75t_L g285 ( .A(n_231), .B(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g314 ( .A(n_231), .B(n_296), .Y(n_314) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
BUFx2_ASAP7_75t_L g278 ( .A(n_232), .Y(n_278) );
INVx2_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
INVx2_ASAP7_75t_L g299 ( .A(n_233), .Y(n_299) );
OAI21x1_ASAP7_75t_SL g233 ( .A1(n_234), .A2(n_236), .B(n_240), .Y(n_233) );
INVx1_ASAP7_75t_L g241 ( .A(n_235), .Y(n_241) );
INVx2_ASAP7_75t_L g286 ( .A(n_242), .Y(n_286) );
HB1xp67_ASAP7_75t_L g346 ( .A(n_242), .Y(n_346) );
AND2x2_ASAP7_75t_L g243 ( .A(n_244), .B(n_245), .Y(n_243) );
INVx1_ASAP7_75t_L g282 ( .A(n_244), .Y(n_282) );
AND2x2_ASAP7_75t_L g361 ( .A(n_244), .B(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g272 ( .A(n_245), .B(n_266), .Y(n_272) );
INVx2_ASAP7_75t_SL g320 ( .A(n_245), .Y(n_320) );
INVx4_ASAP7_75t_L g251 ( .A(n_246), .Y(n_251) );
AND2x2_ASAP7_75t_L g349 ( .A(n_246), .B(n_292), .Y(n_349) );
AND2x2_ASAP7_75t_SL g367 ( .A(n_246), .B(n_362), .Y(n_367) );
NAND2x1p5_ASAP7_75t_L g384 ( .A(n_246), .B(n_260), .Y(n_384) );
INVx1_ASAP7_75t_L g390 ( .A(n_248), .Y(n_390) );
OR2x2_ASAP7_75t_L g248 ( .A(n_249), .B(n_252), .Y(n_248) );
INVx1_ASAP7_75t_L g309 ( .A(n_249), .Y(n_309) );
OR2x2_ASAP7_75t_L g322 ( .A(n_249), .B(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_250), .B(n_251), .Y(n_249) );
OR2x2_ASAP7_75t_L g374 ( .A(n_250), .B(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g404 ( .A(n_250), .B(n_292), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_251), .B(n_254), .Y(n_280) );
AND2x2_ASAP7_75t_L g372 ( .A(n_251), .B(n_362), .Y(n_372) );
AND2x4_ASAP7_75t_L g434 ( .A(n_251), .B(n_313), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_253), .B(n_255), .Y(n_252) );
INVx2_ASAP7_75t_L g258 ( .A(n_253), .Y(n_258) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
NOR2xp67_ASAP7_75t_SL g257 ( .A(n_258), .B(n_259), .Y(n_257) );
OAI322xp33_ASAP7_75t_SL g270 ( .A1(n_258), .A2(n_271), .A3(n_273), .B1(n_276), .B2(n_279), .C1(n_281), .C2(n_283), .Y(n_270) );
INVx1_ASAP7_75t_L g428 ( .A(n_258), .Y(n_428) );
OR2x2_ASAP7_75t_L g281 ( .A(n_259), .B(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g307 ( .A(n_260), .B(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_260), .B(n_308), .Y(n_323) );
INVx2_ASAP7_75t_L g350 ( .A(n_260), .Y(n_350) );
AND2x4_ASAP7_75t_L g362 ( .A(n_260), .B(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_SL g365 ( .A(n_262), .B(n_278), .Y(n_365) );
AOI21xp5_ASAP7_75t_L g263 ( .A1(n_264), .A2(n_268), .B(n_270), .Y(n_263) );
AND2x2_ASAP7_75t_L g331 ( .A(n_265), .B(n_298), .Y(n_331) );
INVx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_266), .B(n_420), .Y(n_419) );
BUFx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVx1_ASAP7_75t_L g289 ( .A(n_267), .Y(n_289) );
AND2x4_ASAP7_75t_SL g371 ( .A(n_267), .B(n_286), .Y(n_371) );
INVx2_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
OR2x2_ASAP7_75t_L g279 ( .A(n_269), .B(n_280), .Y(n_279) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_272), .B(n_356), .Y(n_355) );
INVx1_ASAP7_75t_SL g273 ( .A(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g407 ( .A(n_274), .B(n_371), .Y(n_407) );
NOR4xp25_ASAP7_75t_L g411 ( .A(n_274), .B(n_288), .C(n_328), .D(n_412), .Y(n_411) );
AND2x2_ASAP7_75t_L g288 ( .A(n_275), .B(n_289), .Y(n_288) );
OR2x2_ASAP7_75t_L g324 ( .A(n_275), .B(n_299), .Y(n_324) );
AND2x4_ASAP7_75t_L g388 ( .A(n_275), .B(n_299), .Y(n_388) );
INVx1_ASAP7_75t_SL g276 ( .A(n_277), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_278), .B(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
NOR2xp33_ASAP7_75t_L g284 ( .A(n_285), .B(n_287), .Y(n_284) );
OR2x2_ASAP7_75t_L g377 ( .A(n_285), .B(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g431 ( .A(n_285), .Y(n_431) );
NAND2xp5_ASAP7_75t_SL g332 ( .A(n_286), .B(n_298), .Y(n_332) );
INVx1_ASAP7_75t_SL g287 ( .A(n_288), .Y(n_287) );
AOI211xp5_ASAP7_75t_SL g290 ( .A1(n_291), .A2(n_293), .B(n_300), .C(n_315), .Y(n_290) );
INVx1_ASAP7_75t_SL g293 ( .A(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_295), .B(n_298), .Y(n_294) );
AND2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_296), .B(n_299), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_297), .B(n_302), .Y(n_301) );
BUFx2_ASAP7_75t_L g379 ( .A(n_297), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_298), .B(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g394 ( .A(n_298), .Y(n_394) );
OAI21xp5_ASAP7_75t_L g306 ( .A1(n_307), .A2(n_309), .B(n_310), .Y(n_306) );
AND2x4_ASAP7_75t_L g343 ( .A(n_307), .B(n_344), .Y(n_343) );
AND2x4_ASAP7_75t_L g437 ( .A(n_307), .B(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_312), .B(n_314), .Y(n_311) );
INVx1_ASAP7_75t_SL g341 ( .A(n_313), .Y(n_341) );
AND2x2_ASAP7_75t_L g400 ( .A(n_314), .B(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g414 ( .A(n_314), .Y(n_414) );
O2A1O1Ixp33_ASAP7_75t_SL g315 ( .A1(n_316), .A2(n_318), .B(n_322), .C(n_324), .Y(n_315) );
NAND2xp5_ASAP7_75t_SL g387 ( .A(n_316), .B(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
OR2x2_ASAP7_75t_L g392 ( .A(n_317), .B(n_393), .Y(n_392) );
OR2x2_ASAP7_75t_L g413 ( .A(n_317), .B(n_414), .Y(n_413) );
INVxp67_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
NOR2xp33_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
OR2x2_ASAP7_75t_L g402 ( .A(n_320), .B(n_344), .Y(n_402) );
OAI22xp5_ASAP7_75t_L g329 ( .A1(n_323), .A2(n_330), .B1(n_332), .B2(n_333), .Y(n_329) );
INVx1_ASAP7_75t_SL g420 ( .A(n_324), .Y(n_420) );
INVx2_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVxp67_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_335), .B(n_337), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_335), .B(n_344), .Y(n_386) );
INVx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVxp67_ASAP7_75t_SL g396 ( .A(n_338), .Y(n_396) );
OAI22xp5_ASAP7_75t_L g339 ( .A1(n_340), .A2(n_342), .B1(n_346), .B2(n_347), .Y(n_339) );
INVx2_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
AOI21xp5_ASAP7_75t_SL g353 ( .A1(n_344), .A2(n_354), .B(n_357), .Y(n_353) );
AND2x2_ASAP7_75t_L g382 ( .A(n_344), .B(n_383), .Y(n_382) );
INVx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
AND3x2_ASAP7_75t_L g348 ( .A(n_345), .B(n_349), .C(n_350), .Y(n_348) );
AND2x2_ASAP7_75t_L g410 ( .A(n_345), .B(n_367), .Y(n_410) );
INVx2_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g395 ( .A(n_350), .B(n_396), .Y(n_395) );
NOR2xp67_ASAP7_75t_L g351 ( .A(n_352), .B(n_408), .Y(n_351) );
NAND4xp25_ASAP7_75t_L g352 ( .A(n_353), .B(n_368), .C(n_389), .D(n_406), .Y(n_352) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
OAI22xp5_ASAP7_75t_L g357 ( .A1(n_358), .A2(n_360), .B1(n_364), .B2(n_366), .Y(n_357) );
INVx1_ASAP7_75t_SL g358 ( .A(n_359), .Y(n_358) );
OAI22xp5_ASAP7_75t_L g432 ( .A1(n_360), .A2(n_374), .B1(n_394), .B2(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx2_ASAP7_75t_L g375 ( .A(n_362), .Y(n_375) );
AOI21xp5_ASAP7_75t_L g435 ( .A1(n_364), .A2(n_387), .B(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx3_ASAP7_75t_SL g366 ( .A(n_367), .Y(n_366) );
AOI221xp5_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_372), .B1(n_373), .B2(n_376), .C(n_380), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx2_ASAP7_75t_SL g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_SL g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
OAI22xp5_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_385), .B1(n_386), .B2(n_387), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_383), .B(n_404), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_383), .B(n_428), .Y(n_427) );
INVx2_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
AOI221xp5_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_391), .B1(n_395), .B2(n_397), .C(n_398), .Y(n_389) );
NAND2xp5_ASAP7_75t_SL g391 ( .A(n_392), .B(n_394), .Y(n_391) );
OAI22xp5_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_402), .B1(n_403), .B2(n_405), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
OAI211xp5_ASAP7_75t_SL g423 ( .A1(n_404), .A2(n_424), .B(n_425), .C(n_427), .Y(n_423) );
OAI211xp5_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_411), .B(n_415), .C(n_422), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_SL g418 ( .A(n_419), .Y(n_418) );
AOI221xp5_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_429), .B1(n_432), .B2(n_434), .C(n_435), .Y(n_422) );
INVx1_ASAP7_75t_SL g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_SL g436 ( .A(n_437), .Y(n_436) );
CKINVDCx20_ASAP7_75t_R g442 ( .A(n_443), .Y(n_442) );
CKINVDCx11_ASAP7_75t_R g443 ( .A(n_444), .Y(n_443) );
CKINVDCx20_ASAP7_75t_R g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
NAND2xp5_ASAP7_75t_SL g813 ( .A(n_448), .B(n_814), .Y(n_813) );
AOI21xp5_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_797), .B(n_809), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_451), .B(n_788), .Y(n_450) );
OAI22xp5_ASAP7_75t_SL g451 ( .A1(n_452), .A2(n_784), .B1(n_785), .B2(n_786), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVxp67_ASAP7_75t_L g802 ( .A(n_454), .Y(n_802) );
NAND4xp75_ASAP7_75t_L g454 ( .A(n_455), .B(n_635), .C(n_701), .D(n_764), .Y(n_454) );
NOR2x1_ASAP7_75t_L g455 ( .A(n_456), .B(n_598), .Y(n_455) );
OR3x1_ASAP7_75t_L g456 ( .A(n_457), .B(n_568), .C(n_595), .Y(n_456) );
AOI21xp5_ASAP7_75t_L g457 ( .A1(n_458), .A2(n_503), .B(n_524), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_460), .B(n_492), .Y(n_459) );
AND2x2_ASAP7_75t_L g698 ( .A(n_460), .B(n_668), .Y(n_698) );
INVx1_ASAP7_75t_L g771 ( .A(n_460), .Y(n_771) );
AND2x2_ASAP7_75t_L g460 ( .A(n_461), .B(n_483), .Y(n_460) );
INVx2_ASAP7_75t_L g523 ( .A(n_461), .Y(n_523) );
HB1xp67_ASAP7_75t_L g586 ( .A(n_461), .Y(n_586) );
AND2x2_ASAP7_75t_L g590 ( .A(n_461), .B(n_506), .Y(n_590) );
AND2x4_ASAP7_75t_L g606 ( .A(n_461), .B(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g610 ( .A(n_461), .Y(n_610) );
AND2x2_ASAP7_75t_L g461 ( .A(n_462), .B(n_471), .Y(n_461) );
NOR3xp33_ASAP7_75t_L g463 ( .A(n_464), .B(n_468), .C(n_470), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
AND2x4_ASAP7_75t_L g491 ( .A(n_465), .B(n_469), .Y(n_491) );
AND2x2_ASAP7_75t_L g465 ( .A(n_466), .B(n_467), .Y(n_465) );
OR2x6_ASAP7_75t_L g481 ( .A(n_466), .B(n_476), .Y(n_481) );
INVxp33_ASAP7_75t_L g532 ( .A(n_466), .Y(n_532) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVxp67_ASAP7_75t_L g565 ( .A(n_472), .Y(n_565) );
NOR2x1p5_ASAP7_75t_L g473 ( .A(n_474), .B(n_475), .Y(n_473) );
INVx1_ASAP7_75t_L g533 ( .A(n_475), .Y(n_533) );
INVx3_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
OAI22xp5_ASAP7_75t_L g509 ( .A1(n_481), .A2(n_510), .B1(n_511), .B2(n_512), .Y(n_509) );
INVxp67_ASAP7_75t_L g556 ( .A(n_481), .Y(n_556) );
AO21x2_ASAP7_75t_L g526 ( .A1(n_482), .A2(n_527), .B(n_535), .Y(n_526) );
AO21x2_ASAP7_75t_L g574 ( .A1(n_482), .A2(n_527), .B(n_535), .Y(n_574) );
AND2x2_ASAP7_75t_L g504 ( .A(n_483), .B(n_505), .Y(n_504) );
INVx4_ASAP7_75t_L g587 ( .A(n_483), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_483), .B(n_577), .Y(n_591) );
INVx2_ASAP7_75t_L g605 ( .A(n_483), .Y(n_605) );
AND2x4_ASAP7_75t_L g609 ( .A(n_483), .B(n_610), .Y(n_609) );
BUFx6f_ASAP7_75t_L g644 ( .A(n_483), .Y(n_644) );
OR2x2_ASAP7_75t_L g650 ( .A(n_483), .B(n_495), .Y(n_650) );
NOR2x1_ASAP7_75t_SL g679 ( .A(n_483), .B(n_506), .Y(n_679) );
NAND2xp5_ASAP7_75t_SL g781 ( .A(n_483), .B(n_753), .Y(n_781) );
OR2x6_ASAP7_75t_L g483 ( .A(n_484), .B(n_485), .Y(n_483) );
INVx1_ASAP7_75t_L g567 ( .A(n_491), .Y(n_567) );
AND2x2_ASAP7_75t_L g678 ( .A(n_492), .B(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
NAND2x1_ASAP7_75t_L g712 ( .A(n_493), .B(n_505), .Y(n_712) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
HB1xp67_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g520 ( .A(n_495), .Y(n_520) );
INVx2_ASAP7_75t_L g578 ( .A(n_495), .Y(n_578) );
AND2x2_ASAP7_75t_L g601 ( .A(n_495), .B(n_506), .Y(n_601) );
HB1xp67_ASAP7_75t_L g628 ( .A(n_495), .Y(n_628) );
INVx1_ASAP7_75t_L g669 ( .A(n_495), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_497), .B(n_498), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_504), .B(n_519), .Y(n_503) );
AND2x2_ASAP7_75t_L g681 ( .A(n_504), .B(n_576), .Y(n_681) );
NOR2xp33_ASAP7_75t_L g595 ( .A(n_505), .B(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g748 ( .A(n_505), .Y(n_748) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx3_ASAP7_75t_L g607 ( .A(n_506), .Y(n_607) );
AND2x4_ASAP7_75t_L g506 ( .A(n_507), .B(n_508), .Y(n_506) );
OAI21xp5_ASAP7_75t_L g508 ( .A1(n_509), .A2(n_513), .B(n_518), .Y(n_508) );
NOR2xp33_ASAP7_75t_L g557 ( .A(n_512), .B(n_558), .Y(n_557) );
OAI22xp5_ASAP7_75t_L g513 ( .A1(n_514), .A2(n_515), .B1(n_516), .B2(n_517), .Y(n_513) );
OAI211xp5_ASAP7_75t_SL g684 ( .A1(n_519), .A2(n_685), .B(n_689), .C(n_695), .Y(n_684) );
NAND2xp5_ASAP7_75t_SL g519 ( .A(n_520), .B(n_521), .Y(n_519) );
AND2x2_ASAP7_75t_SL g600 ( .A(n_521), .B(n_601), .Y(n_600) );
INVx2_ASAP7_75t_SL g731 ( .A(n_521), .Y(n_731) );
INVx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
AND2x2_ASAP7_75t_L g653 ( .A(n_523), .B(n_607), .Y(n_653) );
OR2x2_ASAP7_75t_L g524 ( .A(n_525), .B(n_544), .Y(n_524) );
AOI32xp33_ASAP7_75t_L g689 ( .A1(n_525), .A2(n_673), .A3(n_690), .B1(n_691), .B2(n_693), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_526), .B(n_536), .Y(n_525) );
INVx2_ASAP7_75t_L g615 ( .A(n_526), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_526), .B(n_547), .Y(n_683) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_528), .B(n_534), .Y(n_527) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx3_ASAP7_75t_L g627 ( .A(n_536), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_536), .B(n_553), .Y(n_658) );
AND2x2_ASAP7_75t_L g663 ( .A(n_536), .B(n_664), .Y(n_663) );
HB1xp67_ASAP7_75t_L g745 ( .A(n_536), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_538), .B(n_539), .Y(n_537) );
OR2x2_ASAP7_75t_L g646 ( .A(n_544), .B(n_647), .Y(n_646) );
INVx3_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
AND2x2_ASAP7_75t_L g597 ( .A(n_545), .B(n_571), .Y(n_597) );
AND2x2_ASAP7_75t_L g746 ( .A(n_545), .B(n_744), .Y(n_746) );
AND2x4_ASAP7_75t_L g545 ( .A(n_546), .B(n_553), .Y(n_545) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx1_ASAP7_75t_L g583 ( .A(n_547), .Y(n_583) );
AND2x4_ASAP7_75t_L g622 ( .A(n_547), .B(n_623), .Y(n_622) );
INVxp67_ASAP7_75t_L g656 ( .A(n_547), .Y(n_656) );
HB1xp67_ASAP7_75t_L g664 ( .A(n_547), .Y(n_664) );
AND2x2_ASAP7_75t_L g673 ( .A(n_547), .B(n_553), .Y(n_673) );
INVx1_ASAP7_75t_L g757 ( .A(n_547), .Y(n_757) );
INVx2_ASAP7_75t_L g594 ( .A(n_553), .Y(n_594) );
INVx1_ASAP7_75t_L g621 ( .A(n_553), .Y(n_621) );
INVx1_ASAP7_75t_L g688 ( .A(n_553), .Y(n_688) );
OR2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_561), .Y(n_553) );
OAI22xp5_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_565), .B1(n_566), .B2(n_567), .Y(n_561) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
OAI32xp33_ASAP7_75t_L g568 ( .A1(n_569), .A2(n_579), .A3(n_584), .B1(n_588), .B2(n_592), .Y(n_568) );
INVx1_ASAP7_75t_SL g569 ( .A(n_570), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_570), .B(n_768), .Y(n_767) );
AND2x2_ASAP7_75t_L g570 ( .A(n_571), .B(n_575), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_571), .B(n_631), .Y(n_630) );
AND2x2_ASAP7_75t_L g672 ( .A(n_571), .B(n_673), .Y(n_672) );
INVxp67_ASAP7_75t_L g697 ( .A(n_571), .Y(n_697) );
AND2x2_ASAP7_75t_L g778 ( .A(n_571), .B(n_620), .Y(n_778) );
AND2x4_ASAP7_75t_L g571 ( .A(n_572), .B(n_574), .Y(n_571) );
INVx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g593 ( .A(n_573), .B(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g692 ( .A(n_573), .B(n_615), .Y(n_692) );
NOR2xp67_ASAP7_75t_L g714 ( .A(n_573), .B(n_594), .Y(n_714) );
NOR2x1_ASAP7_75t_L g756 ( .A(n_573), .B(n_757), .Y(n_756) );
INVx2_ASAP7_75t_L g623 ( .A(n_574), .Y(n_623) );
INVx1_ASAP7_75t_L g647 ( .A(n_574), .Y(n_647) );
AND2x2_ASAP7_75t_L g662 ( .A(n_574), .B(n_594), .Y(n_662) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g690 ( .A(n_576), .B(n_679), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_576), .B(n_609), .Y(n_760) );
INVx3_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
HB1xp67_ASAP7_75t_L g729 ( .A(n_577), .Y(n_729) );
INVx2_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
HB1xp67_ASAP7_75t_L g711 ( .A(n_578), .Y(n_711) );
INVxp67_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
OR2x2_ASAP7_75t_L g612 ( .A(n_581), .B(n_613), .Y(n_612) );
NOR2xp67_ASAP7_75t_L g696 ( .A(n_581), .B(n_697), .Y(n_696) );
NOR2xp67_ASAP7_75t_SL g783 ( .A(n_581), .B(n_721), .Y(n_783) );
INVx3_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
BUFx3_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g640 ( .A(n_583), .B(n_594), .Y(n_640) );
NAND2xp5_ASAP7_75t_SL g708 ( .A(n_584), .B(n_650), .Y(n_708) );
INVx2_ASAP7_75t_SL g584 ( .A(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_SL g674 ( .A(n_585), .B(n_601), .Y(n_674) );
AND2x4_ASAP7_75t_SL g585 ( .A(n_586), .B(n_587), .Y(n_585) );
NOR2x1_ASAP7_75t_L g633 ( .A(n_587), .B(n_634), .Y(n_633) );
AND2x4_ASAP7_75t_L g739 ( .A(n_587), .B(n_610), .Y(n_739) );
HB1xp67_ASAP7_75t_L g768 ( .A(n_587), .Y(n_768) );
NAND2xp5_ASAP7_75t_SL g759 ( .A(n_588), .B(n_760), .Y(n_759) );
OR2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_591), .Y(n_588) );
OR2x2_ASAP7_75t_L g710 ( .A(n_589), .B(n_711), .Y(n_710) );
NOR2x1_ASAP7_75t_L g775 ( .A(n_589), .B(n_776), .Y(n_775) );
INVx2_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g699 ( .A(n_590), .B(n_644), .Y(n_699) );
INVxp33_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
NAND2x1p5_ASAP7_75t_L g613 ( .A(n_593), .B(n_614), .Y(n_613) );
AND2x2_ASAP7_75t_L g773 ( .A(n_593), .B(n_655), .Y(n_773) );
INVx2_ASAP7_75t_SL g596 ( .A(n_597), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_599), .B(n_616), .Y(n_598) );
OAI21xp33_ASAP7_75t_L g599 ( .A1(n_600), .A2(n_602), .B(n_611), .Y(n_599) );
AND2x2_ASAP7_75t_L g734 ( .A(n_601), .B(n_609), .Y(n_734) );
NAND2xp33_ASAP7_75t_R g602 ( .A(n_603), .B(n_608), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_605), .B(n_606), .Y(n_604) );
INVx1_ASAP7_75t_L g776 ( .A(n_605), .Y(n_776) );
INVx4_ASAP7_75t_L g634 ( .A(n_606), .Y(n_634) );
INVx1_ASAP7_75t_L g753 ( .A(n_607), .Y(n_753) );
INVx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g747 ( .A(n_609), .B(n_748), .Y(n_747) );
AND2x2_ASAP7_75t_SL g751 ( .A(n_609), .B(n_752), .Y(n_751) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
OAI22xp5_ASAP7_75t_L g780 ( .A1(n_612), .A2(n_677), .B1(n_781), .B2(n_782), .Y(n_780) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
AND2x4_ASAP7_75t_L g641 ( .A(n_615), .B(n_627), .Y(n_641) );
AND2x2_ASAP7_75t_L g655 ( .A(n_615), .B(n_656), .Y(n_655) );
A2O1A1Ixp33_ASAP7_75t_SL g616 ( .A1(n_617), .A2(n_624), .B(n_629), .C(n_632), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx3_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g703 ( .A(n_619), .B(n_704), .Y(n_703) );
AND2x2_ASAP7_75t_L g619 ( .A(n_620), .B(n_622), .Y(n_619) );
INVx1_ASAP7_75t_L g631 ( .A(n_620), .Y(n_631) );
INVx2_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g691 ( .A(n_621), .B(n_692), .Y(n_691) );
AND2x2_ASAP7_75t_L g700 ( .A(n_621), .B(n_622), .Y(n_700) );
INVx1_ASAP7_75t_L g732 ( .A(n_621), .Y(n_732) );
AND2x4_ASAP7_75t_L g713 ( .A(n_622), .B(n_714), .Y(n_713) );
AND2x2_ASAP7_75t_L g735 ( .A(n_622), .B(n_626), .Y(n_735) );
AND2x2_ASAP7_75t_L g743 ( .A(n_622), .B(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_626), .B(n_628), .Y(n_625) );
INVx1_ASAP7_75t_L g718 ( .A(n_626), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_626), .B(n_640), .Y(n_720) );
AND2x2_ASAP7_75t_L g723 ( .A(n_626), .B(n_673), .Y(n_723) );
INVx3_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_627), .B(n_688), .Y(n_737) );
AND2x2_ASAP7_75t_L g665 ( .A(n_628), .B(n_653), .Y(n_665) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g761 ( .A(n_631), .B(n_641), .Y(n_761) );
BUFx2_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_633), .B(n_668), .Y(n_667) );
INVx2_ASAP7_75t_L g645 ( .A(n_634), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_634), .B(n_649), .Y(n_648) );
AND2x2_ASAP7_75t_L g635 ( .A(n_636), .B(n_675), .Y(n_635) );
NOR2xp33_ASAP7_75t_L g636 ( .A(n_637), .B(n_659), .Y(n_636) );
OAI222xp33_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_642), .B1(n_646), .B2(n_648), .C1(n_651), .C2(n_654), .Y(n_637) );
INVx1_ASAP7_75t_SL g638 ( .A(n_639), .Y(n_638) );
AND2x2_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .Y(n_639) );
NOR2xp33_ASAP7_75t_L g642 ( .A(n_643), .B(n_645), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_SL g652 ( .A(n_644), .B(n_653), .Y(n_652) );
OR2x6_ASAP7_75t_L g724 ( .A(n_644), .B(n_694), .Y(n_724) );
NAND5xp2_ASAP7_75t_L g727 ( .A(n_644), .B(n_647), .C(n_663), .D(n_728), .E(n_730), .Y(n_727) );
NAND2x1_ASAP7_75t_L g763 ( .A(n_645), .B(n_649), .Y(n_763) );
INVx2_ASAP7_75t_SL g649 ( .A(n_650), .Y(n_649) );
NOR2x1_ASAP7_75t_L g693 ( .A(n_650), .B(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
AOI22xp5_ASAP7_75t_L g742 ( .A1(n_652), .A2(n_743), .B1(n_746), .B2(n_747), .Y(n_742) );
INVx2_ASAP7_75t_L g694 ( .A(n_653), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_653), .B(n_669), .Y(n_706) );
INVx3_ASAP7_75t_L g741 ( .A(n_654), .Y(n_741) );
NAND2x1p5_ASAP7_75t_L g654 ( .A(n_655), .B(n_657), .Y(n_654) );
AND2x2_ASAP7_75t_L g686 ( .A(n_655), .B(n_687), .Y(n_686) );
BUFx2_ASAP7_75t_L g719 ( .A(n_655), .Y(n_719) );
INVx2_ASAP7_75t_SL g657 ( .A(n_658), .Y(n_657) );
OR2x2_ASAP7_75t_L g682 ( .A(n_658), .B(n_683), .Y(n_682) );
NAND2xp5_ASAP7_75t_SL g659 ( .A(n_660), .B(n_671), .Y(n_659) );
AOI21xp5_ASAP7_75t_L g660 ( .A1(n_661), .A2(n_665), .B(n_666), .Y(n_660) );
AND2x4_ASAP7_75t_L g661 ( .A(n_662), .B(n_663), .Y(n_661) );
INVx1_ASAP7_75t_L g670 ( .A(n_662), .Y(n_670) );
AOI22xp5_ASAP7_75t_L g671 ( .A1(n_665), .A2(n_672), .B1(n_673), .B2(n_674), .Y(n_671) );
NOR2xp33_ASAP7_75t_L g666 ( .A(n_667), .B(n_670), .Y(n_666) );
HB1xp67_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
AND2x4_ASAP7_75t_SL g752 ( .A(n_669), .B(n_753), .Y(n_752) );
NOR2xp33_ASAP7_75t_L g675 ( .A(n_676), .B(n_684), .Y(n_675) );
AOI21xp33_ASAP7_75t_L g676 ( .A1(n_677), .A2(n_680), .B(n_682), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
BUFx2_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g721 ( .A(n_692), .Y(n_721) );
AOI22xp5_ASAP7_75t_L g695 ( .A1(n_696), .A2(n_698), .B1(n_699), .B2(n_700), .Y(n_695) );
AND2x2_ASAP7_75t_L g701 ( .A(n_702), .B(n_725), .Y(n_701) );
NOR3xp33_ASAP7_75t_L g702 ( .A(n_703), .B(n_707), .C(n_715), .Y(n_702) );
INVx2_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
BUFx2_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
OA21x2_ASAP7_75t_SL g707 ( .A1(n_708), .A2(n_709), .B(n_713), .Y(n_707) );
NAND2xp33_ASAP7_75t_SL g709 ( .A(n_710), .B(n_712), .Y(n_709) );
AOI21xp33_ASAP7_75t_L g715 ( .A1(n_716), .A2(n_722), .B(n_724), .Y(n_715) );
OAI211xp5_ASAP7_75t_L g716 ( .A1(n_717), .A2(n_719), .B(n_720), .C(n_721), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
AOI22xp5_ASAP7_75t_L g758 ( .A1(n_719), .A2(n_759), .B1(n_761), .B2(n_762), .Y(n_758) );
INVx1_ASAP7_75t_SL g722 ( .A(n_723), .Y(n_722) );
NOR2xp33_ASAP7_75t_L g725 ( .A(n_726), .B(n_749), .Y(n_725) );
NAND4xp25_ASAP7_75t_L g726 ( .A(n_727), .B(n_733), .C(n_740), .D(n_742), .Y(n_726) );
HB1xp67_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
AND2x2_ASAP7_75t_L g738 ( .A(n_729), .B(n_739), .Y(n_738) );
NOR2xp33_ASAP7_75t_L g730 ( .A(n_731), .B(n_732), .Y(n_730) );
INVx1_ASAP7_75t_L g769 ( .A(n_732), .Y(n_769) );
AOI22xp5_ASAP7_75t_L g733 ( .A1(n_734), .A2(n_735), .B1(n_736), .B2(n_738), .Y(n_733) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_738), .B(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
OAI21xp5_ASAP7_75t_SL g749 ( .A1(n_750), .A2(n_754), .B(n_758), .Y(n_749) );
INVx1_ASAP7_75t_SL g750 ( .A(n_751), .Y(n_750) );
INVxp67_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
HB1xp67_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
AND2x2_ASAP7_75t_L g764 ( .A(n_765), .B(n_779), .Y(n_764) );
AOI21xp5_ASAP7_75t_L g765 ( .A1(n_766), .A2(n_769), .B(n_770), .Y(n_765) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
OAI22xp5_ASAP7_75t_L g770 ( .A1(n_771), .A2(n_772), .B1(n_774), .B2(n_777), .Y(n_770) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
INVx1_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
INVx1_ASAP7_75t_SL g777 ( .A(n_778), .Y(n_777) );
INVx1_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
CKINVDCx11_ASAP7_75t_R g801 ( .A(n_784), .Y(n_801) );
CKINVDCx11_ASAP7_75t_R g786 ( .A(n_787), .Y(n_786) );
CKINVDCx5p33_ASAP7_75t_R g805 ( .A(n_787), .Y(n_805) );
INVx1_ASAP7_75t_L g798 ( .A(n_788), .Y(n_798) );
INVx1_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
INVx1_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
AOI21xp5_ASAP7_75t_L g797 ( .A1(n_798), .A2(n_799), .B(n_806), .Y(n_797) );
INVx1_ASAP7_75t_SL g800 ( .A(n_801), .Y(n_800) );
INVx4_ASAP7_75t_SL g803 ( .A(n_804), .Y(n_803) );
INVx3_ASAP7_75t_SL g804 ( .A(n_805), .Y(n_804) );
NOR2xp33_ASAP7_75t_L g806 ( .A(n_807), .B(n_808), .Y(n_806) );
CKINVDCx20_ASAP7_75t_R g809 ( .A(n_810), .Y(n_809) );
BUFx2_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
INVxp67_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
endmodule