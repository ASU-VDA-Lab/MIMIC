module real_aes_11347_n_249 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_246, n_248, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_249);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_249;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_254;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_260;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1441;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_1382;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1346;
wire n_1383;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_411;
wire n_498;
wire n_1397;
wire n_765;
wire n_648;
wire n_1487;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1510;
wire n_1495;
wire n_712;
wire n_266;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_258;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_877;
wire n_424;
wire n_802;
wire n_1488;
wire n_337;
wire n_264;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_1392;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1500;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1386;
wire n_406;
wire n_1493;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_255;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_261;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_1462;
wire n_701;
wire n_809;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_689;
wire n_1483;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1474;
wire n_1032;
wire n_721;
wire n_1431;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1162;
wire n_1463;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_253;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_257;
wire n_285;
wire n_1377;
wire n_800;
wire n_1175;
wire n_778;
wire n_1170;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_856;
wire n_594;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1373;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_263;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_267;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_769;
wire n_434;
wire n_250;
wire n_1455;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_251;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_273;
wire n_1482;
wire n_1038;
wire n_276;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_1494;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_262;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_252;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_1496;
wire n_524;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_1457;
wire n_719;
wire n_465;
wire n_1343;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_640;
wire n_1176;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1420;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_892;
wire n_372;
wire n_578;
wire n_938;
wire n_327;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1290;
wire n_1318;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_969;
wire n_256;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_269;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_275;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_1481;
wire n_907;
wire n_1430;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_516;
wire n_335;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1436;
wire n_793;
wire n_1390;
wire n_272;
wire n_1412;
wire n_757;
wire n_803;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_1097;
wire n_703;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_259;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AOI22xp33_ASAP7_75t_L g936 ( .A1(n_0), .A2(n_64), .B1(n_813), .B2(n_886), .Y(n_936) );
INVx1_ASAP7_75t_L g972 ( .A(n_0), .Y(n_972) );
AO22x2_ASAP7_75t_L g645 ( .A1(n_1), .A2(n_646), .B1(n_700), .B2(n_701), .Y(n_645) );
INVxp67_ASAP7_75t_L g700 ( .A(n_1), .Y(n_700) );
AOI22xp5_ASAP7_75t_L g1185 ( .A1(n_1), .A2(n_6), .B1(n_1169), .B2(n_1186), .Y(n_1185) );
OAI22xp5_ASAP7_75t_L g285 ( .A1(n_2), .A2(n_201), .B1(n_286), .B2(n_294), .Y(n_285) );
INVx1_ASAP7_75t_L g408 ( .A(n_2), .Y(n_408) );
AOI22xp33_ASAP7_75t_L g814 ( .A1(n_3), .A2(n_214), .B1(n_690), .B2(n_815), .Y(n_814) );
INVx1_ASAP7_75t_L g824 ( .A(n_3), .Y(n_824) );
CKINVDCx5p33_ASAP7_75t_R g1036 ( .A(n_4), .Y(n_1036) );
HB1xp67_ASAP7_75t_L g263 ( .A(n_5), .Y(n_263) );
INVx1_ASAP7_75t_L g452 ( .A(n_5), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_5), .B(n_179), .Y(n_494) );
AND2x2_ASAP7_75t_L g498 ( .A(n_5), .B(n_290), .Y(n_498) );
INVxp67_ASAP7_75t_SL g1377 ( .A(n_7), .Y(n_1377) );
AOI22xp33_ASAP7_75t_L g1415 ( .A1(n_7), .A2(n_189), .B1(n_690), .B2(n_1416), .Y(n_1415) );
AOI22xp5_ASAP7_75t_L g1189 ( .A1(n_8), .A2(n_213), .B1(n_1175), .B2(n_1178), .Y(n_1189) );
INVx1_ASAP7_75t_L g595 ( .A(n_9), .Y(n_595) );
OAI22xp33_ASAP7_75t_L g630 ( .A1(n_9), .A2(n_130), .B1(n_631), .B2(n_634), .Y(n_630) );
CKINVDCx5p33_ASAP7_75t_R g326 ( .A(n_10), .Y(n_326) );
INVx1_ASAP7_75t_L g778 ( .A(n_11), .Y(n_778) );
OAI22xp5_ASAP7_75t_L g820 ( .A1(n_11), .A2(n_71), .B1(n_821), .B2(n_822), .Y(n_820) );
CKINVDCx14_ASAP7_75t_R g1194 ( .A(n_12), .Y(n_1194) );
INVxp67_ASAP7_75t_L g1375 ( .A(n_13), .Y(n_1375) );
AOI221xp5_ASAP7_75t_L g1412 ( .A1(n_13), .A2(n_151), .B1(n_816), .B2(n_915), .C(n_1413), .Y(n_1412) );
XNOR2x2_ASAP7_75t_L g455 ( .A(n_14), .B(n_456), .Y(n_455) );
CKINVDCx5p33_ASAP7_75t_R g1001 ( .A(n_15), .Y(n_1001) );
AOI21xp33_ASAP7_75t_L g479 ( .A1(n_16), .A2(n_480), .B(n_481), .Y(n_479) );
INVx1_ASAP7_75t_L g559 ( .A(n_16), .Y(n_559) );
INVxp67_ASAP7_75t_SL g580 ( .A(n_17), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g624 ( .A1(n_17), .A2(n_223), .B1(n_615), .B2(n_625), .Y(n_624) );
AO22x2_ASAP7_75t_L g1082 ( .A1(n_18), .A2(n_1083), .B1(n_1084), .B2(n_1134), .Y(n_1082) );
INVxp67_ASAP7_75t_SL g1083 ( .A(n_18), .Y(n_1083) );
XNOR2xp5_ASAP7_75t_L g834 ( .A(n_19), .B(n_835), .Y(n_834) );
OAI22xp5_ASAP7_75t_L g338 ( .A1(n_20), .A2(n_43), .B1(n_339), .B2(n_347), .Y(n_338) );
INVx1_ASAP7_75t_L g440 ( .A(n_20), .Y(n_440) );
INVxp33_ASAP7_75t_L g1405 ( .A(n_21), .Y(n_1405) );
AOI22xp33_ASAP7_75t_L g1420 ( .A1(n_21), .A2(n_98), .B1(n_561), .B2(n_1116), .Y(n_1420) );
INVx2_ASAP7_75t_L g333 ( .A(n_22), .Y(n_333) );
OR2x2_ASAP7_75t_L g558 ( .A(n_22), .B(n_543), .Y(n_558) );
OAI22xp5_ASAP7_75t_L g495 ( .A1(n_23), .A2(n_146), .B1(n_496), .B2(n_502), .Y(n_495) );
INVx1_ASAP7_75t_L g534 ( .A(n_23), .Y(n_534) );
CKINVDCx5p33_ASAP7_75t_R g483 ( .A(n_24), .Y(n_483) );
AOI22xp33_ASAP7_75t_SL g607 ( .A1(n_25), .A2(n_74), .B1(n_604), .B2(n_608), .Y(n_607) );
INVxp33_ASAP7_75t_L g641 ( .A(n_25), .Y(n_641) );
AOI22xp33_ASAP7_75t_L g938 ( .A1(n_26), .A2(n_193), .B1(n_815), .B2(n_917), .Y(n_938) );
OAI22xp5_ASAP7_75t_L g980 ( .A1(n_26), .A2(n_193), .B1(n_502), .B2(n_981), .Y(n_980) );
AOI22xp33_ASAP7_75t_L g789 ( .A1(n_27), .A2(n_93), .B1(n_790), .B2(n_791), .Y(n_789) );
AOI22xp33_ASAP7_75t_L g805 ( .A1(n_27), .A2(n_93), .B1(n_806), .B2(n_808), .Y(n_805) );
BUFx2_ASAP7_75t_L g281 ( .A(n_28), .Y(n_281) );
BUFx2_ASAP7_75t_L g379 ( .A(n_28), .Y(n_379) );
INVx1_ASAP7_75t_L g450 ( .A(n_28), .Y(n_450) );
OR2x2_ASAP7_75t_L g1010 ( .A(n_28), .B(n_494), .Y(n_1010) );
AOI22xp33_ASAP7_75t_SL g904 ( .A1(n_29), .A2(n_172), .B1(n_793), .B2(n_856), .Y(n_904) );
AOI22xp33_ASAP7_75t_L g908 ( .A1(n_29), .A2(n_172), .B1(n_909), .B2(n_910), .Y(n_908) );
INVx1_ASAP7_75t_L g847 ( .A(n_30), .Y(n_847) );
AOI22xp33_ASAP7_75t_L g855 ( .A1(n_30), .A2(n_171), .B1(n_604), .B2(n_856), .Y(n_855) );
INVxp33_ASAP7_75t_L g1404 ( .A(n_31), .Y(n_1404) );
AOI21xp33_ASAP7_75t_L g1423 ( .A1(n_31), .A2(n_618), .B(n_1424), .Y(n_1423) );
INVx1_ASAP7_75t_L g588 ( .A(n_32), .Y(n_588) );
AOI22xp33_ASAP7_75t_L g620 ( .A1(n_32), .A2(n_58), .B1(n_621), .B2(n_622), .Y(n_620) );
OAI221xp5_ASAP7_75t_L g655 ( .A1(n_33), .A2(n_209), .B1(n_634), .B2(n_656), .C(n_657), .Y(n_655) );
INVx1_ASAP7_75t_L g667 ( .A(n_33), .Y(n_667) );
OAI22xp33_ASAP7_75t_L g898 ( .A1(n_34), .A2(n_53), .B1(n_264), .B2(n_586), .Y(n_898) );
AOI22xp33_ASAP7_75t_L g913 ( .A1(n_34), .A2(n_155), .B1(n_914), .B2(n_915), .Y(n_913) );
INVx1_ASAP7_75t_L g1389 ( .A(n_35), .Y(n_1389) );
OAI22xp33_ASAP7_75t_L g506 ( .A1(n_36), .A2(n_41), .B1(n_507), .B2(n_509), .Y(n_506) );
AOI221xp5_ASAP7_75t_L g527 ( .A1(n_36), .A2(n_41), .B1(n_516), .B2(n_528), .C(n_530), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g1121 ( .A1(n_37), .A2(n_60), .B1(n_1119), .B2(n_1122), .Y(n_1121) );
INVxp67_ASAP7_75t_SL g1127 ( .A(n_37), .Y(n_1127) );
INVx1_ASAP7_75t_L g1477 ( .A(n_38), .Y(n_1477) );
OAI22xp5_ASAP7_75t_L g1501 ( .A1(n_38), .A2(n_51), .B1(n_1502), .B2(n_1504), .Y(n_1501) );
AOI22xp33_ASAP7_75t_L g850 ( .A1(n_39), .A2(n_202), .B1(n_516), .B2(n_618), .Y(n_850) );
AOI22xp33_ASAP7_75t_SL g862 ( .A1(n_39), .A2(n_202), .B1(n_601), .B2(n_863), .Y(n_862) );
XNOR2xp5_ASAP7_75t_L g924 ( .A(n_40), .B(n_925), .Y(n_924) );
CKINVDCx5p33_ASAP7_75t_R g462 ( .A(n_42), .Y(n_462) );
INVx1_ASAP7_75t_L g318 ( .A(n_43), .Y(n_318) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_44), .A2(n_75), .B1(n_604), .B2(n_606), .Y(n_603) );
AOI22xp33_ASAP7_75t_SL g614 ( .A1(n_44), .A2(n_75), .B1(n_615), .B2(n_616), .Y(n_614) );
INVx1_ASAP7_75t_L g784 ( .A(n_45), .Y(n_784) );
AOI22xp33_ASAP7_75t_L g797 ( .A1(n_45), .A2(n_224), .B1(n_798), .B2(n_801), .Y(n_797) );
CKINVDCx5p33_ASAP7_75t_R g387 ( .A(n_46), .Y(n_387) );
OAI22xp5_ASAP7_75t_L g840 ( .A1(n_47), .A2(n_207), .B1(n_634), .B2(n_841), .Y(n_840) );
OAI22xp33_ASAP7_75t_L g873 ( .A1(n_47), .A2(n_207), .B1(n_594), .B2(n_874), .Y(n_873) );
AOI221xp5_ASAP7_75t_L g738 ( .A1(n_48), .A2(n_69), .B1(n_418), .B2(n_484), .C(n_591), .Y(n_738) );
AOI22xp33_ASAP7_75t_L g748 ( .A1(n_48), .A2(n_69), .B1(n_621), .B2(n_749), .Y(n_748) );
CKINVDCx5p33_ASAP7_75t_R g465 ( .A(n_49), .Y(n_465) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_50), .A2(n_85), .B1(n_601), .B2(n_610), .Y(n_609) );
INVxp67_ASAP7_75t_SL g629 ( .A(n_50), .Y(n_629) );
AOI221xp5_ASAP7_75t_L g1480 ( .A1(n_51), .A2(n_65), .B1(n_601), .B2(n_610), .C(n_961), .Y(n_1480) );
AOI22xp33_ASAP7_75t_L g1457 ( .A1(n_52), .A2(n_136), .B1(n_815), .B2(n_917), .Y(n_1457) );
INVx1_ASAP7_75t_L g1491 ( .A(n_52), .Y(n_1491) );
OAI22xp33_ASAP7_75t_L g893 ( .A1(n_53), .A2(n_199), .B1(n_339), .B2(n_347), .Y(n_893) );
INVxp33_ASAP7_75t_L g1402 ( .A(n_54), .Y(n_1402) );
NAND2xp33_ASAP7_75t_SL g1421 ( .A(n_54), .B(n_1422), .Y(n_1421) );
AOI22xp33_ASAP7_75t_SL g1107 ( .A1(n_55), .A2(n_108), .B1(n_591), .B2(n_1108), .Y(n_1107) );
AOI22xp33_ASAP7_75t_L g1118 ( .A1(n_55), .A2(n_108), .B1(n_1119), .B2(n_1120), .Y(n_1118) );
CKINVDCx5p33_ASAP7_75t_R g473 ( .A(n_56), .Y(n_473) );
XNOR2xp5_ASAP7_75t_L g1443 ( .A(n_57), .B(n_1444), .Y(n_1443) );
INVxp33_ASAP7_75t_L g583 ( .A(n_58), .Y(n_583) );
AO22x2_ASAP7_75t_L g768 ( .A1(n_59), .A2(n_769), .B1(n_829), .B2(n_830), .Y(n_768) );
INVxp67_ASAP7_75t_SL g829 ( .A(n_59), .Y(n_829) );
AOI22xp5_ASAP7_75t_L g1190 ( .A1(n_59), .A2(n_88), .B1(n_1169), .B2(n_1186), .Y(n_1190) );
INVxp33_ASAP7_75t_L g1133 ( .A(n_60), .Y(n_1133) );
CKINVDCx5p33_ASAP7_75t_R g946 ( .A(n_61), .Y(n_946) );
INVx1_ASAP7_75t_L g992 ( .A(n_62), .Y(n_992) );
AOI221xp5_ASAP7_75t_L g1053 ( .A1(n_62), .A2(n_123), .B1(n_811), .B2(n_1054), .C(n_1056), .Y(n_1053) );
AOI22xp5_ASAP7_75t_SL g1180 ( .A1(n_63), .A2(n_80), .B1(n_1163), .B2(n_1169), .Y(n_1180) );
INVx1_ASAP7_75t_L g969 ( .A(n_64), .Y(n_969) );
OAI22xp5_ASAP7_75t_L g1499 ( .A1(n_65), .A2(n_177), .B1(n_569), .B2(n_1500), .Y(n_1499) );
AOI22xp33_ASAP7_75t_L g937 ( .A1(n_66), .A2(n_217), .B1(n_554), .B2(n_912), .Y(n_937) );
OAI211xp5_ASAP7_75t_SL g950 ( .A1(n_66), .A2(n_509), .B(n_951), .C(n_962), .Y(n_950) );
INVx1_ASAP7_75t_L g665 ( .A(n_67), .Y(n_665) );
AOI22xp33_ASAP7_75t_L g699 ( .A1(n_67), .A2(n_185), .B1(n_561), .B2(n_690), .Y(n_699) );
INVx1_ASAP7_75t_L g1430 ( .A(n_68), .Y(n_1430) );
INVxp67_ASAP7_75t_SL g1093 ( .A(n_70), .Y(n_1093) );
AOI22xp33_ASAP7_75t_SL g1111 ( .A1(n_70), .A2(n_105), .B1(n_791), .B2(n_1108), .Y(n_1111) );
INVx1_ASAP7_75t_L g781 ( .A(n_71), .Y(n_781) );
CKINVDCx16_ASAP7_75t_R g1167 ( .A(n_72), .Y(n_1167) );
AOI22xp33_ASAP7_75t_L g677 ( .A1(n_73), .A2(n_196), .B1(n_604), .B2(n_678), .Y(n_677) );
AOI22xp33_ASAP7_75t_L g689 ( .A1(n_73), .A2(n_196), .B1(n_615), .B2(n_690), .Y(n_689) );
INVxp67_ASAP7_75t_SL g642 ( .A(n_74), .Y(n_642) );
OAI22xp5_ASAP7_75t_L g891 ( .A1(n_76), .A2(n_116), .B1(n_329), .B2(n_892), .Y(n_891) );
AOI22xp33_ASAP7_75t_SL g905 ( .A1(n_76), .A2(n_116), .B1(n_856), .B2(n_860), .Y(n_905) );
INVx1_ASAP7_75t_L g890 ( .A(n_77), .Y(n_890) );
OAI222xp33_ASAP7_75t_L g896 ( .A1(n_77), .A2(n_155), .B1(n_167), .B2(n_478), .C1(n_822), .C2(n_897), .Y(n_896) );
AOI22xp33_ASAP7_75t_L g1124 ( .A1(n_78), .A2(n_109), .B1(n_815), .B2(n_917), .Y(n_1124) );
INVxp33_ASAP7_75t_SL g1130 ( .A(n_78), .Y(n_1130) );
OAI221xp5_ASAP7_75t_L g1396 ( .A1(n_79), .A2(n_157), .B1(n_1011), .B2(n_1397), .C(n_1398), .Y(n_1396) );
INVx1_ASAP7_75t_L g1425 ( .A(n_79), .Y(n_1425) );
INVx1_ASAP7_75t_L g943 ( .A(n_81), .Y(n_943) );
AOI221xp5_ASAP7_75t_L g957 ( .A1(n_81), .A2(n_163), .B1(n_611), .B2(n_958), .C(n_961), .Y(n_957) );
AOI221xp5_ASAP7_75t_L g720 ( .A1(n_82), .A2(n_94), .B1(n_721), .B2(n_722), .C(n_724), .Y(n_720) );
INVx1_ASAP7_75t_L g754 ( .A(n_82), .Y(n_754) );
CKINVDCx5p33_ASAP7_75t_R g399 ( .A(n_83), .Y(n_399) );
INVx1_ASAP7_75t_L g1020 ( .A(n_84), .Y(n_1020) );
AOI22xp33_ASAP7_75t_L g1070 ( .A1(n_84), .A2(n_244), .B1(n_747), .B2(n_1071), .Y(n_1070) );
INVxp33_ASAP7_75t_L g636 ( .A(n_85), .Y(n_636) );
INVx1_ASAP7_75t_L g377 ( .A(n_86), .Y(n_377) );
INVx1_ASAP7_75t_L g543 ( .A(n_86), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g865 ( .A1(n_87), .A2(n_144), .B1(n_516), .B2(n_866), .Y(n_865) );
INVx1_ASAP7_75t_L g879 ( .A(n_87), .Y(n_879) );
OAI22xp5_ASAP7_75t_L g1448 ( .A1(n_89), .A2(n_91), .B1(n_545), .B2(n_1449), .Y(n_1448) );
INVx1_ASAP7_75t_L g1482 ( .A(n_89), .Y(n_1482) );
AOI22xp33_ASAP7_75t_SL g851 ( .A1(n_90), .A2(n_125), .B1(n_852), .B2(n_853), .Y(n_851) );
AOI22xp33_ASAP7_75t_L g859 ( .A1(n_90), .A2(n_125), .B1(n_860), .B2(n_861), .Y(n_859) );
INVx1_ASAP7_75t_L g1483 ( .A(n_91), .Y(n_1483) );
CKINVDCx5p33_ASAP7_75t_R g396 ( .A(n_92), .Y(n_396) );
INVx1_ASAP7_75t_L g756 ( .A(n_94), .Y(n_756) );
AOI22xp33_ASAP7_75t_L g1226 ( .A1(n_95), .A2(n_218), .B1(n_1175), .B2(n_1227), .Y(n_1226) );
CKINVDCx20_ASAP7_75t_R g1258 ( .A(n_96), .Y(n_1258) );
CKINVDCx5p33_ASAP7_75t_R g931 ( .A(n_97), .Y(n_931) );
INVxp33_ASAP7_75t_L g1401 ( .A(n_98), .Y(n_1401) );
CKINVDCx5p33_ASAP7_75t_R g929 ( .A(n_99), .Y(n_929) );
INVx1_ASAP7_75t_L g734 ( .A(n_100), .Y(n_734) );
AOI22xp33_ASAP7_75t_L g751 ( .A1(n_100), .A2(n_216), .B1(n_523), .B2(n_691), .Y(n_751) );
AOI22xp33_ASAP7_75t_L g933 ( .A1(n_101), .A2(n_162), .B1(n_909), .B2(n_934), .Y(n_933) );
INVx1_ASAP7_75t_L g975 ( .A(n_101), .Y(n_975) );
AOI22xp33_ASAP7_75t_L g739 ( .A1(n_102), .A2(n_194), .B1(n_718), .B2(n_740), .Y(n_739) );
AOI22xp33_ASAP7_75t_L g746 ( .A1(n_102), .A2(n_194), .B1(n_523), .B2(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g838 ( .A(n_103), .Y(n_838) );
AOI22xp33_ASAP7_75t_L g857 ( .A1(n_103), .A2(n_169), .B1(n_591), .B2(n_601), .Y(n_857) );
NOR2xp33_ASAP7_75t_L g328 ( .A(n_104), .B(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g438 ( .A(n_104), .Y(n_438) );
INVxp33_ASAP7_75t_SL g1087 ( .A(n_105), .Y(n_1087) );
AOI22xp33_ASAP7_75t_L g600 ( .A1(n_106), .A2(n_240), .B1(n_601), .B2(n_602), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g617 ( .A1(n_106), .A2(n_240), .B1(n_358), .B2(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g1462 ( .A(n_107), .Y(n_1462) );
OAI221xp5_ASAP7_75t_L g1484 ( .A1(n_107), .A2(n_507), .B1(n_979), .B2(n_1485), .C(n_1487), .Y(n_1484) );
INVxp67_ASAP7_75t_SL g1131 ( .A(n_109), .Y(n_1131) );
AOI22xp33_ASAP7_75t_L g792 ( .A1(n_110), .A2(n_222), .B1(n_793), .B2(n_794), .Y(n_792) );
AOI22xp33_ASAP7_75t_L g810 ( .A1(n_110), .A2(n_222), .B1(n_690), .B2(n_811), .Y(n_810) );
INVx1_ASAP7_75t_L g255 ( .A(n_111), .Y(n_255) );
OA22x2_ASAP7_75t_L g278 ( .A1(n_112), .A2(n_279), .B1(n_453), .B2(n_454), .Y(n_278) );
INVxp67_ASAP7_75t_SL g454 ( .A(n_112), .Y(n_454) );
INVx1_ASAP7_75t_L g1390 ( .A(n_113), .Y(n_1390) );
CKINVDCx5p33_ASAP7_75t_R g844 ( .A(n_114), .Y(n_844) );
CKINVDCx5p33_ASAP7_75t_R g773 ( .A(n_115), .Y(n_773) );
INVx1_ASAP7_75t_L g658 ( .A(n_117), .Y(n_658) );
AOI22xp33_ASAP7_75t_L g686 ( .A1(n_117), .A2(n_135), .B1(n_601), .B2(n_681), .Y(n_686) );
CKINVDCx5p33_ASAP7_75t_R g1042 ( .A(n_118), .Y(n_1042) );
AOI22xp33_ASAP7_75t_L g717 ( .A1(n_119), .A2(n_198), .B1(n_718), .B2(n_719), .Y(n_717) );
INVx1_ASAP7_75t_L g757 ( .A(n_119), .Y(n_757) );
CKINVDCx5p33_ASAP7_75t_R g1030 ( .A(n_120), .Y(n_1030) );
AOI22xp5_ASAP7_75t_L g1174 ( .A1(n_121), .A2(n_195), .B1(n_1175), .B2(n_1178), .Y(n_1174) );
AOI22xp33_ASAP7_75t_L g812 ( .A1(n_122), .A2(n_227), .B1(n_808), .B2(n_813), .Y(n_812) );
INVx1_ASAP7_75t_L g827 ( .A(n_122), .Y(n_827) );
INVx1_ASAP7_75t_L g1003 ( .A(n_123), .Y(n_1003) );
CKINVDCx5p33_ASAP7_75t_R g488 ( .A(n_124), .Y(n_488) );
OAI221xp5_ASAP7_75t_L g535 ( .A1(n_124), .A2(n_536), .B1(n_544), .B2(n_545), .C(n_548), .Y(n_535) );
CKINVDCx5p33_ASAP7_75t_R g1034 ( .A(n_126), .Y(n_1034) );
AOI22xp33_ASAP7_75t_L g1228 ( .A1(n_127), .A2(n_128), .B1(n_1163), .B2(n_1229), .Y(n_1228) );
INVx1_ASAP7_75t_L g1393 ( .A(n_129), .Y(n_1393) );
INVxp67_ASAP7_75t_SL g592 ( .A(n_130), .Y(n_592) );
CKINVDCx14_ASAP7_75t_R g1195 ( .A(n_131), .Y(n_1195) );
INVx1_ASAP7_75t_L g674 ( .A(n_132), .Y(n_674) );
AOI22xp33_ASAP7_75t_SL g697 ( .A1(n_132), .A2(n_137), .B1(n_516), .B2(n_698), .Y(n_697) );
AOI22xp5_ASAP7_75t_L g1184 ( .A1(n_133), .A2(n_150), .B1(n_1175), .B2(n_1178), .Y(n_1184) );
OAI22xp5_ASAP7_75t_L g727 ( .A1(n_134), .A2(n_190), .B1(n_728), .B2(n_732), .Y(n_727) );
INVx1_ASAP7_75t_L g762 ( .A(n_134), .Y(n_762) );
INVx1_ASAP7_75t_L g650 ( .A(n_135), .Y(n_650) );
INVx1_ASAP7_75t_L g1494 ( .A(n_136), .Y(n_1494) );
INVx1_ASAP7_75t_L g669 ( .A(n_137), .Y(n_669) );
INVx1_ASAP7_75t_L g766 ( .A(n_138), .Y(n_766) );
AOI22xp33_ASAP7_75t_L g867 ( .A1(n_139), .A2(n_210), .B1(n_868), .B2(n_869), .Y(n_867) );
INVx1_ASAP7_75t_L g876 ( .A(n_139), .Y(n_876) );
INVx1_ASAP7_75t_L g900 ( .A(n_140), .Y(n_900) );
AOI22xp33_ASAP7_75t_L g916 ( .A1(n_140), .A2(n_143), .B1(n_815), .B2(n_917), .Y(n_916) );
AOI22xp33_ASAP7_75t_L g679 ( .A1(n_141), .A2(n_165), .B1(n_680), .B2(n_681), .Y(n_679) );
AOI22xp33_ASAP7_75t_L g692 ( .A1(n_141), .A2(n_165), .B1(n_516), .B2(n_618), .Y(n_692) );
CKINVDCx5p33_ASAP7_75t_R g475 ( .A(n_142), .Y(n_475) );
INVx1_ASAP7_75t_L g901 ( .A(n_143), .Y(n_901) );
INVx1_ASAP7_75t_L g872 ( .A(n_144), .Y(n_872) );
INVxp33_ASAP7_75t_SL g1088 ( .A(n_145), .Y(n_1088) );
AOI22xp33_ASAP7_75t_SL g1109 ( .A1(n_145), .A2(n_178), .B1(n_1103), .B2(n_1110), .Y(n_1109) );
INVx1_ASAP7_75t_L g531 ( .A(n_146), .Y(n_531) );
AOI22x1_ASAP7_75t_SL g880 ( .A1(n_147), .A2(n_881), .B1(n_918), .B2(n_919), .Y(n_880) );
INVx1_ASAP7_75t_L g918 ( .A(n_147), .Y(n_918) );
AO221x2_ASAP7_75t_L g1192 ( .A1(n_147), .A2(n_230), .B1(n_1169), .B2(n_1186), .C(n_1193), .Y(n_1192) );
INVx1_ASAP7_75t_L g948 ( .A(n_148), .Y(n_948) );
CKINVDCx16_ASAP7_75t_R g1170 ( .A(n_149), .Y(n_1170) );
INVxp33_ASAP7_75t_L g1383 ( .A(n_151), .Y(n_1383) );
CKINVDCx5p33_ASAP7_75t_R g997 ( .A(n_152), .Y(n_997) );
INVx1_ASAP7_75t_L g885 ( .A(n_153), .Y(n_885) );
AOI22xp33_ASAP7_75t_L g906 ( .A1(n_153), .A2(n_199), .B1(n_681), .B2(n_790), .Y(n_906) );
HB1xp67_ASAP7_75t_L g257 ( .A(n_154), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g1150 ( .A(n_154), .B(n_255), .Y(n_1150) );
AND3x2_ASAP7_75t_L g1166 ( .A(n_154), .B(n_255), .C(n_1153), .Y(n_1166) );
AOI22xp5_ASAP7_75t_SL g1202 ( .A1(n_156), .A2(n_166), .B1(n_1163), .B2(n_1169), .Y(n_1202) );
INVx1_ASAP7_75t_L g1427 ( .A(n_157), .Y(n_1427) );
CKINVDCx5p33_ASAP7_75t_R g319 ( .A(n_158), .Y(n_319) );
INVx2_ASAP7_75t_L g268 ( .A(n_159), .Y(n_268) );
AOI22xp5_ASAP7_75t_SL g1201 ( .A1(n_160), .A2(n_225), .B1(n_1175), .B2(n_1178), .Y(n_1201) );
CKINVDCx5p33_ASAP7_75t_R g653 ( .A(n_161), .Y(n_653) );
INVx1_ASAP7_75t_L g977 ( .A(n_162), .Y(n_977) );
INVx1_ASAP7_75t_L g945 ( .A(n_163), .Y(n_945) );
AOI22xp33_ASAP7_75t_L g1102 ( .A1(n_164), .A2(n_181), .B1(n_1103), .B2(n_1105), .Y(n_1102) );
AOI22xp33_ASAP7_75t_L g1113 ( .A1(n_164), .A2(n_181), .B1(n_1114), .B2(n_1116), .Y(n_1113) );
CKINVDCx5p33_ASAP7_75t_R g889 ( .A(n_167), .Y(n_889) );
INVx1_ASAP7_75t_L g1153 ( .A(n_168), .Y(n_1153) );
INVx1_ASAP7_75t_L g843 ( .A(n_169), .Y(n_843) );
CKINVDCx16_ASAP7_75t_R g572 ( .A(n_170), .Y(n_572) );
INVx1_ASAP7_75t_L g846 ( .A(n_171), .Y(n_846) );
AO221x2_ASAP7_75t_L g1255 ( .A1(n_173), .A2(n_248), .B1(n_1229), .B2(n_1256), .C(n_1257), .Y(n_1255) );
AOI22x1_ASAP7_75t_L g1369 ( .A1(n_173), .A2(n_1370), .B1(n_1371), .B2(n_1432), .Y(n_1369) );
INVx1_ASAP7_75t_L g1432 ( .A(n_173), .Y(n_1432) );
AOI22xp33_ASAP7_75t_L g1437 ( .A1(n_173), .A2(n_1438), .B1(n_1442), .B2(n_1506), .Y(n_1437) );
INVx1_ASAP7_75t_L g1471 ( .A(n_174), .Y(n_1471) );
AOI22xp33_ASAP7_75t_SL g903 ( .A1(n_175), .A2(n_220), .B1(n_484), .B2(n_681), .Y(n_903) );
AOI22xp33_ASAP7_75t_L g911 ( .A1(n_175), .A2(n_220), .B1(n_813), .B2(n_912), .Y(n_911) );
INVx1_ASAP7_75t_L g1023 ( .A(n_176), .Y(n_1023) );
AOI221xp5_ASAP7_75t_L g1066 ( .A1(n_176), .A2(n_241), .B1(n_811), .B2(n_1067), .C(n_1069), .Y(n_1066) );
INVx1_ASAP7_75t_L g1479 ( .A(n_177), .Y(n_1479) );
INVxp33_ASAP7_75t_L g1091 ( .A(n_178), .Y(n_1091) );
INVx1_ASAP7_75t_L g270 ( .A(n_179), .Y(n_270) );
INVx2_ASAP7_75t_L g290 ( .A(n_179), .Y(n_290) );
AOI22xp33_ASAP7_75t_L g1466 ( .A1(n_180), .A2(n_208), .B1(n_1467), .B2(n_1469), .Y(n_1466) );
OAI22xp5_ASAP7_75t_L g1495 ( .A1(n_180), .A2(n_208), .B1(n_981), .B2(n_1496), .Y(n_1495) );
CKINVDCx14_ASAP7_75t_R g1260 ( .A(n_182), .Y(n_1260) );
CKINVDCx5p33_ASAP7_75t_R g1455 ( .A(n_183), .Y(n_1455) );
INVx1_ASAP7_75t_L g467 ( .A(n_184), .Y(n_467) );
AOI221xp5_ASAP7_75t_L g515 ( .A1(n_184), .A2(n_211), .B1(n_516), .B2(n_518), .C(n_521), .Y(n_515) );
INVx1_ASAP7_75t_L g664 ( .A(n_185), .Y(n_664) );
CKINVDCx5p33_ASAP7_75t_R g284 ( .A(n_186), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g709 ( .A(n_187), .B(n_710), .Y(n_709) );
XNOR2xp5_ASAP7_75t_L g987 ( .A(n_188), .B(n_988), .Y(n_987) );
XNOR2x1_ASAP7_75t_L g1137 ( .A(n_188), .B(n_988), .Y(n_1137) );
INVxp33_ASAP7_75t_L g1380 ( .A(n_189), .Y(n_1380) );
INVx1_ASAP7_75t_L g760 ( .A(n_190), .Y(n_760) );
CKINVDCx16_ASAP7_75t_R g1160 ( .A(n_191), .Y(n_1160) );
INVx1_ASAP7_75t_L g783 ( .A(n_192), .Y(n_783) );
AOI22xp33_ASAP7_75t_L g802 ( .A1(n_192), .A2(n_203), .B1(n_790), .B2(n_791), .Y(n_802) );
INVx1_ASAP7_75t_L g1465 ( .A(n_197), .Y(n_1465) );
OAI211xp5_ASAP7_75t_SL g1473 ( .A1(n_197), .A2(n_509), .B(n_1474), .C(n_1481), .Y(n_1473) );
INVx1_ASAP7_75t_L g753 ( .A(n_198), .Y(n_753) );
CKINVDCx5p33_ASAP7_75t_R g477 ( .A(n_200), .Y(n_477) );
INVx1_ASAP7_75t_L g410 ( .A(n_201), .Y(n_410) );
INVx1_ASAP7_75t_L g776 ( .A(n_203), .Y(n_776) );
INVx1_ASAP7_75t_L g487 ( .A(n_204), .Y(n_487) );
HB1xp67_ASAP7_75t_L g544 ( .A(n_204), .Y(n_544) );
OAI211xp5_ASAP7_75t_L g355 ( .A1(n_205), .A2(n_356), .B(n_361), .C(n_372), .Y(n_355) );
INVx1_ASAP7_75t_L g445 ( .A(n_205), .Y(n_445) );
INVx1_ASAP7_75t_L g584 ( .A(n_206), .Y(n_584) );
INVx1_ASAP7_75t_L g668 ( .A(n_209), .Y(n_668) );
INVx1_ASAP7_75t_L g877 ( .A(n_210), .Y(n_877) );
AOI21xp33_ASAP7_75t_L g469 ( .A1(n_211), .A2(n_418), .B(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g1154 ( .A(n_212), .Y(n_1154) );
NAND2xp5_ASAP7_75t_L g1159 ( .A(n_212), .B(n_1152), .Y(n_1159) );
INVx1_ASAP7_75t_L g825 ( .A(n_214), .Y(n_825) );
INVx1_ASAP7_75t_L g1094 ( .A(n_215), .Y(n_1094) );
OAI22xp5_ASAP7_75t_L g1128 ( .A1(n_215), .A2(n_234), .B1(n_594), .B2(n_822), .Y(n_1128) );
INVx1_ASAP7_75t_L g735 ( .A(n_216), .Y(n_735) );
OAI221xp5_ASAP7_75t_L g966 ( .A1(n_217), .A2(n_507), .B1(n_967), .B2(n_974), .C(n_979), .Y(n_966) );
INVx1_ASAP7_75t_L g1090 ( .A(n_219), .Y(n_1090) );
OAI211xp5_ASAP7_75t_L g300 ( .A1(n_221), .A2(n_301), .B(n_306), .C(n_313), .Y(n_300) );
INVx1_ASAP7_75t_L g406 ( .A(n_221), .Y(n_406) );
INVx1_ASAP7_75t_L g578 ( .A(n_223), .Y(n_578) );
INVx1_ASAP7_75t_L g774 ( .A(n_224), .Y(n_774) );
CKINVDCx5p33_ASAP7_75t_R g1456 ( .A(n_226), .Y(n_1456) );
INVx1_ASAP7_75t_L g819 ( .A(n_227), .Y(n_819) );
INVx1_ASAP7_75t_L g1395 ( .A(n_228), .Y(n_1395) );
INVx2_ASAP7_75t_L g267 ( .A(n_229), .Y(n_267) );
CKINVDCx5p33_ASAP7_75t_R g1032 ( .A(n_231), .Y(n_1032) );
OAI221xp5_ASAP7_75t_L g1005 ( .A1(n_232), .A2(n_233), .B1(n_1006), .B2(n_1011), .C(n_1013), .Y(n_1005) );
OAI22xp5_ASAP7_75t_L g1047 ( .A1(n_232), .A2(n_233), .B1(n_1048), .B2(n_1051), .Y(n_1047) );
INVx1_ASAP7_75t_L g1095 ( .A(n_234), .Y(n_1095) );
INVx1_ASAP7_75t_L g654 ( .A(n_235), .Y(n_654) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_235), .A2(n_237), .B1(n_604), .B2(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g726 ( .A(n_236), .Y(n_726) );
AOI22xp33_ASAP7_75t_L g750 ( .A1(n_236), .A2(n_245), .B1(n_549), .B2(n_554), .Y(n_750) );
INVx1_ASAP7_75t_L g651 ( .A(n_237), .Y(n_651) );
CKINVDCx20_ASAP7_75t_R g1155 ( .A(n_238), .Y(n_1155) );
CKINVDCx5p33_ASAP7_75t_R g391 ( .A(n_239), .Y(n_391) );
INVx1_ASAP7_75t_L g1025 ( .A(n_241), .Y(n_1025) );
INVx1_ASAP7_75t_L g337 ( .A(n_242), .Y(n_337) );
BUFx3_ASAP7_75t_L g353 ( .A(n_242), .Y(n_353) );
BUFx3_ASAP7_75t_L g336 ( .A(n_243), .Y(n_336) );
INVx1_ASAP7_75t_L g346 ( .A(n_243), .Y(n_346) );
INVx1_ASAP7_75t_L g1027 ( .A(n_244), .Y(n_1027) );
INVx1_ASAP7_75t_L g737 ( .A(n_245), .Y(n_737) );
CKINVDCx5p33_ASAP7_75t_R g942 ( .A(n_246), .Y(n_942) );
CKINVDCx5p33_ASAP7_75t_R g365 ( .A(n_247), .Y(n_365) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_271), .B(n_1140), .Y(n_249) );
INVx2_ASAP7_75t_SL g250 ( .A(n_251), .Y(n_250) );
INVx1_ASAP7_75t_SL g251 ( .A(n_252), .Y(n_251) );
AND2x4_ASAP7_75t_L g252 ( .A(n_253), .B(n_258), .Y(n_252) );
AND2x4_ASAP7_75t_L g1436 ( .A(n_253), .B(n_259), .Y(n_1436) );
NOR2xp33_ASAP7_75t_SL g253 ( .A(n_254), .B(n_256), .Y(n_253) );
INVx1_ASAP7_75t_SL g1441 ( .A(n_254), .Y(n_1441) );
NAND2xp5_ASAP7_75t_L g1512 ( .A(n_254), .B(n_256), .Y(n_1512) );
HB1xp67_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g1440 ( .A(n_256), .B(n_1441), .Y(n_1440) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_260), .B(n_264), .Y(n_259) );
INVxp67_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
OR2x2_ASAP7_75t_L g280 ( .A(n_261), .B(n_281), .Y(n_280) );
OR2x6_ASAP7_75t_L g575 ( .A(n_261), .B(n_281), .Y(n_575) );
HB1xp67_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g599 ( .A(n_262), .B(n_270), .Y(n_599) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
OR2x2_ASAP7_75t_L g418 ( .A(n_263), .B(n_289), .Y(n_418) );
INVx8_ASAP7_75t_L g283 ( .A(n_264), .Y(n_283) );
OR2x6_ASAP7_75t_L g264 ( .A(n_265), .B(n_269), .Y(n_264) );
BUFx6f_ASAP7_75t_L g420 ( .A(n_265), .Y(n_420) );
OR2x6_ASAP7_75t_L g586 ( .A(n_265), .B(n_288), .Y(n_586) );
INVx1_ASAP7_75t_L g971 ( .A(n_265), .Y(n_971) );
INVx2_ASAP7_75t_SL g1019 ( .A(n_265), .Y(n_1019) );
OR2x2_ASAP7_75t_L g1040 ( .A(n_265), .B(n_1010), .Y(n_1040) );
BUFx6f_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_267), .B(n_268), .Y(n_266) );
INVx2_ASAP7_75t_L g293 ( .A(n_267), .Y(n_293) );
AND2x4_ASAP7_75t_L g298 ( .A(n_267), .B(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g305 ( .A(n_267), .Y(n_305) );
INVx1_ASAP7_75t_L g312 ( .A(n_267), .Y(n_312) );
AND2x2_ASAP7_75t_L g317 ( .A(n_267), .B(n_268), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_268), .B(n_293), .Y(n_292) );
INVx2_ASAP7_75t_L g299 ( .A(n_268), .Y(n_299) );
INVx1_ASAP7_75t_L g304 ( .A(n_268), .Y(n_304) );
INVx1_ASAP7_75t_L g321 ( .A(n_268), .Y(n_321) );
INVx1_ASAP7_75t_L g501 ( .A(n_268), .Y(n_501) );
AND2x4_ASAP7_75t_L g320 ( .A(n_269), .B(n_321), .Y(n_320) );
INVx2_ASAP7_75t_SL g269 ( .A(n_270), .Y(n_269) );
OR2x2_ASAP7_75t_L g822 ( .A(n_270), .B(n_324), .Y(n_822) );
OR2x2_ASAP7_75t_L g874 ( .A(n_270), .B(n_324), .Y(n_874) );
OAI22xp33_ASAP7_75t_L g271 ( .A1(n_272), .A2(n_273), .B1(n_921), .B2(n_1139), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
XNOR2xp5_ASAP7_75t_L g273 ( .A(n_274), .B(n_703), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
XNOR2x1_ASAP7_75t_L g276 ( .A(n_277), .B(n_570), .Y(n_276) );
XNOR2x1_ASAP7_75t_L g277 ( .A(n_278), .B(n_455), .Y(n_277) );
INVx1_ASAP7_75t_L g453 ( .A(n_279), .Y(n_453) );
OAI211xp5_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_282), .B(n_327), .C(n_380), .Y(n_279) );
AOI31xp33_ASAP7_75t_L g817 ( .A1(n_280), .A2(n_818), .A3(n_823), .B(n_826), .Y(n_817) );
AOI31xp33_ASAP7_75t_L g1125 ( .A1(n_280), .A2(n_1126), .A3(n_1129), .B(n_1132), .Y(n_1125) );
AND2x4_ASAP7_75t_L g413 ( .A(n_281), .B(n_414), .Y(n_413) );
AND2x4_ASAP7_75t_L g562 ( .A(n_281), .B(n_563), .Y(n_562) );
AND2x4_ASAP7_75t_L g626 ( .A(n_281), .B(n_414), .Y(n_626) );
AOI211xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_284), .B(n_285), .C(n_300), .Y(n_282) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_283), .A2(n_583), .B1(n_584), .B2(n_585), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g673 ( .A1(n_283), .A2(n_585), .B1(n_653), .B2(n_674), .Y(n_673) );
AOI22xp33_ASAP7_75t_L g826 ( .A1(n_283), .A2(n_773), .B1(n_827), .B2(n_828), .Y(n_826) );
AOI22xp33_ASAP7_75t_SL g878 ( .A1(n_283), .A2(n_828), .B1(n_844), .B2(n_879), .Y(n_878) );
AOI22xp33_ASAP7_75t_SL g1132 ( .A1(n_283), .A2(n_828), .B1(n_1090), .B2(n_1133), .Y(n_1132) );
OAI22xp33_ASAP7_75t_L g403 ( .A1(n_284), .A2(n_397), .B1(n_404), .B2(n_406), .Y(n_403) );
OR2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_291), .Y(n_286) );
AOI322xp5_ASAP7_75t_L g313 ( .A1(n_287), .A2(n_314), .A3(n_318), .B1(n_319), .B2(n_320), .C1(n_322), .C2(n_326), .Y(n_313) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x4_ASAP7_75t_L g295 ( .A(n_288), .B(n_296), .Y(n_295) );
AND2x4_ASAP7_75t_L g579 ( .A(n_288), .B(n_499), .Y(n_579) );
AND2x4_ASAP7_75t_L g581 ( .A(n_288), .B(n_296), .Y(n_581) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g310 ( .A(n_290), .Y(n_310) );
INVx2_ASAP7_75t_L g426 ( .A(n_291), .Y(n_426) );
BUFx2_ASAP7_75t_L g1026 ( .A(n_291), .Y(n_1026) );
BUFx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
INVx1_ASAP7_75t_L g433 ( .A(n_292), .Y(n_433) );
INVx1_ASAP7_75t_L g461 ( .A(n_292), .Y(n_461) );
INVx1_ASAP7_75t_L g490 ( .A(n_293), .Y(n_490) );
AND2x4_ASAP7_75t_L g499 ( .A(n_293), .B(n_500), .Y(n_499) );
INVx5_ASAP7_75t_SL g294 ( .A(n_295), .Y(n_294) );
AOI22xp33_ASAP7_75t_L g823 ( .A1(n_295), .A2(n_579), .B1(n_824), .B2(n_825), .Y(n_823) );
AOI22xp33_ASAP7_75t_SL g875 ( .A1(n_295), .A2(n_579), .B1(n_876), .B2(n_877), .Y(n_875) );
AOI22xp5_ASAP7_75t_L g899 ( .A1(n_295), .A2(n_579), .B1(n_900), .B2(n_901), .Y(n_899) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g429 ( .A(n_298), .Y(n_429) );
INVx3_ASAP7_75t_L g437 ( .A(n_298), .Y(n_437) );
BUFx6f_ASAP7_75t_L g796 ( .A(n_298), .Y(n_796) );
AND2x4_ASAP7_75t_L g311 ( .A(n_299), .B(n_312), .Y(n_311) );
OAI22xp33_ASAP7_75t_L g1386 ( .A1(n_301), .A2(n_1387), .B1(n_1389), .B2(n_1390), .Y(n_1386) );
OAI221xp5_ASAP7_75t_L g1485 ( .A1(n_301), .A2(n_973), .B1(n_1455), .B2(n_1456), .C(n_1486), .Y(n_1485) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
BUFx2_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVx2_ASAP7_75t_L g423 ( .A(n_303), .Y(n_423) );
INVx3_ASAP7_75t_L g468 ( .A(n_303), .Y(n_468) );
INVx2_ASAP7_75t_L g478 ( .A(n_303), .Y(n_478) );
AND2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_305), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_304), .B(n_305), .Y(n_444) );
INVx1_ASAP7_75t_L g324 ( .A(n_305), .Y(n_324) );
NAND4xp25_ASAP7_75t_SL g576 ( .A(n_306), .B(n_577), .C(n_582), .D(n_587), .Y(n_576) );
NAND4xp25_ASAP7_75t_SL g662 ( .A(n_306), .B(n_663), .C(n_666), .D(n_673), .Y(n_662) );
CKINVDCx11_ASAP7_75t_R g306 ( .A(n_307), .Y(n_306) );
AOI211xp5_ASAP7_75t_L g818 ( .A1(n_307), .A2(n_722), .B(n_819), .C(n_820), .Y(n_818) );
AOI211xp5_ASAP7_75t_L g871 ( .A1(n_307), .A2(n_791), .B(n_872), .C(n_873), .Y(n_871) );
NOR3xp33_ASAP7_75t_L g895 ( .A(n_307), .B(n_896), .C(n_898), .Y(n_895) );
AOI211xp5_ASAP7_75t_L g1126 ( .A1(n_307), .A2(n_722), .B(n_1127), .C(n_1128), .Y(n_1126) );
AND2x4_ASAP7_75t_L g307 ( .A(n_308), .B(n_311), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVxp67_ASAP7_75t_L g325 ( .A(n_309), .Y(n_325) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
NAND2x1p5_ASAP7_75t_L g451 ( .A(n_310), .B(n_452), .Y(n_451) );
BUFx3_ASAP7_75t_L g511 ( .A(n_311), .Y(n_511) );
BUFx6f_ASAP7_75t_L g591 ( .A(n_311), .Y(n_591) );
BUFx6f_ASAP7_75t_L g611 ( .A(n_311), .Y(n_611) );
BUFx2_ASAP7_75t_L g672 ( .A(n_311), .Y(n_672) );
BUFx3_ASAP7_75t_L g999 ( .A(n_311), .Y(n_999) );
INVx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx2_ASAP7_75t_L g680 ( .A(n_315), .Y(n_680) );
INVx3_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
BUFx6f_ASAP7_75t_L g484 ( .A(n_316), .Y(n_484) );
AND2x4_ASAP7_75t_L g508 ( .A(n_316), .B(n_498), .Y(n_508) );
BUFx2_ASAP7_75t_L g721 ( .A(n_316), .Y(n_721) );
BUFx6f_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx3_ASAP7_75t_L g471 ( .A(n_317), .Y(n_471) );
AOI322xp5_ASAP7_75t_L g361 ( .A1(n_319), .A2(n_326), .A3(n_362), .B1(n_364), .B2(n_365), .C1(n_366), .C2(n_370), .Y(n_361) );
INVx2_ASAP7_75t_L g594 ( .A(n_320), .Y(n_594) );
AOI222xp33_ASAP7_75t_L g666 ( .A1(n_320), .A2(n_322), .B1(n_667), .B2(n_668), .C1(n_669), .C2(n_670), .Y(n_666) );
INVx2_ASAP7_75t_L g821 ( .A(n_320), .Y(n_821) );
INVx2_ASAP7_75t_L g897 ( .A(n_320), .Y(n_897) );
AOI22xp5_ASAP7_75t_L g486 ( .A1(n_321), .A2(n_487), .B1(n_488), .B2(n_489), .Y(n_486) );
INVx1_ASAP7_75t_L g730 ( .A(n_321), .Y(n_730) );
HB1xp67_ASAP7_75t_L g964 ( .A(n_321), .Y(n_964) );
AOI222xp33_ASAP7_75t_L g587 ( .A1(n_322), .A2(n_588), .B1(n_589), .B2(n_592), .C1(n_593), .C2(n_595), .Y(n_587) );
AND2x4_ASAP7_75t_L g322 ( .A(n_323), .B(n_325), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
OAI31xp33_ASAP7_75t_SL g327 ( .A1(n_328), .A2(n_338), .A3(n_355), .B(n_375), .Y(n_327) );
INVx4_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
AOI22xp33_ASAP7_75t_L g639 ( .A1(n_330), .A2(n_640), .B1(n_641), .B2(n_642), .Y(n_639) );
AOI22xp33_ASAP7_75t_L g648 ( .A1(n_330), .A2(n_649), .B1(n_650), .B2(n_651), .Y(n_648) );
AOI22xp33_ASAP7_75t_L g772 ( .A1(n_330), .A2(n_348), .B1(n_773), .B2(n_774), .Y(n_772) );
AOI22xp33_ASAP7_75t_L g845 ( .A1(n_330), .A2(n_640), .B1(n_846), .B2(n_847), .Y(n_845) );
AOI22xp33_ASAP7_75t_L g1089 ( .A1(n_330), .A2(n_348), .B1(n_1090), .B2(n_1091), .Y(n_1089) );
AND2x6_ASAP7_75t_L g330 ( .A(n_331), .B(n_334), .Y(n_330) );
AND2x4_ASAP7_75t_L g637 ( .A(n_331), .B(n_638), .Y(n_637) );
AND2x4_ASAP7_75t_L g649 ( .A(n_331), .B(n_638), .Y(n_649) );
INVx1_ASAP7_75t_SL g331 ( .A(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g632 ( .A(n_332), .B(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g342 ( .A(n_333), .Y(n_342) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_333), .Y(n_350) );
AND2x2_ASAP7_75t_L g384 ( .A(n_333), .B(n_377), .Y(n_384) );
INVx2_ASAP7_75t_L g415 ( .A(n_333), .Y(n_415) );
INVx1_ASAP7_75t_L g411 ( .A(n_334), .Y(n_411) );
HB1xp67_ASAP7_75t_L g616 ( .A(n_334), .Y(n_616) );
BUFx6f_ASAP7_75t_L g625 ( .A(n_334), .Y(n_625) );
INVx2_ASAP7_75t_L g935 ( .A(n_334), .Y(n_935) );
INVx1_ASAP7_75t_L g1117 ( .A(n_334), .Y(n_1117) );
BUFx6f_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx2_ASAP7_75t_L g394 ( .A(n_335), .Y(n_394) );
INVx1_ASAP7_75t_L g524 ( .A(n_335), .Y(n_524) );
INVx1_ASAP7_75t_L g567 ( .A(n_335), .Y(n_567) );
BUFx6f_ASAP7_75t_L g691 ( .A(n_335), .Y(n_691) );
AND2x4_ASAP7_75t_L g335 ( .A(n_336), .B(n_337), .Y(n_335) );
INVx2_ASAP7_75t_L g354 ( .A(n_336), .Y(n_354) );
AND2x2_ASAP7_75t_L g360 ( .A(n_336), .B(n_353), .Y(n_360) );
INVx1_ASAP7_75t_L g344 ( .A(n_337), .Y(n_344) );
OR2x2_ASAP7_75t_L g339 ( .A(n_340), .B(n_343), .Y(n_339) );
INVx1_ASAP7_75t_L g364 ( .A(n_340), .Y(n_364) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
AND2x2_ASAP7_75t_L g357 ( .A(n_341), .B(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g374 ( .A(n_341), .Y(n_374) );
AND2x6_ASAP7_75t_L g640 ( .A(n_341), .B(n_363), .Y(n_640) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
AND2x6_ASAP7_75t_L g370 ( .A(n_342), .B(n_371), .Y(n_370) );
INVx2_ASAP7_75t_L g398 ( .A(n_343), .Y(n_398) );
BUFx2_ASAP7_75t_L g1059 ( .A(n_343), .Y(n_1059) );
OR2x2_ASAP7_75t_L g1077 ( .A(n_343), .B(n_558), .Y(n_1077) );
INVx1_ASAP7_75t_L g1454 ( .A(n_343), .Y(n_1454) );
OR2x2_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
AND2x2_ASAP7_75t_L g402 ( .A(n_344), .B(n_345), .Y(n_402) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
AND2x4_ASAP7_75t_L g363 ( .A(n_346), .B(n_353), .Y(n_363) );
INVx4_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
AOI22xp33_ASAP7_75t_L g635 ( .A1(n_348), .A2(n_584), .B1(n_636), .B2(n_637), .Y(n_635) );
AOI221xp5_ASAP7_75t_L g652 ( .A1(n_348), .A2(n_640), .B1(n_653), .B2(n_654), .C(n_655), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g842 ( .A1(n_348), .A2(n_649), .B1(n_843), .B2(n_844), .Y(n_842) );
AND2x4_ASAP7_75t_L g348 ( .A(n_349), .B(n_351), .Y(n_348) );
AND2x2_ASAP7_75t_SL g366 ( .A(n_349), .B(n_367), .Y(n_366) );
AND2x4_ASAP7_75t_L g780 ( .A(n_349), .B(n_367), .Y(n_780) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx6_ASAP7_75t_L g520 ( .A(n_351), .Y(n_520) );
INVx2_ASAP7_75t_L g555 ( .A(n_351), .Y(n_555) );
AND2x2_ASAP7_75t_L g563 ( .A(n_351), .B(n_541), .Y(n_563) );
BUFx2_ASAP7_75t_L g621 ( .A(n_351), .Y(n_621) );
AND2x4_ASAP7_75t_L g351 ( .A(n_352), .B(n_354), .Y(n_351) );
INVx1_ASAP7_75t_L g371 ( .A(n_352), .Y(n_371) );
INVx2_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g369 ( .A(n_354), .Y(n_369) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AOI211xp5_ASAP7_75t_L g628 ( .A1(n_357), .A2(n_373), .B(n_629), .C(n_630), .Y(n_628) );
HB1xp67_ASAP7_75t_L g777 ( .A(n_358), .Y(n_777) );
HB1xp67_ASAP7_75t_L g839 ( .A(n_358), .Y(n_839) );
HB1xp67_ASAP7_75t_L g1120 ( .A(n_358), .Y(n_1120) );
BUFx6f_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
AND2x4_ASAP7_75t_L g373 ( .A(n_359), .B(n_374), .Y(n_373) );
INVx2_ASAP7_75t_L g517 ( .A(n_359), .Y(n_517) );
BUFx6f_ASAP7_75t_L g659 ( .A(n_359), .Y(n_659) );
INVx1_ASAP7_75t_L g765 ( .A(n_359), .Y(n_765) );
BUFx6f_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
BUFx6f_ASAP7_75t_L g550 ( .A(n_360), .Y(n_550) );
INVx2_ASAP7_75t_L g390 ( .A(n_362), .Y(n_390) );
BUFx6f_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx2_ASAP7_75t_SL g409 ( .A(n_363), .Y(n_409) );
BUFx6f_ASAP7_75t_L g523 ( .A(n_363), .Y(n_523) );
BUFx2_ASAP7_75t_L g615 ( .A(n_363), .Y(n_615) );
BUFx6f_ASAP7_75t_L g816 ( .A(n_363), .Y(n_816) );
BUFx3_ASAP7_75t_L g1115 ( .A(n_363), .Y(n_1115) );
BUFx6f_ASAP7_75t_L g1468 ( .A(n_363), .Y(n_1468) );
OAI22xp5_ASAP7_75t_L g430 ( .A1(n_365), .A2(n_431), .B1(n_434), .B2(n_438), .Y(n_430) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g633 ( .A(n_368), .Y(n_633) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g538 ( .A(n_369), .Y(n_538) );
INVx3_ASAP7_75t_L g634 ( .A(n_370), .Y(n_634) );
AOI222xp33_ASAP7_75t_L g775 ( .A1(n_370), .A2(n_776), .B1(n_777), .B2(n_778), .C1(n_779), .C2(n_781), .Y(n_775) );
AOI22xp33_ASAP7_75t_L g888 ( .A1(n_370), .A2(n_780), .B1(n_889), .B2(n_890), .Y(n_888) );
AOI222xp33_ASAP7_75t_L g1092 ( .A1(n_370), .A2(n_780), .B1(n_912), .B2(n_1093), .C1(n_1094), .C2(n_1095), .Y(n_1092) );
BUFx3_ASAP7_75t_L g547 ( .A(n_371), .Y(n_547) );
NAND3xp33_ASAP7_75t_L g883 ( .A(n_372), .B(n_884), .C(n_888), .Y(n_883) );
CKINVDCx8_ASAP7_75t_R g372 ( .A(n_373), .Y(n_372) );
INVx5_ASAP7_75t_L g771 ( .A(n_373), .Y(n_771) );
AOI211xp5_ASAP7_75t_L g837 ( .A1(n_373), .A2(n_838), .B(n_839), .C(n_840), .Y(n_837) );
OAI21xp33_ASAP7_75t_L g657 ( .A1(n_374), .A2(n_658), .B(n_659), .Y(n_657) );
INVx1_ASAP7_75t_SL g643 ( .A(n_375), .Y(n_643) );
OAI31xp33_ASAP7_75t_L g882 ( .A1(n_375), .A2(n_883), .A3(n_891), .B(n_893), .Y(n_882) );
AND2x4_ASAP7_75t_L g375 ( .A(n_376), .B(n_378), .Y(n_375) );
AND2x4_ASAP7_75t_L g661 ( .A(n_376), .B(n_378), .Y(n_661) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
AND2x4_ASAP7_75t_L g414 ( .A(n_377), .B(n_415), .Y(n_414) );
INVx2_ASAP7_75t_L g983 ( .A(n_378), .Y(n_983) );
BUFx2_ASAP7_75t_L g1081 ( .A(n_378), .Y(n_1081) );
BUFx2_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx2_ASAP7_75t_L g385 ( .A(n_379), .Y(n_385) );
OR2x6_ASAP7_75t_L g417 ( .A(n_379), .B(n_418), .Y(n_417) );
NOR2xp33_ASAP7_75t_L g380 ( .A(n_381), .B(n_416), .Y(n_380) );
OAI33xp33_ASAP7_75t_L g381 ( .A1(n_382), .A2(n_386), .A3(n_395), .B1(n_403), .B2(n_407), .B3(n_412), .Y(n_381) );
INVx1_ASAP7_75t_SL g613 ( .A(n_382), .Y(n_613) );
OR2x2_ASAP7_75t_L g382 ( .A(n_383), .B(n_385), .Y(n_382) );
OR2x6_ASAP7_75t_L g526 ( .A(n_383), .B(n_385), .Y(n_526) );
INVx2_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g695 ( .A(n_384), .Y(n_695) );
INVx2_ASAP7_75t_SL g1069 ( .A(n_384), .Y(n_1069) );
BUFx3_ASAP7_75t_L g1414 ( .A(n_384), .Y(n_1414) );
INVx2_ASAP7_75t_L g513 ( .A(n_385), .Y(n_513) );
AND2x4_ASAP7_75t_L g598 ( .A(n_385), .B(n_599), .Y(n_598) );
OR2x2_ASAP7_75t_L g694 ( .A(n_385), .B(n_695), .Y(n_694) );
AND2x4_ASAP7_75t_L g788 ( .A(n_385), .B(n_599), .Y(n_788) );
BUFx2_ASAP7_75t_L g1497 ( .A(n_385), .Y(n_1497) );
OAI22xp5_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_388), .B1(n_391), .B2(n_392), .Y(n_386) );
OAI22xp5_ASAP7_75t_L g424 ( .A1(n_387), .A2(n_391), .B1(n_425), .B2(n_427), .Y(n_424) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
OAI22xp5_ASAP7_75t_L g530 ( .A1(n_390), .A2(n_531), .B1(n_532), .B2(n_534), .Y(n_530) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx2_ASAP7_75t_L g533 ( .A(n_394), .Y(n_533) );
OR2x2_ASAP7_75t_L g1079 ( .A(n_394), .B(n_558), .Y(n_1079) );
OAI22xp33_ASAP7_75t_SL g395 ( .A1(n_396), .A2(n_397), .B1(n_399), .B2(n_400), .Y(n_395) );
OAI22xp33_ASAP7_75t_L g419 ( .A1(n_396), .A2(n_399), .B1(n_420), .B2(n_421), .Y(n_419) );
INVx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx2_ASAP7_75t_L g1461 ( .A(n_398), .Y(n_1461) );
INVx1_ASAP7_75t_L g1503 ( .A(n_398), .Y(n_1503) );
BUFx2_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx2_ASAP7_75t_L g405 ( .A(n_402), .Y(n_405) );
BUFx4f_ASAP7_75t_L g1058 ( .A(n_402), .Y(n_1058) );
BUFx3_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
OR2x6_ASAP7_75t_L g569 ( .A(n_405), .B(n_557), .Y(n_569) );
OAI221xp5_ASAP7_75t_L g1451 ( .A1(n_405), .A2(n_1452), .B1(n_1455), .B2(n_1456), .C(n_1457), .Y(n_1451) );
OAI22xp5_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_409), .B1(n_410), .B2(n_411), .Y(n_407) );
INVx2_ASAP7_75t_L g561 ( .A(n_409), .Y(n_561) );
INVx1_ASAP7_75t_L g868 ( .A(n_409), .Y(n_868) );
INVx4_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
AOI221xp5_ASAP7_75t_L g514 ( .A1(n_413), .A2(n_515), .B1(n_525), .B2(n_527), .C(n_535), .Y(n_514) );
AOI33xp33_ASAP7_75t_L g803 ( .A1(n_413), .A2(n_804), .A3(n_805), .B1(n_810), .B2(n_812), .B3(n_814), .Y(n_803) );
AOI33xp33_ASAP7_75t_L g907 ( .A1(n_413), .A2(n_804), .A3(n_908), .B1(n_911), .B2(n_913), .B3(n_916), .Y(n_907) );
BUFx4f_ASAP7_75t_L g939 ( .A(n_413), .Y(n_939) );
AOI33xp33_ASAP7_75t_L g1112 ( .A1(n_413), .A2(n_804), .A3(n_1113), .B1(n_1118), .B2(n_1121), .B3(n_1124), .Y(n_1112) );
BUFx4f_ASAP7_75t_L g1459 ( .A(n_413), .Y(n_1459) );
INVx2_ASAP7_75t_L g1061 ( .A(n_414), .Y(n_1061) );
AND2x4_ASAP7_75t_L g541 ( .A(n_415), .B(n_542), .Y(n_541) );
OAI33xp33_ASAP7_75t_L g416 ( .A1(n_417), .A2(n_419), .A3(n_424), .B1(n_430), .B2(n_439), .B3(n_446), .Y(n_416) );
OAI33xp33_ASAP7_75t_L g1015 ( .A1(n_417), .A2(n_446), .A3(n_1016), .B1(n_1024), .B2(n_1029), .B3(n_1033), .Y(n_1015) );
OAI33xp33_ASAP7_75t_L g1373 ( .A1(n_417), .A2(n_1374), .A3(n_1379), .B1(n_1385), .B2(n_1386), .B3(n_1391), .Y(n_1373) );
OAI22xp33_ASAP7_75t_L g439 ( .A1(n_420), .A2(n_440), .B1(n_441), .B2(n_445), .Y(n_439) );
INVx1_ASAP7_75t_L g1382 ( .A(n_420), .Y(n_1382) );
INVx1_ASAP7_75t_L g1388 ( .A(n_420), .Y(n_1388) );
BUFx2_ASAP7_75t_L g1486 ( .A(n_420), .Y(n_1486) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_423), .B(n_486), .Y(n_485) );
OR2x6_ASAP7_75t_L g742 ( .A(n_423), .B(n_492), .Y(n_742) );
OR2x2_ASAP7_75t_L g979 ( .A(n_423), .B(n_492), .Y(n_979) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g861 ( .A(n_427), .Y(n_861) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
AND2x4_ASAP7_75t_L g503 ( .A(n_428), .B(n_504), .Y(n_503) );
INVx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g740 ( .A(n_429), .Y(n_740) );
INVx2_ASAP7_75t_SL g431 ( .A(n_432), .Y(n_431) );
INVx2_ASAP7_75t_L g976 ( .A(n_432), .Y(n_976) );
INVx2_ASAP7_75t_L g1392 ( .A(n_432), .Y(n_1392) );
BUFx3_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g953 ( .A(n_433), .Y(n_953) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx2_ASAP7_75t_SL g435 ( .A(n_436), .Y(n_435) );
INVx2_ASAP7_75t_L g685 ( .A(n_436), .Y(n_685) );
INVx2_ASAP7_75t_L g1106 ( .A(n_436), .Y(n_1106) );
BUFx6f_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx3_ASAP7_75t_L g464 ( .A(n_437), .Y(n_464) );
INVx3_ASAP7_75t_L g995 ( .A(n_437), .Y(n_995) );
INVx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g1384 ( .A(n_442), .Y(n_1384) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
BUFx6f_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
AOI33xp33_ASAP7_75t_L g597 ( .A1(n_447), .A2(n_598), .A3(n_600), .B1(n_603), .B2(n_607), .B3(n_609), .Y(n_597) );
AOI33xp33_ASAP7_75t_L g786 ( .A1(n_447), .A2(n_787), .A3(n_789), .B1(n_792), .B2(n_797), .B3(n_802), .Y(n_786) );
AOI33xp33_ASAP7_75t_L g902 ( .A1(n_447), .A2(n_598), .A3(n_903), .B1(n_904), .B2(n_905), .B3(n_906), .Y(n_902) );
INVx6_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx5_ASAP7_75t_L g687 ( .A(n_448), .Y(n_687) );
OR2x6_ASAP7_75t_L g448 ( .A(n_449), .B(n_451), .Y(n_448) );
NAND2x1p5_ASAP7_75t_L g540 ( .A(n_449), .B(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
OR2x2_ASAP7_75t_L g557 ( .A(n_450), .B(n_558), .Y(n_557) );
AND2x4_ASAP7_75t_L g996 ( .A(n_450), .B(n_498), .Y(n_996) );
BUFx2_ASAP7_75t_L g481 ( .A(n_451), .Y(n_481) );
INVx2_ASAP7_75t_L g725 ( .A(n_451), .Y(n_725) );
NAND4xp25_ASAP7_75t_L g456 ( .A(n_457), .B(n_514), .C(n_552), .D(n_564), .Y(n_456) );
OAI31xp33_ASAP7_75t_L g457 ( .A1(n_458), .A2(n_495), .A3(n_506), .B(n_512), .Y(n_457) );
OAI221xp5_ASAP7_75t_L g458 ( .A1(n_459), .A2(n_466), .B1(n_472), .B2(n_476), .C(n_482), .Y(n_458) );
OAI22xp5_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_462), .B1(n_463), .B2(n_465), .Y(n_459) );
OAI22xp5_ASAP7_75t_L g472 ( .A1(n_460), .A2(n_473), .B1(n_474), .B2(n_475), .Y(n_472) );
BUFx2_ASAP7_75t_L g1376 ( .A(n_460), .Y(n_1376) );
INVx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g1490 ( .A(n_461), .Y(n_1490) );
OAI22xp5_ASAP7_75t_L g521 ( .A1(n_462), .A2(n_465), .B1(n_522), .B2(n_524), .Y(n_521) );
INVx2_ASAP7_75t_L g608 ( .A(n_463), .Y(n_608) );
INVx2_ASAP7_75t_SL g678 ( .A(n_463), .Y(n_678) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx2_ASAP7_75t_L g474 ( .A(n_464), .Y(n_474) );
HB1xp67_ASAP7_75t_L g719 ( .A(n_464), .Y(n_719) );
INVx2_ASAP7_75t_L g1378 ( .A(n_464), .Y(n_1378) );
OAI21xp5_ASAP7_75t_L g466 ( .A1(n_467), .A2(n_468), .B(n_469), .Y(n_466) );
BUFx2_ASAP7_75t_L g968 ( .A(n_468), .Y(n_968) );
INVx1_ASAP7_75t_L g1022 ( .A(n_468), .Y(n_1022) );
BUFx2_ASAP7_75t_L g601 ( .A(n_470), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_470), .B(n_714), .Y(n_713) );
INVx2_ASAP7_75t_SL g470 ( .A(n_471), .Y(n_470) );
INVx2_ASAP7_75t_L g480 ( .A(n_471), .Y(n_480) );
INVx2_ASAP7_75t_SL g960 ( .A(n_471), .Y(n_960) );
AOI222xp33_ASAP7_75t_L g552 ( .A1(n_473), .A2(n_483), .B1(n_553), .B2(n_559), .C1(n_560), .C2(n_562), .Y(n_552) );
INVx1_ASAP7_75t_L g606 ( .A(n_474), .Y(n_606) );
INVx2_ASAP7_75t_L g856 ( .A(n_474), .Y(n_856) );
AOI22xp5_ASAP7_75t_L g564 ( .A1(n_475), .A2(n_477), .B1(n_565), .B2(n_568), .Y(n_564) );
OAI21xp33_ASAP7_75t_L g476 ( .A1(n_477), .A2(n_478), .B(n_479), .Y(n_476) );
BUFx3_ASAP7_75t_L g790 ( .A(n_480), .Y(n_790) );
A2O1A1Ixp33_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_484), .B(n_485), .C(n_491), .Y(n_482) );
NAND2x1p5_ASAP7_75t_L g1012 ( .A(n_489), .B(n_1009), .Y(n_1012) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
OR2x6_ASAP7_75t_L g732 ( .A(n_490), .B(n_492), .Y(n_732) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g714 ( .A(n_492), .Y(n_714) );
INVx1_ASAP7_75t_L g731 ( .A(n_492), .Y(n_731) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx3_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
AOI22xp33_ASAP7_75t_L g733 ( .A1(n_497), .A2(n_503), .B1(n_734), .B2(n_735), .Y(n_733) );
INVx3_ASAP7_75t_L g981 ( .A(n_497), .Y(n_981) );
AND2x2_ASAP7_75t_L g497 ( .A(n_498), .B(n_499), .Y(n_497) );
INVx2_ASAP7_75t_L g505 ( .A(n_498), .Y(n_505) );
INVx1_ASAP7_75t_L g605 ( .A(n_499), .Y(n_605) );
BUFx6f_ASAP7_75t_L g718 ( .A(n_499), .Y(n_718) );
BUFx2_ASAP7_75t_L g793 ( .A(n_499), .Y(n_793) );
BUFx6f_ASAP7_75t_L g800 ( .A(n_499), .Y(n_800) );
BUFx2_ASAP7_75t_L g860 ( .A(n_499), .Y(n_860) );
BUFx6f_ASAP7_75t_L g1104 ( .A(n_499), .Y(n_1104) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx3_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx3_ASAP7_75t_L g1496 ( .A(n_503), .Y(n_1496) );
AND2x4_ASAP7_75t_L g510 ( .A(n_504), .B(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
CKINVDCx6p67_ASAP7_75t_R g507 ( .A(n_508), .Y(n_507) );
AOI221xp5_ASAP7_75t_L g736 ( .A1(n_508), .A2(n_737), .B1(n_738), .B2(n_739), .C(n_741), .Y(n_736) );
INVx8_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
AOI221xp5_ASAP7_75t_SL g716 ( .A1(n_510), .A2(n_717), .B1(n_720), .B2(n_726), .C(n_727), .Y(n_716) );
INVx1_ASAP7_75t_L g723 ( .A(n_511), .Y(n_723) );
INVx1_ASAP7_75t_L g743 ( .A(n_512), .Y(n_743) );
INVx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
NOR2xp67_ASAP7_75t_L g712 ( .A(n_513), .B(n_713), .Y(n_712) );
INVx3_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx2_ASAP7_75t_L g749 ( .A(n_517), .Y(n_749) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
HB1xp67_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
BUFx6f_ASAP7_75t_L g529 ( .A(n_520), .Y(n_529) );
INVx2_ASAP7_75t_L g619 ( .A(n_520), .Y(n_619) );
INVx2_ASAP7_75t_L g638 ( .A(n_520), .Y(n_638) );
INVx1_ASAP7_75t_L g698 ( .A(n_520), .Y(n_698) );
INVx2_ASAP7_75t_L g807 ( .A(n_520), .Y(n_807) );
INVx2_ASAP7_75t_SL g1418 ( .A(n_520), .Y(n_1418) );
INVx1_ASAP7_75t_L g909 ( .A(n_522), .Y(n_909) );
INVx2_ASAP7_75t_SL g522 ( .A(n_523), .Y(n_522) );
BUFx3_ASAP7_75t_L g811 ( .A(n_523), .Y(n_811) );
AND2x4_ASAP7_75t_L g1045 ( .A(n_523), .B(n_1046), .Y(n_1045) );
INVx1_ASAP7_75t_L g910 ( .A(n_524), .Y(n_910) );
INVx1_ASAP7_75t_L g917 ( .A(n_524), .Y(n_917) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
CKINVDCx5p33_ASAP7_75t_R g804 ( .A(n_526), .Y(n_804) );
OAI22xp5_ASAP7_75t_SL g1450 ( .A1(n_526), .A2(n_1451), .B1(n_1458), .B2(n_1460), .Y(n_1450) );
INVx4_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx2_ASAP7_75t_L g866 ( .A(n_529), .Y(n_866) );
INVx1_ASAP7_75t_L g853 ( .A(n_532), .Y(n_853) );
INVx1_ASAP7_75t_L g869 ( .A(n_532), .Y(n_869) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx2_ASAP7_75t_L g761 ( .A(n_536), .Y(n_761) );
INVx1_ASAP7_75t_L g930 ( .A(n_536), .Y(n_930) );
NAND2x1p5_ASAP7_75t_L g536 ( .A(n_537), .B(n_539), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx2_ASAP7_75t_L g1050 ( .A(n_538), .Y(n_1050) );
INVx2_ASAP7_75t_SL g539 ( .A(n_540), .Y(n_539) );
OR2x6_ASAP7_75t_L g545 ( .A(n_540), .B(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g551 ( .A(n_540), .Y(n_551) );
AND2x4_ASAP7_75t_L g1049 ( .A(n_541), .B(n_1050), .Y(n_1049) );
INVx1_ASAP7_75t_L g1052 ( .A(n_541), .Y(n_1052) );
AND2x2_ASAP7_75t_L g1426 ( .A(n_541), .B(n_547), .Y(n_1426) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx2_ASAP7_75t_L g759 ( .A(n_545), .Y(n_759) );
OR2x2_ASAP7_75t_L g1051 ( .A(n_546), .B(n_1052), .Y(n_1051) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
NAND3xp33_ASAP7_75t_SL g927 ( .A(n_548), .B(n_928), .C(n_932), .Y(n_927) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_549), .B(n_551), .Y(n_548) );
INVx1_ASAP7_75t_L g1123 ( .A(n_549), .Y(n_1123) );
BUFx6f_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g623 ( .A(n_550), .Y(n_623) );
INVx2_ASAP7_75t_SL g887 ( .A(n_550), .Y(n_887) );
BUFx3_ASAP7_75t_L g912 ( .A(n_550), .Y(n_912) );
AND2x4_ASAP7_75t_L g1065 ( .A(n_550), .B(n_1046), .Y(n_1065) );
INVx1_ASAP7_75t_L g1068 ( .A(n_550), .Y(n_1068) );
AND2x2_ASAP7_75t_L g763 ( .A(n_551), .B(n_764), .Y(n_763) );
AOI22xp5_ASAP7_75t_L g755 ( .A1(n_553), .A2(n_560), .B1(n_756), .B2(n_757), .Y(n_755) );
AOI22xp33_ASAP7_75t_L g944 ( .A1(n_553), .A2(n_560), .B1(n_945), .B2(n_946), .Y(n_944) );
AND2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_556), .Y(n_553) );
BUFx2_ASAP7_75t_L g1119 ( .A(n_554), .Y(n_1119) );
INVx2_ASAP7_75t_SL g554 ( .A(n_555), .Y(n_554) );
INVx1_ASAP7_75t_L g813 ( .A(n_555), .Y(n_813) );
AND2x2_ASAP7_75t_L g560 ( .A(n_556), .B(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
OR2x6_ASAP7_75t_L g566 ( .A(n_557), .B(n_567), .Y(n_566) );
OR2x2_ASAP7_75t_L g1500 ( .A(n_557), .B(n_567), .Y(n_1500) );
OR2x2_ASAP7_75t_L g1502 ( .A(n_557), .B(n_1503), .Y(n_1502) );
OR2x2_ASAP7_75t_L g1504 ( .A(n_557), .B(n_1505), .Y(n_1504) );
INVx2_ASAP7_75t_L g1046 ( .A(n_558), .Y(n_1046) );
OR2x6_ASAP7_75t_L g711 ( .A(n_562), .B(n_712), .Y(n_711) );
INVx2_ASAP7_75t_L g1041 ( .A(n_562), .Y(n_1041) );
AOI22xp5_ASAP7_75t_L g752 ( .A1(n_565), .A2(n_568), .B1(n_753), .B2(n_754), .Y(n_752) );
AOI22xp33_ASAP7_75t_L g941 ( .A1(n_565), .A2(n_568), .B1(n_942), .B2(n_943), .Y(n_941) );
CKINVDCx6p67_ASAP7_75t_R g565 ( .A(n_566), .Y(n_565) );
INVx2_ASAP7_75t_L g747 ( .A(n_567), .Y(n_747) );
CKINVDCx6p67_ASAP7_75t_R g568 ( .A(n_569), .Y(n_568) );
OA22x2_ASAP7_75t_L g570 ( .A1(n_571), .A2(n_644), .B1(n_645), .B2(n_702), .Y(n_570) );
INVx1_ASAP7_75t_L g702 ( .A(n_571), .Y(n_702) );
XNOR2xp5_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .Y(n_571) );
AOI211xp5_ASAP7_75t_L g573 ( .A1(n_574), .A2(n_576), .B(n_596), .C(n_627), .Y(n_573) );
AOI221x1_ASAP7_75t_L g646 ( .A1(n_574), .A2(n_647), .B1(n_660), .B2(n_662), .C(n_675), .Y(n_646) );
CKINVDCx16_ASAP7_75t_R g574 ( .A(n_575), .Y(n_574) );
AOI31xp33_ASAP7_75t_L g870 ( .A1(n_575), .A2(n_871), .A3(n_875), .B(n_878), .Y(n_870) );
AO21x1_ASAP7_75t_SL g894 ( .A1(n_575), .A2(n_895), .B(n_899), .Y(n_894) );
AOI22xp5_ASAP7_75t_L g577 ( .A1(n_578), .A2(n_579), .B1(n_580), .B2(n_581), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_579), .A2(n_581), .B1(n_664), .B2(n_665), .Y(n_663) );
AOI22xp33_ASAP7_75t_SL g1129 ( .A1(n_579), .A2(n_581), .B1(n_1130), .B2(n_1131), .Y(n_1129) );
INVx4_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx5_ASAP7_75t_L g828 ( .A(n_586), .Y(n_828) );
INVx2_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx2_ASAP7_75t_SL g791 ( .A(n_590), .Y(n_791) );
INVx2_ASAP7_75t_SL g590 ( .A(n_591), .Y(n_590) );
BUFx6f_ASAP7_75t_L g602 ( .A(n_591), .Y(n_602) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_SL g596 ( .A(n_597), .B(n_612), .Y(n_596) );
NAND3xp33_ASAP7_75t_L g676 ( .A(n_598), .B(n_677), .C(n_679), .Y(n_676) );
BUFx2_ASAP7_75t_SL g973 ( .A(n_599), .Y(n_973) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
BUFx2_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx2_ASAP7_75t_SL g682 ( .A(n_611), .Y(n_682) );
HB1xp67_ASAP7_75t_L g863 ( .A(n_611), .Y(n_863) );
AOI33xp33_ASAP7_75t_L g612 ( .A1(n_613), .A2(n_614), .A3(n_617), .B1(n_620), .B2(n_624), .B3(n_626), .Y(n_612) );
BUFx6f_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g1072 ( .A(n_619), .Y(n_1072) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
NAND3xp33_ASAP7_75t_L g696 ( .A(n_626), .B(n_697), .C(n_699), .Y(n_696) );
AOI33xp33_ASAP7_75t_L g745 ( .A1(n_626), .A2(n_693), .A3(n_746), .B1(n_748), .B2(n_750), .B3(n_751), .Y(n_745) );
NAND3xp33_ASAP7_75t_L g864 ( .A(n_626), .B(n_865), .C(n_867), .Y(n_864) );
AOI31xp33_ASAP7_75t_SL g627 ( .A1(n_628), .A2(n_635), .A3(n_639), .B(n_643), .Y(n_627) );
INVx2_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g656 ( .A(n_632), .Y(n_656) );
AOI22xp33_ASAP7_75t_L g1086 ( .A1(n_637), .A2(n_640), .B1(n_1087), .B2(n_1088), .Y(n_1086) );
AOI22xp33_ASAP7_75t_L g782 ( .A1(n_640), .A2(n_649), .B1(n_783), .B2(n_784), .Y(n_782) );
CKINVDCx6p67_ASAP7_75t_R g892 ( .A(n_640), .Y(n_892) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g701 ( .A(n_646), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_648), .B(n_652), .Y(n_647) );
INVx1_ASAP7_75t_L g809 ( .A(n_659), .Y(n_809) );
BUFx6f_ASAP7_75t_L g915 ( .A(n_659), .Y(n_915) );
AND2x4_ASAP7_75t_L g1073 ( .A(n_659), .B(n_1074), .Y(n_1073) );
BUFx6f_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
AOI211x1_ASAP7_75t_SL g769 ( .A1(n_661), .A2(n_770), .B(n_785), .C(n_817), .Y(n_769) );
AO211x2_ASAP7_75t_L g835 ( .A1(n_661), .A2(n_836), .B(n_848), .C(n_870), .Y(n_835) );
INVx1_ASAP7_75t_L g1097 ( .A(n_661), .Y(n_1097) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
NAND4xp25_ASAP7_75t_L g675 ( .A(n_676), .B(n_683), .C(n_688), .D(n_696), .Y(n_675) );
INVx2_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
NAND3xp33_ASAP7_75t_L g683 ( .A(n_684), .B(n_686), .C(n_687), .Y(n_683) );
NAND3xp33_ASAP7_75t_L g854 ( .A(n_687), .B(n_855), .C(n_857), .Y(n_854) );
AOI33xp33_ASAP7_75t_L g1099 ( .A1(n_687), .A2(n_1100), .A3(n_1102), .B1(n_1107), .B2(n_1109), .B3(n_1111), .Y(n_1099) );
CKINVDCx8_ASAP7_75t_R g1385 ( .A(n_687), .Y(n_1385) );
NAND3xp33_ASAP7_75t_L g688 ( .A(n_689), .B(n_692), .C(n_693), .Y(n_688) );
BUFx6f_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g1055 ( .A(n_691), .Y(n_1055) );
NAND3xp33_ASAP7_75t_L g849 ( .A(n_693), .B(n_850), .C(n_851), .Y(n_849) );
INVx3_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
OAI22xp5_ASAP7_75t_L g703 ( .A1(n_704), .A2(n_705), .B1(n_832), .B2(n_920), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
AOI21x1_ASAP7_75t_L g705 ( .A1(n_706), .A2(n_767), .B(n_831), .Y(n_705) );
INVx2_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
AND2x2_ASAP7_75t_L g831 ( .A(n_707), .B(n_768), .Y(n_831) );
XOR2x2_ASAP7_75t_L g707 ( .A(n_708), .B(n_766), .Y(n_707) );
NOR3xp33_ASAP7_75t_L g708 ( .A(n_709), .B(n_715), .C(n_744), .Y(n_708) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g947 ( .A(n_711), .B(n_948), .Y(n_947) );
NAND2xp5_ASAP7_75t_L g1470 ( .A(n_711), .B(n_1471), .Y(n_1470) );
AND2x2_ASAP7_75t_L g963 ( .A(n_714), .B(n_964), .Y(n_963) );
AOI31xp33_ASAP7_75t_L g715 ( .A1(n_716), .A2(n_733), .A3(n_736), .B(n_743), .Y(n_715) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx2_ASAP7_75t_SL g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g961 ( .A(n_725), .Y(n_961) );
NAND2x1p5_ASAP7_75t_L g728 ( .A(n_729), .B(n_731), .Y(n_728) );
NAND2x1_ASAP7_75t_SL g1008 ( .A(n_729), .B(n_1009), .Y(n_1008) );
INVx2_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
CKINVDCx11_ASAP7_75t_R g965 ( .A(n_732), .Y(n_965) );
INVx1_ASAP7_75t_L g956 ( .A(n_740), .Y(n_956) );
INVx2_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
NAND4xp25_ASAP7_75t_L g744 ( .A(n_745), .B(n_752), .C(n_755), .D(n_758), .Y(n_744) );
AOI221xp5_ASAP7_75t_L g758 ( .A1(n_759), .A2(n_760), .B1(n_761), .B2(n_762), .C(n_763), .Y(n_758) );
AOI22xp33_ASAP7_75t_L g928 ( .A1(n_759), .A2(n_929), .B1(n_930), .B2(n_931), .Y(n_928) );
BUFx2_ASAP7_75t_L g1447 ( .A(n_763), .Y(n_1447) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
INVx2_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
INVx1_ASAP7_75t_L g830 ( .A(n_769), .Y(n_830) );
NAND4xp25_ASAP7_75t_L g770 ( .A(n_771), .B(n_772), .C(n_775), .D(n_782), .Y(n_770) );
NAND4xp25_ASAP7_75t_L g1085 ( .A(n_771), .B(n_1086), .C(n_1089), .D(n_1092), .Y(n_1085) );
BUFx4f_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
INVx1_ASAP7_75t_L g841 ( .A(n_780), .Y(n_841) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_786), .B(n_803), .Y(n_785) );
BUFx3_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
NAND3xp33_ASAP7_75t_L g858 ( .A(n_788), .B(n_859), .C(n_862), .Y(n_858) );
INVx2_ASAP7_75t_L g1101 ( .A(n_788), .Y(n_1101) );
INVx2_ASAP7_75t_SL g794 ( .A(n_795), .Y(n_794) );
INVx4_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
BUFx3_ASAP7_75t_L g801 ( .A(n_796), .Y(n_801) );
INVx2_ASAP7_75t_SL g1028 ( .A(n_796), .Y(n_1028) );
INVx2_ASAP7_75t_SL g1031 ( .A(n_796), .Y(n_1031) );
INVx3_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
INVx2_ASAP7_75t_SL g799 ( .A(n_800), .Y(n_799) );
AND2x2_ASAP7_75t_L g1004 ( .A(n_800), .B(n_996), .Y(n_1004) );
INVx1_ASAP7_75t_L g978 ( .A(n_801), .Y(n_978) );
INVx1_ASAP7_75t_L g1394 ( .A(n_801), .Y(n_1394) );
AOI33xp33_ASAP7_75t_L g932 ( .A1(n_804), .A2(n_933), .A3(n_936), .B1(n_937), .B2(n_938), .B3(n_939), .Y(n_932) );
BUFx3_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
HB1xp67_ASAP7_75t_L g914 ( .A(n_807), .Y(n_914) );
INVx1_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
BUFx2_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
BUFx4f_ASAP7_75t_L g852 ( .A(n_816), .Y(n_852) );
INVx1_ASAP7_75t_L g1505 ( .A(n_816), .Y(n_1505) );
INVx1_ASAP7_75t_L g920 ( .A(n_832), .Y(n_920) );
INVx1_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
XNOR2x1_ASAP7_75t_L g833 ( .A(n_834), .B(n_880), .Y(n_833) );
NAND3xp33_ASAP7_75t_L g836 ( .A(n_837), .B(n_842), .C(n_845), .Y(n_836) );
NAND4xp25_ASAP7_75t_L g848 ( .A(n_849), .B(n_854), .C(n_858), .D(n_864), .Y(n_848) );
INVx1_ASAP7_75t_L g1478 ( .A(n_861), .Y(n_1478) );
AND4x1_ASAP7_75t_L g881 ( .A(n_882), .B(n_894), .C(n_902), .D(n_907), .Y(n_881) );
NAND4xp25_ASAP7_75t_L g919 ( .A(n_882), .B(n_894), .C(n_902), .D(n_907), .Y(n_919) );
NAND2xp5_ASAP7_75t_L g884 ( .A(n_885), .B(n_886), .Y(n_884) );
INVx2_ASAP7_75t_L g886 ( .A(n_887), .Y(n_886) );
INVx1_ASAP7_75t_L g1422 ( .A(n_887), .Y(n_1422) );
INVxp67_ASAP7_75t_SL g1139 ( .A(n_921), .Y(n_1139) );
AOI22xp33_ASAP7_75t_L g921 ( .A1(n_922), .A2(n_984), .B1(n_985), .B2(n_1138), .Y(n_921) );
INVx1_ASAP7_75t_L g1138 ( .A(n_922), .Y(n_1138) );
HB1xp67_ASAP7_75t_L g922 ( .A(n_923), .Y(n_922) );
INVx1_ASAP7_75t_L g923 ( .A(n_924), .Y(n_923) );
AND3x1_ASAP7_75t_L g925 ( .A(n_926), .B(n_947), .C(n_949), .Y(n_925) );
NOR2xp33_ASAP7_75t_L g926 ( .A(n_927), .B(n_940), .Y(n_926) );
AOI22xp33_ASAP7_75t_L g962 ( .A1(n_929), .A2(n_931), .B1(n_963), .B2(n_965), .Y(n_962) );
INVx1_ASAP7_75t_L g1449 ( .A(n_930), .Y(n_1449) );
INVx1_ASAP7_75t_L g934 ( .A(n_935), .Y(n_934) );
INVx1_ASAP7_75t_L g1469 ( .A(n_935), .Y(n_1469) );
NAND2xp5_ASAP7_75t_L g940 ( .A(n_941), .B(n_944), .Y(n_940) );
OAI221xp5_ASAP7_75t_L g951 ( .A1(n_942), .A2(n_946), .B1(n_952), .B2(n_954), .C(n_957), .Y(n_951) );
OAI31xp33_ASAP7_75t_L g949 ( .A1(n_950), .A2(n_966), .A3(n_980), .B(n_982), .Y(n_949) );
BUFx2_ASAP7_75t_L g952 ( .A(n_953), .Y(n_952) );
INVx2_ASAP7_75t_L g1476 ( .A(n_953), .Y(n_1476) );
INVx1_ASAP7_75t_L g954 ( .A(n_955), .Y(n_954) );
INVx1_ASAP7_75t_L g955 ( .A(n_956), .Y(n_955) );
INVx1_ASAP7_75t_L g958 ( .A(n_959), .Y(n_958) );
INVx1_ASAP7_75t_L g959 ( .A(n_960), .Y(n_959) );
AND2x4_ASAP7_75t_L g1002 ( .A(n_960), .B(n_996), .Y(n_1002) );
BUFx3_ASAP7_75t_L g1108 ( .A(n_960), .Y(n_1108) );
AOI22xp33_ASAP7_75t_L g1481 ( .A1(n_963), .A2(n_965), .B1(n_1482), .B2(n_1483), .Y(n_1481) );
OAI221xp5_ASAP7_75t_L g967 ( .A1(n_968), .A2(n_969), .B1(n_970), .B2(n_972), .C(n_973), .Y(n_967) );
INVx1_ASAP7_75t_L g970 ( .A(n_971), .Y(n_970) );
OAI22xp5_ASAP7_75t_L g974 ( .A1(n_975), .A2(n_976), .B1(n_977), .B2(n_978), .Y(n_974) );
BUFx8_ASAP7_75t_SL g982 ( .A(n_983), .Y(n_982) );
INVx2_ASAP7_75t_L g1407 ( .A(n_983), .Y(n_1407) );
INVx1_ASAP7_75t_L g984 ( .A(n_985), .Y(n_984) );
INVxp67_ASAP7_75t_L g985 ( .A(n_986), .Y(n_985) );
AOI22x1_ASAP7_75t_L g986 ( .A1(n_987), .A2(n_1082), .B1(n_1135), .B2(n_1136), .Y(n_986) );
AND2x2_ASAP7_75t_L g988 ( .A(n_989), .B(n_1037), .Y(n_988) );
NOR3xp33_ASAP7_75t_L g989 ( .A(n_990), .B(n_1005), .C(n_1015), .Y(n_989) );
NAND2xp5_ASAP7_75t_L g990 ( .A(n_991), .B(n_1000), .Y(n_990) );
AOI22xp33_ASAP7_75t_L g991 ( .A1(n_992), .A2(n_993), .B1(n_997), .B2(n_998), .Y(n_991) );
AOI22xp33_ASAP7_75t_L g1400 ( .A1(n_993), .A2(n_998), .B1(n_1401), .B2(n_1402), .Y(n_1400) );
BUFx2_ASAP7_75t_L g993 ( .A(n_994), .Y(n_993) );
AND2x4_ASAP7_75t_L g994 ( .A(n_995), .B(n_996), .Y(n_994) );
BUFx3_ASAP7_75t_L g1493 ( .A(n_995), .Y(n_1493) );
AND2x6_ASAP7_75t_L g998 ( .A(n_996), .B(n_999), .Y(n_998) );
OAI221xp5_ASAP7_75t_L g1056 ( .A1(n_997), .A2(n_1001), .B1(n_1057), .B2(n_1059), .C(n_1060), .Y(n_1056) );
NAND2x1p5_ASAP7_75t_L g1014 ( .A(n_999), .B(n_1009), .Y(n_1014) );
AOI22xp33_ASAP7_75t_L g1000 ( .A1(n_1001), .A2(n_1002), .B1(n_1003), .B2(n_1004), .Y(n_1000) );
AOI22xp33_ASAP7_75t_L g1403 ( .A1(n_1002), .A2(n_1004), .B1(n_1404), .B2(n_1405), .Y(n_1403) );
INVx2_ASAP7_75t_L g1006 ( .A(n_1007), .Y(n_1006) );
INVx2_ASAP7_75t_SL g1397 ( .A(n_1007), .Y(n_1397) );
INVx2_ASAP7_75t_L g1007 ( .A(n_1008), .Y(n_1007) );
INVx3_ASAP7_75t_L g1009 ( .A(n_1010), .Y(n_1009) );
BUFx4f_ASAP7_75t_L g1011 ( .A(n_1012), .Y(n_1011) );
BUFx2_ASAP7_75t_L g1013 ( .A(n_1014), .Y(n_1013) );
BUFx3_ASAP7_75t_L g1398 ( .A(n_1014), .Y(n_1398) );
OAI22xp33_ASAP7_75t_L g1016 ( .A1(n_1017), .A2(n_1020), .B1(n_1021), .B2(n_1023), .Y(n_1016) );
OAI22xp33_ASAP7_75t_L g1033 ( .A1(n_1017), .A2(n_1034), .B1(n_1035), .B2(n_1036), .Y(n_1033) );
BUFx2_ASAP7_75t_L g1017 ( .A(n_1018), .Y(n_1017) );
INVx2_ASAP7_75t_L g1018 ( .A(n_1019), .Y(n_1018) );
INVx1_ASAP7_75t_L g1021 ( .A(n_1022), .Y(n_1021) );
INVx1_ASAP7_75t_L g1035 ( .A(n_1022), .Y(n_1035) );
OAI22xp5_ASAP7_75t_L g1024 ( .A1(n_1025), .A2(n_1026), .B1(n_1027), .B2(n_1028), .Y(n_1024) );
OAI22xp5_ASAP7_75t_L g1029 ( .A1(n_1026), .A2(n_1030), .B1(n_1031), .B2(n_1032), .Y(n_1029) );
AOI211xp5_ASAP7_75t_L g1044 ( .A1(n_1030), .A2(n_1045), .B(n_1047), .C(n_1053), .Y(n_1044) );
INVx1_ASAP7_75t_L g1110 ( .A(n_1031), .Y(n_1110) );
AOI22xp33_ASAP7_75t_L g1075 ( .A1(n_1032), .A2(n_1034), .B1(n_1076), .B2(n_1078), .Y(n_1075) );
AOI221xp5_ASAP7_75t_L g1062 ( .A1(n_1036), .A2(n_1063), .B1(n_1066), .B2(n_1070), .C(n_1073), .Y(n_1062) );
AOI21xp5_ASAP7_75t_L g1037 ( .A1(n_1038), .A2(n_1042), .B(n_1043), .Y(n_1037) );
INVx1_ASAP7_75t_L g1038 ( .A(n_1039), .Y(n_1038) );
INVx5_ASAP7_75t_L g1431 ( .A(n_1039), .Y(n_1431) );
AND2x4_ASAP7_75t_L g1039 ( .A(n_1040), .B(n_1041), .Y(n_1039) );
AOI31xp33_ASAP7_75t_L g1043 ( .A1(n_1044), .A2(n_1062), .A3(n_1075), .B(n_1080), .Y(n_1043) );
AOI22xp33_ASAP7_75t_L g1428 ( .A1(n_1045), .A2(n_1076), .B1(n_1389), .B2(n_1393), .Y(n_1428) );
INVx2_ASAP7_75t_SL g1048 ( .A(n_1049), .Y(n_1048) );
AOI322xp5_ASAP7_75t_L g1419 ( .A1(n_1049), .A2(n_1420), .A3(n_1421), .B1(n_1423), .B2(n_1425), .C1(n_1426), .C2(n_1427), .Y(n_1419) );
INVx1_ASAP7_75t_SL g1074 ( .A(n_1052), .Y(n_1074) );
INVx1_ASAP7_75t_L g1054 ( .A(n_1055), .Y(n_1054) );
INVx1_ASAP7_75t_L g1057 ( .A(n_1058), .Y(n_1057) );
INVx1_ASAP7_75t_L g1464 ( .A(n_1058), .Y(n_1464) );
INVx1_ASAP7_75t_L g1060 ( .A(n_1061), .Y(n_1060) );
BUFx2_ASAP7_75t_L g1424 ( .A(n_1061), .Y(n_1424) );
INVx1_ASAP7_75t_L g1063 ( .A(n_1064), .Y(n_1063) );
INVx1_ASAP7_75t_L g1064 ( .A(n_1065), .Y(n_1064) );
INVx1_ASAP7_75t_L g1411 ( .A(n_1065), .Y(n_1411) );
INVx1_ASAP7_75t_L g1067 ( .A(n_1068), .Y(n_1067) );
INVx2_ASAP7_75t_L g1071 ( .A(n_1072), .Y(n_1071) );
AOI221xp5_ASAP7_75t_L g1409 ( .A1(n_1073), .A2(n_1390), .B1(n_1410), .B2(n_1412), .C(n_1415), .Y(n_1409) );
INVx6_ASAP7_75t_L g1076 ( .A(n_1077), .Y(n_1076) );
NAND2xp5_ASAP7_75t_L g1429 ( .A(n_1078), .B(n_1395), .Y(n_1429) );
INVx4_ASAP7_75t_L g1078 ( .A(n_1079), .Y(n_1078) );
INVx2_ASAP7_75t_L g1080 ( .A(n_1081), .Y(n_1080) );
INVx2_ASAP7_75t_L g1135 ( .A(n_1082), .Y(n_1135) );
INVx1_ASAP7_75t_L g1134 ( .A(n_1084), .Y(n_1134) );
AOI211x1_ASAP7_75t_L g1084 ( .A1(n_1085), .A2(n_1096), .B(n_1098), .C(n_1125), .Y(n_1084) );
INVx1_ASAP7_75t_L g1096 ( .A(n_1097), .Y(n_1096) );
NAND2xp5_ASAP7_75t_L g1098 ( .A(n_1099), .B(n_1112), .Y(n_1098) );
INVx2_ASAP7_75t_L g1100 ( .A(n_1101), .Y(n_1100) );
BUFx3_ASAP7_75t_L g1103 ( .A(n_1104), .Y(n_1103) );
HB1xp67_ASAP7_75t_L g1105 ( .A(n_1106), .Y(n_1105) );
BUFx3_ASAP7_75t_L g1114 ( .A(n_1115), .Y(n_1114) );
INVx1_ASAP7_75t_L g1116 ( .A(n_1117), .Y(n_1116) );
INVx1_ASAP7_75t_L g1122 ( .A(n_1123), .Y(n_1122) );
INVx3_ASAP7_75t_SL g1136 ( .A(n_1137), .Y(n_1136) );
OAI221xp5_ASAP7_75t_L g1140 ( .A1(n_1141), .A2(n_1363), .B1(n_1367), .B2(n_1433), .C(n_1437), .Y(n_1140) );
AOI221xp5_ASAP7_75t_L g1141 ( .A1(n_1142), .A2(n_1253), .B1(n_1254), .B2(n_1262), .C(n_1302), .Y(n_1141) );
A2O1A1Ixp33_ASAP7_75t_L g1142 ( .A1(n_1143), .A2(n_1196), .B(n_1222), .C(n_1230), .Y(n_1142) );
NAND2xp5_ASAP7_75t_L g1143 ( .A(n_1144), .B(n_1171), .Y(n_1143) );
INVxp67_ASAP7_75t_L g1207 ( .A(n_1144), .Y(n_1207) );
HB1xp67_ASAP7_75t_L g1144 ( .A(n_1145), .Y(n_1144) );
AND2x2_ASAP7_75t_L g1199 ( .A(n_1145), .B(n_1200), .Y(n_1199) );
INVx2_ASAP7_75t_SL g1219 ( .A(n_1145), .Y(n_1219) );
INVx1_ASAP7_75t_L g1233 ( .A(n_1145), .Y(n_1233) );
NAND2xp5_ASAP7_75t_L g1266 ( .A(n_1145), .B(n_1173), .Y(n_1266) );
AND2x2_ASAP7_75t_L g1279 ( .A(n_1145), .B(n_1172), .Y(n_1279) );
NOR2xp33_ASAP7_75t_L g1310 ( .A(n_1145), .B(n_1172), .Y(n_1310) );
AND2x4_ASAP7_75t_L g1322 ( .A(n_1145), .B(n_1216), .Y(n_1322) );
CKINVDCx5p33_ASAP7_75t_R g1145 ( .A(n_1146), .Y(n_1145) );
AND2x2_ASAP7_75t_L g1215 ( .A(n_1146), .B(n_1216), .Y(n_1215) );
AND2x2_ASAP7_75t_L g1285 ( .A(n_1146), .B(n_1200), .Y(n_1285) );
OR2x2_ASAP7_75t_L g1146 ( .A(n_1147), .B(n_1161), .Y(n_1146) );
OAI22xp5_ASAP7_75t_L g1147 ( .A1(n_1148), .A2(n_1155), .B1(n_1156), .B2(n_1160), .Y(n_1147) );
BUFx3_ASAP7_75t_L g1259 ( .A(n_1148), .Y(n_1259) );
BUFx6f_ASAP7_75t_L g1148 ( .A(n_1149), .Y(n_1148) );
OAI22xp5_ASAP7_75t_L g1193 ( .A1(n_1149), .A2(n_1158), .B1(n_1194), .B2(n_1195), .Y(n_1193) );
OR2x2_ASAP7_75t_L g1149 ( .A(n_1150), .B(n_1151), .Y(n_1149) );
OR2x2_ASAP7_75t_L g1158 ( .A(n_1150), .B(n_1159), .Y(n_1158) );
INVx1_ASAP7_75t_L g1177 ( .A(n_1150), .Y(n_1177) );
INVx1_ASAP7_75t_L g1176 ( .A(n_1151), .Y(n_1176) );
NAND2xp5_ASAP7_75t_L g1151 ( .A(n_1152), .B(n_1154), .Y(n_1151) );
HB1xp67_ASAP7_75t_L g1511 ( .A(n_1152), .Y(n_1511) );
INVx1_ASAP7_75t_L g1152 ( .A(n_1153), .Y(n_1152) );
INVx1_ASAP7_75t_L g1165 ( .A(n_1154), .Y(n_1165) );
HB1xp67_ASAP7_75t_L g1261 ( .A(n_1156), .Y(n_1261) );
INVx1_ASAP7_75t_L g1156 ( .A(n_1157), .Y(n_1156) );
INVx1_ASAP7_75t_L g1157 ( .A(n_1158), .Y(n_1157) );
INVx1_ASAP7_75t_L g1179 ( .A(n_1159), .Y(n_1179) );
OAI22xp5_ASAP7_75t_L g1161 ( .A1(n_1162), .A2(n_1167), .B1(n_1168), .B2(n_1170), .Y(n_1161) );
INVx1_ASAP7_75t_L g1162 ( .A(n_1163), .Y(n_1162) );
BUFx3_ASAP7_75t_L g1256 ( .A(n_1163), .Y(n_1256) );
AND2x4_ASAP7_75t_L g1163 ( .A(n_1164), .B(n_1166), .Y(n_1163) );
AND2x2_ASAP7_75t_L g1186 ( .A(n_1164), .B(n_1166), .Y(n_1186) );
HB1xp67_ASAP7_75t_L g1509 ( .A(n_1164), .Y(n_1509) );
INVx1_ASAP7_75t_L g1164 ( .A(n_1165), .Y(n_1164) );
AND2x4_ASAP7_75t_L g1169 ( .A(n_1165), .B(n_1166), .Y(n_1169) );
INVx2_ASAP7_75t_L g1229 ( .A(n_1168), .Y(n_1229) );
INVx1_ASAP7_75t_L g1366 ( .A(n_1168), .Y(n_1366) );
INVx2_ASAP7_75t_L g1168 ( .A(n_1169), .Y(n_1168) );
AND2x2_ASAP7_75t_L g1304 ( .A(n_1171), .B(n_1296), .Y(n_1304) );
AND2x2_ASAP7_75t_L g1171 ( .A(n_1172), .B(n_1181), .Y(n_1171) );
NAND2xp5_ASAP7_75t_L g1209 ( .A(n_1172), .B(n_1210), .Y(n_1209) );
NAND3xp33_ASAP7_75t_L g1308 ( .A(n_1172), .B(n_1192), .C(n_1255), .Y(n_1308) );
AND2x2_ASAP7_75t_L g1341 ( .A(n_1172), .B(n_1203), .Y(n_1341) );
INVx2_ASAP7_75t_L g1172 ( .A(n_1173), .Y(n_1172) );
BUFx2_ASAP7_75t_L g1198 ( .A(n_1173), .Y(n_1198) );
INVx2_ASAP7_75t_L g1220 ( .A(n_1173), .Y(n_1220) );
NAND2xp5_ASAP7_75t_L g1268 ( .A(n_1173), .B(n_1203), .Y(n_1268) );
NAND2xp5_ASAP7_75t_L g1307 ( .A(n_1173), .B(n_1215), .Y(n_1307) );
AND2x2_ASAP7_75t_L g1319 ( .A(n_1173), .B(n_1211), .Y(n_1319) );
AND2x2_ASAP7_75t_L g1332 ( .A(n_1173), .B(n_1247), .Y(n_1332) );
OR2x2_ASAP7_75t_L g1356 ( .A(n_1173), .B(n_1182), .Y(n_1356) );
AND2x2_ASAP7_75t_L g1173 ( .A(n_1174), .B(n_1180), .Y(n_1173) );
AND2x4_ASAP7_75t_L g1175 ( .A(n_1176), .B(n_1177), .Y(n_1175) );
AND2x4_ASAP7_75t_L g1178 ( .A(n_1177), .B(n_1179), .Y(n_1178) );
BUFx2_ASAP7_75t_L g1227 ( .A(n_1178), .Y(n_1227) );
INVx1_ASAP7_75t_L g1298 ( .A(n_1181), .Y(n_1298) );
NOR2xp33_ASAP7_75t_L g1306 ( .A(n_1181), .B(n_1203), .Y(n_1306) );
AND2x2_ASAP7_75t_L g1181 ( .A(n_1182), .B(n_1187), .Y(n_1181) );
OR2x2_ASAP7_75t_L g1251 ( .A(n_1182), .B(n_1212), .Y(n_1251) );
AND2x2_ASAP7_75t_L g1280 ( .A(n_1182), .B(n_1281), .Y(n_1280) );
AND2x2_ASAP7_75t_L g1290 ( .A(n_1182), .B(n_1191), .Y(n_1290) );
AND2x2_ASAP7_75t_L g1350 ( .A(n_1182), .B(n_1192), .Y(n_1350) );
BUFx3_ASAP7_75t_L g1182 ( .A(n_1183), .Y(n_1182) );
INVxp67_ASAP7_75t_L g1204 ( .A(n_1183), .Y(n_1204) );
BUFx2_ASAP7_75t_L g1211 ( .A(n_1183), .Y(n_1211) );
AND2x2_ASAP7_75t_L g1323 ( .A(n_1183), .B(n_1243), .Y(n_1323) );
OR2x2_ASAP7_75t_L g1330 ( .A(n_1183), .B(n_1192), .Y(n_1330) );
AND2x2_ASAP7_75t_L g1183 ( .A(n_1184), .B(n_1185), .Y(n_1183) );
INVx1_ASAP7_75t_L g1272 ( .A(n_1187), .Y(n_1272) );
NAND2xp5_ASAP7_75t_L g1327 ( .A(n_1187), .B(n_1204), .Y(n_1327) );
AND2x2_ASAP7_75t_L g1187 ( .A(n_1188), .B(n_1191), .Y(n_1187) );
INVx2_ASAP7_75t_L g1206 ( .A(n_1188), .Y(n_1206) );
AND2x2_ASAP7_75t_L g1213 ( .A(n_1188), .B(n_1192), .Y(n_1213) );
OR2x2_ASAP7_75t_L g1244 ( .A(n_1188), .B(n_1192), .Y(n_1244) );
AND2x2_ASAP7_75t_L g1188 ( .A(n_1189), .B(n_1190), .Y(n_1188) );
AOI221xp5_ASAP7_75t_L g1196 ( .A1(n_1191), .A2(n_1197), .B1(n_1203), .B2(n_1207), .C(n_1208), .Y(n_1196) );
NOR2x1_ASAP7_75t_L g1264 ( .A(n_1191), .B(n_1211), .Y(n_1264) );
INVx2_ASAP7_75t_SL g1191 ( .A(n_1192), .Y(n_1191) );
AND2x2_ASAP7_75t_L g1205 ( .A(n_1192), .B(n_1206), .Y(n_1205) );
INVx1_ASAP7_75t_L g1313 ( .A(n_1197), .Y(n_1313) );
AND2x2_ASAP7_75t_L g1197 ( .A(n_1198), .B(n_1199), .Y(n_1197) );
INVx2_ASAP7_75t_L g1250 ( .A(n_1198), .Y(n_1250) );
NAND2xp5_ASAP7_75t_L g1284 ( .A(n_1198), .B(n_1285), .Y(n_1284) );
AND2x2_ASAP7_75t_L g1300 ( .A(n_1198), .B(n_1210), .Y(n_1300) );
INVx1_ASAP7_75t_L g1240 ( .A(n_1199), .Y(n_1240) );
OAI221xp5_ASAP7_75t_L g1208 ( .A1(n_1200), .A2(n_1209), .B1(n_1212), .B2(n_1214), .C(n_1217), .Y(n_1208) );
INVx3_ASAP7_75t_L g1216 ( .A(n_1200), .Y(n_1216) );
AND2x2_ASAP7_75t_L g1234 ( .A(n_1200), .B(n_1224), .Y(n_1234) );
OR2x2_ASAP7_75t_L g1275 ( .A(n_1200), .B(n_1225), .Y(n_1275) );
AND2x2_ASAP7_75t_L g1200 ( .A(n_1201), .B(n_1202), .Y(n_1200) );
O2A1O1Ixp33_ASAP7_75t_L g1338 ( .A1(n_1203), .A2(n_1265), .B(n_1323), .C(n_1339), .Y(n_1338) );
AND2x2_ASAP7_75t_L g1203 ( .A(n_1204), .B(n_1205), .Y(n_1203) );
AND2x2_ASAP7_75t_L g1242 ( .A(n_1204), .B(n_1243), .Y(n_1242) );
AOI322xp5_ASAP7_75t_L g1269 ( .A1(n_1204), .A2(n_1216), .A3(n_1270), .B1(n_1274), .B2(n_1276), .C1(n_1277), .C2(n_1280), .Y(n_1269) );
AND2x2_ASAP7_75t_L g1334 ( .A(n_1204), .B(n_1335), .Y(n_1334) );
AND2x2_ASAP7_75t_L g1221 ( .A(n_1205), .B(n_1220), .Y(n_1221) );
AND2x2_ASAP7_75t_L g1238 ( .A(n_1205), .B(n_1211), .Y(n_1238) );
OAI21xp33_ASAP7_75t_L g1252 ( .A1(n_1205), .A2(n_1210), .B(n_1218), .Y(n_1252) );
INVx1_ASAP7_75t_L g1273 ( .A(n_1205), .Y(n_1273) );
AND2x2_ASAP7_75t_L g1318 ( .A(n_1205), .B(n_1319), .Y(n_1318) );
NOR2xp33_ASAP7_75t_L g1210 ( .A(n_1206), .B(n_1211), .Y(n_1210) );
AOI21xp5_ASAP7_75t_L g1217 ( .A1(n_1206), .A2(n_1218), .B(n_1221), .Y(n_1217) );
NAND4xp25_ASAP7_75t_L g1309 ( .A(n_1206), .B(n_1255), .C(n_1296), .D(n_1310), .Y(n_1309) );
INVx1_ASAP7_75t_L g1235 ( .A(n_1210), .Y(n_1235) );
AND2x2_ASAP7_75t_L g1360 ( .A(n_1211), .B(n_1213), .Y(n_1360) );
INVx1_ASAP7_75t_L g1212 ( .A(n_1213), .Y(n_1212) );
AND2x2_ASAP7_75t_L g1281 ( .A(n_1213), .B(n_1220), .Y(n_1281) );
NAND2xp5_ASAP7_75t_L g1361 ( .A(n_1213), .B(n_1362), .Y(n_1361) );
OAI222xp33_ASAP7_75t_SL g1354 ( .A1(n_1214), .A2(n_1294), .B1(n_1355), .B2(n_1357), .C1(n_1359), .C2(n_1361), .Y(n_1354) );
INVx1_ASAP7_75t_L g1214 ( .A(n_1215), .Y(n_1214) );
INVx1_ASAP7_75t_L g1276 ( .A(n_1216), .Y(n_1276) );
OR2x2_ASAP7_75t_L g1316 ( .A(n_1216), .B(n_1317), .Y(n_1316) );
AND2x2_ASAP7_75t_L g1358 ( .A(n_1216), .B(n_1225), .Y(n_1358) );
NAND2xp5_ASAP7_75t_L g1287 ( .A(n_1218), .B(n_1288), .Y(n_1287) );
AND2x2_ASAP7_75t_L g1218 ( .A(n_1219), .B(n_1220), .Y(n_1218) );
INVx2_ASAP7_75t_L g1237 ( .A(n_1219), .Y(n_1237) );
NOR2xp33_ASAP7_75t_L g1274 ( .A(n_1219), .B(n_1275), .Y(n_1274) );
NOR2xp33_ASAP7_75t_L g1315 ( .A(n_1219), .B(n_1316), .Y(n_1315) );
NAND2xp5_ASAP7_75t_L g1351 ( .A(n_1219), .B(n_1352), .Y(n_1351) );
NOR2xp33_ASAP7_75t_L g1335 ( .A(n_1220), .B(n_1244), .Y(n_1335) );
NAND2xp5_ASAP7_75t_L g1346 ( .A(n_1220), .B(n_1322), .Y(n_1346) );
AND2x2_ASAP7_75t_L g1349 ( .A(n_1220), .B(n_1350), .Y(n_1349) );
O2A1O1Ixp33_ASAP7_75t_L g1347 ( .A1(n_1222), .A2(n_1276), .B(n_1348), .C(n_1351), .Y(n_1347) );
INVx2_ASAP7_75t_L g1222 ( .A(n_1223), .Y(n_1222) );
AND2x2_ASAP7_75t_L g1301 ( .A(n_1223), .B(n_1233), .Y(n_1301) );
AND2x2_ASAP7_75t_L g1321 ( .A(n_1223), .B(n_1322), .Y(n_1321) );
INVx1_ASAP7_75t_L g1223 ( .A(n_1224), .Y(n_1223) );
INVx1_ASAP7_75t_L g1289 ( .A(n_1224), .Y(n_1289) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1225), .Y(n_1224) );
INVx1_ASAP7_75t_L g1247 ( .A(n_1225), .Y(n_1247) );
INVx1_ASAP7_75t_L g1317 ( .A(n_1225), .Y(n_1317) );
AND2x2_ASAP7_75t_L g1225 ( .A(n_1226), .B(n_1228), .Y(n_1225) );
NOR3xp33_ASAP7_75t_L g1230 ( .A(n_1231), .B(n_1239), .C(n_1248), .Y(n_1230) );
OAI21xp33_ASAP7_75t_L g1231 ( .A1(n_1232), .A2(n_1235), .B(n_1236), .Y(n_1231) );
INVx1_ASAP7_75t_L g1328 ( .A(n_1232), .Y(n_1328) );
NAND2xp5_ASAP7_75t_L g1232 ( .A(n_1233), .B(n_1234), .Y(n_1232) );
NAND2xp5_ASAP7_75t_L g1357 ( .A(n_1233), .B(n_1358), .Y(n_1357) );
NAND2xp5_ASAP7_75t_L g1249 ( .A(n_1234), .B(n_1250), .Y(n_1249) );
INVx1_ASAP7_75t_L g1337 ( .A(n_1234), .Y(n_1337) );
NAND2xp5_ASAP7_75t_L g1236 ( .A(n_1237), .B(n_1238), .Y(n_1236) );
INVx1_ASAP7_75t_L g1245 ( .A(n_1238), .Y(n_1245) );
AOI22xp5_ASAP7_75t_L g1295 ( .A1(n_1238), .A2(n_1296), .B1(n_1297), .B2(n_1301), .Y(n_1295) );
AND2x2_ASAP7_75t_L g1339 ( .A(n_1238), .B(n_1279), .Y(n_1339) );
O2A1O1Ixp33_ASAP7_75t_L g1239 ( .A1(n_1240), .A2(n_1241), .B(n_1245), .C(n_1246), .Y(n_1239) );
INVx1_ASAP7_75t_L g1241 ( .A(n_1242), .Y(n_1241) );
INVx1_ASAP7_75t_L g1243 ( .A(n_1244), .Y(n_1243) );
A2O1A1Ixp33_ASAP7_75t_L g1329 ( .A1(n_1245), .A2(n_1330), .B(n_1331), .C(n_1333), .Y(n_1329) );
NOR3xp33_ASAP7_75t_L g1277 ( .A(n_1246), .B(n_1272), .C(n_1278), .Y(n_1277) );
INVx1_ASAP7_75t_L g1246 ( .A(n_1247), .Y(n_1246) );
A2O1A1Ixp33_ASAP7_75t_L g1263 ( .A1(n_1247), .A2(n_1264), .B(n_1265), .C(n_1267), .Y(n_1263) );
OAI21xp33_ASAP7_75t_L g1248 ( .A1(n_1249), .A2(n_1251), .B(n_1252), .Y(n_1248) );
OR2x2_ASAP7_75t_L g1326 ( .A(n_1250), .B(n_1327), .Y(n_1326) );
NAND2xp5_ASAP7_75t_L g1353 ( .A(n_1250), .B(n_1264), .Y(n_1353) );
NOR2xp33_ASAP7_75t_L g1291 ( .A(n_1251), .B(n_1292), .Y(n_1291) );
INVx2_ASAP7_75t_L g1253 ( .A(n_1254), .Y(n_1253) );
INVx3_ASAP7_75t_L g1254 ( .A(n_1255), .Y(n_1254) );
NAND2xp5_ASAP7_75t_L g1312 ( .A(n_1255), .B(n_1290), .Y(n_1312) );
OAI22xp33_ASAP7_75t_L g1257 ( .A1(n_1258), .A2(n_1259), .B1(n_1260), .B2(n_1261), .Y(n_1257) );
NAND4xp25_ASAP7_75t_SL g1262 ( .A(n_1263), .B(n_1269), .C(n_1282), .D(n_1295), .Y(n_1262) );
INVx1_ASAP7_75t_L g1265 ( .A(n_1266), .Y(n_1265) );
INVx1_ASAP7_75t_L g1267 ( .A(n_1268), .Y(n_1267) );
INVx1_ASAP7_75t_L g1270 ( .A(n_1271), .Y(n_1270) );
NAND2xp5_ASAP7_75t_L g1271 ( .A(n_1272), .B(n_1273), .Y(n_1271) );
OR2x2_ASAP7_75t_L g1355 ( .A(n_1272), .B(n_1356), .Y(n_1355) );
INVx1_ASAP7_75t_L g1296 ( .A(n_1275), .Y(n_1296) );
INVx1_ASAP7_75t_L g1278 ( .A(n_1279), .Y(n_1278) );
O2A1O1Ixp33_ASAP7_75t_L g1282 ( .A1(n_1283), .A2(n_1286), .B(n_1290), .C(n_1291), .Y(n_1282) );
INVx1_ASAP7_75t_L g1283 ( .A(n_1284), .Y(n_1283) );
CKINVDCx5p33_ASAP7_75t_R g1294 ( .A(n_1285), .Y(n_1294) );
INVx1_ASAP7_75t_L g1286 ( .A(n_1287), .Y(n_1286) );
INVx1_ASAP7_75t_L g1288 ( .A(n_1289), .Y(n_1288) );
INVx1_ASAP7_75t_L g1293 ( .A(n_1289), .Y(n_1293) );
INVx1_ASAP7_75t_L g1345 ( .A(n_1290), .Y(n_1345) );
OR2x2_ASAP7_75t_L g1292 ( .A(n_1293), .B(n_1294), .Y(n_1292) );
OAI221xp5_ASAP7_75t_SL g1305 ( .A1(n_1294), .A2(n_1306), .B1(n_1307), .B2(n_1308), .C(n_1309), .Y(n_1305) );
NAND2xp5_ASAP7_75t_L g1297 ( .A(n_1298), .B(n_1299), .Y(n_1297) );
INVx1_ASAP7_75t_L g1299 ( .A(n_1300), .Y(n_1299) );
NAND3xp33_ASAP7_75t_L g1302 ( .A(n_1303), .B(n_1324), .C(n_1343), .Y(n_1302) );
NOR4xp25_ASAP7_75t_SL g1303 ( .A(n_1304), .B(n_1305), .C(n_1311), .D(n_1320), .Y(n_1303) );
OAI21xp33_ASAP7_75t_L g1311 ( .A1(n_1312), .A2(n_1313), .B(n_1314), .Y(n_1311) );
NAND2xp5_ASAP7_75t_L g1314 ( .A(n_1315), .B(n_1318), .Y(n_1314) );
INVx1_ASAP7_75t_L g1342 ( .A(n_1316), .Y(n_1342) );
AND2x2_ASAP7_75t_L g1320 ( .A(n_1321), .B(n_1323), .Y(n_1320) );
AOI221xp5_ASAP7_75t_L g1324 ( .A1(n_1322), .A2(n_1325), .B1(n_1328), .B2(n_1329), .C(n_1336), .Y(n_1324) );
INVx1_ASAP7_75t_L g1325 ( .A(n_1326), .Y(n_1325) );
INVx1_ASAP7_75t_L g1331 ( .A(n_1332), .Y(n_1331) );
INVx1_ASAP7_75t_L g1333 ( .A(n_1334), .Y(n_1333) );
OAI21xp5_ASAP7_75t_L g1340 ( .A1(n_1334), .A2(n_1341), .B(n_1342), .Y(n_1340) );
OAI21xp5_ASAP7_75t_L g1336 ( .A1(n_1337), .A2(n_1338), .B(n_1340), .Y(n_1336) );
NOR3xp33_ASAP7_75t_SL g1343 ( .A(n_1344), .B(n_1347), .C(n_1354), .Y(n_1343) );
NOR2xp33_ASAP7_75t_L g1344 ( .A(n_1345), .B(n_1346), .Y(n_1344) );
INVx1_ASAP7_75t_L g1348 ( .A(n_1349), .Y(n_1348) );
INVx1_ASAP7_75t_L g1352 ( .A(n_1353), .Y(n_1352) );
INVx1_ASAP7_75t_L g1362 ( .A(n_1356), .Y(n_1362) );
INVx1_ASAP7_75t_L g1359 ( .A(n_1360), .Y(n_1359) );
CKINVDCx5p33_ASAP7_75t_R g1363 ( .A(n_1364), .Y(n_1363) );
INVx1_ASAP7_75t_L g1364 ( .A(n_1365), .Y(n_1364) );
INVx1_ASAP7_75t_L g1365 ( .A(n_1366), .Y(n_1365) );
INVx1_ASAP7_75t_L g1367 ( .A(n_1368), .Y(n_1367) );
INVx1_ASAP7_75t_L g1368 ( .A(n_1369), .Y(n_1368) );
INVx1_ASAP7_75t_L g1370 ( .A(n_1371), .Y(n_1370) );
NAND2xp5_ASAP7_75t_L g1371 ( .A(n_1372), .B(n_1406), .Y(n_1371) );
NOR3xp33_ASAP7_75t_L g1372 ( .A(n_1373), .B(n_1396), .C(n_1399), .Y(n_1372) );
OAI22xp5_ASAP7_75t_L g1374 ( .A1(n_1375), .A2(n_1376), .B1(n_1377), .B2(n_1378), .Y(n_1374) );
OAI22xp33_ASAP7_75t_L g1379 ( .A1(n_1380), .A2(n_1381), .B1(n_1383), .B2(n_1384), .Y(n_1379) );
INVx1_ASAP7_75t_L g1381 ( .A(n_1382), .Y(n_1381) );
INVx1_ASAP7_75t_L g1387 ( .A(n_1388), .Y(n_1387) );
OAI22xp5_ASAP7_75t_L g1391 ( .A1(n_1392), .A2(n_1393), .B1(n_1394), .B2(n_1395), .Y(n_1391) );
NAND2xp5_ASAP7_75t_L g1399 ( .A(n_1400), .B(n_1403), .Y(n_1399) );
AOI22xp5_ASAP7_75t_L g1406 ( .A1(n_1407), .A2(n_1408), .B1(n_1430), .B2(n_1431), .Y(n_1406) );
NAND4xp25_ASAP7_75t_L g1408 ( .A(n_1409), .B(n_1419), .C(n_1428), .D(n_1429), .Y(n_1408) );
INVx1_ASAP7_75t_L g1410 ( .A(n_1411), .Y(n_1410) );
INVx3_ASAP7_75t_L g1413 ( .A(n_1414), .Y(n_1413) );
INVx2_ASAP7_75t_L g1416 ( .A(n_1417), .Y(n_1416) );
INVx1_ASAP7_75t_L g1417 ( .A(n_1418), .Y(n_1417) );
INVx2_ASAP7_75t_L g1433 ( .A(n_1434), .Y(n_1433) );
INVx1_ASAP7_75t_L g1434 ( .A(n_1435), .Y(n_1434) );
INVx1_ASAP7_75t_L g1435 ( .A(n_1436), .Y(n_1435) );
INVx1_ASAP7_75t_L g1438 ( .A(n_1439), .Y(n_1438) );
CKINVDCx5p33_ASAP7_75t_R g1439 ( .A(n_1440), .Y(n_1439) );
A2O1A1Ixp33_ASAP7_75t_L g1507 ( .A1(n_1441), .A2(n_1508), .B(n_1510), .C(n_1512), .Y(n_1507) );
INVxp33_ASAP7_75t_SL g1442 ( .A(n_1443), .Y(n_1442) );
HB1xp67_ASAP7_75t_L g1444 ( .A(n_1445), .Y(n_1444) );
AND4x1_ASAP7_75t_L g1445 ( .A(n_1446), .B(n_1470), .C(n_1472), .D(n_1498), .Y(n_1445) );
NOR3xp33_ASAP7_75t_SL g1446 ( .A(n_1447), .B(n_1448), .C(n_1450), .Y(n_1446) );
BUFx2_ASAP7_75t_L g1452 ( .A(n_1453), .Y(n_1452) );
INVx2_ASAP7_75t_L g1453 ( .A(n_1454), .Y(n_1453) );
CKINVDCx5p33_ASAP7_75t_R g1458 ( .A(n_1459), .Y(n_1458) );
OAI221xp5_ASAP7_75t_L g1460 ( .A1(n_1461), .A2(n_1462), .B1(n_1463), .B2(n_1465), .C(n_1466), .Y(n_1460) );
BUFx2_ASAP7_75t_L g1463 ( .A(n_1464), .Y(n_1463) );
BUFx3_ASAP7_75t_L g1467 ( .A(n_1468), .Y(n_1467) );
OAI31xp33_ASAP7_75t_L g1472 ( .A1(n_1473), .A2(n_1484), .A3(n_1495), .B(n_1497), .Y(n_1472) );
OAI221xp5_ASAP7_75t_L g1474 ( .A1(n_1475), .A2(n_1477), .B1(n_1478), .B2(n_1479), .C(n_1480), .Y(n_1474) );
INVx1_ASAP7_75t_L g1475 ( .A(n_1476), .Y(n_1475) );
OAI22xp5_ASAP7_75t_L g1487 ( .A1(n_1488), .A2(n_1491), .B1(n_1492), .B2(n_1494), .Y(n_1487) );
INVx1_ASAP7_75t_L g1488 ( .A(n_1489), .Y(n_1488) );
INVx1_ASAP7_75t_L g1489 ( .A(n_1490), .Y(n_1489) );
CKINVDCx5p33_ASAP7_75t_R g1492 ( .A(n_1493), .Y(n_1492) );
NOR2xp33_ASAP7_75t_L g1498 ( .A(n_1499), .B(n_1501), .Y(n_1498) );
HB1xp67_ASAP7_75t_L g1506 ( .A(n_1507), .Y(n_1506) );
INVx1_ASAP7_75t_L g1508 ( .A(n_1509), .Y(n_1508) );
INVx1_ASAP7_75t_L g1510 ( .A(n_1511), .Y(n_1510) );
endmodule