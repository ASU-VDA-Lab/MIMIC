module fake_jpeg_4343_n_327 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_327);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_327;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx8_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx4f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_8),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_34),
.B(n_36),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_33),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_42),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_18),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_57),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_42),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_58),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_34),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_59),
.Y(n_77)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_61),
.A2(n_29),
.B1(n_16),
.B2(n_23),
.Y(n_87)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_63),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_20),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_64),
.B(n_22),
.Y(n_81)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_24),
.Y(n_79)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_64),
.B(n_20),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_69),
.B(n_92),
.Y(n_100)
);

O2A1O1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_60),
.A2(n_30),
.B(n_21),
.C(n_29),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_75),
.Y(n_103)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_81),
.B(n_93),
.Y(n_95)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_84),
.Y(n_99)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_48),
.A2(n_32),
.B(n_36),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_54),
.B(n_32),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_28),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_87),
.A2(n_90),
.B1(n_25),
.B2(n_23),
.Y(n_108)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_88),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_52),
.A2(n_29),
.B1(n_25),
.B2(n_16),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_89),
.A2(n_16),
.B1(n_32),
.B2(n_25),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_46),
.Y(n_90)
);

CKINVDCx12_ASAP7_75t_R g91 ( 
.A(n_56),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_91),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_62),
.B(n_28),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_53),
.B(n_18),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_94),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_97),
.B(n_101),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_65),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_77),
.A2(n_53),
.B1(n_61),
.B2(n_51),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_102),
.A2(n_106),
.B1(n_112),
.B2(n_71),
.Y(n_136)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_104),
.B(n_105),
.Y(n_131)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_69),
.A2(n_51),
.B1(n_52),
.B2(n_55),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_107),
.A2(n_116),
.B1(n_71),
.B2(n_74),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_108),
.Y(n_137)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_73),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_109),
.B(n_117),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_77),
.B(n_68),
.Y(n_110)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_110),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_90),
.A2(n_50),
.B1(n_23),
.B2(n_31),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_111),
.A2(n_71),
.B1(n_74),
.B2(n_82),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_81),
.A2(n_50),
.B1(n_63),
.B2(n_57),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_69),
.B(n_93),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_113),
.B(n_20),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_72),
.B(n_17),
.Y(n_114)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_114),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_85),
.A2(n_31),
.B1(n_17),
.B2(n_26),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_73),
.Y(n_117)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_92),
.Y(n_119)
);

INVx13_ASAP7_75t_L g126 ( 
.A(n_119),
.Y(n_126)
);

AOI32xp33_ASAP7_75t_L g121 ( 
.A1(n_72),
.A2(n_19),
.A3(n_47),
.B1(n_66),
.B2(n_21),
.Y(n_121)
);

CKINVDCx12_ASAP7_75t_R g146 ( 
.A(n_121),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_78),
.B(n_26),
.Y(n_122)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_122),
.Y(n_138)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_120),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_124),
.B(n_136),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_95),
.B(n_93),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_125),
.B(n_140),
.Y(n_156)
);

AND2x6_ASAP7_75t_L g128 ( 
.A(n_96),
.B(n_75),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_128),
.B(n_102),
.Y(n_161)
);

BUFx12f_ASAP7_75t_L g129 ( 
.A(n_115),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_129),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_132),
.A2(n_134),
.B1(n_105),
.B2(n_76),
.Y(n_169)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_103),
.B(n_75),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_133),
.A2(n_135),
.B(n_139),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_96),
.A2(n_79),
.B(n_70),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_101),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_113),
.A2(n_74),
.B1(n_84),
.B2(n_76),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_141),
.A2(n_137),
.B(n_106),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_95),
.B(n_113),
.Y(n_142)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_142),
.Y(n_163)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_120),
.Y(n_143)
);

INVxp67_ASAP7_75t_SL g154 ( 
.A(n_143),
.Y(n_154)
);

INVx13_ASAP7_75t_L g144 ( 
.A(n_109),
.Y(n_144)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_144),
.Y(n_171)
);

INVx13_ASAP7_75t_L g145 ( 
.A(n_117),
.Y(n_145)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_145),
.Y(n_172)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_97),
.Y(n_147)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_147),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_128),
.A2(n_142),
.B(n_139),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_149),
.A2(n_144),
.B1(n_126),
.B2(n_104),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_140),
.A2(n_98),
.B(n_110),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_150),
.B(n_152),
.C(n_162),
.Y(n_190)
);

MAJx2_ASAP7_75t_L g152 ( 
.A(n_135),
.B(n_125),
.C(n_123),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_137),
.A2(n_95),
.B1(n_119),
.B2(n_100),
.Y(n_153)
);

OAI21xp33_ASAP7_75t_SL g185 ( 
.A1(n_153),
.A2(n_159),
.B(n_166),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_131),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_155),
.B(n_161),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_157),
.A2(n_168),
.B1(n_169),
.B2(n_175),
.Y(n_196)
);

INVx2_ASAP7_75t_SL g158 ( 
.A(n_131),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_158),
.B(n_174),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_135),
.A2(n_100),
.B1(n_98),
.B2(n_112),
.Y(n_159)
);

MAJx2_ASAP7_75t_L g162 ( 
.A(n_123),
.B(n_114),
.C(n_122),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_136),
.B(n_99),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_164),
.B(n_167),
.Y(n_177)
);

OAI21xp33_ASAP7_75t_SL g166 ( 
.A1(n_141),
.A2(n_78),
.B(n_70),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_146),
.B(n_91),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_146),
.A2(n_133),
.B1(n_147),
.B2(n_127),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_127),
.B(n_115),
.C(n_80),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_170),
.B(n_176),
.Y(n_184)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_148),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_148),
.A2(n_80),
.B(n_2),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_133),
.B(n_120),
.Y(n_176)
);

INVx13_ASAP7_75t_L g178 ( 
.A(n_154),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_178),
.B(n_182),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_156),
.B(n_130),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_180),
.B(n_193),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_161),
.A2(n_130),
.B1(n_138),
.B2(n_76),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_181),
.A2(n_157),
.B1(n_168),
.B2(n_152),
.Y(n_212)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_170),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_158),
.A2(n_124),
.B1(n_143),
.B2(n_138),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_183),
.A2(n_203),
.B(n_27),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_150),
.B(n_129),
.Y(n_186)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_186),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_160),
.B(n_126),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_187),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_172),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_188),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_163),
.B(n_129),
.Y(n_189)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_189),
.Y(n_207)
);

INVx13_ASAP7_75t_L g191 ( 
.A(n_172),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_191),
.B(n_194),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_153),
.B(n_145),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_192),
.B(n_197),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_173),
.B(n_145),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_171),
.Y(n_194)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_165),
.Y(n_197)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_171),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_198),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_164),
.B(n_129),
.Y(n_199)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_199),
.Y(n_208)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_175),
.Y(n_200)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_200),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_159),
.B(n_144),
.Y(n_201)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_201),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_202),
.B(n_151),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_158),
.A2(n_82),
.B1(n_126),
.B2(n_94),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_195),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_205),
.B(n_213),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_212),
.A2(n_201),
.B1(n_196),
.B2(n_179),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_189),
.B(n_162),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_190),
.B(n_149),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_214),
.B(n_178),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_184),
.B(n_176),
.C(n_151),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_216),
.B(n_225),
.C(n_208),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_217),
.A2(n_224),
.B(n_226),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_221),
.B(n_190),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_177),
.B(n_167),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_222),
.B(n_177),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_191),
.Y(n_223)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_223),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_195),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_184),
.B(n_118),
.C(n_94),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_186),
.A2(n_94),
.B(n_118),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_188),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_228),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g263 ( 
.A(n_229),
.B(n_210),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_212),
.B(n_199),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_SL g259 ( 
.A(n_230),
.B(n_247),
.C(n_250),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_231),
.B(n_236),
.C(n_245),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_232),
.B(n_233),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_216),
.B(n_182),
.C(n_181),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_211),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_237),
.B(n_239),
.Y(n_251)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_218),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_206),
.A2(n_196),
.B1(n_197),
.B2(n_185),
.Y(n_240)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_240),
.Y(n_252)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_218),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_241),
.B(n_207),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_206),
.A2(n_192),
.B1(n_202),
.B2(n_200),
.Y(n_242)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_242),
.Y(n_255)
);

OR2x2_ASAP7_75t_L g243 ( 
.A(n_224),
.B(n_180),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_243),
.B(n_249),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_225),
.B(n_193),
.C(n_194),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_227),
.A2(n_198),
.B1(n_178),
.B2(n_191),
.Y(n_246)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_246),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_221),
.B(n_118),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_248),
.B(n_226),
.Y(n_254)
);

OR2x2_ASAP7_75t_L g249 ( 
.A(n_228),
.B(n_24),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_222),
.B(n_24),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_253),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_254),
.B(n_250),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_238),
.B(n_207),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_256),
.A2(n_258),
.B(n_265),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_235),
.A2(n_227),
.B1(n_208),
.B2(n_215),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_257),
.A2(n_229),
.B1(n_236),
.B2(n_245),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_244),
.B(n_219),
.Y(n_258)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_234),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_262),
.B(n_243),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_263),
.B(n_230),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_235),
.A2(n_209),
.B(n_220),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_240),
.A2(n_215),
.B1(n_219),
.B2(n_220),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_266),
.A2(n_233),
.B1(n_2),
.B2(n_3),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_231),
.B(n_217),
.C(n_204),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_268),
.B(n_248),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_269),
.A2(n_270),
.B(n_275),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_261),
.B(n_246),
.Y(n_270)
);

BUFx2_ASAP7_75t_L g271 ( 
.A(n_262),
.Y(n_271)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_271),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_272),
.B(n_276),
.Y(n_285)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_273),
.Y(n_294)
);

BUFx24_ASAP7_75t_SL g274 ( 
.A(n_255),
.Y(n_274)
);

NOR2xp67_ASAP7_75t_SL g287 ( 
.A(n_274),
.B(n_259),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_257),
.B(n_249),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_277),
.B(n_280),
.C(n_260),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_263),
.B(n_232),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_278),
.B(n_264),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_279),
.A2(n_282),
.B1(n_261),
.B2(n_252),
.Y(n_286)
);

BUFx12_ASAP7_75t_L g280 ( 
.A(n_266),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_9),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_284),
.B(n_292),
.C(n_293),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_286),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_287),
.B(n_272),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_281),
.A2(n_268),
.B1(n_260),
.B2(n_251),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_288),
.B(n_291),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_283),
.A2(n_254),
.B1(n_264),
.B2(n_10),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_277),
.B(n_1),
.C(n_3),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_278),
.B(n_9),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_295),
.B(n_8),
.C(n_14),
.Y(n_304)
);

NOR2x1_ASAP7_75t_SL g296 ( 
.A(n_280),
.B(n_9),
.Y(n_296)
);

OR2x2_ASAP7_75t_L g299 ( 
.A(n_296),
.B(n_8),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_297),
.B(n_299),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_294),
.A2(n_280),
.B(n_271),
.Y(n_298)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_298),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_289),
.B(n_1),
.Y(n_300)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_300),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_290),
.B(n_1),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_301),
.B(n_1),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_304),
.B(n_305),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_284),
.B(n_10),
.C(n_14),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_301),
.B(n_295),
.Y(n_310)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_310),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_306),
.B(n_285),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_311),
.B(n_302),
.C(n_292),
.Y(n_315)
);

AOI322xp5_ASAP7_75t_L g317 ( 
.A1(n_312),
.A2(n_314),
.A3(n_10),
.B1(n_13),
.B2(n_12),
.C1(n_11),
.C2(n_15),
.Y(n_317)
);

AOI21x1_ASAP7_75t_L g314 ( 
.A1(n_303),
.A2(n_285),
.B(n_293),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_315),
.B(n_317),
.Y(n_320)
);

NOR2x1_ASAP7_75t_L g318 ( 
.A(n_307),
.B(n_12),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_318),
.B(n_319),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_308),
.A2(n_15),
.B(n_12),
.Y(n_319)
);

AOI322xp5_ASAP7_75t_L g322 ( 
.A1(n_320),
.A2(n_316),
.A3(n_313),
.B1(n_309),
.B2(n_312),
.C1(n_3),
.C2(n_6),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_321),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_323),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_324),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_325),
.A2(n_5),
.B1(n_7),
.B2(n_321),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_7),
.Y(n_327)
);


endmodule