module fake_netlist_5_911_n_1920 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1920);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1920;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_164;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1891;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_759;
wire n_1892;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_1916;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_252;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_448;
wire n_259;
wire n_1851;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_1874;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_1902;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1875;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_174;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_968;
wire n_912;
wire n_315;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_753;
wire n_621;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1363;
wire n_1301;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1400;
wire n_1342;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_990;
wire n_836;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1834;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_172;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_1904;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_177;
wire n_421;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1898;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_242;
wire n_1032;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

BUFx2_ASAP7_75t_L g158 ( 
.A(n_156),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_40),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_1),
.Y(n_160)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_50),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_124),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_64),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_132),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_114),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_22),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_39),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_90),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_29),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_121),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_99),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_42),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_92),
.Y(n_173)
);

INVx2_ASAP7_75t_SL g174 ( 
.A(n_98),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_57),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_26),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_103),
.Y(n_177)
);

BUFx8_ASAP7_75t_SL g178 ( 
.A(n_80),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_110),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_106),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_43),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_113),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_53),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_24),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_157),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_86),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_7),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_84),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_11),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_37),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_72),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_153),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_68),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_45),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_149),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_37),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_14),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_32),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_130),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_141),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_137),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_9),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_111),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_19),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_31),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_46),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_144),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_129),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_76),
.Y(n_209)
);

INVx2_ASAP7_75t_SL g210 ( 
.A(n_126),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_96),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_29),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_33),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_22),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_117),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_54),
.Y(n_216)
);

INVx2_ASAP7_75t_SL g217 ( 
.A(n_105),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_27),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_52),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_101),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_63),
.Y(n_221)
);

BUFx8_ASAP7_75t_SL g222 ( 
.A(n_85),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_21),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_28),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_30),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_44),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_5),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_151),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_83),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_78),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_71),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_27),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_10),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_34),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_135),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_2),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_10),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_66),
.Y(n_238)
);

BUFx2_ASAP7_75t_L g239 ( 
.A(n_139),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_94),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_60),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_81),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_75),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_5),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_6),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_134),
.Y(n_246)
);

BUFx8_ASAP7_75t_SL g247 ( 
.A(n_79),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_35),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_109),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_19),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_11),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_56),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_2),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_128),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_120),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_118),
.Y(n_256)
);

INVx2_ASAP7_75t_SL g257 ( 
.A(n_3),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_145),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_93),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_89),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_3),
.Y(n_261)
);

BUFx5_ASAP7_75t_L g262 ( 
.A(n_112),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_67),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_108),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_147),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_16),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_51),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_87),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_123),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_70),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_9),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_48),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_31),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_150),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_133),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_58),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_6),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_125),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_119),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_8),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_32),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_47),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_14),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_74),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_91),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_17),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_136),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_138),
.Y(n_288)
);

HB1xp67_ASAP7_75t_L g289 ( 
.A(n_49),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_34),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_13),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_115),
.Y(n_292)
);

INVx1_ASAP7_75t_SL g293 ( 
.A(n_8),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_77),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_143),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_7),
.Y(n_296)
);

BUFx10_ASAP7_75t_L g297 ( 
.A(n_116),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_88),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_142),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_30),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_62),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_33),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_100),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_12),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_28),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_104),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_0),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_127),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_41),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_1),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_0),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_18),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_82),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_311),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_204),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_311),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_311),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_204),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_170),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_271),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_170),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_311),
.Y(n_322)
);

INVxp67_ASAP7_75t_SL g323 ( 
.A(n_161),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_250),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_225),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_166),
.Y(n_326)
);

INVxp67_ASAP7_75t_SL g327 ( 
.A(n_289),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_187),
.Y(n_328)
);

INVxp33_ASAP7_75t_SL g329 ( 
.A(n_169),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_311),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_160),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_185),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_160),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_169),
.Y(n_334)
);

INVxp67_ASAP7_75t_SL g335 ( 
.A(n_158),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_226),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_271),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_184),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_213),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_197),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_185),
.Y(n_341)
);

INVxp33_ASAP7_75t_SL g342 ( 
.A(n_176),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_227),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_234),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_236),
.Y(n_345)
);

CKINVDCx16_ASAP7_75t_R g346 ( 
.A(n_216),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_189),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_240),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_248),
.Y(n_349)
);

INVxp67_ASAP7_75t_SL g350 ( 
.A(n_239),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_190),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_226),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_251),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_196),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_266),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_277),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_198),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_280),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_290),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_202),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_302),
.Y(n_361)
);

INVxp67_ASAP7_75t_SL g362 ( 
.A(n_241),
.Y(n_362)
);

INVx2_ASAP7_75t_SL g363 ( 
.A(n_213),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_205),
.Y(n_364)
);

INVxp67_ASAP7_75t_SL g365 ( 
.A(n_241),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_212),
.Y(n_366)
);

CKINVDCx14_ASAP7_75t_R g367 ( 
.A(n_297),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_304),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_159),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_240),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_171),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_214),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_223),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_175),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_300),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_287),
.Y(n_376)
);

CKINVDCx16_ASAP7_75t_R g377 ( 
.A(n_287),
.Y(n_377)
);

HB1xp67_ASAP7_75t_L g378 ( 
.A(n_176),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_300),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_195),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_199),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_224),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_200),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_178),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_203),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_233),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_211),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_215),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_220),
.Y(n_389)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_336),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_330),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_330),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_314),
.Y(n_393)
);

INVx4_ASAP7_75t_L g394 ( 
.A(n_336),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_314),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_336),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_362),
.B(n_257),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_335),
.B(n_174),
.Y(n_398)
);

AND2x4_ASAP7_75t_L g399 ( 
.A(n_369),
.B(n_174),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_316),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_316),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_317),
.Y(n_402)
);

AND2x4_ASAP7_75t_L g403 ( 
.A(n_371),
.B(n_210),
.Y(n_403)
);

INVx5_ASAP7_75t_L g404 ( 
.A(n_336),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_317),
.Y(n_405)
);

AND2x4_ASAP7_75t_L g406 ( 
.A(n_374),
.B(n_380),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_SL g407 ( 
.A(n_329),
.B(n_218),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_322),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_322),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_336),
.Y(n_410)
);

INVx2_ASAP7_75t_SL g411 ( 
.A(n_315),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_352),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_352),
.Y(n_413)
);

NAND2xp33_ASAP7_75t_L g414 ( 
.A(n_326),
.B(n_305),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_350),
.B(n_210),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_323),
.B(n_327),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_331),
.Y(n_417)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_352),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_352),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_331),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_381),
.B(n_217),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_352),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_333),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_383),
.B(n_217),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_333),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g426 ( 
.A(n_334),
.Y(n_426)
);

AND2x4_ASAP7_75t_L g427 ( 
.A(n_385),
.B(n_167),
.Y(n_427)
);

AND2x6_ASAP7_75t_L g428 ( 
.A(n_387),
.B(n_226),
.Y(n_428)
);

BUFx8_ASAP7_75t_L g429 ( 
.A(n_318),
.Y(n_429)
);

INVx5_ASAP7_75t_L g430 ( 
.A(n_363),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_339),
.Y(n_431)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_339),
.Y(n_432)
);

BUFx3_ASAP7_75t_L g433 ( 
.A(n_388),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_375),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_319),
.Y(n_435)
);

AND2x4_ASAP7_75t_L g436 ( 
.A(n_389),
.B(n_167),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_375),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_379),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_329),
.A2(n_232),
.B1(n_312),
.B2(n_218),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_379),
.Y(n_440)
);

HB1xp67_ASAP7_75t_L g441 ( 
.A(n_378),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_338),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_340),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_343),
.Y(n_444)
);

AND2x6_ASAP7_75t_L g445 ( 
.A(n_320),
.B(n_226),
.Y(n_445)
);

INVx3_ASAP7_75t_L g446 ( 
.A(n_363),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_344),
.Y(n_447)
);

INVxp67_ASAP7_75t_L g448 ( 
.A(n_325),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_345),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_353),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_355),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_356),
.Y(n_452)
);

NAND2xp33_ASAP7_75t_SL g453 ( 
.A(n_324),
.B(n_257),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_365),
.B(n_297),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_358),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_337),
.B(n_297),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_321),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_359),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_393),
.Y(n_459)
);

BUFx6f_ASAP7_75t_SL g460 ( 
.A(n_406),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_435),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_393),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_397),
.B(n_367),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_442),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_397),
.B(n_326),
.Y(n_465)
);

AND2x4_ASAP7_75t_L g466 ( 
.A(n_399),
.B(n_361),
.Y(n_466)
);

BUFx2_ASAP7_75t_L g467 ( 
.A(n_448),
.Y(n_467)
);

BUFx6f_ASAP7_75t_L g468 ( 
.A(n_396),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_442),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_396),
.Y(n_470)
);

INVx2_ASAP7_75t_SL g471 ( 
.A(n_454),
.Y(n_471)
);

INVx3_ASAP7_75t_L g472 ( 
.A(n_396),
.Y(n_472)
);

OR2x6_ASAP7_75t_L g473 ( 
.A(n_454),
.B(n_349),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_443),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_393),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_398),
.B(n_226),
.Y(n_476)
);

INVx4_ASAP7_75t_L g477 ( 
.A(n_396),
.Y(n_477)
);

INVx1_ASAP7_75t_SL g478 ( 
.A(n_457),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_429),
.Y(n_479)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_396),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_443),
.Y(n_481)
);

INVx2_ASAP7_75t_SL g482 ( 
.A(n_456),
.Y(n_482)
);

BUFx10_ASAP7_75t_L g483 ( 
.A(n_416),
.Y(n_483)
);

AND3x1_ASAP7_75t_L g484 ( 
.A(n_407),
.B(n_368),
.C(n_342),
.Y(n_484)
);

INVx4_ASAP7_75t_L g485 ( 
.A(n_396),
.Y(n_485)
);

OR2x2_ASAP7_75t_L g486 ( 
.A(n_426),
.B(n_346),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_395),
.Y(n_487)
);

AOI22x1_ASAP7_75t_L g488 ( 
.A1(n_399),
.A2(n_386),
.B1(n_382),
.B2(n_373),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_444),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_415),
.B(n_256),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_444),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_395),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_395),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_414),
.B(n_342),
.Y(n_494)
);

INVx1_ASAP7_75t_SL g495 ( 
.A(n_426),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_453),
.B(n_328),
.Y(n_496)
);

NAND2xp33_ASAP7_75t_R g497 ( 
.A(n_456),
.B(n_324),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_448),
.B(n_328),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_400),
.Y(n_499)
);

BUFx2_ASAP7_75t_L g500 ( 
.A(n_441),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_400),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_441),
.B(n_347),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_447),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_406),
.B(n_256),
.Y(n_504)
);

NOR3xp33_ASAP7_75t_L g505 ( 
.A(n_439),
.B(n_377),
.C(n_351),
.Y(n_505)
);

INVx3_ASAP7_75t_L g506 ( 
.A(n_413),
.Y(n_506)
);

INVx3_ASAP7_75t_L g507 ( 
.A(n_413),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_400),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_409),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_447),
.Y(n_510)
);

AOI22xp33_ASAP7_75t_L g511 ( 
.A1(n_427),
.A2(n_256),
.B1(n_272),
.B2(n_221),
.Y(n_511)
);

INVx4_ASAP7_75t_L g512 ( 
.A(n_413),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_409),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_449),
.Y(n_514)
);

AOI22xp33_ASAP7_75t_L g515 ( 
.A1(n_427),
.A2(n_256),
.B1(n_272),
.B2(n_229),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_409),
.Y(n_516)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_413),
.Y(n_517)
);

BUFx6f_ASAP7_75t_SL g518 ( 
.A(n_406),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_449),
.Y(n_519)
);

OAI22xp33_ASAP7_75t_SL g520 ( 
.A1(n_407),
.A2(n_386),
.B1(n_382),
.B2(n_373),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_451),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_433),
.B(n_347),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_433),
.B(n_351),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_L g524 ( 
.A1(n_406),
.A2(n_354),
.B1(n_372),
.B2(n_366),
.Y(n_524)
);

OR2x2_ASAP7_75t_L g525 ( 
.A(n_411),
.B(n_354),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_451),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_452),
.Y(n_527)
);

BUFx4f_ASAP7_75t_L g528 ( 
.A(n_450),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_452),
.Y(n_529)
);

INVx2_ASAP7_75t_SL g530 ( 
.A(n_399),
.Y(n_530)
);

INVx4_ASAP7_75t_L g531 ( 
.A(n_413),
.Y(n_531)
);

BUFx6f_ASAP7_75t_SL g532 ( 
.A(n_399),
.Y(n_532)
);

INVx2_ASAP7_75t_SL g533 ( 
.A(n_403),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_430),
.B(n_357),
.Y(n_534)
);

AOI21x1_ASAP7_75t_L g535 ( 
.A1(n_391),
.A2(n_259),
.B(n_243),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_401),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_401),
.Y(n_537)
);

INVx2_ASAP7_75t_SL g538 ( 
.A(n_403),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_433),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_402),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_402),
.Y(n_541)
);

INVx3_ASAP7_75t_L g542 ( 
.A(n_413),
.Y(n_542)
);

OAI21xp5_ASAP7_75t_L g543 ( 
.A1(n_421),
.A2(n_263),
.B(n_260),
.Y(n_543)
);

INVx3_ASAP7_75t_L g544 ( 
.A(n_394),
.Y(n_544)
);

INVx2_ASAP7_75t_SL g545 ( 
.A(n_403),
.Y(n_545)
);

OR2x2_ASAP7_75t_L g546 ( 
.A(n_411),
.B(n_357),
.Y(n_546)
);

INVx4_ASAP7_75t_L g547 ( 
.A(n_394),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_405),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_405),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_403),
.B(n_256),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_450),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_408),
.Y(n_552)
);

INVx2_ASAP7_75t_SL g553 ( 
.A(n_427),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_430),
.B(n_360),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_408),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_391),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_392),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_450),
.Y(n_558)
);

INVx3_ASAP7_75t_L g559 ( 
.A(n_394),
.Y(n_559)
);

BUFx4f_ASAP7_75t_L g560 ( 
.A(n_450),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_392),
.Y(n_561)
);

BUFx3_ASAP7_75t_L g562 ( 
.A(n_430),
.Y(n_562)
);

INVx3_ASAP7_75t_L g563 ( 
.A(n_394),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_450),
.Y(n_564)
);

AND2x4_ASAP7_75t_L g565 ( 
.A(n_411),
.B(n_265),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_450),
.Y(n_566)
);

BUFx6f_ASAP7_75t_L g567 ( 
.A(n_458),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_429),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_458),
.Y(n_569)
);

BUFx8_ASAP7_75t_SL g570 ( 
.A(n_439),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_458),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_432),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_432),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_432),
.Y(n_574)
);

XNOR2xp5_ASAP7_75t_L g575 ( 
.A(n_427),
.B(n_332),
.Y(n_575)
);

INVxp67_ASAP7_75t_SL g576 ( 
.A(n_390),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_458),
.B(n_272),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_432),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_458),
.Y(n_579)
);

INVx3_ASAP7_75t_L g580 ( 
.A(n_390),
.Y(n_580)
);

INVxp67_ASAP7_75t_L g581 ( 
.A(n_421),
.Y(n_581)
);

INVxp33_ASAP7_75t_L g582 ( 
.A(n_424),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_430),
.B(n_360),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_390),
.Y(n_584)
);

BUFx3_ASAP7_75t_L g585 ( 
.A(n_430),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_446),
.B(n_364),
.Y(n_586)
);

NAND3xp33_ASAP7_75t_L g587 ( 
.A(n_424),
.B(n_364),
.C(n_372),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_458),
.Y(n_588)
);

AND2x4_ASAP7_75t_L g589 ( 
.A(n_436),
.B(n_278),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_390),
.Y(n_590)
);

AOI22xp33_ASAP7_75t_SL g591 ( 
.A1(n_429),
.A2(n_232),
.B1(n_312),
.B2(n_370),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_423),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_455),
.Y(n_593)
);

INVx6_ASAP7_75t_L g594 ( 
.A(n_430),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_423),
.Y(n_595)
);

OR2x6_ASAP7_75t_L g596 ( 
.A(n_436),
.B(n_279),
.Y(n_596)
);

HB1xp67_ASAP7_75t_L g597 ( 
.A(n_446),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_436),
.B(n_272),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_455),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_455),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_417),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_430),
.B(n_366),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_418),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_423),
.Y(n_604)
);

OAI22xp5_ASAP7_75t_L g605 ( 
.A1(n_436),
.A2(n_286),
.B1(n_261),
.B2(n_253),
.Y(n_605)
);

AOI22xp33_ASAP7_75t_L g606 ( 
.A1(n_417),
.A2(n_272),
.B1(n_294),
.B2(n_284),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_425),
.Y(n_607)
);

INVx2_ASAP7_75t_SL g608 ( 
.A(n_446),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_582),
.B(n_446),
.Y(n_609)
);

BUFx6f_ASAP7_75t_L g610 ( 
.A(n_553),
.Y(n_610)
);

AND2x4_ASAP7_75t_L g611 ( 
.A(n_539),
.B(n_420),
.Y(n_611)
);

AND2x4_ASAP7_75t_L g612 ( 
.A(n_464),
.B(n_420),
.Y(n_612)
);

INVx4_ASAP7_75t_L g613 ( 
.A(n_566),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_582),
.B(n_341),
.Y(n_614)
);

INVx1_ASAP7_75t_SL g615 ( 
.A(n_495),
.Y(n_615)
);

INVxp67_ASAP7_75t_L g616 ( 
.A(n_467),
.Y(n_616)
);

INVx4_ASAP7_75t_SL g617 ( 
.A(n_460),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_469),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_474),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_481),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_459),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_489),
.Y(n_622)
);

OR2x6_ASAP7_75t_L g623 ( 
.A(n_500),
.B(n_308),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_581),
.B(n_418),
.Y(n_624)
);

AND2x4_ASAP7_75t_L g625 ( 
.A(n_491),
.B(n_425),
.Y(n_625)
);

NAND2x1p5_ASAP7_75t_L g626 ( 
.A(n_553),
.B(n_238),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_459),
.Y(n_627)
);

OR2x2_ASAP7_75t_L g628 ( 
.A(n_486),
.B(n_293),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_503),
.Y(n_629)
);

INVx3_ASAP7_75t_L g630 ( 
.A(n_580),
.Y(n_630)
);

INVxp67_ASAP7_75t_SL g631 ( 
.A(n_544),
.Y(n_631)
);

INVx3_ASAP7_75t_L g632 ( 
.A(n_580),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_462),
.Y(n_633)
);

BUFx6f_ASAP7_75t_L g634 ( 
.A(n_590),
.Y(n_634)
);

BUFx3_ASAP7_75t_L g635 ( 
.A(n_461),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_471),
.B(n_418),
.Y(n_636)
);

AO22x2_ASAP7_75t_L g637 ( 
.A1(n_505),
.A2(n_306),
.B1(n_12),
.B2(n_13),
.Y(n_637)
);

AND2x4_ASAP7_75t_L g638 ( 
.A(n_510),
.B(n_425),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_514),
.Y(n_639)
);

AND2x4_ASAP7_75t_L g640 ( 
.A(n_519),
.B(n_431),
.Y(n_640)
);

HB1xp67_ASAP7_75t_L g641 ( 
.A(n_471),
.Y(n_641)
);

BUFx10_ASAP7_75t_L g642 ( 
.A(n_498),
.Y(n_642)
);

AND2x4_ASAP7_75t_L g643 ( 
.A(n_521),
.B(n_526),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_527),
.Y(n_644)
);

INVx2_ASAP7_75t_SL g645 ( 
.A(n_586),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_572),
.B(n_418),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_586),
.B(n_348),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_462),
.Y(n_648)
);

NAND3xp33_ASAP7_75t_L g649 ( 
.A(n_543),
.B(n_177),
.C(n_173),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_529),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_601),
.Y(n_651)
);

HB1xp67_ASAP7_75t_L g652 ( 
.A(n_473),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_482),
.B(n_376),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_597),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_556),
.Y(n_655)
);

BUFx6f_ASAP7_75t_L g656 ( 
.A(n_590),
.Y(n_656)
);

AND2x4_ASAP7_75t_L g657 ( 
.A(n_530),
.B(n_431),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_556),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_557),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_465),
.B(n_525),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_557),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_475),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_561),
.Y(n_663)
);

AOI22xp5_ASAP7_75t_L g664 ( 
.A1(n_482),
.A2(n_179),
.B1(n_270),
.B2(n_269),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_572),
.B(n_410),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_561),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_573),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_530),
.B(n_262),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_533),
.B(n_262),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_573),
.Y(n_670)
);

NAND2x1p5_ASAP7_75t_L g671 ( 
.A(n_533),
.B(n_431),
.Y(n_671)
);

INVxp67_ASAP7_75t_SL g672 ( 
.A(n_544),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_574),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_574),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_475),
.Y(n_675)
);

BUFx3_ASAP7_75t_L g676 ( 
.A(n_461),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_479),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_578),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_487),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_502),
.B(n_384),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_578),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_487),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_536),
.Y(n_683)
);

OR2x2_ASAP7_75t_L g684 ( 
.A(n_486),
.B(n_525),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_538),
.B(n_410),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_536),
.Y(n_686)
);

INVxp67_ASAP7_75t_L g687 ( 
.A(n_463),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_546),
.B(n_168),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_492),
.Y(n_689)
);

BUFx6f_ASAP7_75t_L g690 ( 
.A(n_590),
.Y(n_690)
);

HAxp5_ASAP7_75t_SL g691 ( 
.A(n_570),
.B(n_222),
.CON(n_691),
.SN(n_691)
);

BUFx3_ASAP7_75t_L g692 ( 
.A(n_608),
.Y(n_692)
);

NAND2x1p5_ASAP7_75t_L g693 ( 
.A(n_538),
.B(n_434),
.Y(n_693)
);

BUFx3_ASAP7_75t_L g694 ( 
.A(n_466),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_537),
.Y(n_695)
);

AOI22xp5_ASAP7_75t_L g696 ( 
.A1(n_545),
.A2(n_209),
.B1(n_208),
.B2(n_313),
.Y(n_696)
);

INVx4_ASAP7_75t_L g697 ( 
.A(n_566),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_537),
.Y(n_698)
);

AOI22xp5_ASAP7_75t_L g699 ( 
.A1(n_545),
.A2(n_494),
.B1(n_484),
.B2(n_496),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_593),
.B(n_410),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_540),
.Y(n_701)
);

AND2x4_ASAP7_75t_L g702 ( 
.A(n_608),
.B(n_434),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_492),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_599),
.B(n_412),
.Y(n_704)
);

AND2x4_ASAP7_75t_L g705 ( 
.A(n_466),
.B(n_434),
.Y(n_705)
);

OAI22xp5_ASAP7_75t_L g706 ( 
.A1(n_473),
.A2(n_305),
.B1(n_307),
.B2(n_237),
.Y(n_706)
);

CKINVDCx14_ASAP7_75t_R g707 ( 
.A(n_479),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_493),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_540),
.Y(n_709)
);

NAND2x1p5_ASAP7_75t_L g710 ( 
.A(n_547),
.B(n_437),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_493),
.Y(n_711)
);

BUFx2_ASAP7_75t_L g712 ( 
.A(n_575),
.Y(n_712)
);

BUFx6f_ASAP7_75t_L g713 ( 
.A(n_590),
.Y(n_713)
);

BUFx3_ASAP7_75t_L g714 ( 
.A(n_466),
.Y(n_714)
);

OR2x2_ASAP7_75t_SL g715 ( 
.A(n_587),
.B(n_429),
.Y(n_715)
);

HB1xp67_ASAP7_75t_L g716 ( 
.A(n_473),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_499),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_473),
.B(n_437),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_522),
.B(n_437),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_568),
.Y(n_720)
);

INVxp67_ASAP7_75t_L g721 ( 
.A(n_523),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_499),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_541),
.Y(n_723)
);

AO22x2_ASAP7_75t_L g724 ( 
.A1(n_476),
.A2(n_4),
.B1(n_15),
.B2(n_16),
.Y(n_724)
);

OAI21xp33_ASAP7_75t_SL g725 ( 
.A1(n_476),
.A2(n_490),
.B(n_511),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_501),
.Y(n_726)
);

NAND3xp33_ASAP7_75t_SL g727 ( 
.A(n_524),
.B(n_303),
.C(n_177),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_541),
.Y(n_728)
);

INVx4_ASAP7_75t_L g729 ( 
.A(n_566),
.Y(n_729)
);

NAND2x1p5_ASAP7_75t_L g730 ( 
.A(n_547),
.B(n_438),
.Y(n_730)
);

INVxp67_ASAP7_75t_L g731 ( 
.A(n_546),
.Y(n_731)
);

INVx3_ASAP7_75t_R g732 ( 
.A(n_565),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_501),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_508),
.Y(n_734)
);

NOR2x1p5_ASAP7_75t_L g735 ( 
.A(n_568),
.B(n_307),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_483),
.B(n_262),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_548),
.Y(n_737)
);

INVx3_ASAP7_75t_L g738 ( 
.A(n_580),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_508),
.Y(n_739)
);

BUFx6f_ASAP7_75t_L g740 ( 
.A(n_589),
.Y(n_740)
);

XOR2x2_ASAP7_75t_L g741 ( 
.A(n_520),
.B(n_4),
.Y(n_741)
);

INVx3_ASAP7_75t_L g742 ( 
.A(n_584),
.Y(n_742)
);

CKINVDCx20_ASAP7_75t_R g743 ( 
.A(n_570),
.Y(n_743)
);

OAI221xp5_ASAP7_75t_L g744 ( 
.A1(n_490),
.A2(n_438),
.B1(n_440),
.B2(n_245),
.C(n_244),
.Y(n_744)
);

NAND2x1p5_ASAP7_75t_L g745 ( 
.A(n_547),
.B(n_544),
.Y(n_745)
);

AND2x6_ASAP7_75t_L g746 ( 
.A(n_589),
.B(n_412),
.Y(n_746)
);

BUFx3_ASAP7_75t_L g747 ( 
.A(n_565),
.Y(n_747)
);

HB1xp67_ASAP7_75t_L g748 ( 
.A(n_596),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_509),
.Y(n_749)
);

INVx3_ASAP7_75t_L g750 ( 
.A(n_584),
.Y(n_750)
);

HB1xp67_ASAP7_75t_L g751 ( 
.A(n_596),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_548),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_549),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_483),
.B(n_438),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_549),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_509),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_552),
.Y(n_757)
);

AND3x4_ASAP7_75t_L g758 ( 
.A(n_591),
.B(n_440),
.C(n_291),
.Y(n_758)
);

AO22x2_ASAP7_75t_L g759 ( 
.A1(n_550),
.A2(n_15),
.B1(n_17),
.B2(n_18),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_552),
.Y(n_760)
);

AOI22xp5_ASAP7_75t_L g761 ( 
.A1(n_532),
.A2(n_201),
.B1(n_309),
.B2(n_228),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_555),
.Y(n_762)
);

BUFx2_ASAP7_75t_L g763 ( 
.A(n_478),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_513),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_555),
.Y(n_765)
);

AND2x4_ASAP7_75t_L g766 ( 
.A(n_589),
.B(n_440),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_513),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_600),
.Y(n_768)
);

AND2x4_ASAP7_75t_L g769 ( 
.A(n_596),
.B(n_168),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_483),
.B(n_605),
.Y(n_770)
);

OAI22xp5_ASAP7_75t_SL g771 ( 
.A1(n_596),
.A2(n_273),
.B1(n_310),
.B2(n_296),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_516),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_592),
.Y(n_773)
);

AOI22xp5_ASAP7_75t_L g774 ( 
.A1(n_532),
.A2(n_192),
.B1(n_207),
.B2(n_301),
.Y(n_774)
);

AO22x2_ASAP7_75t_L g775 ( 
.A1(n_550),
.A2(n_20),
.B1(n_21),
.B2(n_23),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_584),
.B(n_262),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_592),
.Y(n_777)
);

AO22x2_ASAP7_75t_L g778 ( 
.A1(n_504),
.A2(n_20),
.B1(n_23),
.B2(n_24),
.Y(n_778)
);

AND2x4_ASAP7_75t_L g779 ( 
.A(n_565),
.B(n_172),
.Y(n_779)
);

AND2x2_ASAP7_75t_L g780 ( 
.A(n_504),
.B(n_281),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_516),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_631),
.B(n_595),
.Y(n_782)
);

NOR2x1_ASAP7_75t_L g783 ( 
.A(n_660),
.B(n_534),
.Y(n_783)
);

BUFx2_ASAP7_75t_L g784 ( 
.A(n_615),
.Y(n_784)
);

INVx2_ASAP7_75t_SL g785 ( 
.A(n_615),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_719),
.B(n_576),
.Y(n_786)
);

HB1xp67_ASAP7_75t_L g787 ( 
.A(n_616),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_657),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_657),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_635),
.Y(n_790)
);

AOI22xp5_ASAP7_75t_L g791 ( 
.A1(n_660),
.A2(n_758),
.B1(n_645),
.B2(n_724),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_702),
.Y(n_792)
);

NAND2x1p5_ASAP7_75t_L g793 ( 
.A(n_610),
.B(n_559),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_631),
.B(n_595),
.Y(n_794)
);

AND2x6_ASAP7_75t_L g795 ( 
.A(n_754),
.B(n_559),
.Y(n_795)
);

INVx3_ASAP7_75t_L g796 ( 
.A(n_610),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_721),
.B(n_532),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_672),
.B(n_721),
.Y(n_798)
);

BUFx6f_ASAP7_75t_L g799 ( 
.A(n_740),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_702),
.Y(n_800)
);

OR2x2_ASAP7_75t_L g801 ( 
.A(n_684),
.B(n_598),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_676),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_705),
.Y(n_803)
);

NOR2x1_ASAP7_75t_L g804 ( 
.A(n_727),
.B(n_554),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_705),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_L g806 ( 
.A(n_687),
.B(n_460),
.Y(n_806)
);

OAI22xp33_ASAP7_75t_L g807 ( 
.A1(n_699),
.A2(n_497),
.B1(n_488),
.B2(n_602),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_655),
.Y(n_808)
);

INVxp67_ASAP7_75t_L g809 ( 
.A(n_614),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_658),
.Y(n_810)
);

CKINVDCx20_ASAP7_75t_R g811 ( 
.A(n_763),
.Y(n_811)
);

BUFx3_ASAP7_75t_L g812 ( 
.A(n_653),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_L g813 ( 
.A(n_687),
.B(n_460),
.Y(n_813)
);

AOI22xp33_ASAP7_75t_L g814 ( 
.A1(n_649),
.A2(n_518),
.B1(n_598),
.B2(n_606),
.Y(n_814)
);

BUFx2_ASAP7_75t_L g815 ( 
.A(n_616),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_659),
.Y(n_816)
);

O2A1O1Ixp5_ASAP7_75t_L g817 ( 
.A1(n_736),
.A2(n_583),
.B(n_577),
.C(n_535),
.Y(n_817)
);

A2O1A1Ixp33_ASAP7_75t_L g818 ( 
.A1(n_688),
.A2(n_603),
.B(n_515),
.C(n_558),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_672),
.B(n_559),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_610),
.B(n_563),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_661),
.Y(n_821)
);

AOI22xp5_ASAP7_75t_L g822 ( 
.A1(n_758),
.A2(n_607),
.B1(n_604),
.B2(n_518),
.Y(n_822)
);

HB1xp67_ASAP7_75t_L g823 ( 
.A(n_641),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_663),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_747),
.B(n_740),
.Y(n_825)
);

OR2x2_ASAP7_75t_L g826 ( 
.A(n_628),
.B(n_283),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_667),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_609),
.B(n_563),
.Y(n_828)
);

INVx4_ASAP7_75t_L g829 ( 
.A(n_740),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_666),
.Y(n_830)
);

AOI22xp5_ASAP7_75t_L g831 ( 
.A1(n_724),
.A2(n_607),
.B1(n_604),
.B2(n_518),
.Y(n_831)
);

INVx2_ASAP7_75t_SL g832 ( 
.A(n_647),
.Y(n_832)
);

BUFx3_ASAP7_75t_L g833 ( 
.A(n_654),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_692),
.B(n_563),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_692),
.B(n_603),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_714),
.B(n_528),
.Y(n_836)
);

INVx4_ASAP7_75t_L g837 ( 
.A(n_714),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_624),
.B(n_603),
.Y(n_838)
);

AND2x4_ASAP7_75t_L g839 ( 
.A(n_617),
.B(n_694),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_683),
.Y(n_840)
);

INVxp67_ASAP7_75t_SL g841 ( 
.A(n_745),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_731),
.B(n_528),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_624),
.B(n_472),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_731),
.B(n_528),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_686),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_688),
.B(n_472),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_670),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_641),
.B(n_560),
.Y(n_848)
);

AOI22xp5_ASAP7_75t_L g849 ( 
.A1(n_724),
.A2(n_649),
.B1(n_778),
.B2(n_775),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_651),
.B(n_472),
.Y(n_850)
);

AOI22xp33_ASAP7_75t_L g851 ( 
.A1(n_727),
.A2(n_564),
.B1(n_588),
.B2(n_551),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_618),
.B(n_480),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_619),
.B(n_620),
.Y(n_853)
);

AOI22xp33_ASAP7_75t_SL g854 ( 
.A1(n_770),
.A2(n_262),
.B1(n_173),
.B2(n_172),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_695),
.Y(n_855)
);

INVx4_ASAP7_75t_L g856 ( 
.A(n_617),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_R g857 ( 
.A(n_707),
.B(n_303),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_SL g858 ( 
.A(n_642),
.B(n_560),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_698),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_701),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_709),
.Y(n_861)
);

AND2x4_ASAP7_75t_L g862 ( 
.A(n_617),
.B(n_569),
.Y(n_862)
);

AOI22xp33_ASAP7_75t_L g863 ( 
.A1(n_744),
.A2(n_579),
.B1(n_571),
.B2(n_262),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_707),
.Y(n_864)
);

AOI22xp33_ASAP7_75t_L g865 ( 
.A1(n_744),
.A2(n_262),
.B1(n_577),
.B2(n_566),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_622),
.B(n_480),
.Y(n_866)
);

INVx2_ASAP7_75t_SL g867 ( 
.A(n_623),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_723),
.Y(n_868)
);

INVx4_ASAP7_75t_L g869 ( 
.A(n_634),
.Y(n_869)
);

NAND2x1p5_ASAP7_75t_L g870 ( 
.A(n_766),
.B(n_567),
.Y(n_870)
);

A2O1A1Ixp33_ASAP7_75t_L g871 ( 
.A1(n_725),
.A2(n_560),
.B(n_506),
.C(n_507),
.Y(n_871)
);

BUFx2_ASAP7_75t_L g872 ( 
.A(n_652),
.Y(n_872)
);

BUFx6f_ASAP7_75t_L g873 ( 
.A(n_746),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_728),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_630),
.B(n_480),
.Y(n_875)
);

HB1xp67_ASAP7_75t_L g876 ( 
.A(n_718),
.Y(n_876)
);

AND2x4_ASAP7_75t_L g877 ( 
.A(n_643),
.B(n_506),
.Y(n_877)
);

INVx5_ASAP7_75t_L g878 ( 
.A(n_746),
.Y(n_878)
);

OR2x6_ASAP7_75t_L g879 ( 
.A(n_652),
.B(n_716),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_673),
.Y(n_880)
);

CKINVDCx8_ASAP7_75t_R g881 ( 
.A(n_677),
.Y(n_881)
);

INVx3_ASAP7_75t_L g882 ( 
.A(n_630),
.Y(n_882)
);

AND2x4_ASAP7_75t_L g883 ( 
.A(n_643),
.B(n_506),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_737),
.Y(n_884)
);

BUFx3_ASAP7_75t_L g885 ( 
.A(n_712),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_SL g886 ( 
.A(n_642),
.B(n_567),
.Y(n_886)
);

BUFx6f_ASAP7_75t_L g887 ( 
.A(n_746),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_752),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_680),
.B(n_477),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_779),
.B(n_780),
.Y(n_890)
);

AND2x6_ASAP7_75t_L g891 ( 
.A(n_632),
.B(n_507),
.Y(n_891)
);

NAND3xp33_ASAP7_75t_SL g892 ( 
.A(n_677),
.B(n_235),
.C(n_252),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_753),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_632),
.B(n_738),
.Y(n_894)
);

BUFx6f_ASAP7_75t_L g895 ( 
.A(n_746),
.Y(n_895)
);

BUFx6f_ASAP7_75t_L g896 ( 
.A(n_746),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_674),
.Y(n_897)
);

BUFx2_ASAP7_75t_L g898 ( 
.A(n_716),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_779),
.B(n_162),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_678),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_755),
.Y(n_901)
);

BUFx2_ASAP7_75t_L g902 ( 
.A(n_623),
.Y(n_902)
);

BUFx3_ASAP7_75t_L g903 ( 
.A(n_720),
.Y(n_903)
);

AND2x4_ASAP7_75t_L g904 ( 
.A(n_612),
.B(n_507),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_681),
.Y(n_905)
);

AOI22xp33_ASAP7_75t_L g906 ( 
.A1(n_766),
.A2(n_567),
.B1(n_517),
.B2(n_542),
.Y(n_906)
);

INVx5_ASAP7_75t_L g907 ( 
.A(n_623),
.Y(n_907)
);

INVx3_ASAP7_75t_L g908 ( 
.A(n_738),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_742),
.B(n_750),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_742),
.Y(n_910)
);

AOI22xp33_ASAP7_75t_L g911 ( 
.A1(n_625),
.A2(n_567),
.B1(n_517),
.B2(n_542),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_750),
.B(n_517),
.Y(n_912)
);

AOI22x1_ASAP7_75t_L g913 ( 
.A1(n_629),
.A2(n_542),
.B1(n_477),
.B2(n_485),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_611),
.Y(n_914)
);

AOI22xp33_ASAP7_75t_L g915 ( 
.A1(n_625),
.A2(n_428),
.B1(n_445),
.B2(n_164),
.Y(n_915)
);

AO21x1_ASAP7_75t_L g916 ( 
.A1(n_736),
.A2(n_669),
.B(n_668),
.Y(n_916)
);

AOI22xp33_ASAP7_75t_L g917 ( 
.A1(n_638),
.A2(n_428),
.B1(n_445),
.B2(n_165),
.Y(n_917)
);

BUFx6f_ASAP7_75t_L g918 ( 
.A(n_634),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_757),
.Y(n_919)
);

BUFx3_ASAP7_75t_L g920 ( 
.A(n_720),
.Y(n_920)
);

OAI22xp5_ASAP7_75t_L g921 ( 
.A1(n_778),
.A2(n_231),
.B1(n_254),
.B2(n_249),
.Y(n_921)
);

BUFx6f_ASAP7_75t_L g922 ( 
.A(n_634),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_639),
.B(n_477),
.Y(n_923)
);

INVx5_ASAP7_75t_L g924 ( 
.A(n_656),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_R g925 ( 
.A(n_743),
.B(n_163),
.Y(n_925)
);

AOI22xp33_ASAP7_75t_L g926 ( 
.A1(n_638),
.A2(n_428),
.B1(n_445),
.B2(n_275),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_611),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_745),
.A2(n_485),
.B(n_531),
.Y(n_928)
);

BUFx4f_ASAP7_75t_L g929 ( 
.A(n_626),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_644),
.B(n_485),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_760),
.Y(n_931)
);

BUFx3_ASAP7_75t_L g932 ( 
.A(n_743),
.Y(n_932)
);

INVx3_ASAP7_75t_L g933 ( 
.A(n_656),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_650),
.B(n_762),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_765),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_626),
.B(n_180),
.Y(n_936)
);

INVx4_ASAP7_75t_L g937 ( 
.A(n_656),
.Y(n_937)
);

AOI22xp5_ASAP7_75t_L g938 ( 
.A1(n_778),
.A2(n_219),
.B1(n_246),
.B2(n_242),
.Y(n_938)
);

INVx3_ASAP7_75t_L g939 ( 
.A(n_690),
.Y(n_939)
);

HB1xp67_ASAP7_75t_L g940 ( 
.A(n_748),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_732),
.B(n_748),
.Y(n_941)
);

BUFx3_ASAP7_75t_L g942 ( 
.A(n_715),
.Y(n_942)
);

INVx3_ASAP7_75t_L g943 ( 
.A(n_690),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_612),
.Y(n_944)
);

OAI22xp5_ASAP7_75t_L g945 ( 
.A1(n_759),
.A2(n_194),
.B1(n_206),
.B2(n_193),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_640),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_621),
.Y(n_947)
);

AOI22xp5_ASAP7_75t_L g948 ( 
.A1(n_759),
.A2(n_230),
.B1(n_255),
.B2(n_191),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_636),
.B(n_531),
.Y(n_949)
);

BUFx3_ASAP7_75t_L g950 ( 
.A(n_769),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_627),
.Y(n_951)
);

OR2x6_ASAP7_75t_L g952 ( 
.A(n_751),
.B(n_512),
.Y(n_952)
);

AND2x2_ASAP7_75t_L g953 ( 
.A(n_769),
.B(n_188),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_633),
.Y(n_954)
);

INVx5_ASAP7_75t_L g955 ( 
.A(n_690),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_640),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_768),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_636),
.B(n_531),
.Y(n_958)
);

OR2x2_ASAP7_75t_L g959 ( 
.A(n_706),
.B(n_751),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_664),
.B(n_186),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_773),
.B(n_512),
.Y(n_961)
);

AOI21xp33_ASAP7_75t_L g962 ( 
.A1(n_759),
.A2(n_181),
.B(n_299),
.Y(n_962)
);

AOI22xp5_ASAP7_75t_L g963 ( 
.A1(n_775),
.A2(n_295),
.B1(n_183),
.B2(n_182),
.Y(n_963)
);

A2O1A1Ixp33_ASAP7_75t_L g964 ( 
.A1(n_668),
.A2(n_669),
.B(n_685),
.C(n_777),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_SL g965 ( 
.A(n_696),
.B(n_288),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_771),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_761),
.B(n_292),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_685),
.Y(n_968)
);

INVxp67_ASAP7_75t_L g969 ( 
.A(n_706),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_SL g970 ( 
.A(n_774),
.B(n_285),
.Y(n_970)
);

INVx3_ASAP7_75t_L g971 ( 
.A(n_713),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_665),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_648),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_735),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_968),
.B(n_662),
.Y(n_975)
);

BUFx12f_ASAP7_75t_L g976 ( 
.A(n_790),
.Y(n_976)
);

OR2x6_ASAP7_75t_L g977 ( 
.A(n_856),
.B(n_637),
.Y(n_977)
);

AOI22xp33_ASAP7_75t_L g978 ( 
.A1(n_962),
.A2(n_775),
.B1(n_637),
.B2(n_741),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_789),
.Y(n_979)
);

BUFx4f_ASAP7_75t_L g980 ( 
.A(n_784),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_934),
.Y(n_981)
);

INVx2_ASAP7_75t_SL g982 ( 
.A(n_785),
.Y(n_982)
);

AND2x4_ASAP7_75t_L g983 ( 
.A(n_839),
.B(n_776),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_798),
.B(n_675),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_SL g985 ( 
.A(n_929),
.B(n_671),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_929),
.B(n_671),
.Y(n_986)
);

HB1xp67_ASAP7_75t_L g987 ( 
.A(n_815),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_934),
.Y(n_988)
);

BUFx2_ASAP7_75t_L g989 ( 
.A(n_811),
.Y(n_989)
);

BUFx12f_ASAP7_75t_L g990 ( 
.A(n_802),
.Y(n_990)
);

OR2x2_ASAP7_75t_L g991 ( 
.A(n_826),
.B(n_776),
.Y(n_991)
);

INVx3_ASAP7_75t_L g992 ( 
.A(n_873),
.Y(n_992)
);

AOI22xp33_ASAP7_75t_L g993 ( 
.A1(n_962),
.A2(n_637),
.B1(n_693),
.B2(n_767),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_946),
.Y(n_994)
);

CKINVDCx20_ASAP7_75t_R g995 ( 
.A(n_864),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_798),
.B(n_679),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_972),
.B(n_682),
.Y(n_997)
);

O2A1O1Ixp33_ASAP7_75t_L g998 ( 
.A1(n_809),
.A2(n_700),
.B(n_704),
.C(n_693),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_956),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_786),
.B(n_689),
.Y(n_1000)
);

AOI22xp33_ASAP7_75t_L g1001 ( 
.A1(n_854),
.A2(n_733),
.B1(n_772),
.B2(n_764),
.Y(n_1001)
);

BUFx6f_ASAP7_75t_L g1002 ( 
.A(n_918),
.Y(n_1002)
);

AO22x1_ASAP7_75t_L g1003 ( 
.A1(n_966),
.A2(n_691),
.B1(n_276),
.B2(n_274),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_828),
.B(n_781),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_788),
.Y(n_1005)
);

AOI22xp33_ASAP7_75t_L g1006 ( 
.A1(n_791),
.A2(n_756),
.B1(n_749),
.B2(n_739),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_783),
.B(n_734),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_957),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_782),
.B(n_703),
.Y(n_1009)
);

AOI21xp33_ASAP7_75t_L g1010 ( 
.A1(n_921),
.A2(n_945),
.B(n_849),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_792),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_782),
.B(n_717),
.Y(n_1012)
);

AND2x2_ASAP7_75t_SL g1013 ( 
.A(n_938),
.B(n_948),
.Y(n_1013)
);

HB1xp67_ASAP7_75t_L g1014 ( 
.A(n_823),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_800),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_827),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_808),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_794),
.B(n_708),
.Y(n_1018)
);

CKINVDCx11_ASAP7_75t_R g1019 ( 
.A(n_881),
.Y(n_1019)
);

AND2x2_ASAP7_75t_SL g1020 ( 
.A(n_938),
.B(n_697),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_810),
.Y(n_1021)
);

BUFx8_ASAP7_75t_L g1022 ( 
.A(n_902),
.Y(n_1022)
);

OR2x6_ASAP7_75t_L g1023 ( 
.A(n_856),
.B(n_730),
.Y(n_1023)
);

CKINVDCx20_ASAP7_75t_R g1024 ( 
.A(n_885),
.Y(n_1024)
);

BUFx2_ASAP7_75t_L g1025 ( 
.A(n_787),
.Y(n_1025)
);

CKINVDCx20_ASAP7_75t_R g1026 ( 
.A(n_925),
.Y(n_1026)
);

BUFx2_ASAP7_75t_L g1027 ( 
.A(n_812),
.Y(n_1027)
);

AND2x4_ASAP7_75t_L g1028 ( 
.A(n_839),
.B(n_713),
.Y(n_1028)
);

INVx3_ASAP7_75t_L g1029 ( 
.A(n_873),
.Y(n_1029)
);

INVxp67_ASAP7_75t_L g1030 ( 
.A(n_940),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_847),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_816),
.Y(n_1032)
);

INVx1_ASAP7_75t_SL g1033 ( 
.A(n_890),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_880),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_794),
.B(n_726),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_889),
.B(n_722),
.Y(n_1036)
);

BUFx2_ASAP7_75t_L g1037 ( 
.A(n_872),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_974),
.Y(n_1038)
);

BUFx6f_ASAP7_75t_L g1039 ( 
.A(n_918),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_L g1040 ( 
.A(n_969),
.B(n_729),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_821),
.Y(n_1041)
);

BUFx6f_ASAP7_75t_L g1042 ( 
.A(n_918),
.Y(n_1042)
);

BUFx2_ASAP7_75t_L g1043 ( 
.A(n_898),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_853),
.B(n_876),
.Y(n_1044)
);

INVx4_ASAP7_75t_L g1045 ( 
.A(n_799),
.Y(n_1045)
);

HB1xp67_ASAP7_75t_L g1046 ( 
.A(n_879),
.Y(n_1046)
);

CKINVDCx20_ASAP7_75t_R g1047 ( 
.A(n_932),
.Y(n_1047)
);

NOR2xp33_ASAP7_75t_L g1048 ( 
.A(n_832),
.B(n_959),
.Y(n_1048)
);

INVx3_ASAP7_75t_SL g1049 ( 
.A(n_903),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_819),
.B(n_711),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_824),
.Y(n_1051)
);

AOI22xp33_ASAP7_75t_L g1052 ( 
.A1(n_791),
.A2(n_646),
.B1(n_700),
.B2(n_704),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_795),
.B(n_665),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_920),
.Y(n_1054)
);

BUFx3_ASAP7_75t_L g1055 ( 
.A(n_833),
.Y(n_1055)
);

INVxp67_ASAP7_75t_SL g1056 ( 
.A(n_841),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_795),
.B(n_646),
.Y(n_1057)
);

INVx4_ASAP7_75t_L g1058 ( 
.A(n_799),
.Y(n_1058)
);

NOR2x1_ASAP7_75t_L g1059 ( 
.A(n_829),
.B(n_729),
.Y(n_1059)
);

AND2x2_ASAP7_75t_L g1060 ( 
.A(n_899),
.B(n_282),
.Y(n_1060)
);

BUFx6f_ASAP7_75t_L g1061 ( 
.A(n_922),
.Y(n_1061)
);

A2O1A1Ixp33_ASAP7_75t_L g1062 ( 
.A1(n_849),
.A2(n_258),
.B(n_264),
.C(n_267),
.Y(n_1062)
);

AOI22xp33_ASAP7_75t_L g1063 ( 
.A1(n_921),
.A2(n_945),
.B1(n_948),
.B2(n_963),
.Y(n_1063)
);

AOI221xp5_ASAP7_75t_L g1064 ( 
.A1(n_963),
.A2(n_268),
.B1(n_298),
.B2(n_713),
.C(n_730),
.Y(n_1064)
);

AOI22xp33_ASAP7_75t_L g1065 ( 
.A1(n_803),
.A2(n_710),
.B1(n_697),
.B2(n_613),
.Y(n_1065)
);

BUFx3_ASAP7_75t_L g1066 ( 
.A(n_879),
.Y(n_1066)
);

CKINVDCx14_ASAP7_75t_R g1067 ( 
.A(n_857),
.Y(n_1067)
);

BUFx2_ASAP7_75t_L g1068 ( 
.A(n_879),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_795),
.B(n_710),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_897),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_799),
.B(n_613),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_942),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_795),
.B(n_512),
.Y(n_1073)
);

AND2x4_ASAP7_75t_L g1074 ( 
.A(n_944),
.B(n_468),
.Y(n_1074)
);

AOI22xp33_ASAP7_75t_L g1075 ( 
.A1(n_805),
.A2(n_247),
.B1(n_445),
.B2(n_428),
.Y(n_1075)
);

INVx4_ASAP7_75t_L g1076 ( 
.A(n_924),
.Y(n_1076)
);

BUFx2_ASAP7_75t_L g1077 ( 
.A(n_950),
.Y(n_1077)
);

INVxp67_ASAP7_75t_SL g1078 ( 
.A(n_870),
.Y(n_1078)
);

INVx4_ASAP7_75t_L g1079 ( 
.A(n_924),
.Y(n_1079)
);

BUFx3_ASAP7_75t_L g1080 ( 
.A(n_867),
.Y(n_1080)
);

O2A1O1Ixp33_ASAP7_75t_L g1081 ( 
.A1(n_807),
.A2(n_412),
.B(n_419),
.C(n_422),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_907),
.Y(n_1082)
);

BUFx6f_ASAP7_75t_L g1083 ( 
.A(n_922),
.Y(n_1083)
);

AND2x2_ASAP7_75t_L g1084 ( 
.A(n_914),
.B(n_25),
.Y(n_1084)
);

OAI22xp5_ASAP7_75t_SL g1085 ( 
.A1(n_907),
.A2(n_941),
.B1(n_797),
.B2(n_813),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_900),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_834),
.B(n_470),
.Y(n_1087)
);

NOR2xp33_ASAP7_75t_L g1088 ( 
.A(n_806),
.B(n_470),
.Y(n_1088)
);

BUFx3_ASAP7_75t_L g1089 ( 
.A(n_907),
.Y(n_1089)
);

INVx5_ASAP7_75t_L g1090 ( 
.A(n_873),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_830),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_840),
.Y(n_1092)
);

HB1xp67_ASAP7_75t_L g1093 ( 
.A(n_927),
.Y(n_1093)
);

NOR2xp33_ASAP7_75t_L g1094 ( 
.A(n_801),
.B(n_470),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_834),
.B(n_470),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_882),
.B(n_908),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_L g1097 ( 
.A(n_822),
.B(n_468),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_892),
.Y(n_1098)
);

OAI22xp5_ASAP7_75t_L g1099 ( 
.A1(n_831),
.A2(n_822),
.B1(n_814),
.B2(n_878),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_SL g1100 ( 
.A(n_837),
.B(n_468),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_882),
.B(n_468),
.Y(n_1101)
);

OR2x6_ASAP7_75t_L g1102 ( 
.A(n_952),
.B(n_594),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_L g1103 ( 
.A(n_842),
.B(n_25),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_845),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_908),
.B(n_422),
.Y(n_1105)
);

AND2x4_ASAP7_75t_L g1106 ( 
.A(n_837),
.B(n_131),
.Y(n_1106)
);

OAI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_871),
.A2(n_445),
.B(n_422),
.Y(n_1107)
);

BUFx3_ASAP7_75t_L g1108 ( 
.A(n_862),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_855),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_905),
.Y(n_1110)
);

BUFx12f_ASAP7_75t_L g1111 ( 
.A(n_862),
.Y(n_1111)
);

BUFx3_ASAP7_75t_L g1112 ( 
.A(n_877),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_931),
.Y(n_1113)
);

NOR2xp33_ASAP7_75t_L g1114 ( 
.A(n_844),
.B(n_26),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_859),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_860),
.Y(n_1116)
);

BUFx2_ASAP7_75t_L g1117 ( 
.A(n_953),
.Y(n_1117)
);

AO22x1_ASAP7_75t_L g1118 ( 
.A1(n_804),
.A2(n_445),
.B1(n_428),
.B2(n_35),
.Y(n_1118)
);

O2A1O1Ixp33_ASAP7_75t_L g1119 ( 
.A1(n_936),
.A2(n_858),
.B(n_960),
.C(n_967),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_861),
.Y(n_1120)
);

INVx5_ASAP7_75t_L g1121 ( 
.A(n_887),
.Y(n_1121)
);

AND2x4_ASAP7_75t_L g1122 ( 
.A(n_829),
.B(n_140),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_935),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_868),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_846),
.B(n_838),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_874),
.B(n_419),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_884),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_947),
.Y(n_1128)
);

CKINVDCx11_ASAP7_75t_R g1129 ( 
.A(n_1019),
.Y(n_1129)
);

CKINVDCx11_ASAP7_75t_R g1130 ( 
.A(n_1024),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_1008),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_1017),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_1021),
.Y(n_1133)
);

INVx2_ASAP7_75t_SL g1134 ( 
.A(n_980),
.Y(n_1134)
);

INVx4_ASAP7_75t_L g1135 ( 
.A(n_1076),
.Y(n_1135)
);

INVx2_ASAP7_75t_SL g1136 ( 
.A(n_980),
.Y(n_1136)
);

BUFx4f_ASAP7_75t_SL g1137 ( 
.A(n_976),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_1032),
.Y(n_1138)
);

BUFx12f_ASAP7_75t_L g1139 ( 
.A(n_990),
.Y(n_1139)
);

BUFx3_ASAP7_75t_L g1140 ( 
.A(n_1049),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1041),
.Y(n_1141)
);

INVx2_ASAP7_75t_SL g1142 ( 
.A(n_1055),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_981),
.B(n_888),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1051),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1091),
.Y(n_1145)
);

INVx4_ASAP7_75t_L g1146 ( 
.A(n_1076),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_1092),
.Y(n_1147)
);

A2O1A1Ixp33_ASAP7_75t_L g1148 ( 
.A1(n_1063),
.A2(n_831),
.B(n_817),
.C(n_964),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_988),
.B(n_893),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1104),
.Y(n_1150)
);

BUFx6f_ASAP7_75t_L g1151 ( 
.A(n_1002),
.Y(n_1151)
);

NOR2xp33_ASAP7_75t_L g1152 ( 
.A(n_1033),
.B(n_970),
.Y(n_1152)
);

INVx3_ASAP7_75t_L g1153 ( 
.A(n_1023),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_984),
.B(n_996),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1109),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_1115),
.Y(n_1156)
);

BUFx2_ASAP7_75t_L g1157 ( 
.A(n_987),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1116),
.Y(n_1158)
);

OR2x2_ASAP7_75t_L g1159 ( 
.A(n_1044),
.B(n_901),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_1120),
.Y(n_1160)
);

HB1xp67_ASAP7_75t_L g1161 ( 
.A(n_1014),
.Y(n_1161)
);

INVx3_ASAP7_75t_L g1162 ( 
.A(n_1023),
.Y(n_1162)
);

AOI22xp33_ASAP7_75t_L g1163 ( 
.A1(n_1013),
.A2(n_1010),
.B1(n_978),
.B2(n_1103),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_1124),
.Y(n_1164)
);

OR2x2_ASAP7_75t_L g1165 ( 
.A(n_1033),
.B(n_919),
.Y(n_1165)
);

OAI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1125),
.A2(n_818),
.B(n_949),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_1125),
.A2(n_958),
.B(n_949),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_984),
.B(n_796),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_1127),
.Y(n_1169)
);

NOR2xp67_ASAP7_75t_SL g1170 ( 
.A(n_1054),
.B(n_878),
.Y(n_1170)
);

BUFx4f_ASAP7_75t_L g1171 ( 
.A(n_1111),
.Y(n_1171)
);

NOR2xp33_ASAP7_75t_L g1172 ( 
.A(n_1048),
.B(n_877),
.Y(n_1172)
);

A2O1A1Ixp33_ASAP7_75t_L g1173 ( 
.A1(n_1010),
.A2(n_848),
.B(n_825),
.C(n_965),
.Y(n_1173)
);

INVx1_ASAP7_75t_SL g1174 ( 
.A(n_1025),
.Y(n_1174)
);

A2O1A1Ixp33_ASAP7_75t_L g1175 ( 
.A1(n_1119),
.A2(n_904),
.B(n_883),
.C(n_930),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_1016),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_1038),
.Y(n_1177)
);

CKINVDCx20_ASAP7_75t_R g1178 ( 
.A(n_995),
.Y(n_1178)
);

NOR2xp33_ASAP7_75t_L g1179 ( 
.A(n_1030),
.B(n_883),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_1031),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_994),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_1034),
.Y(n_1182)
);

AND2x4_ASAP7_75t_L g1183 ( 
.A(n_1108),
.B(n_904),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_999),
.Y(n_1184)
);

BUFx3_ASAP7_75t_L g1185 ( 
.A(n_1037),
.Y(n_1185)
);

BUFx6f_ASAP7_75t_L g1186 ( 
.A(n_1002),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1070),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1036),
.A2(n_1056),
.B(n_998),
.Y(n_1188)
);

O2A1O1Ixp33_ASAP7_75t_SL g1189 ( 
.A1(n_1062),
.A2(n_836),
.B(n_886),
.C(n_894),
.Y(n_1189)
);

BUFx6f_ASAP7_75t_L g1190 ( 
.A(n_1002),
.Y(n_1190)
);

BUFx6f_ASAP7_75t_L g1191 ( 
.A(n_1039),
.Y(n_1191)
);

BUFx3_ASAP7_75t_L g1192 ( 
.A(n_1043),
.Y(n_1192)
);

AND2x2_ASAP7_75t_L g1193 ( 
.A(n_1117),
.B(n_951),
.Y(n_1193)
);

O2A1O1Ixp5_ASAP7_75t_L g1194 ( 
.A1(n_1099),
.A2(n_916),
.B(n_958),
.C(n_820),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1086),
.Y(n_1195)
);

OR2x6_ASAP7_75t_L g1196 ( 
.A(n_1023),
.B(n_952),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1110),
.Y(n_1197)
);

BUFx3_ASAP7_75t_L g1198 ( 
.A(n_1027),
.Y(n_1198)
);

AND2x2_ASAP7_75t_L g1199 ( 
.A(n_1060),
.B(n_954),
.Y(n_1199)
);

BUFx2_ASAP7_75t_L g1200 ( 
.A(n_989),
.Y(n_1200)
);

AOI22xp33_ASAP7_75t_L g1201 ( 
.A1(n_1114),
.A2(n_973),
.B1(n_796),
.B2(n_865),
.Y(n_1201)
);

AND2x2_ASAP7_75t_SL g1202 ( 
.A(n_1020),
.B(n_887),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_SL g1203 ( 
.A(n_982),
.B(n_878),
.Y(n_1203)
);

AO21x2_ASAP7_75t_L g1204 ( 
.A1(n_1107),
.A2(n_843),
.B(n_928),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1113),
.Y(n_1205)
);

BUFx16f_ASAP7_75t_R g1206 ( 
.A(n_1022),
.Y(n_1206)
);

BUFx6f_ASAP7_75t_L g1207 ( 
.A(n_1039),
.Y(n_1207)
);

HB1xp67_ASAP7_75t_L g1208 ( 
.A(n_1093),
.Y(n_1208)
);

INVx1_ASAP7_75t_SL g1209 ( 
.A(n_1047),
.Y(n_1209)
);

AND2x4_ASAP7_75t_L g1210 ( 
.A(n_1112),
.B(n_952),
.Y(n_1210)
);

BUFx6f_ASAP7_75t_L g1211 ( 
.A(n_1039),
.Y(n_1211)
);

AOI22xp33_ASAP7_75t_SL g1212 ( 
.A1(n_977),
.A2(n_896),
.B1(n_887),
.B2(n_895),
.Y(n_1212)
);

NAND2x1_ASAP7_75t_L g1213 ( 
.A(n_1079),
.B(n_869),
.Y(n_1213)
);

AND2x2_ASAP7_75t_L g1214 ( 
.A(n_1084),
.B(n_910),
.Y(n_1214)
);

INVx1_ASAP7_75t_SL g1215 ( 
.A(n_1068),
.Y(n_1215)
);

INVx1_ASAP7_75t_SL g1216 ( 
.A(n_1077),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1123),
.Y(n_1217)
);

AND2x4_ASAP7_75t_L g1218 ( 
.A(n_1066),
.B(n_895),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1011),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_996),
.B(n_894),
.Y(n_1220)
);

OAI221xp5_ASAP7_75t_L g1221 ( 
.A1(n_993),
.A2(n_863),
.B1(n_851),
.B2(n_930),
.C(n_923),
.Y(n_1221)
);

BUFx6f_ASAP7_75t_L g1222 ( 
.A(n_1042),
.Y(n_1222)
);

AND2x4_ASAP7_75t_L g1223 ( 
.A(n_1028),
.B(n_895),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_1128),
.Y(n_1224)
);

NOR2x1_ASAP7_75t_SL g1225 ( 
.A(n_1102),
.B(n_924),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_1005),
.Y(n_1226)
);

OAI21x1_ASAP7_75t_L g1227 ( 
.A1(n_1107),
.A2(n_913),
.B(n_875),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1015),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_975),
.B(n_909),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_975),
.B(n_909),
.Y(n_1230)
);

BUFx3_ASAP7_75t_L g1231 ( 
.A(n_1089),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_SL g1232 ( 
.A(n_1098),
.B(n_955),
.Y(n_1232)
);

INVx3_ASAP7_75t_L g1233 ( 
.A(n_1090),
.Y(n_1233)
);

AOI22xp33_ASAP7_75t_L g1234 ( 
.A1(n_977),
.A2(n_896),
.B1(n_923),
.B2(n_852),
.Y(n_1234)
);

INVx1_ASAP7_75t_SL g1235 ( 
.A(n_991),
.Y(n_1235)
);

NOR2x1_ASAP7_75t_SL g1236 ( 
.A(n_1102),
.B(n_955),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1009),
.B(n_835),
.Y(n_1237)
);

INVx3_ASAP7_75t_L g1238 ( 
.A(n_1090),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1000),
.A2(n_1012),
.B(n_1035),
.Y(n_1239)
);

AND2x4_ASAP7_75t_L g1240 ( 
.A(n_1028),
.B(n_1046),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_979),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1000),
.A2(n_961),
.B(n_793),
.Y(n_1242)
);

AOI22xp5_ASAP7_75t_L g1243 ( 
.A1(n_1085),
.A2(n_896),
.B1(n_850),
.B2(n_866),
.Y(n_1243)
);

CKINVDCx8_ASAP7_75t_R g1244 ( 
.A(n_1082),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_997),
.Y(n_1245)
);

BUFx2_ASAP7_75t_L g1246 ( 
.A(n_1022),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_997),
.Y(n_1247)
);

INVx2_ASAP7_75t_L g1248 ( 
.A(n_1126),
.Y(n_1248)
);

AND3x1_ASAP7_75t_SL g1249 ( 
.A(n_1064),
.B(n_36),
.C(n_38),
.Y(n_1249)
);

BUFx2_ASAP7_75t_L g1250 ( 
.A(n_1072),
.Y(n_1250)
);

AOI22xp5_ASAP7_75t_L g1251 ( 
.A1(n_1026),
.A2(n_891),
.B1(n_870),
.B2(n_971),
.Y(n_1251)
);

INVx2_ASAP7_75t_SL g1252 ( 
.A(n_1080),
.Y(n_1252)
);

BUFx8_ASAP7_75t_L g1253 ( 
.A(n_1042),
.Y(n_1253)
);

AOI22xp5_ASAP7_75t_L g1254 ( 
.A1(n_1099),
.A2(n_1067),
.B1(n_983),
.B2(n_1040),
.Y(n_1254)
);

A2O1A1Ixp33_ASAP7_75t_L g1255 ( 
.A1(n_1097),
.A2(n_961),
.B(n_912),
.C(n_875),
.Y(n_1255)
);

AOI221x1_ASAP7_75t_L g1256 ( 
.A1(n_1088),
.A2(n_912),
.B1(n_971),
.B2(n_943),
.C(n_939),
.Y(n_1256)
);

INVx4_ASAP7_75t_L g1257 ( 
.A(n_1079),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1126),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1007),
.Y(n_1259)
);

HB1xp67_ASAP7_75t_L g1260 ( 
.A(n_1042),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1007),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1009),
.A2(n_793),
.B(n_955),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1012),
.A2(n_906),
.B(n_911),
.Y(n_1263)
);

INVx3_ASAP7_75t_L g1264 ( 
.A(n_1090),
.Y(n_1264)
);

NOR2xp67_ASAP7_75t_L g1265 ( 
.A(n_1045),
.B(n_943),
.Y(n_1265)
);

OAI22xp5_ASAP7_75t_L g1266 ( 
.A1(n_977),
.A2(n_922),
.B1(n_933),
.B2(n_939),
.Y(n_1266)
);

INVx1_ASAP7_75t_SL g1267 ( 
.A(n_1061),
.Y(n_1267)
);

BUFx3_ASAP7_75t_L g1268 ( 
.A(n_1061),
.Y(n_1268)
);

BUFx6f_ASAP7_75t_L g1269 ( 
.A(n_1061),
.Y(n_1269)
);

BUFx6f_ASAP7_75t_L g1270 ( 
.A(n_1083),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1105),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1105),
.Y(n_1272)
);

INVx3_ASAP7_75t_SL g1273 ( 
.A(n_1106),
.Y(n_1273)
);

AOI22xp33_ASAP7_75t_L g1274 ( 
.A1(n_1052),
.A2(n_933),
.B1(n_891),
.B2(n_937),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_1074),
.Y(n_1275)
);

BUFx12f_ASAP7_75t_L g1276 ( 
.A(n_1083),
.Y(n_1276)
);

AOI22xp33_ASAP7_75t_L g1277 ( 
.A1(n_983),
.A2(n_891),
.B1(n_937),
.B2(n_869),
.Y(n_1277)
);

AND2x2_ASAP7_75t_SL g1278 ( 
.A(n_1106),
.B(n_926),
.Y(n_1278)
);

BUFx6f_ASAP7_75t_L g1279 ( 
.A(n_1083),
.Y(n_1279)
);

BUFx2_ASAP7_75t_L g1280 ( 
.A(n_1045),
.Y(n_1280)
);

INVx1_ASAP7_75t_SL g1281 ( 
.A(n_1122),
.Y(n_1281)
);

INVx3_ASAP7_75t_L g1282 ( 
.A(n_1090),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1096),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1167),
.A2(n_1069),
.B(n_1073),
.Y(n_1284)
);

AOI22xp33_ASAP7_75t_L g1285 ( 
.A1(n_1163),
.A2(n_985),
.B1(n_986),
.B2(n_1094),
.Y(n_1285)
);

AND2x2_ASAP7_75t_L g1286 ( 
.A(n_1235),
.B(n_1074),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1235),
.B(n_1122),
.Y(n_1287)
);

INVx3_ASAP7_75t_L g1288 ( 
.A(n_1233),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1131),
.Y(n_1289)
);

HB1xp67_ASAP7_75t_L g1290 ( 
.A(n_1161),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1132),
.Y(n_1291)
);

AO21x2_ASAP7_75t_L g1292 ( 
.A1(n_1188),
.A2(n_1069),
.B(n_1087),
.Y(n_1292)
);

OAI21x1_ASAP7_75t_L g1293 ( 
.A1(n_1227),
.A2(n_1081),
.B(n_1087),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_L g1294 ( 
.A1(n_1163),
.A2(n_1006),
.B1(n_1004),
.B2(n_1035),
.Y(n_1294)
);

OR2x2_ASAP7_75t_L g1295 ( 
.A(n_1159),
.B(n_1096),
.Y(n_1295)
);

OAI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1254),
.A2(n_1018),
.B1(n_1004),
.B2(n_1050),
.Y(n_1296)
);

AOI222xp33_ASAP7_75t_L g1297 ( 
.A1(n_1278),
.A2(n_1003),
.B1(n_1118),
.B2(n_1018),
.C1(n_1075),
.C2(n_1078),
.Y(n_1297)
);

INVx3_ASAP7_75t_L g1298 ( 
.A(n_1233),
.Y(n_1298)
);

BUFx2_ASAP7_75t_R g1299 ( 
.A(n_1177),
.Y(n_1299)
);

BUFx6f_ASAP7_75t_L g1300 ( 
.A(n_1151),
.Y(n_1300)
);

OA21x2_ASAP7_75t_L g1301 ( 
.A1(n_1256),
.A2(n_1095),
.B(n_1053),
.Y(n_1301)
);

AOI221xp5_ASAP7_75t_L g1302 ( 
.A1(n_1148),
.A2(n_1001),
.B1(n_1053),
.B2(n_1057),
.C(n_1065),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1138),
.Y(n_1303)
);

OR2x6_ASAP7_75t_L g1304 ( 
.A(n_1196),
.B(n_1102),
.Y(n_1304)
);

INVx3_ASAP7_75t_L g1305 ( 
.A(n_1238),
.Y(n_1305)
);

OAI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1173),
.A2(n_1073),
.B(n_1059),
.Y(n_1306)
);

OAI21x1_ASAP7_75t_SL g1307 ( 
.A1(n_1225),
.A2(n_1101),
.B(n_1058),
.Y(n_1307)
);

NAND2x1p5_ASAP7_75t_L g1308 ( 
.A(n_1153),
.B(n_1121),
.Y(n_1308)
);

INVx1_ASAP7_75t_SL g1309 ( 
.A(n_1174),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1147),
.Y(n_1310)
);

OR2x6_ASAP7_75t_L g1311 ( 
.A(n_1196),
.B(n_1153),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1156),
.Y(n_1312)
);

AO21x1_ASAP7_75t_L g1313 ( 
.A1(n_1188),
.A2(n_1100),
.B(n_1071),
.Y(n_1313)
);

BUFx3_ASAP7_75t_L g1314 ( 
.A(n_1253),
.Y(n_1314)
);

BUFx2_ASAP7_75t_L g1315 ( 
.A(n_1185),
.Y(n_1315)
);

OAI21x1_ASAP7_75t_L g1316 ( 
.A1(n_1262),
.A2(n_1101),
.B(n_992),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1160),
.Y(n_1317)
);

OAI21x1_ASAP7_75t_L g1318 ( 
.A1(n_1242),
.A2(n_1029),
.B(n_992),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1164),
.Y(n_1319)
);

OAI21x1_ASAP7_75t_L g1320 ( 
.A1(n_1242),
.A2(n_1029),
.B(n_917),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1193),
.B(n_1058),
.Y(n_1321)
);

NAND3xp33_ASAP7_75t_L g1322 ( 
.A(n_1152),
.B(n_915),
.C(n_1121),
.Y(n_1322)
);

INVx1_ASAP7_75t_SL g1323 ( 
.A(n_1174),
.Y(n_1323)
);

OAI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1165),
.A2(n_1121),
.B1(n_36),
.B2(n_419),
.Y(n_1324)
);

OAI21x1_ASAP7_75t_L g1325 ( 
.A1(n_1167),
.A2(n_891),
.B(n_1121),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1169),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1214),
.B(n_55),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1133),
.Y(n_1328)
);

AOI221xp5_ASAP7_75t_SL g1329 ( 
.A1(n_1266),
.A2(n_59),
.B1(n_61),
.B2(n_65),
.C(n_69),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1245),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1199),
.B(n_73),
.Y(n_1331)
);

BUFx6f_ASAP7_75t_L g1332 ( 
.A(n_1151),
.Y(n_1332)
);

AOI22xp33_ASAP7_75t_SL g1333 ( 
.A1(n_1202),
.A2(n_428),
.B1(n_445),
.B2(n_102),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1141),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1144),
.Y(n_1335)
);

AOI21xp5_ASAP7_75t_L g1336 ( 
.A1(n_1239),
.A2(n_585),
.B(n_562),
.Y(n_1336)
);

OAI21x1_ASAP7_75t_L g1337 ( 
.A1(n_1239),
.A2(n_95),
.B(n_97),
.Y(n_1337)
);

HB1xp67_ASAP7_75t_L g1338 ( 
.A(n_1161),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1247),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_1145),
.Y(n_1340)
);

INVx3_ASAP7_75t_L g1341 ( 
.A(n_1238),
.Y(n_1341)
);

HB1xp67_ASAP7_75t_L g1342 ( 
.A(n_1208),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1172),
.B(n_107),
.Y(n_1343)
);

OAI21x1_ASAP7_75t_L g1344 ( 
.A1(n_1166),
.A2(n_122),
.B(n_146),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1150),
.Y(n_1345)
);

OAI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1281),
.A2(n_585),
.B1(n_562),
.B2(n_594),
.Y(n_1346)
);

OAI21x1_ASAP7_75t_L g1347 ( 
.A1(n_1166),
.A2(n_148),
.B(n_152),
.Y(n_1347)
);

AOI22xp33_ASAP7_75t_L g1348 ( 
.A1(n_1259),
.A2(n_428),
.B1(n_445),
.B2(n_154),
.Y(n_1348)
);

OAI21x1_ASAP7_75t_SL g1349 ( 
.A1(n_1236),
.A2(n_155),
.B(n_428),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1240),
.B(n_404),
.Y(n_1350)
);

OR2x2_ASAP7_75t_L g1351 ( 
.A(n_1200),
.B(n_404),
.Y(n_1351)
);

AOI22xp5_ASAP7_75t_L g1352 ( 
.A1(n_1281),
.A2(n_404),
.B1(n_594),
.B2(n_1249),
.Y(n_1352)
);

AOI22xp33_ASAP7_75t_L g1353 ( 
.A1(n_1261),
.A2(n_404),
.B1(n_1221),
.B2(n_1143),
.Y(n_1353)
);

O2A1O1Ixp33_ASAP7_75t_SL g1354 ( 
.A1(n_1175),
.A2(n_404),
.B(n_1255),
.C(n_1154),
.Y(n_1354)
);

O2A1O1Ixp5_ASAP7_75t_SL g1355 ( 
.A1(n_1283),
.A2(n_404),
.B(n_1266),
.C(n_1162),
.Y(n_1355)
);

OA21x2_ASAP7_75t_L g1356 ( 
.A1(n_1194),
.A2(n_404),
.B(n_1154),
.Y(n_1356)
);

OA21x2_ASAP7_75t_L g1357 ( 
.A1(n_1194),
.A2(n_1263),
.B(n_1237),
.Y(n_1357)
);

XNOR2xp5_ASAP7_75t_L g1358 ( 
.A(n_1178),
.B(n_1209),
.Y(n_1358)
);

AOI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1221),
.A2(n_1237),
.B(n_1220),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1155),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1158),
.Y(n_1361)
);

OA21x2_ASAP7_75t_L g1362 ( 
.A1(n_1168),
.A2(n_1229),
.B(n_1230),
.Y(n_1362)
);

OAI21x1_ASAP7_75t_L g1363 ( 
.A1(n_1229),
.A2(n_1230),
.B(n_1248),
.Y(n_1363)
);

OAI21xp5_ASAP7_75t_L g1364 ( 
.A1(n_1201),
.A2(n_1243),
.B(n_1189),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_1258),
.Y(n_1365)
);

BUFx2_ASAP7_75t_L g1366 ( 
.A(n_1192),
.Y(n_1366)
);

BUFx3_ASAP7_75t_L g1367 ( 
.A(n_1253),
.Y(n_1367)
);

BUFx6f_ASAP7_75t_L g1368 ( 
.A(n_1151),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1143),
.B(n_1149),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1181),
.Y(n_1370)
);

AOI21xp5_ASAP7_75t_L g1371 ( 
.A1(n_1204),
.A2(n_1149),
.B(n_1274),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1184),
.Y(n_1372)
);

OR2x2_ASAP7_75t_L g1373 ( 
.A(n_1209),
.B(n_1208),
.Y(n_1373)
);

NAND2x1p5_ASAP7_75t_L g1374 ( 
.A(n_1162),
.B(n_1170),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1219),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1273),
.B(n_1179),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1271),
.Y(n_1377)
);

BUFx12f_ASAP7_75t_L g1378 ( 
.A(n_1129),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1228),
.Y(n_1379)
);

AOI21xp5_ASAP7_75t_L g1380 ( 
.A1(n_1204),
.A2(n_1274),
.B(n_1201),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1187),
.Y(n_1381)
);

OAI21x1_ASAP7_75t_L g1382 ( 
.A1(n_1272),
.A2(n_1234),
.B(n_1264),
.Y(n_1382)
);

OA21x2_ASAP7_75t_L g1383 ( 
.A1(n_1195),
.A2(n_1205),
.B(n_1197),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1226),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1217),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1176),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1157),
.B(n_1215),
.Y(n_1387)
);

AOI22xp33_ASAP7_75t_L g1388 ( 
.A1(n_1241),
.A2(n_1182),
.B1(n_1180),
.B2(n_1224),
.Y(n_1388)
);

OA21x2_ASAP7_75t_L g1389 ( 
.A1(n_1251),
.A2(n_1277),
.B(n_1203),
.Y(n_1389)
);

INVx6_ASAP7_75t_L g1390 ( 
.A(n_1276),
.Y(n_1390)
);

O2A1O1Ixp33_ASAP7_75t_L g1391 ( 
.A1(n_1232),
.A2(n_1215),
.B(n_1216),
.C(n_1134),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1260),
.Y(n_1392)
);

OA21x2_ASAP7_75t_L g1393 ( 
.A1(n_1275),
.A2(n_1249),
.B(n_1265),
.Y(n_1393)
);

AO21x2_ASAP7_75t_L g1394 ( 
.A1(n_1260),
.A2(n_1210),
.B(n_1218),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1240),
.B(n_1216),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1267),
.Y(n_1396)
);

AND2x2_ASAP7_75t_SL g1397 ( 
.A(n_1171),
.B(n_1246),
.Y(n_1397)
);

NAND2x1p5_ASAP7_75t_L g1398 ( 
.A(n_1264),
.B(n_1282),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1282),
.Y(n_1399)
);

BUFx3_ASAP7_75t_L g1400 ( 
.A(n_1198),
.Y(n_1400)
);

OAI22xp5_ASAP7_75t_L g1401 ( 
.A1(n_1212),
.A2(n_1196),
.B1(n_1136),
.B2(n_1210),
.Y(n_1401)
);

OAI21x1_ASAP7_75t_L g1402 ( 
.A1(n_1213),
.A2(n_1212),
.B(n_1206),
.Y(n_1402)
);

BUFx3_ASAP7_75t_L g1403 ( 
.A(n_1140),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1267),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1186),
.Y(n_1405)
);

OAI21x1_ASAP7_75t_L g1406 ( 
.A1(n_1206),
.A2(n_1257),
.B(n_1135),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1186),
.Y(n_1407)
);

NOR4xp25_ASAP7_75t_L g1408 ( 
.A(n_1252),
.B(n_1142),
.C(n_1244),
.D(n_1280),
.Y(n_1408)
);

O2A1O1Ixp33_ASAP7_75t_L g1409 ( 
.A1(n_1231),
.A2(n_1218),
.B(n_1250),
.C(n_1183),
.Y(n_1409)
);

BUFx12f_ASAP7_75t_L g1410 ( 
.A(n_1130),
.Y(n_1410)
);

OAI21xp5_ASAP7_75t_L g1411 ( 
.A1(n_1183),
.A2(n_1223),
.B(n_1257),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_1186),
.Y(n_1412)
);

O2A1O1Ixp33_ASAP7_75t_SL g1413 ( 
.A1(n_1190),
.A2(n_1211),
.B(n_1270),
.C(n_1269),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1190),
.Y(n_1414)
);

BUFx2_ASAP7_75t_L g1415 ( 
.A(n_1268),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_1190),
.Y(n_1416)
);

AOI21xp5_ASAP7_75t_SL g1417 ( 
.A1(n_1223),
.A2(n_1135),
.B(n_1146),
.Y(n_1417)
);

OAI21x1_ASAP7_75t_L g1418 ( 
.A1(n_1146),
.A2(n_1211),
.B(n_1270),
.Y(n_1418)
);

OA21x2_ASAP7_75t_L g1419 ( 
.A1(n_1191),
.A2(n_1211),
.B(n_1270),
.Y(n_1419)
);

OAI21x1_ASAP7_75t_L g1420 ( 
.A1(n_1191),
.A2(n_1207),
.B(n_1222),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1191),
.Y(n_1421)
);

CKINVDCx6p67_ASAP7_75t_R g1422 ( 
.A(n_1139),
.Y(n_1422)
);

AOI22xp33_ASAP7_75t_L g1423 ( 
.A1(n_1137),
.A2(n_1171),
.B1(n_1207),
.B2(n_1222),
.Y(n_1423)
);

HB1xp67_ASAP7_75t_L g1424 ( 
.A(n_1207),
.Y(n_1424)
);

CKINVDCx5p33_ASAP7_75t_R g1425 ( 
.A(n_1137),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1222),
.Y(n_1426)
);

OR2x6_ASAP7_75t_L g1427 ( 
.A(n_1269),
.B(n_1279),
.Y(n_1427)
);

INVx3_ASAP7_75t_L g1428 ( 
.A(n_1269),
.Y(n_1428)
);

OAI21x1_ASAP7_75t_L g1429 ( 
.A1(n_1279),
.A2(n_1227),
.B(n_1262),
.Y(n_1429)
);

INVx3_ASAP7_75t_L g1430 ( 
.A(n_1300),
.Y(n_1430)
);

OAI22xp33_ASAP7_75t_L g1431 ( 
.A1(n_1352),
.A2(n_1279),
.B1(n_1324),
.B2(n_1376),
.Y(n_1431)
);

AND2x4_ASAP7_75t_L g1432 ( 
.A(n_1304),
.B(n_1311),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1369),
.B(n_1295),
.Y(n_1433)
);

HB1xp67_ASAP7_75t_L g1434 ( 
.A(n_1290),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1340),
.Y(n_1435)
);

AOI22xp33_ASAP7_75t_L g1436 ( 
.A1(n_1297),
.A2(n_1324),
.B1(n_1364),
.B2(n_1322),
.Y(n_1436)
);

OR2x6_ASAP7_75t_L g1437 ( 
.A(n_1410),
.B(n_1417),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1340),
.Y(n_1438)
);

AND2x4_ASAP7_75t_L g1439 ( 
.A(n_1304),
.B(n_1311),
.Y(n_1439)
);

BUFx2_ASAP7_75t_L g1440 ( 
.A(n_1400),
.Y(n_1440)
);

OAI22xp5_ASAP7_75t_L g1441 ( 
.A1(n_1285),
.A2(n_1423),
.B1(n_1294),
.B2(n_1309),
.Y(n_1441)
);

AOI221xp5_ASAP7_75t_L g1442 ( 
.A1(n_1296),
.A2(n_1408),
.B1(n_1380),
.B2(n_1359),
.C(n_1354),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1345),
.Y(n_1443)
);

OAI21x1_ASAP7_75t_L g1444 ( 
.A1(n_1429),
.A2(n_1337),
.B(n_1293),
.Y(n_1444)
);

BUFx2_ASAP7_75t_L g1445 ( 
.A(n_1400),
.Y(n_1445)
);

INVx4_ASAP7_75t_L g1446 ( 
.A(n_1390),
.Y(n_1446)
);

AOI22xp5_ASAP7_75t_L g1447 ( 
.A1(n_1401),
.A2(n_1397),
.B1(n_1287),
.B2(n_1343),
.Y(n_1447)
);

CKINVDCx5p33_ASAP7_75t_R g1448 ( 
.A(n_1378),
.Y(n_1448)
);

INVx6_ASAP7_75t_L g1449 ( 
.A(n_1390),
.Y(n_1449)
);

OR2x2_ASAP7_75t_L g1450 ( 
.A(n_1373),
.B(n_1290),
.Y(n_1450)
);

NAND3x1_ASAP7_75t_L g1451 ( 
.A(n_1387),
.B(n_1395),
.C(n_1411),
.Y(n_1451)
);

INVx3_ASAP7_75t_L g1452 ( 
.A(n_1300),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1345),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1370),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1286),
.B(n_1321),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1370),
.Y(n_1456)
);

OAI22xp33_ASAP7_75t_L g1457 ( 
.A1(n_1304),
.A2(n_1311),
.B1(n_1410),
.B2(n_1323),
.Y(n_1457)
);

INVx1_ASAP7_75t_SL g1458 ( 
.A(n_1315),
.Y(n_1458)
);

AND2x6_ASAP7_75t_L g1459 ( 
.A(n_1377),
.B(n_1330),
.Y(n_1459)
);

INVx4_ASAP7_75t_L g1460 ( 
.A(n_1390),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1372),
.Y(n_1461)
);

AOI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1389),
.A2(n_1296),
.B1(n_1285),
.B2(n_1331),
.Y(n_1462)
);

BUFx6f_ASAP7_75t_L g1463 ( 
.A(n_1300),
.Y(n_1463)
);

AOI21xp5_ASAP7_75t_L g1464 ( 
.A1(n_1354),
.A2(n_1284),
.B(n_1371),
.Y(n_1464)
);

AOI22xp33_ASAP7_75t_L g1465 ( 
.A1(n_1389),
.A2(n_1302),
.B1(n_1327),
.B2(n_1393),
.Y(n_1465)
);

BUFx3_ASAP7_75t_L g1466 ( 
.A(n_1403),
.Y(n_1466)
);

AND2x4_ASAP7_75t_L g1467 ( 
.A(n_1394),
.B(n_1392),
.Y(n_1467)
);

AOI22xp33_ASAP7_75t_L g1468 ( 
.A1(n_1389),
.A2(n_1393),
.B1(n_1397),
.B2(n_1294),
.Y(n_1468)
);

OAI211xp5_ASAP7_75t_L g1469 ( 
.A1(n_1391),
.A2(n_1329),
.B(n_1409),
.C(n_1338),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1383),
.Y(n_1470)
);

INVx3_ASAP7_75t_L g1471 ( 
.A(n_1300),
.Y(n_1471)
);

OR2x6_ASAP7_75t_L g1472 ( 
.A(n_1402),
.B(n_1314),
.Y(n_1472)
);

OR2x2_ASAP7_75t_L g1473 ( 
.A(n_1338),
.B(n_1342),
.Y(n_1473)
);

BUFx2_ASAP7_75t_L g1474 ( 
.A(n_1366),
.Y(n_1474)
);

NAND3xp33_ASAP7_75t_L g1475 ( 
.A(n_1388),
.B(n_1306),
.C(n_1393),
.Y(n_1475)
);

OR2x2_ASAP7_75t_L g1476 ( 
.A(n_1342),
.B(n_1372),
.Y(n_1476)
);

AOI221xp5_ASAP7_75t_L g1477 ( 
.A1(n_1353),
.A2(n_1326),
.B1(n_1317),
.B2(n_1291),
.C(n_1312),
.Y(n_1477)
);

NOR2xp33_ASAP7_75t_L g1478 ( 
.A(n_1358),
.B(n_1299),
.Y(n_1478)
);

OAI221xp5_ASAP7_75t_L g1479 ( 
.A1(n_1333),
.A2(n_1423),
.B1(n_1353),
.B2(n_1348),
.C(n_1403),
.Y(n_1479)
);

CKINVDCx5p33_ASAP7_75t_R g1480 ( 
.A(n_1378),
.Y(n_1480)
);

INVx2_ASAP7_75t_SL g1481 ( 
.A(n_1314),
.Y(n_1481)
);

NAND3xp33_ASAP7_75t_L g1482 ( 
.A(n_1388),
.B(n_1333),
.C(n_1355),
.Y(n_1482)
);

OAI22xp33_ASAP7_75t_L g1483 ( 
.A1(n_1367),
.A2(n_1422),
.B1(n_1374),
.B2(n_1415),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1289),
.Y(n_1484)
);

AOI22xp33_ASAP7_75t_L g1485 ( 
.A1(n_1394),
.A2(n_1289),
.B1(n_1319),
.B2(n_1384),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1328),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1330),
.B(n_1339),
.Y(n_1487)
);

AOI22xp33_ASAP7_75t_L g1488 ( 
.A1(n_1319),
.A2(n_1384),
.B1(n_1367),
.B2(n_1339),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1334),
.Y(n_1489)
);

AOI222xp33_ASAP7_75t_L g1490 ( 
.A1(n_1303),
.A2(n_1310),
.B1(n_1335),
.B2(n_1361),
.C1(n_1360),
.C2(n_1375),
.Y(n_1490)
);

AOI22xp33_ASAP7_75t_L g1491 ( 
.A1(n_1313),
.A2(n_1386),
.B1(n_1365),
.B2(n_1381),
.Y(n_1491)
);

INVx3_ASAP7_75t_L g1492 ( 
.A(n_1332),
.Y(n_1492)
);

AND2x4_ASAP7_75t_L g1493 ( 
.A(n_1402),
.B(n_1404),
.Y(n_1493)
);

NOR2xp33_ASAP7_75t_L g1494 ( 
.A(n_1425),
.B(n_1351),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1365),
.B(n_1377),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_SL g1496 ( 
.A1(n_1344),
.A2(n_1347),
.B1(n_1374),
.B2(n_1349),
.Y(n_1496)
);

BUFx6f_ASAP7_75t_L g1497 ( 
.A(n_1332),
.Y(n_1497)
);

AOI22xp33_ASAP7_75t_SL g1498 ( 
.A1(n_1357),
.A2(n_1379),
.B1(n_1307),
.B2(n_1362),
.Y(n_1498)
);

NAND2xp33_ASAP7_75t_SL g1499 ( 
.A(n_1425),
.B(n_1332),
.Y(n_1499)
);

AND2x4_ASAP7_75t_L g1500 ( 
.A(n_1396),
.B(n_1399),
.Y(n_1500)
);

OAI22xp5_ASAP7_75t_SL g1501 ( 
.A1(n_1398),
.A2(n_1385),
.B1(n_1427),
.B2(n_1308),
.Y(n_1501)
);

AND2x4_ASAP7_75t_L g1502 ( 
.A(n_1399),
.B(n_1288),
.Y(n_1502)
);

INVx3_ASAP7_75t_L g1503 ( 
.A(n_1332),
.Y(n_1503)
);

BUFx2_ASAP7_75t_SL g1504 ( 
.A(n_1405),
.Y(n_1504)
);

OAI22xp5_ASAP7_75t_L g1505 ( 
.A1(n_1308),
.A2(n_1348),
.B1(n_1398),
.B2(n_1414),
.Y(n_1505)
);

CKINVDCx6p67_ASAP7_75t_R g1506 ( 
.A(n_1427),
.Y(n_1506)
);

OAI21x1_ASAP7_75t_L g1507 ( 
.A1(n_1316),
.A2(n_1325),
.B(n_1318),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1383),
.Y(n_1508)
);

OR2x6_ASAP7_75t_L g1509 ( 
.A(n_1406),
.B(n_1382),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1363),
.B(n_1362),
.Y(n_1510)
);

OAI22xp33_ASAP7_75t_L g1511 ( 
.A1(n_1362),
.A2(n_1288),
.B1(n_1341),
.B2(n_1298),
.Y(n_1511)
);

OAI21xp5_ASAP7_75t_L g1512 ( 
.A1(n_1382),
.A2(n_1320),
.B(n_1336),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1424),
.B(n_1416),
.Y(n_1513)
);

AOI22xp33_ASAP7_75t_L g1514 ( 
.A1(n_1298),
.A2(n_1305),
.B1(n_1341),
.B2(n_1350),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1424),
.B(n_1412),
.Y(n_1515)
);

INVx3_ASAP7_75t_L g1516 ( 
.A(n_1368),
.Y(n_1516)
);

AND2x4_ASAP7_75t_L g1517 ( 
.A(n_1305),
.B(n_1406),
.Y(n_1517)
);

OA21x2_ASAP7_75t_L g1518 ( 
.A1(n_1420),
.A2(n_1418),
.B(n_1356),
.Y(n_1518)
);

INVx2_ASAP7_75t_SL g1519 ( 
.A(n_1368),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1292),
.Y(n_1520)
);

OAI211xp5_ASAP7_75t_SL g1521 ( 
.A1(n_1407),
.A2(n_1426),
.B(n_1421),
.C(n_1416),
.Y(n_1521)
);

CKINVDCx20_ASAP7_75t_R g1522 ( 
.A(n_1368),
.Y(n_1522)
);

OR2x6_ASAP7_75t_L g1523 ( 
.A(n_1418),
.B(n_1427),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1419),
.Y(n_1524)
);

AOI221xp5_ASAP7_75t_SL g1525 ( 
.A1(n_1405),
.A2(n_1412),
.B1(n_1368),
.B2(n_1428),
.C(n_1346),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1357),
.B(n_1428),
.Y(n_1526)
);

AOI21xp33_ASAP7_75t_L g1527 ( 
.A1(n_1292),
.A2(n_1301),
.B(n_1356),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1301),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1419),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_SL g1530 ( 
.A(n_1420),
.B(n_1413),
.Y(n_1530)
);

AOI22xp33_ASAP7_75t_L g1531 ( 
.A1(n_1419),
.A2(n_1413),
.B1(n_1013),
.B2(n_1163),
.Y(n_1531)
);

CKINVDCx8_ASAP7_75t_R g1532 ( 
.A(n_1425),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1340),
.Y(n_1533)
);

AOI222xp33_ASAP7_75t_L g1534 ( 
.A1(n_1324),
.A2(n_1013),
.B1(n_1163),
.B2(n_978),
.C1(n_741),
.C2(n_407),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1369),
.B(n_1235),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1286),
.B(n_1287),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1286),
.B(n_1287),
.Y(n_1537)
);

CKINVDCx5p33_ASAP7_75t_R g1538 ( 
.A(n_1378),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1340),
.Y(n_1539)
);

A2O1A1Ixp33_ASAP7_75t_L g1540 ( 
.A1(n_1364),
.A2(n_1163),
.B(n_1063),
.C(n_1013),
.Y(n_1540)
);

INVxp67_ASAP7_75t_SL g1541 ( 
.A(n_1342),
.Y(n_1541)
);

INVx4_ASAP7_75t_L g1542 ( 
.A(n_1390),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1369),
.B(n_1235),
.Y(n_1543)
);

OAI22xp33_ASAP7_75t_SL g1544 ( 
.A1(n_1369),
.A2(n_407),
.B1(n_948),
.B2(n_938),
.Y(n_1544)
);

AO21x2_ASAP7_75t_L g1545 ( 
.A1(n_1284),
.A2(n_1380),
.B(n_1371),
.Y(n_1545)
);

CKINVDCx20_ASAP7_75t_R g1546 ( 
.A(n_1425),
.Y(n_1546)
);

CKINVDCx11_ASAP7_75t_R g1547 ( 
.A(n_1378),
.Y(n_1547)
);

AND2x2_ASAP7_75t_SL g1548 ( 
.A(n_1442),
.B(n_1436),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1433),
.B(n_1535),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1543),
.B(n_1450),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1455),
.B(n_1536),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1537),
.B(n_1513),
.Y(n_1552)
);

OAI22xp5_ASAP7_75t_L g1553 ( 
.A1(n_1540),
.A2(n_1479),
.B1(n_1462),
.B2(n_1447),
.Y(n_1553)
);

AND2x4_ASAP7_75t_L g1554 ( 
.A(n_1493),
.B(n_1432),
.Y(n_1554)
);

OR2x2_ASAP7_75t_L g1555 ( 
.A(n_1473),
.B(n_1476),
.Y(n_1555)
);

AND2x4_ASAP7_75t_L g1556 ( 
.A(n_1493),
.B(n_1432),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1434),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1541),
.B(n_1490),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1470),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1439),
.B(n_1467),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1500),
.B(n_1438),
.Y(n_1561)
);

CKINVDCx5p33_ASAP7_75t_R g1562 ( 
.A(n_1547),
.Y(n_1562)
);

AND2x2_ASAP7_75t_SL g1563 ( 
.A(n_1468),
.B(n_1439),
.Y(n_1563)
);

CKINVDCx20_ASAP7_75t_R g1564 ( 
.A(n_1546),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1486),
.Y(n_1565)
);

AOI22xp33_ASAP7_75t_L g1566 ( 
.A1(n_1534),
.A2(n_1544),
.B1(n_1441),
.B2(n_1431),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1489),
.Y(n_1567)
);

HB1xp67_ASAP7_75t_L g1568 ( 
.A(n_1524),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1435),
.Y(n_1569)
);

NAND2xp33_ASAP7_75t_SL g1570 ( 
.A(n_1501),
.B(n_1446),
.Y(n_1570)
);

CKINVDCx16_ASAP7_75t_R g1571 ( 
.A(n_1522),
.Y(n_1571)
);

CKINVDCx16_ASAP7_75t_R g1572 ( 
.A(n_1478),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1467),
.B(n_1500),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1443),
.Y(n_1574)
);

CKINVDCx20_ASAP7_75t_R g1575 ( 
.A(n_1448),
.Y(n_1575)
);

INVxp67_ASAP7_75t_L g1576 ( 
.A(n_1474),
.Y(n_1576)
);

AOI221xp5_ASAP7_75t_L g1577 ( 
.A1(n_1475),
.A2(n_1469),
.B1(n_1465),
.B2(n_1457),
.C(n_1477),
.Y(n_1577)
);

INVx4_ASAP7_75t_L g1578 ( 
.A(n_1437),
.Y(n_1578)
);

AND2x6_ASAP7_75t_L g1579 ( 
.A(n_1517),
.B(n_1453),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_1454),
.Y(n_1580)
);

O2A1O1Ixp33_ASAP7_75t_L g1581 ( 
.A1(n_1483),
.A2(n_1505),
.B(n_1437),
.C(n_1464),
.Y(n_1581)
);

INVx3_ASAP7_75t_L g1582 ( 
.A(n_1502),
.Y(n_1582)
);

OR2x6_ASAP7_75t_L g1583 ( 
.A(n_1509),
.B(n_1472),
.Y(n_1583)
);

NOR3xp33_ASAP7_75t_SL g1584 ( 
.A(n_1480),
.B(n_1538),
.C(n_1521),
.Y(n_1584)
);

OR2x2_ASAP7_75t_L g1585 ( 
.A(n_1533),
.B(n_1539),
.Y(n_1585)
);

OR2x6_ASAP7_75t_L g1586 ( 
.A(n_1509),
.B(n_1472),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1456),
.B(n_1461),
.Y(n_1587)
);

INVx2_ASAP7_75t_SL g1588 ( 
.A(n_1449),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_1508),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1529),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1515),
.B(n_1440),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1495),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1445),
.B(n_1458),
.Y(n_1593)
);

CKINVDCx8_ASAP7_75t_R g1594 ( 
.A(n_1504),
.Y(n_1594)
);

CKINVDCx20_ASAP7_75t_R g1595 ( 
.A(n_1532),
.Y(n_1595)
);

BUFx8_ASAP7_75t_SL g1596 ( 
.A(n_1466),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1487),
.B(n_1484),
.Y(n_1597)
);

HB1xp67_ASAP7_75t_L g1598 ( 
.A(n_1526),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1510),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1528),
.Y(n_1600)
);

BUFx3_ASAP7_75t_L g1601 ( 
.A(n_1449),
.Y(n_1601)
);

INVxp67_ASAP7_75t_SL g1602 ( 
.A(n_1520),
.Y(n_1602)
);

AND2x4_ASAP7_75t_L g1603 ( 
.A(n_1517),
.B(n_1523),
.Y(n_1603)
);

CKINVDCx5p33_ASAP7_75t_R g1604 ( 
.A(n_1481),
.Y(n_1604)
);

OAI21x1_ASAP7_75t_SL g1605 ( 
.A1(n_1531),
.A2(n_1491),
.B(n_1542),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1528),
.Y(n_1606)
);

NOR3xp33_ASAP7_75t_SL g1607 ( 
.A(n_1499),
.B(n_1494),
.C(n_1511),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1518),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1502),
.B(n_1485),
.Y(n_1609)
);

BUFx2_ASAP7_75t_L g1610 ( 
.A(n_1523),
.Y(n_1610)
);

NOR3xp33_ASAP7_75t_SL g1611 ( 
.A(n_1530),
.B(n_1482),
.C(n_1512),
.Y(n_1611)
);

CKINVDCx20_ASAP7_75t_R g1612 ( 
.A(n_1506),
.Y(n_1612)
);

CKINVDCx5p33_ASAP7_75t_R g1613 ( 
.A(n_1446),
.Y(n_1613)
);

OAI21xp5_ASAP7_75t_L g1614 ( 
.A1(n_1451),
.A2(n_1496),
.B(n_1525),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_1518),
.Y(n_1615)
);

AOI21xp33_ASAP7_75t_L g1616 ( 
.A1(n_1545),
.A2(n_1488),
.B(n_1514),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1459),
.B(n_1430),
.Y(n_1617)
);

AOI22xp33_ASAP7_75t_L g1618 ( 
.A1(n_1545),
.A2(n_1542),
.B1(n_1460),
.B2(n_1459),
.Y(n_1618)
);

CKINVDCx5p33_ASAP7_75t_R g1619 ( 
.A(n_1460),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1430),
.B(n_1516),
.Y(n_1620)
);

OR2x2_ASAP7_75t_L g1621 ( 
.A(n_1520),
.B(n_1498),
.Y(n_1621)
);

BUFx3_ASAP7_75t_L g1622 ( 
.A(n_1579),
.Y(n_1622)
);

HB1xp67_ASAP7_75t_L g1623 ( 
.A(n_1568),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1559),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1598),
.B(n_1527),
.Y(n_1625)
);

AOI22xp33_ASAP7_75t_L g1626 ( 
.A1(n_1548),
.A2(n_1459),
.B1(n_1503),
.B2(n_1452),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1590),
.Y(n_1627)
);

OR2x2_ASAP7_75t_L g1628 ( 
.A(n_1598),
.B(n_1507),
.Y(n_1628)
);

AND2x4_ASAP7_75t_L g1629 ( 
.A(n_1603),
.B(n_1444),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1600),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1589),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1600),
.Y(n_1632)
);

HB1xp67_ASAP7_75t_L g1633 ( 
.A(n_1568),
.Y(n_1633)
);

OR2x2_ASAP7_75t_L g1634 ( 
.A(n_1621),
.B(n_1452),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1606),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1606),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1580),
.Y(n_1637)
);

INVx2_ASAP7_75t_SL g1638 ( 
.A(n_1603),
.Y(n_1638)
);

AND2x4_ASAP7_75t_L g1639 ( 
.A(n_1603),
.B(n_1471),
.Y(n_1639)
);

INVx2_ASAP7_75t_SL g1640 ( 
.A(n_1579),
.Y(n_1640)
);

BUFx4_ASAP7_75t_SL g1641 ( 
.A(n_1575),
.Y(n_1641)
);

HB1xp67_ASAP7_75t_L g1642 ( 
.A(n_1599),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1608),
.B(n_1471),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1615),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1565),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1615),
.B(n_1492),
.Y(n_1646)
);

OR2x2_ASAP7_75t_L g1647 ( 
.A(n_1555),
.B(n_1492),
.Y(n_1647)
);

BUFx2_ASAP7_75t_L g1648 ( 
.A(n_1583),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1580),
.Y(n_1649)
);

BUFx3_ASAP7_75t_L g1650 ( 
.A(n_1579),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1583),
.B(n_1503),
.Y(n_1651)
);

OR2x2_ASAP7_75t_L g1652 ( 
.A(n_1557),
.B(n_1516),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1569),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1574),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1567),
.Y(n_1655)
);

HB1xp67_ASAP7_75t_L g1656 ( 
.A(n_1602),
.Y(n_1656)
);

INVx3_ASAP7_75t_L g1657 ( 
.A(n_1579),
.Y(n_1657)
);

INVx2_ASAP7_75t_SL g1658 ( 
.A(n_1579),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1583),
.B(n_1463),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1586),
.B(n_1463),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1585),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1586),
.B(n_1463),
.Y(n_1662)
);

NOR2xp33_ASAP7_75t_L g1663 ( 
.A(n_1634),
.B(n_1548),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1647),
.B(n_1591),
.Y(n_1664)
);

OAI21xp5_ASAP7_75t_SL g1665 ( 
.A1(n_1626),
.A2(n_1566),
.B(n_1553),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1638),
.B(n_1560),
.Y(n_1666)
);

NAND2xp33_ASAP7_75t_SL g1667 ( 
.A(n_1641),
.B(n_1584),
.Y(n_1667)
);

OAI221xp5_ASAP7_75t_L g1668 ( 
.A1(n_1648),
.A2(n_1566),
.B1(n_1577),
.B2(n_1614),
.C(n_1607),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1638),
.B(n_1610),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1647),
.B(n_1550),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1647),
.B(n_1558),
.Y(n_1671)
);

NAND3xp33_ASAP7_75t_L g1672 ( 
.A(n_1625),
.B(n_1611),
.C(n_1581),
.Y(n_1672)
);

AOI221xp5_ASAP7_75t_L g1673 ( 
.A1(n_1625),
.A2(n_1576),
.B1(n_1616),
.B2(n_1549),
.C(n_1592),
.Y(n_1673)
);

NAND2xp33_ASAP7_75t_SL g1674 ( 
.A(n_1641),
.B(n_1612),
.Y(n_1674)
);

AOI22xp33_ASAP7_75t_L g1675 ( 
.A1(n_1648),
.A2(n_1563),
.B1(n_1605),
.B2(n_1578),
.Y(n_1675)
);

OAI22xp5_ASAP7_75t_L g1676 ( 
.A1(n_1626),
.A2(n_1594),
.B1(n_1563),
.B2(n_1613),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1638),
.B(n_1556),
.Y(n_1677)
);

OAI22xp5_ASAP7_75t_L g1678 ( 
.A1(n_1634),
.A2(n_1613),
.B1(n_1612),
.B2(n_1604),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1639),
.B(n_1651),
.Y(n_1679)
);

OAI22xp5_ASAP7_75t_L g1680 ( 
.A1(n_1634),
.A2(n_1604),
.B1(n_1578),
.B2(n_1618),
.Y(n_1680)
);

NAND3xp33_ASAP7_75t_L g1681 ( 
.A(n_1628),
.B(n_1618),
.C(n_1609),
.Y(n_1681)
);

NOR3xp33_ASAP7_75t_L g1682 ( 
.A(n_1648),
.B(n_1570),
.C(n_1572),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1642),
.B(n_1552),
.Y(n_1683)
);

NOR3xp33_ASAP7_75t_L g1684 ( 
.A(n_1628),
.B(n_1570),
.C(n_1571),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1642),
.B(n_1573),
.Y(n_1685)
);

NAND2xp33_ASAP7_75t_SL g1686 ( 
.A(n_1640),
.B(n_1595),
.Y(n_1686)
);

NAND3xp33_ASAP7_75t_L g1687 ( 
.A(n_1628),
.B(n_1561),
.C(n_1617),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1661),
.B(n_1593),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1661),
.B(n_1645),
.Y(n_1689)
);

NOR3xp33_ASAP7_75t_L g1690 ( 
.A(n_1651),
.B(n_1588),
.C(n_1562),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1661),
.B(n_1551),
.Y(n_1691)
);

OAI21xp33_ASAP7_75t_SL g1692 ( 
.A1(n_1640),
.A2(n_1586),
.B(n_1587),
.Y(n_1692)
);

NAND3xp33_ASAP7_75t_L g1693 ( 
.A(n_1656),
.B(n_1597),
.C(n_1582),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1639),
.B(n_1554),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_SL g1695 ( 
.A(n_1622),
.B(n_1554),
.Y(n_1695)
);

OAI221xp5_ASAP7_75t_L g1696 ( 
.A1(n_1640),
.A2(n_1601),
.B1(n_1619),
.B2(n_1582),
.C(n_1519),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1645),
.B(n_1554),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1652),
.B(n_1556),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1639),
.B(n_1556),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1652),
.B(n_1620),
.Y(n_1700)
);

NAND2xp33_ASAP7_75t_SL g1701 ( 
.A(n_1658),
.B(n_1595),
.Y(n_1701)
);

NAND3xp33_ASAP7_75t_L g1702 ( 
.A(n_1656),
.B(n_1652),
.C(n_1653),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1651),
.B(n_1601),
.Y(n_1703)
);

OAI221xp5_ASAP7_75t_L g1704 ( 
.A1(n_1658),
.A2(n_1497),
.B1(n_1596),
.B2(n_1575),
.C(n_1564),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1655),
.B(n_1596),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1643),
.B(n_1497),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1671),
.B(n_1623),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1679),
.B(n_1629),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1689),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1702),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1691),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1697),
.Y(n_1712)
);

INVx3_ASAP7_75t_L g1713 ( 
.A(n_1669),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1694),
.B(n_1629),
.Y(n_1714)
);

HB1xp67_ASAP7_75t_L g1715 ( 
.A(n_1693),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1669),
.B(n_1629),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1706),
.B(n_1629),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1663),
.B(n_1673),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1670),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1663),
.B(n_1623),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1706),
.B(n_1629),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1700),
.Y(n_1722)
);

OAI221xp5_ASAP7_75t_SL g1723 ( 
.A1(n_1665),
.A2(n_1650),
.B1(n_1622),
.B2(n_1658),
.C(n_1633),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1699),
.B(n_1629),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1687),
.B(n_1633),
.Y(n_1725)
);

OR2x2_ASAP7_75t_L g1726 ( 
.A(n_1683),
.B(n_1681),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1677),
.B(n_1657),
.Y(n_1727)
);

INVx3_ASAP7_75t_L g1728 ( 
.A(n_1703),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1688),
.Y(n_1729)
);

OR2x2_ASAP7_75t_L g1730 ( 
.A(n_1664),
.B(n_1655),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1685),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1698),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1672),
.B(n_1655),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1695),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1703),
.B(n_1657),
.Y(n_1735)
);

INVx1_ASAP7_75t_SL g1736 ( 
.A(n_1674),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1695),
.Y(n_1737)
);

NOR2xp33_ASAP7_75t_L g1738 ( 
.A(n_1674),
.B(n_1564),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1666),
.B(n_1646),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1692),
.B(n_1655),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_SL g1741 ( 
.A(n_1682),
.B(n_1639),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1705),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1684),
.B(n_1657),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1730),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1733),
.B(n_1678),
.Y(n_1745)
);

INVx2_ASAP7_75t_L g1746 ( 
.A(n_1739),
.Y(n_1746)
);

OR2x2_ASAP7_75t_L g1747 ( 
.A(n_1733),
.B(n_1654),
.Y(n_1747)
);

OR2x2_ASAP7_75t_L g1748 ( 
.A(n_1710),
.B(n_1654),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1730),
.Y(n_1749)
);

OR2x2_ASAP7_75t_L g1750 ( 
.A(n_1710),
.B(n_1654),
.Y(n_1750)
);

AND2x4_ASAP7_75t_L g1751 ( 
.A(n_1728),
.B(n_1743),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1739),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1718),
.B(n_1675),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1718),
.B(n_1668),
.Y(n_1754)
);

INVx3_ASAP7_75t_L g1755 ( 
.A(n_1713),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1709),
.Y(n_1756)
);

INVx2_ASAP7_75t_L g1757 ( 
.A(n_1739),
.Y(n_1757)
);

INVx2_ASAP7_75t_L g1758 ( 
.A(n_1713),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1742),
.B(n_1690),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1713),
.Y(n_1760)
);

INVxp67_ASAP7_75t_SL g1761 ( 
.A(n_1715),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1717),
.B(n_1657),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1709),
.Y(n_1763)
);

NOR2xp67_ASAP7_75t_L g1764 ( 
.A(n_1715),
.B(n_1704),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1742),
.B(n_1680),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1709),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1711),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1717),
.B(n_1721),
.Y(n_1768)
);

OR2x2_ASAP7_75t_L g1769 ( 
.A(n_1710),
.B(n_1654),
.Y(n_1769)
);

INVx3_ASAP7_75t_L g1770 ( 
.A(n_1713),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1717),
.B(n_1657),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1719),
.B(n_1653),
.Y(n_1772)
);

NOR2xp33_ASAP7_75t_L g1773 ( 
.A(n_1738),
.B(n_1696),
.Y(n_1773)
);

OR2x2_ASAP7_75t_L g1774 ( 
.A(n_1731),
.B(n_1637),
.Y(n_1774)
);

NOR2x1_ASAP7_75t_L g1775 ( 
.A(n_1736),
.B(n_1676),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1719),
.B(n_1653),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1711),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1721),
.B(n_1650),
.Y(n_1778)
);

INVx2_ASAP7_75t_L g1779 ( 
.A(n_1712),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1721),
.B(n_1650),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1712),
.B(n_1639),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1714),
.B(n_1650),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1729),
.Y(n_1783)
);

INVx1_ASAP7_75t_SL g1784 ( 
.A(n_1736),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1729),
.B(n_1639),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1748),
.Y(n_1786)
);

INVxp67_ASAP7_75t_SL g1787 ( 
.A(n_1764),
.Y(n_1787)
);

INVx2_ASAP7_75t_L g1788 ( 
.A(n_1755),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1748),
.Y(n_1789)
);

AOI21x1_ASAP7_75t_L g1790 ( 
.A1(n_1754),
.A2(n_1741),
.B(n_1725),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1784),
.B(n_1726),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1750),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_1755),
.Y(n_1793)
);

OAI33xp33_ASAP7_75t_L g1794 ( 
.A1(n_1753),
.A2(n_1745),
.A3(n_1767),
.B1(n_1783),
.B2(n_1777),
.B3(n_1765),
.Y(n_1794)
);

AOI32xp33_ASAP7_75t_L g1795 ( 
.A1(n_1775),
.A2(n_1743),
.A3(n_1737),
.B1(n_1734),
.B2(n_1726),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1778),
.B(n_1780),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1778),
.B(n_1728),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1755),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1750),
.Y(n_1799)
);

OA222x2_ASAP7_75t_L g1800 ( 
.A1(n_1770),
.A2(n_1725),
.B1(n_1728),
.B2(n_1737),
.C1(n_1734),
.C2(n_1622),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1761),
.B(n_1732),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1780),
.B(n_1728),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1768),
.B(n_1724),
.Y(n_1803)
);

NOR2xp33_ASAP7_75t_SL g1804 ( 
.A(n_1775),
.B(n_1723),
.Y(n_1804)
);

OR2x6_ASAP7_75t_L g1805 ( 
.A(n_1751),
.B(n_1740),
.Y(n_1805)
);

INVx3_ASAP7_75t_L g1806 ( 
.A(n_1770),
.Y(n_1806)
);

AOI22xp33_ASAP7_75t_L g1807 ( 
.A1(n_1773),
.A2(n_1667),
.B1(n_1701),
.B2(n_1686),
.Y(n_1807)
);

A2O1A1Ixp33_ASAP7_75t_L g1808 ( 
.A1(n_1759),
.A2(n_1723),
.B(n_1667),
.C(n_1686),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1767),
.B(n_1732),
.Y(n_1809)
);

NOR2xp33_ASAP7_75t_L g1810 ( 
.A(n_1751),
.B(n_1720),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1769),
.Y(n_1811)
);

NAND4xp25_ASAP7_75t_L g1812 ( 
.A(n_1751),
.B(n_1777),
.C(n_1783),
.D(n_1720),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1768),
.B(n_1724),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1769),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1779),
.B(n_1731),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1779),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1782),
.B(n_1724),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1772),
.Y(n_1818)
);

OAI211xp5_ASAP7_75t_L g1819 ( 
.A1(n_1758),
.A2(n_1740),
.B(n_1701),
.C(n_1707),
.Y(n_1819)
);

NAND2x1_ASAP7_75t_L g1820 ( 
.A(n_1770),
.B(n_1735),
.Y(n_1820)
);

AOI21xp33_ASAP7_75t_L g1821 ( 
.A1(n_1804),
.A2(n_1744),
.B(n_1749),
.Y(n_1821)
);

AOI21xp5_ASAP7_75t_L g1822 ( 
.A1(n_1787),
.A2(n_1776),
.B(n_1747),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1816),
.Y(n_1823)
);

OAI21xp5_ASAP7_75t_L g1824 ( 
.A1(n_1808),
.A2(n_1747),
.B(n_1758),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1795),
.B(n_1731),
.Y(n_1825)
);

INVx1_ASAP7_75t_SL g1826 ( 
.A(n_1791),
.Y(n_1826)
);

AOI221xp5_ASAP7_75t_L g1827 ( 
.A1(n_1794),
.A2(n_1744),
.B1(n_1749),
.B2(n_1760),
.C(n_1756),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1796),
.B(n_1782),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1786),
.Y(n_1829)
);

INVx1_ASAP7_75t_SL g1830 ( 
.A(n_1801),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1789),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1792),
.Y(n_1832)
);

HB1xp67_ASAP7_75t_L g1833 ( 
.A(n_1799),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1811),
.Y(n_1834)
);

NAND2xp33_ASAP7_75t_SL g1835 ( 
.A(n_1807),
.B(n_1760),
.Y(n_1835)
);

OAI21xp33_ASAP7_75t_L g1836 ( 
.A1(n_1808),
.A2(n_1746),
.B(n_1752),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1814),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1809),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1806),
.Y(n_1839)
);

OR2x2_ASAP7_75t_L g1840 ( 
.A(n_1812),
.B(n_1746),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1815),
.Y(n_1841)
);

OR2x2_ASAP7_75t_L g1842 ( 
.A(n_1805),
.B(n_1752),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1810),
.B(n_1757),
.Y(n_1843)
);

INVx2_ASAP7_75t_L g1844 ( 
.A(n_1806),
.Y(n_1844)
);

NAND2xp33_ASAP7_75t_R g1845 ( 
.A(n_1805),
.B(n_1762),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1833),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1828),
.B(n_1796),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1839),
.Y(n_1848)
);

BUFx3_ASAP7_75t_L g1849 ( 
.A(n_1829),
.Y(n_1849)
);

O2A1O1Ixp33_ASAP7_75t_SL g1850 ( 
.A1(n_1821),
.A2(n_1819),
.B(n_1820),
.C(n_1800),
.Y(n_1850)
);

OAI32xp33_ASAP7_75t_L g1851 ( 
.A1(n_1845),
.A2(n_1810),
.A3(n_1806),
.B1(n_1790),
.B2(n_1793),
.Y(n_1851)
);

OR2x2_ASAP7_75t_L g1852 ( 
.A(n_1826),
.B(n_1805),
.Y(n_1852)
);

NOR2x1p5_ASAP7_75t_L g1853 ( 
.A(n_1840),
.B(n_1790),
.Y(n_1853)
);

NOR2xp33_ASAP7_75t_L g1854 ( 
.A(n_1830),
.B(n_1805),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1843),
.B(n_1797),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1833),
.Y(n_1856)
);

AOI21xp5_ASAP7_75t_L g1857 ( 
.A1(n_1835),
.A2(n_1818),
.B(n_1793),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_L g1858 ( 
.A(n_1831),
.B(n_1832),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1823),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1834),
.B(n_1757),
.Y(n_1860)
);

OAI22xp5_ASAP7_75t_L g1861 ( 
.A1(n_1825),
.A2(n_1802),
.B1(n_1797),
.B2(n_1798),
.Y(n_1861)
);

OR2x2_ASAP7_75t_L g1862 ( 
.A(n_1842),
.B(n_1817),
.Y(n_1862)
);

NOR2xp33_ASAP7_75t_L g1863 ( 
.A(n_1838),
.B(n_1802),
.Y(n_1863)
);

AND2x4_ASAP7_75t_L g1864 ( 
.A(n_1839),
.B(n_1817),
.Y(n_1864)
);

OR2x2_ASAP7_75t_L g1865 ( 
.A(n_1862),
.B(n_1837),
.Y(n_1865)
);

NOR2xp33_ASAP7_75t_L g1866 ( 
.A(n_1852),
.B(n_1835),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1855),
.B(n_1841),
.Y(n_1867)
);

AOI21xp5_ASAP7_75t_L g1868 ( 
.A1(n_1850),
.A2(n_1824),
.B(n_1822),
.Y(n_1868)
);

INVxp67_ASAP7_75t_L g1869 ( 
.A(n_1854),
.Y(n_1869)
);

INVx2_ASAP7_75t_SL g1870 ( 
.A(n_1864),
.Y(n_1870)
);

AOI22xp5_ASAP7_75t_L g1871 ( 
.A1(n_1853),
.A2(n_1845),
.B1(n_1836),
.B2(n_1827),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1846),
.Y(n_1872)
);

AOI22xp5_ASAP7_75t_L g1873 ( 
.A1(n_1847),
.A2(n_1844),
.B1(n_1798),
.B2(n_1788),
.Y(n_1873)
);

OAI211xp5_ASAP7_75t_L g1874 ( 
.A1(n_1851),
.A2(n_1844),
.B(n_1788),
.C(n_1803),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1856),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1848),
.Y(n_1876)
);

INVx2_ASAP7_75t_SL g1877 ( 
.A(n_1870),
.Y(n_1877)
);

OAI21xp5_ASAP7_75t_L g1878 ( 
.A1(n_1868),
.A2(n_1857),
.B(n_1861),
.Y(n_1878)
);

AOI21xp5_ASAP7_75t_L g1879 ( 
.A1(n_1871),
.A2(n_1858),
.B(n_1861),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1866),
.B(n_1849),
.Y(n_1880)
);

AND2x2_ASAP7_75t_L g1881 ( 
.A(n_1869),
.B(n_1863),
.Y(n_1881)
);

OA33x2_ASAP7_75t_L g1882 ( 
.A1(n_1867),
.A2(n_1858),
.A3(n_1860),
.B1(n_1859),
.B2(n_1864),
.B3(n_1707),
.Y(n_1882)
);

O2A1O1Ixp33_ASAP7_75t_L g1883 ( 
.A1(n_1872),
.A2(n_1860),
.B(n_1756),
.C(n_1766),
.Y(n_1883)
);

NAND3xp33_ASAP7_75t_SL g1884 ( 
.A(n_1874),
.B(n_1813),
.C(n_1803),
.Y(n_1884)
);

AOI22xp33_ASAP7_75t_L g1885 ( 
.A1(n_1875),
.A2(n_1813),
.B1(n_1763),
.B2(n_1766),
.Y(n_1885)
);

OAI221xp5_ASAP7_75t_L g1886 ( 
.A1(n_1865),
.A2(n_1763),
.B1(n_1785),
.B2(n_1781),
.C(n_1722),
.Y(n_1886)
);

NAND4xp25_ASAP7_75t_L g1887 ( 
.A(n_1878),
.B(n_1876),
.C(n_1873),
.D(n_1771),
.Y(n_1887)
);

AOI211x1_ASAP7_75t_L g1888 ( 
.A1(n_1879),
.A2(n_1771),
.B(n_1762),
.C(n_1735),
.Y(n_1888)
);

AOI22xp5_ASAP7_75t_L g1889 ( 
.A1(n_1884),
.A2(n_1722),
.B1(n_1716),
.B2(n_1659),
.Y(n_1889)
);

NOR3xp33_ASAP7_75t_L g1890 ( 
.A(n_1880),
.B(n_1722),
.C(n_1774),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1877),
.Y(n_1891)
);

NOR2xp33_ASAP7_75t_L g1892 ( 
.A(n_1887),
.B(n_1881),
.Y(n_1892)
);

NOR3xp33_ASAP7_75t_L g1893 ( 
.A(n_1891),
.B(n_1883),
.C(n_1886),
.Y(n_1893)
);

AOI211x1_ASAP7_75t_L g1894 ( 
.A1(n_1888),
.A2(n_1882),
.B(n_1885),
.C(n_1716),
.Y(n_1894)
);

NOR3xp33_ASAP7_75t_SL g1895 ( 
.A(n_1890),
.B(n_1627),
.C(n_1637),
.Y(n_1895)
);

OAI21xp5_ASAP7_75t_SL g1896 ( 
.A1(n_1889),
.A2(n_1660),
.B(n_1662),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_SL g1897 ( 
.A(n_1891),
.B(n_1774),
.Y(n_1897)
);

OAI22xp5_ASAP7_75t_SL g1898 ( 
.A1(n_1892),
.A2(n_1622),
.B1(n_1497),
.B2(n_1627),
.Y(n_1898)
);

AOI22x1_ASAP7_75t_L g1899 ( 
.A1(n_1893),
.A2(n_1897),
.B1(n_1894),
.B2(n_1895),
.Y(n_1899)
);

AND2x2_ASAP7_75t_L g1900 ( 
.A(n_1896),
.B(n_1708),
.Y(n_1900)
);

OAI211xp5_ASAP7_75t_SL g1901 ( 
.A1(n_1892),
.A2(n_1637),
.B(n_1649),
.C(n_1631),
.Y(n_1901)
);

NAND3xp33_ASAP7_75t_SL g1902 ( 
.A(n_1893),
.B(n_1716),
.C(n_1727),
.Y(n_1902)
);

AND2x4_ASAP7_75t_L g1903 ( 
.A(n_1900),
.B(n_1727),
.Y(n_1903)
);

AOI22xp5_ASAP7_75t_L g1904 ( 
.A1(n_1902),
.A2(n_1898),
.B1(n_1901),
.B2(n_1899),
.Y(n_1904)
);

AND2x2_ASAP7_75t_L g1905 ( 
.A(n_1900),
.B(n_1708),
.Y(n_1905)
);

AOI22xp5_ASAP7_75t_L g1906 ( 
.A1(n_1903),
.A2(n_1714),
.B1(n_1662),
.B2(n_1660),
.Y(n_1906)
);

HB1xp67_ASAP7_75t_L g1907 ( 
.A(n_1906),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1907),
.B(n_1904),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1907),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1909),
.Y(n_1910)
);

INVx2_ASAP7_75t_L g1911 ( 
.A(n_1908),
.Y(n_1911)
);

AOI22xp5_ASAP7_75t_L g1912 ( 
.A1(n_1910),
.A2(n_1905),
.B1(n_1662),
.B2(n_1660),
.Y(n_1912)
);

OAI22xp5_ASAP7_75t_SL g1913 ( 
.A1(n_1911),
.A2(n_1649),
.B1(n_1631),
.B2(n_1644),
.Y(n_1913)
);

INVx2_ASAP7_75t_L g1914 ( 
.A(n_1912),
.Y(n_1914)
);

OAI22xp5_ASAP7_75t_SL g1915 ( 
.A1(n_1914),
.A2(n_1913),
.B1(n_1649),
.B2(n_1624),
.Y(n_1915)
);

AND2x4_ASAP7_75t_L g1916 ( 
.A(n_1915),
.B(n_1659),
.Y(n_1916)
);

OAI21x1_ASAP7_75t_SL g1917 ( 
.A1(n_1916),
.A2(n_1630),
.B(n_1632),
.Y(n_1917)
);

AOI22xp33_ASAP7_75t_L g1918 ( 
.A1(n_1917),
.A2(n_1659),
.B1(n_1646),
.B2(n_1643),
.Y(n_1918)
);

OAI22xp5_ASAP7_75t_L g1919 ( 
.A1(n_1918),
.A2(n_1644),
.B1(n_1646),
.B2(n_1643),
.Y(n_1919)
);

AOI211xp5_ASAP7_75t_L g1920 ( 
.A1(n_1919),
.A2(n_1624),
.B(n_1636),
.C(n_1635),
.Y(n_1920)
);


endmodule