module fake_jpeg_3342_n_178 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_178);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_178;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_37),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_28),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_1),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_9),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_30),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_11),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

BUFx10_ASAP7_75t_L g63 ( 
.A(n_4),
.Y(n_63)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_2),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_7),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_31),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_26),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_17),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_73),
.Y(n_78)
);

BUFx24_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

NAND2xp67_ASAP7_75t_L g80 ( 
.A(n_74),
.B(n_77),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_76),
.B(n_56),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_75),
.A2(n_53),
.B1(n_49),
.B2(n_59),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_79),
.A2(n_63),
.B1(n_68),
.B2(n_51),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_77),
.A2(n_53),
.B1(n_65),
.B2(n_54),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_81),
.A2(n_86),
.B1(n_87),
.B2(n_74),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_61),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_88),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_72),
.A2(n_64),
.B1(n_55),
.B2(n_66),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_71),
.A2(n_64),
.B1(n_66),
.B2(n_52),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_74),
.B(n_69),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_85),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

CKINVDCx5p33_ASAP7_75t_R g92 ( 
.A(n_84),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_100),
.Y(n_107)
);

A2O1A1Ixp33_ASAP7_75t_L g93 ( 
.A1(n_89),
.A2(n_50),
.B(n_60),
.C(n_67),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_93),
.B(n_97),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_102),
.Y(n_113)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_95),
.Y(n_120)
);

BUFx2_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_96),
.Y(n_116)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_84),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_98),
.B(n_99),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_84),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_101),
.A2(n_51),
.B1(n_63),
.B2(n_48),
.Y(n_109)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_104),
.B(n_5),
.Y(n_118)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_105),
.B(n_22),
.Y(n_110)
);

OA22x2_ASAP7_75t_L g108 ( 
.A1(n_102),
.A2(n_76),
.B1(n_63),
.B2(n_57),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_108),
.B(n_118),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_109),
.A2(n_111),
.B1(n_10),
.B2(n_12),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_110),
.B(n_117),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_101),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_SL g115 ( 
.A(n_94),
.B(n_24),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_SL g123 ( 
.A(n_115),
.B(n_8),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_103),
.B(n_3),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_90),
.B(n_5),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_91),
.A2(n_6),
.B(n_7),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_121),
.B(n_122),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_96),
.B(n_6),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_123),
.B(n_127),
.Y(n_143)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_120),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_125),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_115),
.B(n_32),
.Y(n_125)
);

OAI21xp33_ASAP7_75t_L g126 ( 
.A1(n_107),
.A2(n_8),
.B(n_10),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_126),
.B(n_130),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_114),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_113),
.A2(n_105),
.B1(n_12),
.B2(n_13),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_128),
.B(n_131),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_113),
.A2(n_118),
.B1(n_112),
.B2(n_111),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_116),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_132),
.B(n_133),
.Y(n_144)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_116),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_108),
.B(n_33),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_135),
.B(n_138),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_108),
.B(n_13),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_136),
.B(n_27),
.Y(n_149)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_106),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_106),
.B(n_14),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_139),
.B(n_140),
.Y(n_151)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_120),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_119),
.B(n_15),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_141),
.B(n_16),
.C(n_18),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_134),
.A2(n_20),
.B1(n_21),
.B2(n_25),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_146),
.A2(n_153),
.B1(n_139),
.B2(n_39),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_137),
.Y(n_147)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_147),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_149),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_134),
.A2(n_47),
.B(n_34),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_152),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_135),
.A2(n_29),
.B(n_36),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_129),
.B(n_125),
.Y(n_154)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_154),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_157),
.B(n_45),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_155),
.A2(n_38),
.B1(n_42),
.B2(n_43),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_160),
.A2(n_146),
.B1(n_153),
.B2(n_148),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_143),
.B(n_44),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_145),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_163),
.A2(n_167),
.B1(n_159),
.B2(n_158),
.Y(n_171)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_164),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_165),
.Y(n_169)
);

OR2x2_ASAP7_75t_L g166 ( 
.A(n_156),
.B(n_142),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_166),
.A2(n_144),
.B(n_150),
.Y(n_170)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_161),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_170),
.A2(n_171),
.B1(n_168),
.B2(n_152),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_172),
.B(n_173),
.Y(n_174)
);

BUFx24_ASAP7_75t_SL g173 ( 
.A(n_169),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_174),
.B(n_151),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_175),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_176),
.A2(n_163),
.B(n_158),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_150),
.Y(n_178)
);


endmodule