module fake_jpeg_31142_n_139 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_139);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_139;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

BUFx12_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_0),
.B(n_9),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_3),
.B(n_2),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_18),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_29),
.B(n_35),
.Y(n_52)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_0),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_36),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_18),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_16),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_15),
.B(n_1),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_39),
.Y(n_61)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_17),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_20),
.B(n_5),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_43),
.Y(n_59)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_22),
.B(n_6),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_31),
.A2(n_23),
.B1(n_25),
.B2(n_19),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_48),
.A2(n_57),
.B1(n_63),
.B2(n_33),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_37),
.B(n_26),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_60),
.Y(n_69)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_17),
.C(n_23),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_50),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_41),
.A2(n_2),
.B1(n_7),
.B2(n_8),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_39),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_32),
.A2(n_25),
.B1(n_14),
.B2(n_21),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_29),
.B(n_14),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_14),
.Y(n_79)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_64),
.Y(n_66)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_35),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_74),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_71),
.A2(n_83),
.B1(n_44),
.B2(n_58),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_72),
.B(n_75),
.Y(n_85)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_73),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_61),
.A2(n_42),
.B(n_25),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_50),
.B(n_41),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_78),
.B(n_79),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_44),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_80),
.B(n_62),
.Y(n_89)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_82),
.Y(n_90)
);

AND2x6_ASAP7_75t_L g82 ( 
.A(n_61),
.B(n_21),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_61),
.A2(n_57),
.B(n_62),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_87),
.B(n_47),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_75),
.Y(n_100)
);

BUFx8_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_93),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_83),
.A2(n_58),
.B1(n_45),
.B2(n_55),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_94),
.A2(n_96),
.B1(n_82),
.B2(n_70),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_69),
.B(n_59),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_95),
.B(n_68),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_67),
.A2(n_75),
.B1(n_72),
.B2(n_80),
.Y(n_96)
);

OA21x2_ASAP7_75t_L g98 ( 
.A1(n_90),
.A2(n_76),
.B(n_74),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_98),
.A2(n_88),
.B(n_92),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_86),
.B(n_72),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_100),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_92),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_101),
.Y(n_111)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_97),
.Y(n_102)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_102),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_103),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_105),
.A2(n_107),
.B1(n_87),
.B2(n_94),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_84),
.B(n_81),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_106),
.Y(n_115)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_108),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_85),
.B(n_66),
.C(n_45),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_109),
.B(n_88),
.C(n_91),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_SL g119 ( 
.A(n_116),
.B(n_118),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_117),
.A2(n_105),
.B(n_107),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_118),
.B(n_109),
.C(n_100),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_120),
.B(n_121),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_114),
.B(n_98),
.Y(n_122)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_122),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_112),
.B(n_98),
.C(n_91),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_123),
.B(n_125),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_111),
.Y(n_124)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_124),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_117),
.A2(n_104),
.B1(n_47),
.B2(n_55),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_119),
.A2(n_115),
.B1(n_113),
.B2(n_110),
.Y(n_127)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_127),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_126),
.B(n_125),
.C(n_113),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_131),
.B(n_133),
.Y(n_134)
);

AOI31xp67_ASAP7_75t_L g133 ( 
.A1(n_129),
.A2(n_110),
.A3(n_104),
.B(n_93),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_132),
.A2(n_130),
.B1(n_128),
.B2(n_126),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_128),
.C(n_93),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_134),
.C(n_56),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_137),
.A2(n_56),
.B1(n_21),
.B2(n_10),
.Y(n_138)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_138),
.Y(n_139)
);


endmodule