module fake_jpeg_31972_n_545 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_545);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_545;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_417;
wire n_362;
wire n_142;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_17),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_17),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_16),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_9),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_12),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_15),
.Y(n_50)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_53),
.Y(n_116)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_54),
.Y(n_115)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

INVx8_ASAP7_75t_L g141 ( 
.A(n_55),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_56),
.Y(n_113)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_57),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_58),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_59),
.Y(n_121)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_60),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_31),
.B(n_15),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_61),
.B(n_62),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g62 ( 
.A(n_21),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_63),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_64),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_65),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_31),
.B(n_14),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_66),
.B(n_80),
.Y(n_110)
);

BUFx24_ASAP7_75t_L g67 ( 
.A(n_28),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g134 ( 
.A(n_67),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_14),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_68),
.B(n_70),
.Y(n_129)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_18),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_69),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_50),
.B(n_0),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_71),
.Y(n_117)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_18),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_72),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_21),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_73),
.B(n_83),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_74),
.Y(n_124)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_34),
.Y(n_75)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_75),
.Y(n_161)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_34),
.Y(n_76)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_76),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_77),
.Y(n_126)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_36),
.Y(n_78)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_78),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_79),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_28),
.B(n_0),
.Y(n_80)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_27),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_81),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_82),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_46),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_84),
.Y(n_166)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_20),
.Y(n_85)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_85),
.Y(n_163)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_25),
.Y(n_86)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_86),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_27),
.Y(n_87)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_87),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_88),
.Y(n_171)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_29),
.Y(n_89)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_89),
.Y(n_142)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_25),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_90),
.B(n_92),
.Y(n_147)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_91),
.Y(n_167)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_27),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_93),
.B(n_94),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_46),
.Y(n_94)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_29),
.Y(n_95)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_95),
.Y(n_174)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_26),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_96),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_26),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_97),
.B(n_100),
.Y(n_157)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_52),
.Y(n_98)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_29),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_99),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_19),
.B(n_0),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_101),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_44),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_102),
.Y(n_145)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_26),
.Y(n_103)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_103),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_19),
.B(n_0),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_104),
.B(n_105),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_28),
.B(n_1),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_24),
.Y(n_106)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_106),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_44),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_107),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_41),
.Y(n_108)
);

INVx2_ASAP7_75t_SL g159 ( 
.A(n_108),
.Y(n_159)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_24),
.Y(n_109)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_109),
.Y(n_150)
);

BUFx12f_ASAP7_75t_L g111 ( 
.A(n_102),
.Y(n_111)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_111),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_98),
.A2(n_23),
.B1(n_33),
.B2(n_39),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_120),
.A2(n_170),
.B1(n_39),
.B2(n_33),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_57),
.A2(n_44),
.B1(n_51),
.B2(n_47),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_125),
.A2(n_64),
.B1(n_56),
.B2(n_74),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_60),
.B(n_23),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_130),
.B(n_172),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_96),
.B(n_45),
.C(n_41),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_143),
.B(n_149),
.C(n_32),
.Y(n_179)
);

AND2x4_ASAP7_75t_SL g149 ( 
.A(n_67),
.B(n_63),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_108),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_151),
.B(n_155),
.Y(n_221)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_75),
.Y(n_154)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_154),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_87),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_76),
.Y(n_156)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_156),
.Y(n_197)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_77),
.Y(n_160)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_160),
.Y(n_208)
);

BUFx12f_ASAP7_75t_L g162 ( 
.A(n_107),
.Y(n_162)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_162),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_67),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_164),
.B(n_51),
.Y(n_224)
);

BUFx12f_ASAP7_75t_L g168 ( 
.A(n_79),
.Y(n_168)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_168),
.Y(n_214)
);

OAI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_82),
.A2(n_41),
.B1(n_47),
.B2(n_37),
.Y(n_170)
);

NAND2x1_ASAP7_75t_SL g172 ( 
.A(n_93),
.B(n_22),
.Y(n_172)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_115),
.Y(n_175)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_175),
.Y(n_243)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_148),
.Y(n_176)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_176),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_131),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_177),
.B(n_186),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_113),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_178),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_179),
.B(n_202),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_112),
.B(n_91),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_180),
.B(n_189),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_126),
.A2(n_88),
.B1(n_84),
.B2(n_58),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g248 ( 
.A1(n_181),
.A2(n_184),
.B1(n_227),
.B2(n_124),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_113),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_182),
.Y(n_271)
);

INVx5_ASAP7_75t_L g183 ( 
.A(n_136),
.Y(n_183)
);

INVx5_ASAP7_75t_L g266 ( 
.A(n_183),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_131),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_119),
.Y(n_187)
);

BUFx2_ASAP7_75t_L g272 ( 
.A(n_187),
.Y(n_272)
);

A2O1A1Ixp33_ASAP7_75t_L g188 ( 
.A1(n_110),
.A2(n_37),
.B(n_35),
.C(n_32),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_188),
.B(n_190),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_112),
.B(n_40),
.Y(n_189)
);

A2O1A1Ixp33_ASAP7_75t_L g190 ( 
.A1(n_139),
.A2(n_35),
.B(n_40),
.C(n_93),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_172),
.A2(n_55),
.B1(n_69),
.B2(n_81),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_191),
.A2(n_194),
.B1(n_216),
.B2(n_226),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_157),
.B(n_42),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_192),
.B(n_210),
.Y(n_242)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_119),
.Y(n_193)
);

BUFx2_ASAP7_75t_L g281 ( 
.A(n_193),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_169),
.A2(n_72),
.B1(n_42),
.B2(n_22),
.Y(n_194)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_116),
.Y(n_195)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_195),
.Y(n_252)
);

INVx6_ASAP7_75t_L g196 ( 
.A(n_121),
.Y(n_196)
);

INVx6_ASAP7_75t_L g276 ( 
.A(n_196),
.Y(n_276)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_140),
.Y(n_199)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_199),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_129),
.B(n_22),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_201),
.B(n_229),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_134),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_121),
.Y(n_203)
);

BUFx5_ASAP7_75t_L g262 ( 
.A(n_203),
.Y(n_262)
);

INVx11_ASAP7_75t_L g204 ( 
.A(n_144),
.Y(n_204)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_204),
.Y(n_277)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_158),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_205),
.Y(n_239)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_150),
.Y(n_206)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_206),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_207),
.B(n_235),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_130),
.A2(n_59),
.B1(n_65),
.B2(n_89),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_209),
.B(n_170),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_157),
.B(n_42),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_118),
.Y(n_211)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_211),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_122),
.Y(n_213)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_213),
.Y(n_256)
);

INVx6_ASAP7_75t_L g215 ( 
.A(n_122),
.Y(n_215)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_215),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_141),
.A2(n_53),
.B1(n_95),
.B2(n_99),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_163),
.Y(n_217)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_217),
.Y(n_275)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_117),
.Y(n_218)
);

CKINVDCx14_ASAP7_75t_R g249 ( 
.A(n_218),
.Y(n_249)
);

INVx11_ASAP7_75t_L g219 ( 
.A(n_145),
.Y(n_219)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_219),
.Y(n_279)
);

BUFx12f_ASAP7_75t_L g220 ( 
.A(n_137),
.Y(n_220)
);

CKINVDCx14_ASAP7_75t_R g263 ( 
.A(n_220),
.Y(n_263)
);

INVx13_ASAP7_75t_L g222 ( 
.A(n_134),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_222),
.Y(n_280)
);

INVx2_ASAP7_75t_SL g223 ( 
.A(n_167),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_223),
.B(n_224),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_129),
.B(n_30),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_225),
.B(n_228),
.Y(n_268)
);

INVx8_ASAP7_75t_L g226 ( 
.A(n_138),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g227 ( 
.A1(n_126),
.A2(n_53),
.B1(n_51),
.B2(n_30),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_135),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_147),
.B(n_1),
.Y(n_229)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_132),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_230),
.B(n_232),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_147),
.B(n_1),
.Y(n_231)
);

NAND3xp33_ASAP7_75t_L g253 ( 
.A(n_231),
.B(n_233),
.C(n_1),
.Y(n_253)
);

INVx6_ASAP7_75t_L g232 ( 
.A(n_123),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_173),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_128),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_234),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_123),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_198),
.B(n_153),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_236),
.B(n_265),
.C(n_159),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_202),
.B(n_149),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_245),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_191),
.B(n_153),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_246),
.A2(n_267),
.B(n_270),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_248),
.B(n_253),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_255),
.A2(n_282),
.B1(n_171),
.B2(n_146),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_221),
.B(n_114),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_259),
.B(n_260),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_188),
.B(n_114),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_190),
.B(n_133),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_185),
.B(n_133),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_197),
.B(n_165),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_208),
.B(n_124),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_274),
.B(n_278),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_205),
.B(n_127),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_L g282 ( 
.A1(n_181),
.A2(n_171),
.B1(n_166),
.B2(n_127),
.Y(n_282)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_252),
.Y(n_284)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_284),
.Y(n_340)
);

AND2x6_ASAP7_75t_L g285 ( 
.A(n_246),
.B(n_222),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_285),
.B(n_288),
.Y(n_332)
);

INVx13_ASAP7_75t_L g286 ( 
.A(n_252),
.Y(n_286)
);

BUFx6f_ASAP7_75t_SL g344 ( 
.A(n_286),
.Y(n_344)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_262),
.Y(n_287)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_287),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_238),
.B(n_223),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_289),
.A2(n_290),
.B1(n_273),
.B2(n_215),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_241),
.A2(n_146),
.B1(n_166),
.B2(n_226),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g291 ( 
.A(n_262),
.Y(n_291)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_291),
.Y(n_331)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_274),
.Y(n_292)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_292),
.Y(n_338)
);

AOI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_250),
.A2(n_183),
.B1(n_220),
.B2(n_174),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_293),
.Y(n_351)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_278),
.Y(n_294)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_294),
.Y(n_339)
);

NAND3xp33_ASAP7_75t_L g297 ( 
.A(n_283),
.B(n_2),
.C(n_3),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_297),
.B(n_302),
.Y(n_348)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_258),
.Y(n_298)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_298),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_246),
.A2(n_194),
.B(n_216),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_300),
.A2(n_311),
.B(n_314),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_259),
.B(n_195),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_237),
.B(n_230),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_303),
.B(n_306),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_304),
.B(n_323),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_260),
.B(n_193),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_305),
.B(n_308),
.Y(n_324)
);

AND2x6_ASAP7_75t_L g306 ( 
.A(n_236),
.B(n_227),
.Y(n_306)
);

INVx6_ASAP7_75t_SL g307 ( 
.A(n_254),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_307),
.B(n_316),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_265),
.B(n_232),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_243),
.Y(n_309)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_309),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_261),
.B(n_161),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_310),
.Y(n_325)
);

OR2x2_ASAP7_75t_SL g311 ( 
.A(n_264),
.B(n_125),
.Y(n_311)
);

INVx11_ASAP7_75t_L g312 ( 
.A(n_266),
.Y(n_312)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_312),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_268),
.B(n_212),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g335 ( 
.A(n_313),
.B(n_315),
.Y(n_335)
);

AND2x6_ASAP7_75t_L g314 ( 
.A(n_240),
.B(n_242),
.Y(n_314)
);

AND2x6_ASAP7_75t_L g315 ( 
.A(n_240),
.B(n_159),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_251),
.Y(n_316)
);

INVx4_ASAP7_75t_L g317 ( 
.A(n_254),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_317),
.B(n_318),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_240),
.B(n_196),
.Y(n_318)
);

BUFx12f_ASAP7_75t_L g320 ( 
.A(n_271),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_320),
.B(n_322),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_247),
.B(n_275),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g341 ( 
.A(n_321),
.B(n_269),
.Y(n_341)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_273),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_245),
.A2(n_214),
.B(n_200),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_294),
.A2(n_241),
.B1(n_245),
.B2(n_255),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_326),
.A2(n_311),
.B1(n_292),
.B2(n_299),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_295),
.A2(n_241),
.B(n_267),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g361 ( 
.A1(n_328),
.A2(n_319),
.B(n_324),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_304),
.B(n_267),
.C(n_244),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_330),
.B(n_342),
.C(n_343),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_333),
.A2(n_337),
.B1(n_272),
.B2(n_281),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_295),
.A2(n_256),
.B1(n_276),
.B2(n_182),
.Y(n_337)
);

CKINVDCx14_ASAP7_75t_R g358 ( 
.A(n_341),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_308),
.B(n_239),
.C(n_270),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_318),
.B(n_270),
.C(n_257),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_296),
.B(n_249),
.C(n_280),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_345),
.B(n_346),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_296),
.B(n_280),
.C(n_263),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_299),
.B(n_256),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_350),
.B(n_298),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_314),
.B(n_279),
.C(n_276),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_354),
.B(n_285),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_319),
.B(n_279),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_356),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_341),
.B(n_305),
.Y(n_359)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_359),
.Y(n_394)
);

AND2x6_ASAP7_75t_L g360 ( 
.A(n_334),
.B(n_315),
.Y(n_360)
);

AO22x1_ASAP7_75t_L g417 ( 
.A1(n_360),
.A2(n_389),
.B1(n_336),
.B2(n_329),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_361),
.A2(n_335),
.B(n_326),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_362),
.A2(n_366),
.B1(n_370),
.B2(n_343),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_325),
.B(n_316),
.Y(n_363)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_363),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_325),
.B(n_352),
.Y(n_364)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_364),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_328),
.B(n_300),
.Y(n_365)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_365),
.A2(n_371),
.B(n_384),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_349),
.A2(n_289),
.B1(n_306),
.B2(n_301),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_SL g367 ( 
.A(n_348),
.B(n_323),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_367),
.B(n_369),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_339),
.A2(n_290),
.B1(n_307),
.B2(n_322),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_332),
.A2(n_287),
.B(n_284),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_372),
.B(n_387),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_350),
.B(n_317),
.Y(n_373)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_373),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_324),
.B(n_281),
.Y(n_374)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_374),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_SL g375 ( 
.A(n_338),
.B(n_312),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_375),
.B(n_388),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_338),
.B(n_320),
.Y(n_376)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_376),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_339),
.B(n_320),
.Y(n_377)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_377),
.Y(n_419)
);

INVx13_ASAP7_75t_L g378 ( 
.A(n_344),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_378),
.B(n_383),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_352),
.B(n_286),
.Y(n_380)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_380),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_381),
.A2(n_353),
.B1(n_340),
.B2(n_266),
.Y(n_420)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_347),
.Y(n_382)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_382),
.Y(n_412)
);

INVxp67_ASAP7_75t_SL g383 ( 
.A(n_344),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_351),
.A2(n_214),
.B1(n_277),
.B2(n_200),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_336),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_385),
.B(n_357),
.Y(n_409)
);

OAI21xp33_ASAP7_75t_L g386 ( 
.A1(n_335),
.A2(n_320),
.B(n_220),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_386),
.A2(n_357),
.B1(n_337),
.B2(n_329),
.Y(n_407)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_347),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_327),
.B(n_272),
.Y(n_388)
);

XNOR2x2_ASAP7_75t_SL g389 ( 
.A(n_334),
.B(n_327),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_379),
.B(n_355),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_391),
.B(n_396),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_L g393 ( 
.A1(n_365),
.A2(n_351),
.B(n_354),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g428 ( 
.A1(n_393),
.A2(n_404),
.B(n_411),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_379),
.B(n_355),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_390),
.B(n_356),
.C(n_330),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_397),
.B(n_398),
.C(n_406),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_361),
.B(n_365),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_369),
.B(n_342),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_407),
.B(n_420),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_409),
.Y(n_433)
);

AOI21xp5_ASAP7_75t_L g411 ( 
.A1(n_371),
.A2(n_357),
.B(n_331),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_413),
.A2(n_418),
.B1(n_381),
.B2(n_374),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_364),
.B(n_331),
.Y(n_414)
);

CKINVDCx16_ASAP7_75t_R g430 ( 
.A(n_414),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_368),
.B(n_345),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_415),
.B(n_416),
.C(n_363),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_368),
.B(n_346),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_417),
.B(n_362),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_366),
.A2(n_353),
.B1(n_340),
.B2(n_271),
.Y(n_418)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_403),
.Y(n_423)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_423),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_402),
.B(n_372),
.Y(n_424)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_424),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_425),
.A2(n_432),
.B1(n_440),
.B2(n_448),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_426),
.B(n_439),
.Y(n_449)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_403),
.Y(n_427)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_427),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_431),
.B(n_397),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_413),
.A2(n_385),
.B1(n_389),
.B2(n_373),
.Y(n_432)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_421),
.Y(n_435)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_435),
.Y(n_467)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_412),
.Y(n_436)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_436),
.Y(n_470)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_405),
.Y(n_437)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_437),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_391),
.B(n_389),
.C(n_359),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_438),
.B(n_441),
.C(n_416),
.Y(n_454)
);

AO22x1_ASAP7_75t_L g439 ( 
.A1(n_417),
.A2(n_360),
.B1(n_370),
.B2(n_388),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_417),
.A2(n_360),
.B1(n_358),
.B2(n_377),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_396),
.B(n_376),
.C(n_375),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_394),
.B(n_410),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_442),
.B(n_443),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_408),
.B(n_387),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_400),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_444),
.B(n_446),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_SL g445 ( 
.A(n_401),
.B(n_367),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g450 ( 
.A1(n_445),
.A2(n_404),
.B1(n_419),
.B2(n_399),
.Y(n_450)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_400),
.Y(n_446)
);

CKINVDCx16_ASAP7_75t_R g447 ( 
.A(n_419),
.Y(n_447)
);

CKINVDCx16_ASAP7_75t_R g466 ( 
.A(n_447),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_418),
.A2(n_384),
.B1(n_382),
.B2(n_380),
.Y(n_448)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_450),
.Y(n_472)
);

INVx3_ASAP7_75t_L g451 ( 
.A(n_433),
.Y(n_451)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_451),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_L g452 ( 
.A1(n_445),
.A2(n_435),
.B1(n_430),
.B2(n_433),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_452),
.B(n_453),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_L g453 ( 
.A1(n_439),
.A2(n_407),
.B1(n_392),
.B2(n_399),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_454),
.B(n_462),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_434),
.B(n_406),
.C(n_415),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_459),
.B(n_465),
.C(n_468),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_441),
.B(n_393),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_463),
.B(n_429),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_434),
.B(n_398),
.C(n_411),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_431),
.B(n_392),
.C(n_395),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_429),
.B(n_212),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_469),
.B(n_443),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_439),
.A2(n_422),
.B1(n_427),
.B2(n_423),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_471),
.A2(n_425),
.B1(n_448),
.B2(n_436),
.Y(n_482)
);

AOI21xp5_ASAP7_75t_SL g473 ( 
.A1(n_449),
.A2(n_428),
.B(n_446),
.Y(n_473)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_473),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_SL g475 ( 
.A1(n_461),
.A2(n_422),
.B1(n_424),
.B2(n_442),
.Y(n_475)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_475),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_476),
.B(n_482),
.Y(n_493)
);

A2O1A1O1Ixp25_ASAP7_75t_L g478 ( 
.A1(n_449),
.A2(n_438),
.B(n_440),
.C(n_428),
.D(n_432),
.Y(n_478)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_478),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_451),
.B(n_437),
.Y(n_479)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_479),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_480),
.B(n_487),
.Y(n_490)
);

AOI21xp5_ASAP7_75t_L g483 ( 
.A1(n_468),
.A2(n_277),
.B(n_378),
.Y(n_483)
);

AOI21xp5_ASAP7_75t_L g491 ( 
.A1(n_483),
.A2(n_457),
.B(n_456),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_471),
.A2(n_378),
.B1(n_235),
.B2(n_187),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_484),
.B(n_486),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_456),
.B(n_203),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_485),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_466),
.B(n_219),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_467),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_458),
.A2(n_213),
.B1(n_178),
.B2(n_204),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_489),
.B(n_470),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g513 ( 
.A(n_491),
.B(n_502),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_L g494 ( 
.A1(n_473),
.A2(n_461),
.B(n_455),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_SL g507 ( 
.A(n_494),
.B(n_503),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_488),
.B(n_454),
.C(n_469),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_498),
.B(n_501),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_SL g510 ( 
.A1(n_500),
.A2(n_482),
.B1(n_484),
.B2(n_457),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_489),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_477),
.B(n_465),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_477),
.B(n_462),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_488),
.B(n_463),
.C(n_459),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_504),
.B(n_474),
.Y(n_511)
);

CKINVDCx16_ASAP7_75t_R g506 ( 
.A(n_495),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_506),
.B(n_508),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_490),
.B(n_475),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_510),
.A2(n_505),
.B1(n_491),
.B2(n_499),
.Y(n_521)
);

OAI21xp5_ASAP7_75t_SL g526 ( 
.A1(n_511),
.A2(n_168),
.B(n_162),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_493),
.B(n_472),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_512),
.B(n_515),
.Y(n_527)
);

NOR2xp67_ASAP7_75t_SL g514 ( 
.A(n_492),
.B(n_478),
.Y(n_514)
);

AOI21xp5_ASAP7_75t_L g520 ( 
.A1(n_514),
.A2(n_517),
.B(n_502),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_493),
.B(n_487),
.Y(n_515)
);

AOI22xp33_ASAP7_75t_L g516 ( 
.A1(n_505),
.A2(n_464),
.B1(n_481),
.B2(n_460),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_L g525 ( 
.A1(n_516),
.A2(n_152),
.B1(n_142),
.B2(n_4),
.Y(n_525)
);

OAI21xp5_ASAP7_75t_SL g517 ( 
.A1(n_496),
.A2(n_504),
.B(n_498),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_SL g518 ( 
.A(n_503),
.B(n_460),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_518),
.B(n_494),
.C(n_497),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_509),
.B(n_496),
.Y(n_519)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_519),
.Y(n_531)
);

XOR2xp5_ASAP7_75t_L g529 ( 
.A(n_520),
.B(n_521),
.Y(n_529)
);

XNOR2x1_ASAP7_75t_L g532 ( 
.A(n_522),
.B(n_525),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_513),
.B(n_497),
.C(n_500),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_523),
.B(n_507),
.C(n_30),
.Y(n_534)
);

AOI322xp5_ASAP7_75t_L g533 ( 
.A1(n_526),
.A2(n_528),
.A3(n_30),
.B1(n_3),
.B2(n_4),
.C1(n_6),
.C2(n_8),
.Y(n_533)
);

OAI21xp5_ASAP7_75t_SL g528 ( 
.A1(n_516),
.A2(n_111),
.B(n_3),
.Y(n_528)
);

AOI322xp5_ASAP7_75t_L g530 ( 
.A1(n_519),
.A2(n_507),
.A3(n_518),
.B1(n_513),
.B2(n_5),
.C1(n_6),
.C2(n_7),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_SL g538 ( 
.A1(n_530),
.A2(n_533),
.B1(n_8),
.B2(n_9),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_534),
.B(n_524),
.C(n_527),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_535),
.B(n_537),
.Y(n_539)
);

O2A1O1Ixp33_ASAP7_75t_SL g536 ( 
.A1(n_529),
.A2(n_527),
.B(n_4),
.C(n_6),
.Y(n_536)
);

OR2x2_ASAP7_75t_L g540 ( 
.A(n_536),
.B(n_538),
.Y(n_540)
);

AOI21xp5_ASAP7_75t_L g537 ( 
.A1(n_531),
.A2(n_2),
.B(n_4),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_540),
.B(n_532),
.Y(n_541)
);

OAI21xp33_ASAP7_75t_L g542 ( 
.A1(n_541),
.A2(n_539),
.B(n_530),
.Y(n_542)
);

AOI22xp5_ASAP7_75t_L g543 ( 
.A1(n_542),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_543)
);

OAI21xp5_ASAP7_75t_L g544 ( 
.A1(n_543),
.A2(n_10),
.B(n_12),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_544),
.B(n_30),
.Y(n_545)
);


endmodule