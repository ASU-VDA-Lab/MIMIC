module real_aes_7199_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_766;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_746;
wire n_153;
wire n_316;
wire n_284;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_505;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_288;
wire n_147;
wire n_756;
wire n_150;
wire n_404;
wire n_598;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_749;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_753;
wire n_283;
wire n_314;
wire n_252;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_762;
wire n_210;
wire n_212;
wire n_325;
wire n_575;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_0), .A2(n_104), .B1(n_117), .B2(n_766), .Y(n_103) );
INVx1_ASAP7_75t_L g112 ( .A(n_1), .Y(n_112) );
INVx1_ASAP7_75t_L g502 ( .A(n_2), .Y(n_502) );
INVx1_ASAP7_75t_L g216 ( .A(n_3), .Y(n_216) );
AOI22xp5_ASAP7_75t_L g760 ( .A1(n_4), .A2(n_80), .B1(n_761), .B2(n_762), .Y(n_760) );
CKINVDCx20_ASAP7_75t_R g762 ( .A(n_4), .Y(n_762) );
AOI22xp33_ASAP7_75t_L g528 ( .A1(n_5), .A2(n_40), .B1(n_172), .B2(n_518), .Y(n_528) );
AOI21xp33_ASAP7_75t_L g196 ( .A1(n_6), .A2(n_153), .B(n_197), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_7), .B(n_146), .Y(n_493) );
AND2x6_ASAP7_75t_L g158 ( .A(n_8), .B(n_159), .Y(n_158) );
AOI21xp5_ASAP7_75t_L g254 ( .A1(n_9), .A2(n_255), .B(n_256), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_10), .B(n_41), .Y(n_109) );
NOR2xp33_ASAP7_75t_L g127 ( .A(n_10), .B(n_41), .Y(n_127) );
INVx1_ASAP7_75t_L g203 ( .A(n_11), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_12), .B(n_247), .Y(n_246) );
INVx1_ASAP7_75t_L g151 ( .A(n_13), .Y(n_151) );
INVx1_ASAP7_75t_L g497 ( .A(n_14), .Y(n_497) );
INVx1_ASAP7_75t_L g261 ( .A(n_15), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_16), .B(n_184), .Y(n_513) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_17), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_18), .B(n_147), .Y(n_474) );
AO32x2_ASAP7_75t_L g526 ( .A1(n_19), .A2(n_146), .A3(n_181), .B1(n_480), .B2(n_527), .Y(n_526) );
NAND2xp5_ASAP7_75t_SL g516 ( .A(n_20), .B(n_172), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_21), .B(n_167), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_22), .B(n_147), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_23), .A2(n_53), .B1(n_172), .B2(n_518), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_24), .B(n_153), .Y(n_227) );
AOI22xp33_ASAP7_75t_SL g524 ( .A1(n_25), .A2(n_77), .B1(n_172), .B2(n_184), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g539 ( .A(n_26), .B(n_172), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_27), .B(n_175), .Y(n_174) );
A2O1A1Ixp33_ASAP7_75t_L g258 ( .A1(n_28), .A2(n_259), .B(n_260), .C(n_262), .Y(n_258) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_29), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_30), .B(n_205), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_31), .B(n_201), .Y(n_218) );
AOI222xp33_ASAP7_75t_SL g129 ( .A1(n_32), .A2(n_130), .B1(n_136), .B2(n_744), .C1(n_745), .C2(n_750), .Y(n_129) );
OAI22xp5_ASAP7_75t_L g131 ( .A1(n_33), .A2(n_44), .B1(n_132), .B2(n_133), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g132 ( .A(n_33), .Y(n_132) );
INVx1_ASAP7_75t_L g190 ( .A(n_34), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_35), .B(n_205), .Y(n_541) );
INVx2_ASAP7_75t_L g156 ( .A(n_36), .Y(n_156) );
NAND2xp5_ASAP7_75t_SL g557 ( .A(n_37), .B(n_172), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_38), .B(n_205), .Y(n_519) );
A2O1A1Ixp33_ASAP7_75t_L g228 ( .A1(n_39), .A2(n_158), .B(n_162), .C(n_229), .Y(n_228) );
INVx1_ASAP7_75t_L g188 ( .A(n_42), .Y(n_188) );
NAND2xp5_ASAP7_75t_SL g271 ( .A(n_43), .B(n_201), .Y(n_271) );
CKINVDCx14_ASAP7_75t_R g133 ( .A(n_44), .Y(n_133) );
NAND2xp5_ASAP7_75t_SL g487 ( .A(n_45), .B(n_172), .Y(n_487) );
OAI22xp5_ASAP7_75t_SL g130 ( .A1(n_46), .A2(n_131), .B1(n_134), .B2(n_135), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g135 ( .A(n_46), .Y(n_135) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_47), .A2(n_88), .B1(n_234), .B2(n_518), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g490 ( .A(n_48), .B(n_172), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_49), .B(n_172), .Y(n_498) );
CKINVDCx16_ASAP7_75t_R g191 ( .A(n_50), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_51), .B(n_492), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_52), .B(n_153), .Y(n_249) );
AOI22xp33_ASAP7_75t_SL g479 ( .A1(n_54), .A2(n_63), .B1(n_172), .B2(n_184), .Y(n_479) );
AOI22xp5_ASAP7_75t_L g183 ( .A1(n_55), .A2(n_162), .B1(n_184), .B2(n_186), .Y(n_183) );
CKINVDCx20_ASAP7_75t_R g237 ( .A(n_56), .Y(n_237) );
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_57), .B(n_172), .Y(n_512) );
CKINVDCx16_ASAP7_75t_R g213 ( .A(n_58), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g561 ( .A(n_59), .B(n_172), .Y(n_561) );
A2O1A1Ixp33_ASAP7_75t_L g199 ( .A1(n_60), .A2(n_171), .B(n_200), .C(n_202), .Y(n_199) );
CKINVDCx20_ASAP7_75t_R g275 ( .A(n_61), .Y(n_275) );
INVx1_ASAP7_75t_L g198 ( .A(n_62), .Y(n_198) );
INVx1_ASAP7_75t_L g159 ( .A(n_64), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_65), .B(n_172), .Y(n_503) );
INVx1_ASAP7_75t_L g150 ( .A(n_66), .Y(n_150) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_67), .Y(n_121) );
AO32x2_ASAP7_75t_L g521 ( .A1(n_68), .A2(n_146), .A3(n_241), .B1(n_480), .B2(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g560 ( .A(n_69), .Y(n_560) );
INVx1_ASAP7_75t_L g536 ( .A(n_70), .Y(n_536) );
A2O1A1Ixp33_ASAP7_75t_SL g166 ( .A1(n_71), .A2(n_167), .B(n_168), .C(n_171), .Y(n_166) );
INVxp67_ASAP7_75t_L g169 ( .A(n_72), .Y(n_169) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_73), .B(n_184), .Y(n_537) );
INVx1_ASAP7_75t_L g116 ( .A(n_74), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g194 ( .A(n_75), .Y(n_194) );
INVx1_ASAP7_75t_L g268 ( .A(n_76), .Y(n_268) );
A2O1A1Ixp33_ASAP7_75t_L g269 ( .A1(n_78), .A2(n_158), .B(n_162), .C(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_79), .B(n_518), .Y(n_517) );
CKINVDCx20_ASAP7_75t_R g761 ( .A(n_80), .Y(n_761) );
NAND2xp5_ASAP7_75t_SL g540 ( .A(n_81), .B(n_184), .Y(n_540) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_82), .B(n_217), .Y(n_230) );
INVx2_ASAP7_75t_L g148 ( .A(n_83), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_84), .B(n_167), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_85), .B(n_184), .Y(n_488) );
A2O1A1Ixp33_ASAP7_75t_L g214 ( .A1(n_86), .A2(n_158), .B(n_162), .C(n_215), .Y(n_214) );
INVx2_ASAP7_75t_L g113 ( .A(n_87), .Y(n_113) );
OR2x2_ASAP7_75t_L g124 ( .A(n_87), .B(n_125), .Y(n_124) );
OR2x2_ASAP7_75t_L g465 ( .A(n_87), .B(n_126), .Y(n_465) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_89), .A2(n_102), .B1(n_184), .B2(n_185), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_90), .B(n_205), .Y(n_204) );
CKINVDCx20_ASAP7_75t_R g221 ( .A(n_91), .Y(n_221) );
A2O1A1Ixp33_ASAP7_75t_L g243 ( .A1(n_92), .A2(n_158), .B(n_162), .C(n_244), .Y(n_243) );
CKINVDCx20_ASAP7_75t_R g251 ( .A(n_93), .Y(n_251) );
INVx1_ASAP7_75t_L g165 ( .A(n_94), .Y(n_165) );
CKINVDCx16_ASAP7_75t_R g257 ( .A(n_95), .Y(n_257) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_96), .B(n_217), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_97), .B(n_184), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_98), .B(n_146), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_99), .B(n_116), .Y(n_115) );
AOI21xp5_ASAP7_75t_L g152 ( .A1(n_100), .A2(n_153), .B(n_160), .Y(n_152) );
OAI22xp5_ASAP7_75t_SL g758 ( .A1(n_101), .A2(n_759), .B1(n_760), .B2(n_763), .Y(n_758) );
CKINVDCx20_ASAP7_75t_R g763 ( .A(n_101), .Y(n_763) );
INVx1_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
CKINVDCx9p33_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g767 ( .A(n_107), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_108), .B(n_110), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
CKINVDCx14_ASAP7_75t_R g110 ( .A(n_111), .Y(n_110) );
NAND3xp33_ASAP7_75t_SL g111 ( .A(n_112), .B(n_113), .C(n_114), .Y(n_111) );
AND2x2_ASAP7_75t_L g126 ( .A(n_112), .B(n_127), .Y(n_126) );
OR2x2_ASAP7_75t_L g466 ( .A(n_113), .B(n_126), .Y(n_466) );
NOR2x2_ASAP7_75t_L g752 ( .A(n_113), .B(n_125), .Y(n_752) );
INVx1_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
AOI22x1_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_129), .B1(n_753), .B2(n_755), .Y(n_117) );
NOR2xp33_ASAP7_75t_L g118 ( .A(n_119), .B(n_122), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
BUFx2_ASAP7_75t_L g754 ( .A(n_120), .Y(n_754) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
AOI21xp5_ASAP7_75t_L g755 ( .A1(n_122), .A2(n_756), .B(n_764), .Y(n_755) );
NOR2xp33_ASAP7_75t_SL g122 ( .A(n_123), .B(n_128), .Y(n_122) );
HB1xp67_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx1_ASAP7_75t_SL g765 ( .A(n_124), .Y(n_765) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
CKINVDCx14_ASAP7_75t_R g744 ( .A(n_130), .Y(n_744) );
INVx1_ASAP7_75t_L g134 ( .A(n_131), .Y(n_134) );
OAI22x1_ASAP7_75t_SL g136 ( .A1(n_137), .A2(n_463), .B1(n_466), .B2(n_467), .Y(n_136) );
OAI22xp5_ASAP7_75t_L g756 ( .A1(n_137), .A2(n_138), .B1(n_757), .B2(n_758), .Y(n_756) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
OAI22xp5_ASAP7_75t_L g745 ( .A1(n_138), .A2(n_746), .B1(n_747), .B2(n_749), .Y(n_745) );
AND2x2_ASAP7_75t_SL g138 ( .A(n_139), .B(n_400), .Y(n_138) );
NOR4xp25_ASAP7_75t_L g139 ( .A(n_140), .B(n_330), .C(n_361), .D(n_380), .Y(n_139) );
NAND4xp25_ASAP7_75t_L g140 ( .A(n_141), .B(n_288), .C(n_303), .D(n_321), .Y(n_140) );
AOI222xp33_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_223), .B1(n_264), .B2(n_276), .C1(n_281), .C2(n_283), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_143), .B(n_206), .Y(n_142) );
INVx1_ASAP7_75t_L g344 ( .A(n_143), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_144), .B(n_177), .Y(n_143) );
AND2x2_ASAP7_75t_L g207 ( .A(n_144), .B(n_195), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_144), .B(n_210), .Y(n_373) );
INVx3_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
OR2x2_ASAP7_75t_L g280 ( .A(n_145), .B(n_179), .Y(n_280) );
AND2x2_ASAP7_75t_L g289 ( .A(n_145), .B(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g315 ( .A(n_145), .Y(n_315) );
AND2x2_ASAP7_75t_L g336 ( .A(n_145), .B(n_179), .Y(n_336) );
BUFx2_ASAP7_75t_L g359 ( .A(n_145), .Y(n_359) );
AND2x2_ASAP7_75t_L g383 ( .A(n_145), .B(n_180), .Y(n_383) );
AND2x2_ASAP7_75t_L g447 ( .A(n_145), .B(n_195), .Y(n_447) );
OA21x2_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_152), .B(n_174), .Y(n_145) );
INVx4_ASAP7_75t_L g176 ( .A(n_146), .Y(n_176) );
OA21x2_ASAP7_75t_L g484 ( .A1(n_146), .A2(n_485), .B(n_493), .Y(n_484) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx1_ASAP7_75t_L g181 ( .A(n_147), .Y(n_181) );
AND2x2_ASAP7_75t_L g147 ( .A(n_148), .B(n_149), .Y(n_147) );
AND2x2_ASAP7_75t_SL g205 ( .A(n_148), .B(n_149), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_150), .B(n_151), .Y(n_149) );
BUFx2_ASAP7_75t_L g255 ( .A(n_153), .Y(n_255) );
AND2x4_ASAP7_75t_L g153 ( .A(n_154), .B(n_158), .Y(n_153) );
NAND2x1p5_ASAP7_75t_L g192 ( .A(n_154), .B(n_158), .Y(n_192) );
AND2x2_ASAP7_75t_L g154 ( .A(n_155), .B(n_157), .Y(n_154) );
INVx1_ASAP7_75t_L g492 ( .A(n_155), .Y(n_492) );
INVx1_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx2_ASAP7_75t_L g163 ( .A(n_156), .Y(n_163) );
INVx1_ASAP7_75t_L g185 ( .A(n_156), .Y(n_185) );
INVx1_ASAP7_75t_L g164 ( .A(n_157), .Y(n_164) );
INVx1_ASAP7_75t_L g167 ( .A(n_157), .Y(n_167) );
INVx3_ASAP7_75t_L g170 ( .A(n_157), .Y(n_170) );
BUFx6f_ASAP7_75t_L g187 ( .A(n_157), .Y(n_187) );
BUFx6f_ASAP7_75t_L g201 ( .A(n_157), .Y(n_201) );
INVx4_ASAP7_75t_SL g173 ( .A(n_158), .Y(n_173) );
BUFx3_ASAP7_75t_L g480 ( .A(n_158), .Y(n_480) );
OAI21xp5_ASAP7_75t_L g485 ( .A1(n_158), .A2(n_486), .B(n_489), .Y(n_485) );
OAI21xp5_ASAP7_75t_L g495 ( .A1(n_158), .A2(n_496), .B(n_500), .Y(n_495) );
OAI21xp5_ASAP7_75t_L g510 ( .A1(n_158), .A2(n_511), .B(n_515), .Y(n_510) );
OAI21xp5_ASAP7_75t_L g534 ( .A1(n_158), .A2(n_535), .B(n_538), .Y(n_534) );
O2A1O1Ixp33_ASAP7_75t_L g160 ( .A1(n_161), .A2(n_165), .B(n_166), .C(n_173), .Y(n_160) );
O2A1O1Ixp33_ASAP7_75t_L g197 ( .A1(n_161), .A2(n_173), .B(n_198), .C(n_199), .Y(n_197) );
O2A1O1Ixp33_ASAP7_75t_L g256 ( .A1(n_161), .A2(n_173), .B(n_257), .C(n_258), .Y(n_256) );
INVx5_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
AND2x6_ASAP7_75t_L g162 ( .A(n_163), .B(n_164), .Y(n_162) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_163), .Y(n_172) );
BUFx3_ASAP7_75t_L g234 ( .A(n_163), .Y(n_234) );
INVx1_ASAP7_75t_L g518 ( .A(n_163), .Y(n_518) );
INVx1_ASAP7_75t_L g514 ( .A(n_167), .Y(n_514) );
NOR2xp33_ASAP7_75t_L g168 ( .A(n_169), .B(n_170), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_170), .B(n_203), .Y(n_202) );
INVx5_ASAP7_75t_L g217 ( .A(n_170), .Y(n_217) );
OAI22xp5_ASAP7_75t_SL g522 ( .A1(n_170), .A2(n_201), .B1(n_523), .B2(n_524), .Y(n_522) );
O2A1O1Ixp5_ASAP7_75t_SL g535 ( .A1(n_171), .A2(n_217), .B(n_536), .C(n_537), .Y(n_535) );
INVx3_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
HB1xp67_ASAP7_75t_L g248 ( .A(n_172), .Y(n_248) );
OAI22xp33_ASAP7_75t_L g182 ( .A1(n_173), .A2(n_183), .B1(n_191), .B2(n_192), .Y(n_182) );
OA21x2_ASAP7_75t_L g195 ( .A1(n_175), .A2(n_196), .B(n_204), .Y(n_195) );
INVx3_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
NOR2xp33_ASAP7_75t_SL g236 ( .A(n_176), .B(n_237), .Y(n_236) );
NAND3xp33_ASAP7_75t_L g475 ( .A(n_176), .B(n_476), .C(n_480), .Y(n_475) );
AO21x1_ASAP7_75t_L g568 ( .A1(n_176), .A2(n_476), .B(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g348 ( .A(n_177), .B(n_279), .Y(n_348) );
INVx1_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g372 ( .A(n_178), .B(n_373), .Y(n_372) );
OR2x2_ASAP7_75t_L g178 ( .A(n_179), .B(n_195), .Y(n_178) );
OR2x2_ASAP7_75t_L g308 ( .A(n_179), .B(n_211), .Y(n_308) );
AND2x2_ASAP7_75t_L g320 ( .A(n_179), .B(n_279), .Y(n_320) );
BUFx2_ASAP7_75t_L g452 ( .A(n_179), .Y(n_452) );
INVx3_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
OR2x2_ASAP7_75t_L g209 ( .A(n_180), .B(n_210), .Y(n_209) );
AND2x2_ASAP7_75t_L g302 ( .A(n_180), .B(n_211), .Y(n_302) );
AND2x2_ASAP7_75t_L g355 ( .A(n_180), .B(n_195), .Y(n_355) );
HB1xp67_ASAP7_75t_L g391 ( .A(n_180), .Y(n_391) );
AO21x2_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_182), .B(n_193), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_181), .B(n_194), .Y(n_193) );
AO21x2_ASAP7_75t_L g211 ( .A1(n_181), .A2(n_212), .B(n_220), .Y(n_211) );
INVx2_ASAP7_75t_L g235 ( .A(n_181), .Y(n_235) );
INVx2_ASAP7_75t_L g219 ( .A(n_184), .Y(n_219) );
INVx3_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
OAI22xp5_ASAP7_75t_SL g186 ( .A1(n_187), .A2(n_188), .B1(n_189), .B2(n_190), .Y(n_186) );
INVx2_ASAP7_75t_L g189 ( .A(n_187), .Y(n_189) );
INVx4_ASAP7_75t_L g259 ( .A(n_187), .Y(n_259) );
OAI21xp5_ASAP7_75t_L g212 ( .A1(n_192), .A2(n_213), .B(n_214), .Y(n_212) );
OAI21xp5_ASAP7_75t_L g267 ( .A1(n_192), .A2(n_268), .B(n_269), .Y(n_267) );
AND2x2_ASAP7_75t_L g278 ( .A(n_195), .B(n_279), .Y(n_278) );
INVx1_ASAP7_75t_SL g290 ( .A(n_195), .Y(n_290) );
INVx2_ASAP7_75t_L g301 ( .A(n_195), .Y(n_301) );
BUFx2_ASAP7_75t_L g325 ( .A(n_195), .Y(n_325) );
AND2x2_ASAP7_75t_SL g382 ( .A(n_195), .B(n_383), .Y(n_382) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_200), .A2(n_516), .B(n_517), .Y(n_515) );
O2A1O1Ixp5_ASAP7_75t_L g559 ( .A1(n_200), .A2(n_501), .B(n_560), .C(n_561), .Y(n_559) );
INVx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
INVx4_ASAP7_75t_L g247 ( .A(n_201), .Y(n_247) );
OAI22xp5_ASAP7_75t_L g476 ( .A1(n_201), .A2(n_477), .B1(n_478), .B2(n_479), .Y(n_476) );
OAI22xp5_ASAP7_75t_L g527 ( .A1(n_201), .A2(n_478), .B1(n_528), .B2(n_529), .Y(n_527) );
INVx1_ASAP7_75t_L g222 ( .A(n_205), .Y(n_222) );
INVx2_ASAP7_75t_L g241 ( .A(n_205), .Y(n_241) );
OA21x2_ASAP7_75t_L g253 ( .A1(n_205), .A2(n_254), .B(n_263), .Y(n_253) );
OA21x2_ASAP7_75t_L g509 ( .A1(n_205), .A2(n_510), .B(n_519), .Y(n_509) );
OA21x2_ASAP7_75t_L g533 ( .A1(n_205), .A2(n_534), .B(n_541), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_207), .B(n_208), .Y(n_206) );
AOI332xp33_ASAP7_75t_L g303 ( .A1(n_207), .A2(n_304), .A3(n_308), .B1(n_309), .B2(n_313), .B3(n_316), .C1(n_317), .C2(n_319), .Y(n_303) );
NAND2x1_ASAP7_75t_L g388 ( .A(n_207), .B(n_279), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_207), .B(n_293), .Y(n_439) );
A2O1A1Ixp33_ASAP7_75t_SL g321 ( .A1(n_208), .A2(n_322), .B(n_325), .C(n_326), .Y(n_321) );
AND2x2_ASAP7_75t_L g460 ( .A(n_208), .B(n_301), .Y(n_460) );
INVx3_ASAP7_75t_SL g208 ( .A(n_209), .Y(n_208) );
OR2x2_ASAP7_75t_L g357 ( .A(n_209), .B(n_358), .Y(n_357) );
OR2x2_ASAP7_75t_L g362 ( .A(n_209), .B(n_359), .Y(n_362) );
INVx1_ASAP7_75t_L g293 ( .A(n_210), .Y(n_293) );
AND2x2_ASAP7_75t_L g396 ( .A(n_210), .B(n_355), .Y(n_396) );
AND2x2_ASAP7_75t_L g397 ( .A(n_210), .B(n_336), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_210), .B(n_407), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_210), .B(n_314), .Y(n_422) );
INVx3_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
INVx3_ASAP7_75t_L g279 ( .A(n_211), .Y(n_279) );
O2A1O1Ixp33_ASAP7_75t_L g215 ( .A1(n_216), .A2(n_217), .B(n_218), .C(n_219), .Y(n_215) );
INVx2_ASAP7_75t_L g478 ( .A(n_217), .Y(n_478) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_217), .A2(n_487), .B(n_488), .Y(n_486) );
AOI21xp5_ASAP7_75t_L g556 ( .A1(n_217), .A2(n_557), .B(n_558), .Y(n_556) );
O2A1O1Ixp33_ASAP7_75t_L g496 ( .A1(n_219), .A2(n_497), .B(n_498), .C(n_499), .Y(n_496) );
NOR2xp33_ASAP7_75t_L g220 ( .A(n_221), .B(n_222), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g250 ( .A(n_222), .B(n_251), .Y(n_250) );
NOR2xp33_ASAP7_75t_L g274 ( .A(n_222), .B(n_275), .Y(n_274) );
OAI31xp33_ASAP7_75t_L g461 ( .A1(n_223), .A2(n_382), .A3(n_389), .B(n_462), .Y(n_461) );
AND2x2_ASAP7_75t_L g223 ( .A(n_224), .B(n_238), .Y(n_223) );
AND2x2_ASAP7_75t_L g264 ( .A(n_224), .B(n_265), .Y(n_264) );
NAND2x1_ASAP7_75t_SL g284 ( .A(n_224), .B(n_285), .Y(n_284) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_224), .Y(n_371) );
AND2x2_ASAP7_75t_L g376 ( .A(n_224), .B(n_287), .Y(n_376) );
INVx3_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
A2O1A1Ixp33_ASAP7_75t_L g288 ( .A1(n_225), .A2(n_289), .B(n_291), .C(n_294), .Y(n_288) );
OR2x2_ASAP7_75t_L g305 ( .A(n_225), .B(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g318 ( .A(n_225), .Y(n_318) );
AND2x2_ASAP7_75t_L g324 ( .A(n_225), .B(n_266), .Y(n_324) );
INVx2_ASAP7_75t_L g342 ( .A(n_225), .Y(n_342) );
AND2x2_ASAP7_75t_L g353 ( .A(n_225), .B(n_307), .Y(n_353) );
AND2x2_ASAP7_75t_L g385 ( .A(n_225), .B(n_343), .Y(n_385) );
AND2x2_ASAP7_75t_L g389 ( .A(n_225), .B(n_312), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_225), .B(n_238), .Y(n_394) );
AND2x2_ASAP7_75t_L g428 ( .A(n_225), .B(n_429), .Y(n_428) );
NOR2xp33_ASAP7_75t_L g462 ( .A(n_225), .B(n_331), .Y(n_462) );
OR2x6_ASAP7_75t_L g225 ( .A(n_226), .B(n_236), .Y(n_225) );
AOI21xp5_ASAP7_75t_SL g226 ( .A1(n_227), .A2(n_228), .B(n_235), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_231), .B(n_232), .Y(n_229) );
AOI21xp5_ASAP7_75t_L g270 ( .A1(n_232), .A2(n_271), .B(n_272), .Y(n_270) );
INVx2_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
INVx1_ASAP7_75t_L g262 ( .A(n_234), .Y(n_262) );
INVx1_ASAP7_75t_L g273 ( .A(n_235), .Y(n_273) );
OA21x2_ASAP7_75t_L g494 ( .A1(n_235), .A2(n_495), .B(n_504), .Y(n_494) );
OA21x2_ASAP7_75t_L g554 ( .A1(n_235), .A2(n_555), .B(n_562), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_238), .B(n_293), .Y(n_292) );
INVx1_ASAP7_75t_L g370 ( .A(n_238), .Y(n_370) );
AND2x2_ASAP7_75t_L g432 ( .A(n_238), .B(n_353), .Y(n_432) );
AND2x2_ASAP7_75t_L g238 ( .A(n_239), .B(n_252), .Y(n_238) );
OR2x2_ASAP7_75t_L g286 ( .A(n_239), .B(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g296 ( .A(n_239), .B(n_297), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_239), .B(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g404 ( .A(n_239), .Y(n_404) );
AND2x2_ASAP7_75t_L g421 ( .A(n_239), .B(n_266), .Y(n_421) );
INVx2_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_L g312 ( .A(n_240), .B(n_252), .Y(n_312) );
AND2x2_ASAP7_75t_L g341 ( .A(n_240), .B(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g352 ( .A(n_240), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_240), .B(n_307), .Y(n_443) );
AO21x2_ASAP7_75t_L g240 ( .A1(n_241), .A2(n_242), .B(n_250), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_243), .B(n_249), .Y(n_242) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_245), .A2(n_246), .B(n_248), .Y(n_244) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g265 ( .A(n_253), .B(n_266), .Y(n_265) );
INVx2_ASAP7_75t_L g287 ( .A(n_253), .Y(n_287) );
AND2x2_ASAP7_75t_L g343 ( .A(n_253), .B(n_307), .Y(n_343) );
NOR2xp33_ASAP7_75t_L g260 ( .A(n_259), .B(n_261), .Y(n_260) );
INVx1_ASAP7_75t_L g499 ( .A(n_259), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_259), .A2(n_539), .B(n_540), .Y(n_538) );
INVx1_ASAP7_75t_L g445 ( .A(n_264), .Y(n_445) );
INVx1_ASAP7_75t_L g449 ( .A(n_265), .Y(n_449) );
INVx2_ASAP7_75t_L g307 ( .A(n_266), .Y(n_307) );
AO21x2_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_273), .B(n_274), .Y(n_266) );
NOR2xp33_ASAP7_75t_L g276 ( .A(n_277), .B(n_280), .Y(n_276) );
INVx1_ASAP7_75t_SL g277 ( .A(n_278), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_278), .B(n_424), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_278), .B(n_383), .Y(n_441) );
OR2x2_ASAP7_75t_L g282 ( .A(n_279), .B(n_280), .Y(n_282) );
INVx1_ASAP7_75t_SL g334 ( .A(n_279), .Y(n_334) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AOI221xp5_ASAP7_75t_L g337 ( .A1(n_285), .A2(n_338), .B1(n_340), .B2(n_344), .C(n_345), .Y(n_337) );
INVx2_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
OR2x2_ASAP7_75t_L g365 ( .A(n_286), .B(n_329), .Y(n_365) );
INVx2_ASAP7_75t_L g297 ( .A(n_287), .Y(n_297) );
INVx1_ASAP7_75t_L g323 ( .A(n_287), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_287), .B(n_307), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_287), .B(n_310), .Y(n_417) );
INVx1_ASAP7_75t_L g425 ( .A(n_287), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_289), .B(n_293), .Y(n_339) );
AND2x4_ASAP7_75t_L g314 ( .A(n_290), .B(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g427 ( .A(n_293), .B(n_383), .Y(n_427) );
NOR2xp33_ASAP7_75t_L g294 ( .A(n_295), .B(n_298), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_296), .B(n_328), .Y(n_327) );
INVxp67_ASAP7_75t_L g435 ( .A(n_297), .Y(n_435) );
INVxp67_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_302), .Y(n_299) );
INVx1_ASAP7_75t_SL g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g335 ( .A(n_301), .B(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g407 ( .A(n_301), .B(n_383), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_301), .B(n_320), .Y(n_413) );
AOI322xp5_ASAP7_75t_L g367 ( .A1(n_302), .A2(n_336), .A3(n_343), .B1(n_368), .B2(n_371), .C1(n_372), .C2(n_374), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_302), .B(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
OR2x2_ASAP7_75t_L g433 ( .A(n_305), .B(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g379 ( .A(n_306), .Y(n_379) );
INVx2_ASAP7_75t_L g310 ( .A(n_307), .Y(n_310) );
INVx1_ASAP7_75t_L g369 ( .A(n_307), .Y(n_369) );
CKINVDCx16_ASAP7_75t_R g316 ( .A(n_308), .Y(n_316) );
NOR2xp33_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
AND2x2_ASAP7_75t_L g405 ( .A(n_310), .B(n_318), .Y(n_405) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g317 ( .A(n_312), .B(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g360 ( .A(n_312), .B(n_353), .Y(n_360) );
AND2x2_ASAP7_75t_L g364 ( .A(n_312), .B(n_324), .Y(n_364) );
OAI21xp33_ASAP7_75t_SL g374 ( .A1(n_313), .A2(n_375), .B(n_377), .Y(n_374) );
OAI22xp33_ASAP7_75t_L g444 ( .A1(n_313), .A2(n_445), .B1(n_446), .B2(n_448), .Y(n_444) );
INVx3_ASAP7_75t_SL g313 ( .A(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g319 ( .A(n_314), .B(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_314), .B(n_334), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_316), .B(n_454), .Y(n_453) );
AND2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
INVx1_ASAP7_75t_L g456 ( .A(n_323), .Y(n_456) );
INVx4_ASAP7_75t_L g329 ( .A(n_324), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_324), .B(n_351), .Y(n_399) );
INVx1_ASAP7_75t_SL g411 ( .A(n_325), .Y(n_411) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
NOR2xp67_ASAP7_75t_L g424 ( .A(n_329), .B(n_425), .Y(n_424) );
OAI211xp5_ASAP7_75t_SL g330 ( .A1(n_331), .A2(n_332), .B(n_337), .C(n_354), .Y(n_330) );
OAI221xp5_ASAP7_75t_SL g450 ( .A1(n_332), .A2(n_370), .B1(n_449), .B2(n_451), .C(n_453), .Y(n_450) );
INVx1_ASAP7_75t_SL g332 ( .A(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_334), .B(n_447), .Y(n_446) );
OAI31xp33_ASAP7_75t_L g426 ( .A1(n_335), .A2(n_412), .A3(n_427), .B(n_428), .Y(n_426) );
INVx1_ASAP7_75t_L g366 ( .A(n_336), .Y(n_366) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g340 ( .A(n_341), .B(n_343), .Y(n_340) );
INVx1_ASAP7_75t_L g416 ( .A(n_341), .Y(n_416) );
AND2x2_ASAP7_75t_L g429 ( .A(n_343), .B(n_352), .Y(n_429) );
AOI21xp33_ASAP7_75t_L g345 ( .A1(n_346), .A2(n_347), .B(n_349), .Y(n_345) );
INVx1_ASAP7_75t_SL g347 ( .A(n_348), .Y(n_347) );
INVxp67_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_351), .B(n_353), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_353), .B(n_456), .Y(n_455) );
OAI21xp33_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_356), .B(n_360), .Y(n_354) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
OAI221xp5_ASAP7_75t_SL g361 ( .A1(n_362), .A2(n_363), .B1(n_365), .B2(n_366), .C(n_367), .Y(n_361) );
A2O1A1Ixp33_ASAP7_75t_L g430 ( .A1(n_362), .A2(n_431), .B(n_433), .C(n_436), .Y(n_430) );
CKINVDCx16_ASAP7_75t_R g363 ( .A(n_364), .Y(n_363) );
NAND2xp5_ASAP7_75t_SL g414 ( .A(n_365), .B(n_415), .Y(n_414) );
NOR2xp33_ASAP7_75t_L g368 ( .A(n_369), .B(n_370), .Y(n_368) );
INVx1_ASAP7_75t_L g392 ( .A(n_373), .Y(n_392) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
AND2x2_ASAP7_75t_L g378 ( .A(n_376), .B(n_379), .Y(n_378) );
AND2x2_ASAP7_75t_L g420 ( .A(n_376), .B(n_421), .Y(n_420) );
INVx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
OAI211xp5_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_384), .B(n_386), .C(n_395), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
OAI221xp5_ASAP7_75t_L g457 ( .A1(n_384), .A2(n_394), .B1(n_458), .B2(n_459), .C(n_461), .Y(n_457) );
INVx1_ASAP7_75t_SL g384 ( .A(n_385), .Y(n_384) );
AOI22xp5_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_389), .B1(n_390), .B2(n_393), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g390 ( .A(n_391), .B(n_392), .Y(n_390) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
OAI21xp5_ASAP7_75t_SL g395 ( .A1(n_396), .A2(n_397), .B(n_398), .Y(n_395) );
INVx1_ASAP7_75t_SL g458 ( .A(n_397), .Y(n_458) );
INVxp67_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
NOR4xp25_ASAP7_75t_L g400 ( .A(n_401), .B(n_430), .C(n_450), .D(n_457), .Y(n_400) );
OAI211xp5_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_406), .B(n_408), .C(n_426), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_403), .B(n_405), .Y(n_402) );
INVxp67_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
O2A1O1Ixp33_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_412), .B(n_414), .C(n_418), .Y(n_408) );
INVx1_ASAP7_75t_SL g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_SL g437 ( .A(n_415), .Y(n_437) );
OR2x2_ASAP7_75t_L g415 ( .A(n_416), .B(n_417), .Y(n_415) );
OR2x2_ASAP7_75t_L g448 ( .A(n_416), .B(n_449), .Y(n_448) );
OAI21xp33_ASAP7_75t_L g418 ( .A1(n_419), .A2(n_422), .B(n_423), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
HB1xp67_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
AOI221xp5_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_438), .B1(n_440), .B2(n_442), .C(n_444), .Y(n_436) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVxp67_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_447), .B(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx2_ASAP7_75t_L g746 ( .A(n_464), .Y(n_746) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g748 ( .A(n_466), .Y(n_748) );
INVx1_ASAP7_75t_L g749 ( .A(n_467), .Y(n_749) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
AND2x2_ASAP7_75t_SL g468 ( .A(n_469), .B(n_678), .Y(n_468) );
NOR5xp2_ASAP7_75t_L g469 ( .A(n_470), .B(n_591), .C(n_637), .D(n_650), .E(n_662), .Y(n_469) );
OAI211xp5_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_505), .B(n_545), .C(n_572), .Y(n_470) );
INVx1_ASAP7_75t_SL g673 ( .A(n_471), .Y(n_673) );
OR2x2_ASAP7_75t_L g471 ( .A(n_472), .B(n_481), .Y(n_471) );
AND2x2_ASAP7_75t_L g597 ( .A(n_472), .B(n_482), .Y(n_597) );
AND2x2_ASAP7_75t_L g625 ( .A(n_472), .B(n_571), .Y(n_625) );
AND2x2_ASAP7_75t_L g633 ( .A(n_472), .B(n_576), .Y(n_633) );
INVx3_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
AND2x2_ASAP7_75t_L g563 ( .A(n_473), .B(n_483), .Y(n_563) );
INVx2_ASAP7_75t_L g575 ( .A(n_473), .Y(n_575) );
AND2x2_ASAP7_75t_L g700 ( .A(n_473), .B(n_642), .Y(n_700) );
OR2x2_ASAP7_75t_L g702 ( .A(n_473), .B(n_703), .Y(n_702) );
AND2x4_ASAP7_75t_L g473 ( .A(n_474), .B(n_475), .Y(n_473) );
INVx1_ASAP7_75t_L g569 ( .A(n_474), .Y(n_569) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_478), .A2(n_490), .B(n_491), .Y(n_489) );
O2A1O1Ixp33_ASAP7_75t_L g500 ( .A1(n_478), .A2(n_501), .B(n_502), .C(n_503), .Y(n_500) );
OAI21xp5_ASAP7_75t_L g555 ( .A1(n_480), .A2(n_556), .B(n_559), .Y(n_555) );
INVx2_ASAP7_75t_SL g481 ( .A(n_482), .Y(n_481) );
AND2x2_ASAP7_75t_L g613 ( .A(n_482), .B(n_585), .Y(n_613) );
NOR2xp33_ASAP7_75t_L g641 ( .A(n_482), .B(n_642), .Y(n_641) );
AND2x2_ASAP7_75t_L g727 ( .A(n_482), .B(n_567), .Y(n_727) );
AND2x2_ASAP7_75t_L g482 ( .A(n_483), .B(n_494), .Y(n_482) );
AND2x2_ASAP7_75t_L g570 ( .A(n_483), .B(n_571), .Y(n_570) );
INVx2_ASAP7_75t_L g617 ( .A(n_483), .Y(n_617) );
AND2x2_ASAP7_75t_L g642 ( .A(n_483), .B(n_554), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_483), .B(n_675), .Y(n_712) );
INVx3_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
AND2x2_ASAP7_75t_L g576 ( .A(n_484), .B(n_554), .Y(n_576) );
AND2x2_ASAP7_75t_L g590 ( .A(n_484), .B(n_553), .Y(n_590) );
AND2x2_ASAP7_75t_L g607 ( .A(n_484), .B(n_494), .Y(n_607) );
AND2x2_ASAP7_75t_L g664 ( .A(n_484), .B(n_665), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_484), .B(n_571), .Y(n_677) );
AND2x2_ASAP7_75t_L g729 ( .A(n_484), .B(n_654), .Y(n_729) );
INVx2_ASAP7_75t_L g501 ( .A(n_492), .Y(n_501) );
AND2x2_ASAP7_75t_L g552 ( .A(n_494), .B(n_553), .Y(n_552) );
INVx2_ASAP7_75t_L g571 ( .A(n_494), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_494), .B(n_554), .Y(n_648) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_506), .A2(n_530), .B(n_542), .Y(n_505) );
INVx1_ASAP7_75t_SL g661 ( .A(n_506), .Y(n_661) );
AND2x4_ASAP7_75t_L g506 ( .A(n_507), .B(n_520), .Y(n_506) );
BUFx3_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
AND2x2_ASAP7_75t_SL g549 ( .A(n_508), .B(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx2_ASAP7_75t_L g544 ( .A(n_509), .Y(n_544) );
INVx1_ASAP7_75t_L g581 ( .A(n_509), .Y(n_581) );
AND2x2_ASAP7_75t_L g602 ( .A(n_509), .B(n_525), .Y(n_602) );
AND2x2_ASAP7_75t_L g636 ( .A(n_509), .B(n_526), .Y(n_636) );
OR2x2_ASAP7_75t_L g655 ( .A(n_509), .B(n_532), .Y(n_655) );
HB1xp67_ASAP7_75t_L g669 ( .A(n_509), .Y(n_669) );
AND2x2_ASAP7_75t_L g682 ( .A(n_509), .B(n_683), .Y(n_682) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_512), .A2(n_513), .B(n_514), .Y(n_511) );
AOI22xp5_ASAP7_75t_L g603 ( .A1(n_520), .A2(n_604), .B1(n_605), .B2(n_614), .Y(n_603) );
AND2x2_ASAP7_75t_L g687 ( .A(n_520), .B(n_688), .Y(n_687) );
AND2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_525), .Y(n_520) );
INVx1_ASAP7_75t_L g548 ( .A(n_521), .Y(n_548) );
BUFx6f_ASAP7_75t_L g585 ( .A(n_521), .Y(n_585) );
INVx1_ASAP7_75t_L g596 ( .A(n_521), .Y(n_596) );
AND2x2_ASAP7_75t_L g611 ( .A(n_521), .B(n_526), .Y(n_611) );
OR2x2_ASAP7_75t_L g565 ( .A(n_525), .B(n_550), .Y(n_565) );
AND2x2_ASAP7_75t_L g595 ( .A(n_525), .B(n_596), .Y(n_595) );
NOR2xp67_ASAP7_75t_L g683 ( .A(n_525), .B(n_684), .Y(n_683) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
AND2x2_ASAP7_75t_L g543 ( .A(n_526), .B(n_544), .Y(n_543) );
BUFx2_ASAP7_75t_L g652 ( .A(n_526), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_530), .B(n_668), .Y(n_667) );
BUFx2_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
AND2x2_ASAP7_75t_L g630 ( .A(n_531), .B(n_596), .Y(n_630) );
INVx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
AND2x2_ASAP7_75t_L g542 ( .A(n_532), .B(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g601 ( .A(n_532), .Y(n_601) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx2_ASAP7_75t_L g550 ( .A(n_533), .Y(n_550) );
OR2x2_ASAP7_75t_L g580 ( .A(n_533), .B(n_581), .Y(n_580) );
HB1xp67_ASAP7_75t_L g635 ( .A(n_533), .Y(n_635) );
AOI32xp33_ASAP7_75t_L g672 ( .A1(n_542), .A2(n_602), .A3(n_673), .B1(n_674), .B2(n_676), .Y(n_672) );
AND2x2_ASAP7_75t_L g598 ( .A(n_543), .B(n_599), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_543), .B(n_697), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_543), .B(n_630), .Y(n_716) );
INVx1_ASAP7_75t_L g721 ( .A(n_543), .Y(n_721) );
AOI22xp5_ASAP7_75t_L g545 ( .A1(n_546), .A2(n_551), .B1(n_564), .B2(n_566), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_547), .B(n_549), .Y(n_546) );
AND2x2_ASAP7_75t_L g651 ( .A(n_547), .B(n_652), .Y(n_651) );
HB1xp67_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_548), .B(n_550), .Y(n_695) );
AOI22xp5_ASAP7_75t_L g572 ( .A1(n_549), .A2(n_573), .B1(n_577), .B2(n_587), .Y(n_572) );
AND2x2_ASAP7_75t_L g594 ( .A(n_549), .B(n_595), .Y(n_594) );
A2O1A1Ixp33_ASAP7_75t_L g645 ( .A1(n_549), .A2(n_563), .B(n_611), .C(n_646), .Y(n_645) );
OAI332xp33_ASAP7_75t_L g650 ( .A1(n_549), .A2(n_651), .A3(n_653), .B1(n_655), .B2(n_656), .B3(n_658), .C1(n_659), .C2(n_661), .Y(n_650) );
INVx2_ASAP7_75t_L g691 ( .A(n_549), .Y(n_691) );
HB1xp67_ASAP7_75t_L g609 ( .A(n_550), .Y(n_609) );
INVx1_ASAP7_75t_L g684 ( .A(n_550), .Y(n_684) );
AND2x2_ASAP7_75t_L g738 ( .A(n_550), .B(n_602), .Y(n_738) );
AND2x2_ASAP7_75t_L g551 ( .A(n_552), .B(n_563), .Y(n_551) );
AND2x2_ASAP7_75t_L g618 ( .A(n_553), .B(n_568), .Y(n_618) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g567 ( .A(n_554), .B(n_568), .Y(n_567) );
OR2x2_ASAP7_75t_L g666 ( .A(n_554), .B(n_568), .Y(n_666) );
INVx1_ASAP7_75t_L g675 ( .A(n_554), .Y(n_675) );
INVx1_ASAP7_75t_L g649 ( .A(n_563), .Y(n_649) );
INVxp67_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
OR2x2_ASAP7_75t_L g733 ( .A(n_565), .B(n_585), .Y(n_733) );
INVx1_ASAP7_75t_SL g644 ( .A(n_566), .Y(n_644) );
AND2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_570), .Y(n_566) );
AND2x2_ASAP7_75t_L g671 ( .A(n_567), .B(n_629), .Y(n_671) );
INVx1_ASAP7_75t_L g690 ( .A(n_567), .Y(n_690) );
NAND2xp5_ASAP7_75t_SL g692 ( .A(n_567), .B(n_657), .Y(n_692) );
INVx1_ASAP7_75t_L g589 ( .A(n_568), .Y(n_589) );
AND2x2_ASAP7_75t_L g593 ( .A(n_570), .B(n_574), .Y(n_593) );
AND2x2_ASAP7_75t_L g660 ( .A(n_570), .B(n_618), .Y(n_660) );
INVx2_ASAP7_75t_L g703 ( .A(n_570), .Y(n_703) );
INVx2_ASAP7_75t_L g586 ( .A(n_571), .Y(n_586) );
AND2x2_ASAP7_75t_L g588 ( .A(n_571), .B(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g573 ( .A(n_574), .B(n_576), .Y(n_573) );
INVx1_ASAP7_75t_L g604 ( .A(n_574), .Y(n_604) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g654 ( .A(n_575), .B(n_648), .Y(n_654) );
OR2x2_ASAP7_75t_L g718 ( .A(n_575), .B(n_677), .Y(n_718) );
INVx1_ASAP7_75t_L g742 ( .A(n_575), .Y(n_742) );
INVx1_ASAP7_75t_L g698 ( .A(n_576), .Y(n_698) );
AND2x2_ASAP7_75t_L g743 ( .A(n_576), .B(n_586), .Y(n_743) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_579), .B(n_582), .Y(n_578) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
OAI22xp5_ASAP7_75t_L g605 ( .A1(n_580), .A2(n_606), .B1(n_608), .B2(n_612), .Y(n_605) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
OAI322xp33_ASAP7_75t_SL g689 ( .A1(n_583), .A2(n_690), .A3(n_691), .B1(n_692), .B2(n_693), .C1(n_696), .C2(n_698), .Y(n_689) );
OR2x2_ASAP7_75t_L g583 ( .A(n_584), .B(n_586), .Y(n_583) );
AND2x2_ASAP7_75t_L g686 ( .A(n_584), .B(n_602), .Y(n_686) );
OR2x2_ASAP7_75t_L g720 ( .A(n_584), .B(n_721), .Y(n_720) );
OR2x2_ASAP7_75t_L g723 ( .A(n_584), .B(n_655), .Y(n_723) );
INVx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g668 ( .A(n_585), .B(n_669), .Y(n_668) );
OR2x2_ASAP7_75t_L g724 ( .A(n_585), .B(n_655), .Y(n_724) );
INVx3_ASAP7_75t_L g657 ( .A(n_586), .Y(n_657) );
AND2x2_ASAP7_75t_L g587 ( .A(n_588), .B(n_590), .Y(n_587) );
INVx1_ASAP7_75t_L g713 ( .A(n_588), .Y(n_713) );
AOI222xp33_ASAP7_75t_L g592 ( .A1(n_590), .A2(n_593), .B1(n_594), .B2(n_597), .C1(n_598), .C2(n_600), .Y(n_592) );
INVx1_ASAP7_75t_L g623 ( .A(n_590), .Y(n_623) );
NAND3xp33_ASAP7_75t_SL g591 ( .A(n_592), .B(n_603), .C(n_620), .Y(n_591) );
AND2x2_ASAP7_75t_L g708 ( .A(n_595), .B(n_609), .Y(n_708) );
BUFx2_ASAP7_75t_L g599 ( .A(n_596), .Y(n_599) );
INVx1_ASAP7_75t_L g640 ( .A(n_596), .Y(n_640) );
AOI221xp5_ASAP7_75t_L g685 ( .A1(n_597), .A2(n_633), .B1(n_686), .B2(n_687), .C(n_689), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_599), .B(n_682), .Y(n_681) );
AND2x2_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
HB1xp67_ASAP7_75t_L g626 ( .A(n_602), .Y(n_626) );
AND2x2_ASAP7_75t_L g639 ( .A(n_602), .B(n_640), .Y(n_639) );
INVx1_ASAP7_75t_SL g606 ( .A(n_607), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_607), .B(n_618), .Y(n_619) );
OR2x2_ASAP7_75t_L g608 ( .A(n_609), .B(n_610), .Y(n_608) );
OAI21xp33_ASAP7_75t_L g614 ( .A1(n_609), .A2(n_615), .B(n_619), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_609), .B(n_639), .Y(n_638) );
INVx1_ASAP7_75t_SL g610 ( .A(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g706 ( .A(n_611), .B(n_688), .Y(n_706) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_617), .B(n_618), .Y(n_616) );
INVx1_ASAP7_75t_L g629 ( .A(n_617), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_618), .B(n_629), .Y(n_628) );
INVx2_ASAP7_75t_L g735 ( .A(n_618), .Y(n_735) );
AOI221xp5_ASAP7_75t_L g620 ( .A1(n_621), .A2(n_626), .B1(n_627), .B2(n_630), .C(n_631), .Y(n_620) );
INVx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
NAND2xp5_ASAP7_75t_SL g710 ( .A(n_622), .B(n_711), .Y(n_710) );
OR2x2_ASAP7_75t_L g622 ( .A(n_623), .B(n_624), .Y(n_622) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g731 ( .A(n_630), .B(n_636), .Y(n_731) );
INVxp67_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_633), .B(n_634), .Y(n_632) );
OAI31xp33_ASAP7_75t_SL g699 ( .A1(n_634), .A2(n_673), .A3(n_700), .B(n_701), .Y(n_699) );
AND2x2_ASAP7_75t_L g634 ( .A(n_635), .B(n_636), .Y(n_634) );
INVx1_ASAP7_75t_L g688 ( .A(n_635), .Y(n_688) );
NAND2xp5_ASAP7_75t_SL g739 ( .A(n_636), .B(n_640), .Y(n_739) );
OAI221xp5_ASAP7_75t_SL g637 ( .A1(n_638), .A2(n_641), .B1(n_643), .B2(n_644), .C(n_645), .Y(n_637) );
INVx1_ASAP7_75t_L g643 ( .A(n_639), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_642), .B(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
OR2x2_ASAP7_75t_L g647 ( .A(n_648), .B(n_649), .Y(n_647) );
INVx1_ASAP7_75t_L g658 ( .A(n_651), .Y(n_658) );
INVx2_ASAP7_75t_L g694 ( .A(n_652), .Y(n_694) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
OR2x2_ASAP7_75t_L g680 ( .A(n_657), .B(n_666), .Y(n_680) );
A2O1A1Ixp33_ASAP7_75t_L g730 ( .A1(n_657), .A2(n_674), .B(n_731), .C(n_732), .Y(n_730) );
OAI221xp5_ASAP7_75t_SL g662 ( .A1(n_658), .A2(n_663), .B1(n_667), .B2(n_670), .C(n_672), .Y(n_662) );
INVx1_ASAP7_75t_SL g659 ( .A(n_660), .Y(n_659) );
A2O1A1Ixp33_ASAP7_75t_L g725 ( .A1(n_661), .A2(n_726), .B(n_728), .C(n_730), .Y(n_725) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
AOI221xp5_ASAP7_75t_L g714 ( .A1(n_664), .A2(n_715), .B1(n_717), .B2(n_719), .C(n_722), .Y(n_714) );
INVx1_ASAP7_75t_SL g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_SL g676 ( .A(n_677), .Y(n_676) );
NOR4xp25_ASAP7_75t_L g678 ( .A(n_679), .B(n_704), .C(n_725), .D(n_736), .Y(n_678) );
OAI211xp5_ASAP7_75t_SL g679 ( .A1(n_680), .A2(n_681), .B(n_685), .C(n_699), .Y(n_679) );
INVx1_ASAP7_75t_SL g734 ( .A(n_686), .Y(n_734) );
OR2x2_ASAP7_75t_L g693 ( .A(n_694), .B(n_695), .Y(n_693) );
INVx1_ASAP7_75t_SL g697 ( .A(n_695), .Y(n_697) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
OAI22xp5_ASAP7_75t_L g722 ( .A1(n_702), .A2(n_711), .B1(n_723), .B2(n_724), .Y(n_722) );
A2O1A1Ixp33_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_707), .B(n_709), .C(n_714), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
AOI31xp33_ASAP7_75t_L g736 ( .A1(n_707), .A2(n_737), .A3(n_739), .B(n_740), .Y(n_736) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVxp67_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
OR2x2_ASAP7_75t_L g711 ( .A(n_712), .B(n_713), .Y(n_711) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_SL g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_SL g728 ( .A(n_729), .Y(n_728) );
AOI21xp5_ASAP7_75t_L g732 ( .A1(n_733), .A2(n_734), .B(n_735), .Y(n_732) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_741), .B(n_743), .Y(n_740) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx2_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx2_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx2_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx1_ASAP7_75t_SL g753 ( .A(n_754), .Y(n_753) );
CKINVDCx20_ASAP7_75t_R g757 ( .A(n_758), .Y(n_757) );
CKINVDCx20_ASAP7_75t_R g759 ( .A(n_760), .Y(n_759) );
INVx1_ASAP7_75t_SL g764 ( .A(n_765), .Y(n_764) );
INVx1_ASAP7_75t_SL g766 ( .A(n_767), .Y(n_766) );
endmodule