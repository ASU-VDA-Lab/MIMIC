module fake_jpeg_28462_n_534 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_534);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_534;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_479;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx11_ASAP7_75t_SL g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_17),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_17),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_8),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_50),
.Y(n_106)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_51),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_52),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_53),
.Y(n_119)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_54),
.Y(n_141)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_55),
.Y(n_124)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_56),
.Y(n_103)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_57),
.Y(n_142)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_58),
.Y(n_107)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_59),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_60),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_61),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_62),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_30),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_63),
.Y(n_149)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_64),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_29),
.B(n_17),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_65),
.B(n_70),
.Y(n_158)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_66),
.Y(n_143)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_67),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_68),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_27),
.B(n_16),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_29),
.B(n_16),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_71),
.B(n_90),
.Y(n_105)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_28),
.Y(n_72)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_72),
.Y(n_102)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_32),
.Y(n_73)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_73),
.Y(n_113)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_74),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_75),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_76),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx3_ASAP7_75t_SL g144 ( 
.A(n_77),
.Y(n_144)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_78),
.Y(n_128)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_27),
.Y(n_79)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_79),
.Y(n_130)
);

BUFx24_ASAP7_75t_L g80 ( 
.A(n_25),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g135 ( 
.A(n_80),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_81),
.Y(n_126)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_31),
.Y(n_82)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_82),
.Y(n_138)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_31),
.Y(n_83)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_83),
.Y(n_140)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_84),
.Y(n_146)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_85),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_86),
.Y(n_160)
);

INVx6_ASAP7_75t_SL g87 ( 
.A(n_41),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_87),
.Y(n_154)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_88),
.Y(n_164)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_19),
.Y(n_89)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_89),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_34),
.B(n_14),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_91),
.Y(n_122)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_28),
.Y(n_92)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_92),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_34),
.B(n_0),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_95),
.Y(n_117)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_94),
.Y(n_156)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_41),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_19),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_96),
.B(n_98),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_39),
.Y(n_97)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_23),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_39),
.Y(n_99)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_99),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_35),
.B(n_21),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_21),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_39),
.Y(n_101)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_101),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_70),
.B(n_35),
.C(n_47),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_109),
.B(n_139),
.C(n_36),
.Y(n_202)
);

BUFx10_ASAP7_75t_L g120 ( 
.A(n_80),
.Y(n_120)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_120),
.Y(n_180)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_51),
.Y(n_125)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_125),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_127),
.B(n_136),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_95),
.B(n_43),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_134),
.B(n_162),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_94),
.B(n_43),
.Y(n_136)
);

HAxp5_ASAP7_75t_SL g137 ( 
.A(n_80),
.B(n_20),
.CON(n_137),
.SN(n_137)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_137),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_60),
.B(n_46),
.C(n_23),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_95),
.A2(n_44),
.B1(n_42),
.B2(n_26),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_145),
.A2(n_152),
.B1(n_161),
.B2(n_63),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_75),
.B(n_46),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_148),
.B(n_153),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_88),
.A2(n_41),
.B1(n_42),
.B2(n_44),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_91),
.B(n_40),
.Y(n_153)
);

INVx6_ASAP7_75t_SL g157 ( 
.A(n_97),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g225 ( 
.A(n_157),
.Y(n_225)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_55),
.Y(n_159)
);

INVx5_ASAP7_75t_L g204 ( 
.A(n_159),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_99),
.A2(n_44),
.B1(n_42),
.B2(n_26),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_72),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_104),
.A2(n_68),
.B1(n_86),
.B2(n_81),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_165),
.A2(n_221),
.B1(n_225),
.B2(n_133),
.Y(n_256)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_160),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_166),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_158),
.B(n_24),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_168),
.B(n_171),
.Y(n_238)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_135),
.Y(n_169)
);

INVx13_ASAP7_75t_L g235 ( 
.A(n_169),
.Y(n_235)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_103),
.Y(n_170)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_170),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_121),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_107),
.Y(n_172)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_172),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_174),
.A2(n_222),
.B1(n_119),
.B2(n_1),
.Y(n_261)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_160),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_175),
.Y(n_267)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_150),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_176),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_121),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_177),
.B(n_188),
.Y(n_229)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_125),
.Y(n_178)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_178),
.Y(n_269)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_135),
.Y(n_179)
);

INVx13_ASAP7_75t_L g247 ( 
.A(n_179),
.Y(n_247)
);

INVx4_ASAP7_75t_SL g181 ( 
.A(n_120),
.Y(n_181)
);

INVx13_ASAP7_75t_L g268 ( 
.A(n_181),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_158),
.B(n_24),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_182),
.B(n_208),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_156),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_183),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_127),
.B(n_40),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_184),
.B(n_142),
.Y(n_249)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_106),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_185),
.Y(n_263)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_113),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_186),
.Y(n_255)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_110),
.Y(n_187)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_187),
.Y(n_272)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_111),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_120),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_189),
.B(n_196),
.Y(n_234)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_138),
.Y(n_191)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_191),
.Y(n_228)
);

BUFx12f_ASAP7_75t_L g192 ( 
.A(n_115),
.Y(n_192)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_192),
.Y(n_270)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_140),
.Y(n_193)
);

CKINVDCx14_ASAP7_75t_R g253 ( 
.A(n_193),
.Y(n_253)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_155),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_194),
.Y(n_237)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_164),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_195),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_136),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_114),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_197),
.B(n_198),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_105),
.B(n_36),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_118),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_199),
.B(n_202),
.Y(n_245)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_116),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_200),
.Y(n_251)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_128),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_201),
.Y(n_266)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_130),
.Y(n_203)
);

INVx11_ASAP7_75t_L g248 ( 
.A(n_203),
.Y(n_248)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_108),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_206),
.B(n_207),
.Y(n_257)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_108),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_105),
.B(n_20),
.Y(n_208)
);

OAI21xp33_ASAP7_75t_L g209 ( 
.A1(n_117),
.A2(n_44),
.B(n_42),
.Y(n_209)
);

O2A1O1Ixp33_ASAP7_75t_L g236 ( 
.A1(n_209),
.A2(n_216),
.B(n_215),
.C(n_214),
.Y(n_236)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_148),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_210),
.B(n_217),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_146),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_211),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_144),
.A2(n_101),
.B1(n_26),
.B2(n_42),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_212),
.A2(n_223),
.B1(n_224),
.B2(n_122),
.Y(n_227)
);

INVx2_ASAP7_75t_SL g213 ( 
.A(n_143),
.Y(n_213)
);

BUFx12f_ASAP7_75t_L g226 ( 
.A(n_213),
.Y(n_226)
);

A2O1A1Ixp33_ASAP7_75t_L g214 ( 
.A1(n_117),
.A2(n_20),
.B(n_44),
.C(n_26),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_214),
.B(n_220),
.Y(n_265)
);

NAND2xp33_ASAP7_75t_SL g216 ( 
.A(n_154),
.B(n_20),
.Y(n_216)
);

OR2x2_ASAP7_75t_L g230 ( 
.A(n_216),
.B(n_218),
.Y(n_230)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_153),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_141),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_112),
.A2(n_62),
.B1(n_77),
.B2(n_76),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_219),
.A2(n_132),
.B1(n_151),
.B2(n_149),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_119),
.B(n_20),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_161),
.A2(n_69),
.B1(n_61),
.B2(n_53),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_145),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_144),
.A2(n_26),
.B1(n_52),
.B2(n_92),
.Y(n_223)
);

INVx8_ASAP7_75t_L g224 ( 
.A(n_124),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_227),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_167),
.B(n_149),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_231),
.B(n_246),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_236),
.B(n_243),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_L g279 ( 
.A1(n_239),
.A2(n_207),
.B1(n_206),
.B2(n_175),
.Y(n_279)
);

OA22x2_ASAP7_75t_L g243 ( 
.A1(n_219),
.A2(n_152),
.B1(n_126),
.B2(n_131),
.Y(n_243)
);

AO22x1_ASAP7_75t_SL g246 ( 
.A1(n_209),
.A2(n_132),
.B1(n_151),
.B2(n_133),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_249),
.B(n_259),
.Y(n_280)
);

AO22x1_ASAP7_75t_L g250 ( 
.A1(n_212),
.A2(n_147),
.B1(n_129),
.B2(n_123),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_250),
.A2(n_204),
.B(n_180),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_205),
.B(n_202),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_254),
.B(n_262),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_256),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_173),
.B(n_0),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_261),
.B(n_169),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_205),
.B(n_124),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_213),
.B(n_170),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_271),
.B(n_180),
.Y(n_286)
);

OAI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_166),
.A2(n_163),
.B1(n_102),
.B2(n_2),
.Y(n_273)
);

OAI22xp33_ASAP7_75t_L g314 ( 
.A1(n_273),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_190),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_274),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_237),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_275),
.B(n_285),
.Y(n_347)
);

A2O1A1Ixp33_ASAP7_75t_L g276 ( 
.A1(n_254),
.A2(n_223),
.B(n_181),
.C(n_172),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_276),
.A2(n_288),
.B(n_319),
.Y(n_323)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_272),
.Y(n_277)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_277),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_279),
.A2(n_253),
.B1(n_266),
.B2(n_260),
.Y(n_328)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_269),
.Y(n_281)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_281),
.Y(n_324)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_269),
.Y(n_282)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_282),
.Y(n_341)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_232),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g333 ( 
.A(n_283),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_245),
.B(n_203),
.C(n_201),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_284),
.B(n_297),
.C(n_238),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_237),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_286),
.B(n_303),
.Y(n_320)
);

XNOR2x1_ASAP7_75t_SL g287 ( 
.A(n_265),
.B(n_195),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_287),
.B(n_240),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_265),
.A2(n_224),
.B1(n_178),
.B2(n_200),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_289),
.A2(n_291),
.B1(n_294),
.B2(n_307),
.Y(n_332)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_272),
.Y(n_290)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_290),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_261),
.A2(n_204),
.B1(n_192),
.B2(n_179),
.Y(n_291)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_257),
.Y(n_293)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_293),
.Y(n_330)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_271),
.Y(n_295)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_295),
.Y(n_335)
);

XOR2x2_ASAP7_75t_L g296 ( 
.A(n_236),
.B(n_192),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_296),
.B(n_268),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_252),
.B(n_2),
.C(n_3),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_230),
.A2(n_13),
.B(n_4),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_298),
.A2(n_304),
.B(n_259),
.Y(n_336)
);

INVx8_ASAP7_75t_L g299 ( 
.A(n_233),
.Y(n_299)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_299),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_234),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_300),
.Y(n_351)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_255),
.Y(n_301)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_301),
.Y(n_337)
);

INVx2_ASAP7_75t_SL g303 ( 
.A(n_243),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_230),
.A2(n_13),
.B(n_4),
.Y(n_304)
);

INVx2_ASAP7_75t_SL g305 ( 
.A(n_243),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_305),
.B(n_308),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_258),
.B(n_3),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_306),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_256),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_229),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_309),
.A2(n_314),
.B1(n_267),
.B2(n_233),
.Y(n_353)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_255),
.Y(n_311)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_311),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_231),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_312),
.B(n_313),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_244),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_249),
.B(n_6),
.Y(n_315)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_315),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_262),
.B(n_230),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_316),
.A2(n_252),
.B(n_246),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_241),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_318),
.B(n_226),
.Y(n_357)
);

AOI22xp33_ASAP7_75t_SL g319 ( 
.A1(n_250),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g393 ( 
.A1(n_321),
.A2(n_329),
.B(n_334),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_327),
.Y(n_363)
);

AOI22xp33_ASAP7_75t_L g371 ( 
.A1(n_328),
.A2(n_353),
.B1(n_295),
.B2(n_309),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_R g329 ( 
.A(n_296),
.B(n_250),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_303),
.A2(n_246),
.B1(n_243),
.B2(n_239),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_331),
.A2(n_342),
.B1(n_354),
.B2(n_356),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_278),
.A2(n_246),
.B(n_260),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_336),
.Y(n_366)
);

OAI32xp33_ASAP7_75t_L g338 ( 
.A1(n_292),
.A2(n_263),
.A3(n_241),
.B1(n_226),
.B2(n_266),
.Y(n_338)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_338),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_316),
.A2(n_240),
.B(n_263),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g362 ( 
.A1(n_339),
.A2(n_358),
.B(n_359),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_340),
.B(n_359),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_303),
.A2(n_267),
.B1(n_233),
.B2(n_242),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_317),
.B(n_251),
.C(n_242),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_345),
.B(n_284),
.C(n_317),
.Y(n_368)
);

AOI32xp33_ASAP7_75t_L g348 ( 
.A1(n_296),
.A2(n_251),
.A3(n_270),
.B1(n_228),
.B2(n_268),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_348),
.B(n_294),
.Y(n_369)
);

OA22x2_ASAP7_75t_L g349 ( 
.A1(n_305),
.A2(n_228),
.B1(n_264),
.B2(n_232),
.Y(n_349)
);

INVx2_ASAP7_75t_SL g360 ( 
.A(n_349),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_305),
.A2(n_267),
.B1(n_264),
.B2(n_248),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_277),
.Y(n_355)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_355),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_292),
.A2(n_248),
.B1(n_226),
.B2(n_270),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_357),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_L g358 ( 
.A1(n_316),
.A2(n_226),
.B(n_268),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_SL g404 ( 
.A(n_361),
.B(n_328),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_322),
.B(n_312),
.Y(n_364)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_364),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_329),
.A2(n_302),
.B(n_278),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_SL g411 ( 
.A1(n_365),
.A2(n_369),
.B(n_341),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_368),
.B(n_373),
.C(n_379),
.Y(n_396)
);

NAND2x1_ASAP7_75t_SL g370 ( 
.A(n_349),
.B(n_287),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_370),
.A2(n_323),
.B(n_342),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_371),
.A2(n_386),
.B1(n_349),
.B2(n_346),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_351),
.B(n_308),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_372),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_340),
.B(n_276),
.C(n_278),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_322),
.B(n_300),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_374),
.B(n_378),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_320),
.A2(n_302),
.B1(n_310),
.B2(n_294),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_375),
.A2(n_381),
.B1(n_389),
.B2(n_344),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_335),
.B(n_313),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_345),
.B(n_327),
.C(n_350),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_334),
.A2(n_321),
.B1(n_350),
.B2(n_332),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_320),
.B(n_357),
.Y(n_382)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_382),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_339),
.B(n_293),
.C(n_289),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_383),
.B(n_390),
.C(n_235),
.Y(n_422)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_325),
.Y(n_384)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_384),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_SL g385 ( 
.A(n_352),
.B(n_280),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_385),
.B(n_346),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_331),
.A2(n_291),
.B1(n_307),
.B2(n_310),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_330),
.B(n_318),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_387),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_347),
.B(n_326),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_388),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_332),
.A2(n_288),
.B1(n_304),
.B2(n_298),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_358),
.B(n_297),
.C(n_290),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_356),
.A2(n_311),
.B1(n_301),
.B2(n_285),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_391),
.B(n_349),
.Y(n_400)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_338),
.Y(n_392)
);

CKINVDCx16_ASAP7_75t_R g403 ( 
.A(n_392),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_394),
.B(n_360),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_SL g442 ( 
.A1(n_395),
.A2(n_398),
.B(n_362),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_365),
.A2(n_323),
.B(n_336),
.Y(n_398)
);

CKINVDCx14_ASAP7_75t_R g437 ( 
.A(n_399),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_400),
.B(n_391),
.Y(n_434)
);

OAI21xp5_ASAP7_75t_L g402 ( 
.A1(n_369),
.A2(n_366),
.B(n_373),
.Y(n_402)
);

AO21x1_ASAP7_75t_L g447 ( 
.A1(n_402),
.A2(n_411),
.B(n_393),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_404),
.B(n_413),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_L g407 ( 
.A1(n_386),
.A2(n_343),
.B1(n_337),
.B2(n_354),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_407),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_408),
.A2(n_410),
.B1(n_414),
.B2(n_377),
.Y(n_443)
);

NOR2xp67_ASAP7_75t_L g409 ( 
.A(n_372),
.B(n_333),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_409),
.B(n_417),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_381),
.A2(n_344),
.B1(n_333),
.B2(n_299),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_379),
.B(n_275),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_360),
.A2(n_299),
.B1(n_341),
.B2(n_324),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_374),
.B(n_324),
.Y(n_416)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_416),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_387),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_385),
.B(n_282),
.Y(n_418)
);

INVxp33_ASAP7_75t_L g444 ( 
.A(n_418),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_361),
.B(n_281),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_419),
.B(n_420),
.C(n_422),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_368),
.B(n_235),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_388),
.B(n_283),
.Y(n_421)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_421),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_378),
.B(n_235),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_424),
.B(n_376),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_426),
.A2(n_450),
.B1(n_377),
.B2(n_403),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_412),
.B(n_364),
.Y(n_429)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_429),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_412),
.B(n_382),
.Y(n_430)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_430),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_396),
.B(n_363),
.C(n_390),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_433),
.B(n_422),
.C(n_396),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_434),
.B(n_435),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_423),
.B(n_376),
.Y(n_435)
);

NOR2x1_ASAP7_75t_L g436 ( 
.A(n_408),
.B(n_389),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_436),
.B(n_443),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g439 ( 
.A1(n_405),
.A2(n_360),
.B1(n_392),
.B2(n_367),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_439),
.A2(n_448),
.B1(n_401),
.B2(n_400),
.Y(n_466)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_416),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_440),
.B(n_441),
.Y(n_451)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_405),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_442),
.B(n_370),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_445),
.B(n_446),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_423),
.B(n_367),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_447),
.B(n_411),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g448 ( 
.A(n_421),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_397),
.B(n_384),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_449),
.Y(n_462)
);

OAI22x1_ASAP7_75t_L g450 ( 
.A1(n_394),
.A2(n_370),
.B1(n_400),
.B2(n_395),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_SL g484 ( 
.A(n_452),
.B(n_469),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_454),
.B(n_456),
.C(n_458),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_433),
.B(n_413),
.C(n_420),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_425),
.B(n_419),
.C(n_402),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_425),
.B(n_383),
.C(n_404),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_459),
.B(n_464),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_427),
.B(n_410),
.C(n_398),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_460),
.B(n_463),
.C(n_467),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_461),
.B(n_443),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_427),
.B(n_397),
.C(n_362),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_447),
.B(n_442),
.Y(n_464)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_466),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_435),
.B(n_393),
.C(n_406),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_447),
.B(n_375),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_468),
.B(n_434),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_441),
.B(n_406),
.C(n_414),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_471),
.B(n_429),
.C(n_448),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_473),
.B(n_476),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_457),
.A2(n_426),
.B1(n_450),
.B2(n_446),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_474),
.A2(n_439),
.B1(n_428),
.B2(n_469),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_L g475 ( 
.A1(n_465),
.A2(n_432),
.B1(n_437),
.B2(n_438),
.Y(n_475)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_475),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_460),
.B(n_434),
.Y(n_476)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_455),
.Y(n_479)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_479),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_481),
.B(n_463),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_482),
.B(n_487),
.C(n_478),
.Y(n_494)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_451),
.Y(n_483)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_483),
.Y(n_502)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_470),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_485),
.B(n_488),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_L g486 ( 
.A1(n_453),
.A2(n_436),
.B(n_430),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_486),
.B(n_449),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_454),
.B(n_428),
.C(n_440),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_462),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_472),
.A2(n_438),
.B1(n_471),
.B2(n_467),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_491),
.B(n_494),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_493),
.B(n_496),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_477),
.B(n_478),
.C(n_487),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_495),
.B(n_497),
.C(n_500),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_477),
.B(n_456),
.C(n_458),
.Y(n_497)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_498),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_486),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_499),
.B(n_484),
.Y(n_510)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_476),
.B(n_431),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_490),
.A2(n_474),
.B1(n_473),
.B2(n_481),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_506),
.B(n_512),
.Y(n_516)
);

NOR2xp67_ASAP7_75t_L g507 ( 
.A(n_495),
.B(n_480),
.Y(n_507)
);

A2O1A1Ixp33_ASAP7_75t_L g514 ( 
.A1(n_507),
.A2(n_511),
.B(n_504),
.C(n_503),
.Y(n_514)
);

AOI21xp5_ASAP7_75t_L g509 ( 
.A1(n_494),
.A2(n_482),
.B(n_484),
.Y(n_509)
);

OAI21xp5_ASAP7_75t_SL g519 ( 
.A1(n_509),
.A2(n_497),
.B(n_505),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_L g515 ( 
.A1(n_510),
.A2(n_513),
.B(n_496),
.Y(n_515)
);

AOI211xp5_ASAP7_75t_L g511 ( 
.A1(n_501),
.A2(n_431),
.B(n_415),
.C(n_444),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_489),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g513 ( 
.A(n_498),
.B(n_415),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_SL g521 ( 
.A1(n_514),
.A2(n_513),
.B(n_380),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_515),
.A2(n_517),
.B1(n_518),
.B2(n_520),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_508),
.B(n_502),
.Y(n_517)
);

BUFx4f_ASAP7_75t_SL g518 ( 
.A(n_508),
.Y(n_518)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_519),
.B(n_492),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_506),
.B(n_500),
.Y(n_520)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_521),
.Y(n_526)
);

XOR2xp5_ASAP7_75t_L g522 ( 
.A(n_516),
.B(n_492),
.Y(n_522)
);

AOI22xp33_ASAP7_75t_SL g525 ( 
.A1(n_522),
.A2(n_524),
.B1(n_493),
.B2(n_518),
.Y(n_525)
);

XOR2xp5_ASAP7_75t_L g528 ( 
.A(n_525),
.B(n_380),
.Y(n_528)
);

OAI21xp5_ASAP7_75t_L g527 ( 
.A1(n_526),
.A2(n_523),
.B(n_522),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_527),
.B(n_528),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_529),
.B(n_247),
.Y(n_530)
);

AO21x1_ASAP7_75t_L g531 ( 
.A1(n_530),
.A2(n_247),
.B(n_11),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_531),
.B(n_247),
.C(n_11),
.Y(n_532)
);

AOI21xp5_ASAP7_75t_SL g533 ( 
.A1(n_532),
.A2(n_9),
.B(n_12),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_533),
.B(n_9),
.Y(n_534)
);


endmodule