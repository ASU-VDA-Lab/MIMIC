module fake_jpeg_18172_n_73 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_73);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_73;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_51;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

INVx2_ASAP7_75t_SL g10 ( 
.A(n_5),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_5),
.Y(n_11)
);

INVx13_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_0),
.B(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_SL g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_24),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_11),
.B(n_20),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_25),
.B(n_26),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_15),
.C(n_20),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_15),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_15),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_SL g43 ( 
.A1(n_32),
.A2(n_12),
.B(n_16),
.Y(n_43)
);

NOR2x1_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_19),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_33),
.B(n_10),
.Y(n_37)
);

OAI21xp33_ASAP7_75t_L g52 ( 
.A1(n_35),
.A2(n_37),
.B(n_45),
.Y(n_52)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_38),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_28),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_17),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_41),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_31),
.A2(n_27),
.B1(n_10),
.B2(n_24),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_31),
.A2(n_13),
.B1(n_18),
.B2(n_9),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_44),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_32),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_27),
.B(n_32),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_46),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_39),
.Y(n_48)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_48),
.B(n_12),
.Y(n_60)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_54),
.Y(n_57)
);

FAx1_ASAP7_75t_SL g55 ( 
.A(n_51),
.B(n_43),
.CI(n_40),
.CON(n_55),
.SN(n_55)
);

A2O1A1O1Ixp25_ASAP7_75t_L g62 ( 
.A1(n_55),
.A2(n_60),
.B(n_52),
.C(n_53),
.D(n_16),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_54),
.B(n_35),
.Y(n_56)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_47),
.A2(n_33),
.B1(n_46),
.B2(n_34),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_58),
.A2(n_59),
.B1(n_49),
.B2(n_47),
.Y(n_61)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_61),
.A2(n_60),
.B1(n_57),
.B2(n_56),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_62),
.B(n_55),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_49),
.C(n_6),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g65 ( 
.A(n_63),
.B(n_58),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_65),
.B(n_67),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_66),
.A2(n_64),
.B1(n_61),
.B2(n_7),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_68),
.B(n_65),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_70),
.A2(n_71),
.B1(n_69),
.B2(n_3),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_68),
.B(n_3),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_7),
.Y(n_73)
);


endmodule