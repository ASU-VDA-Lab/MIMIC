module real_jpeg_33323_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_595;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_620;
wire n_578;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_605;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_601;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_288;
wire n_78;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_611;
wire n_104;
wire n_153;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_615;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_589;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_515;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_596;
wire n_312;
wire n_617;
wire n_325;
wire n_307;
wire n_316;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_604;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_572;
wire n_586;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_613;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_616;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_534;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_608;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_597;
wire n_618;
wire n_609;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_625;
wire n_85;
wire n_591;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx2_ASAP7_75t_L g189 ( 
.A(n_0),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_0),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_0),
.Y(n_234)
);

BUFx12f_ASAP7_75t_L g255 ( 
.A(n_0),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_1),
.A2(n_66),
.B1(n_71),
.B2(n_72),
.Y(n_65)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_1),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_1),
.A2(n_71),
.B1(n_223),
.B2(n_228),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_1),
.A2(n_71),
.B1(n_387),
.B2(n_481),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_SL g533 ( 
.A1(n_1),
.A2(n_71),
.B1(n_534),
.B2(n_535),
.Y(n_533)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_2),
.A2(n_141),
.B1(n_142),
.B2(n_144),
.Y(n_140)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_2),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_2),
.A2(n_144),
.B1(n_281),
.B2(n_284),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_L g514 ( 
.A1(n_2),
.A2(n_144),
.B1(n_481),
.B2(n_515),
.Y(n_514)
);

AOI22xp33_ASAP7_75t_SL g522 ( 
.A1(n_2),
.A2(n_144),
.B1(n_523),
.B2(n_524),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_4),
.A2(n_149),
.B1(n_152),
.B2(n_157),
.Y(n_148)
);

INVx2_ASAP7_75t_R g157 ( 
.A(n_4),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_4),
.A2(n_157),
.B1(n_329),
.B2(n_333),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g432 ( 
.A1(n_4),
.A2(n_157),
.B1(n_433),
.B2(n_436),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_4),
.A2(n_157),
.B1(n_498),
.B2(n_502),
.Y(n_497)
);

AOI21x1_ASAP7_75t_L g75 ( 
.A1(n_5),
.A2(n_76),
.B(n_82),
.Y(n_75)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_5),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_5),
.A2(n_83),
.B1(n_237),
.B2(n_238),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_5),
.A2(n_83),
.B1(n_320),
.B2(n_324),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_5),
.A2(n_83),
.B1(n_160),
.B2(n_398),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g54 ( 
.A1(n_6),
.A2(n_55),
.B(n_59),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_6),
.B(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_6),
.B(n_242),
.Y(n_241)
);

OAI32xp33_ASAP7_75t_L g441 ( 
.A1(n_6),
.A2(n_122),
.A3(n_442),
.B1(n_445),
.B2(n_451),
.Y(n_441)
);

INVx1_ASAP7_75t_SL g452 ( 
.A(n_6),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_6),
.B(n_146),
.Y(n_511)
);

OAI22xp33_ASAP7_75t_SL g540 ( 
.A1(n_6),
.A2(n_298),
.B1(n_533),
.B2(n_541),
.Y(n_540)
);

AOI22xp33_ASAP7_75t_L g558 ( 
.A1(n_6),
.A2(n_452),
.B1(n_559),
.B2(n_564),
.Y(n_558)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_7),
.A2(n_99),
.B1(n_102),
.B2(n_106),
.Y(n_98)
);

INVx2_ASAP7_75t_R g106 ( 
.A(n_7),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_7),
.A2(n_106),
.B1(n_271),
.B2(n_276),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_7),
.A2(n_106),
.B1(n_338),
.B2(n_340),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_7),
.A2(n_106),
.B1(n_459),
.B2(n_463),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_8),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_9),
.Y(n_127)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_9),
.Y(n_131)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_10),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_10),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_10),
.Y(n_466)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_11),
.Y(n_625)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_12),
.Y(n_94)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_12),
.Y(n_97)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_12),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_13),
.A2(n_304),
.B1(n_305),
.B2(n_307),
.Y(n_303)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_13),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_13),
.A2(n_307),
.B1(n_383),
.B2(n_386),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_14),
.A2(n_192),
.B1(n_193),
.B2(n_196),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_14),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_14),
.A2(n_192),
.B1(n_258),
.B2(n_262),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_14),
.A2(n_192),
.B1(n_276),
.B2(n_317),
.Y(n_316)
);

OAI22xp33_ASAP7_75t_SL g597 ( 
.A1(n_14),
.A2(n_192),
.B1(n_338),
.B2(n_598),
.Y(n_597)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_15),
.A2(n_21),
.B(n_624),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_15),
.B(n_625),
.Y(n_624)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_16),
.A2(n_249),
.B1(n_250),
.B2(n_251),
.Y(n_248)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_16),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_L g347 ( 
.A1(n_16),
.A2(n_251),
.B1(n_348),
.B2(n_350),
.Y(n_347)
);

AOI22xp33_ASAP7_75t_L g607 ( 
.A1(n_16),
.A2(n_251),
.B1(n_608),
.B2(n_613),
.Y(n_607)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_17),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_17),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_17),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_17),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_18),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_18),
.Y(n_134)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_18),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_19),
.A2(n_205),
.B1(n_207),
.B2(n_208),
.Y(n_204)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_19),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_19),
.A2(n_207),
.B1(n_310),
.B2(n_311),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_19),
.A2(n_207),
.B1(n_317),
.B2(n_373),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_584),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_422),
.B(n_579),
.Y(n_23)
);

NAND4xp25_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_292),
.C(n_402),
.D(n_415),
.Y(n_24)
);

OR2x2_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_243),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_26),
.B(n_243),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_158),
.C(n_218),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_SL g424 ( 
.A(n_27),
.B(n_425),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_73),
.Y(n_27)
);

HB1xp67_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_29),
.B(n_74),
.C(n_118),
.Y(n_245)
);

OAI22xp33_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_54),
.B1(n_63),
.B2(n_65),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_30),
.A2(n_328),
.B1(n_334),
.B2(n_336),
.Y(n_327)
);

OAI22x1_ASAP7_75t_L g362 ( 
.A1(n_30),
.A2(n_63),
.B1(n_280),
.B2(n_328),
.Y(n_362)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_31),
.A2(n_279),
.B1(n_286),
.B2(n_288),
.Y(n_278)
);

NAND2x1p5_ASAP7_75t_L g400 ( 
.A(n_31),
.B(n_337),
.Y(n_400)
);

NAND2xp33_ASAP7_75t_SL g601 ( 
.A(n_31),
.B(n_397),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_43),
.Y(n_31)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_36),
.B1(n_39),
.B2(n_41),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_34),
.Y(n_326)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_35),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_35),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_35),
.Y(n_563)
);

BUFx12f_ASAP7_75t_L g615 ( 
.A(n_35),
.Y(n_615)
);

INVx2_ASAP7_75t_SL g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_38),
.Y(n_168)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_38),
.Y(n_178)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g151 ( 
.A(n_40),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_40),
.Y(n_277)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_47),
.B1(n_50),
.B2(n_52),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx3_ASAP7_75t_L g399 ( 
.A(n_45),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_46),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_46),
.Y(n_600)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_51),
.Y(n_339)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_57),
.Y(n_216)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_59),
.Y(n_182)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_61),
.Y(n_333)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_62),
.Y(n_163)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_62),
.Y(n_285)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_62),
.Y(n_332)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_63),
.Y(n_242)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_64),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g335 ( 
.A(n_64),
.Y(n_335)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_65),
.Y(n_288)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_68),
.Y(n_341)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_69),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_118),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_87),
.B1(n_98),
.B2(n_107),
.Y(n_74)
);

OAI22x1_ASAP7_75t_SL g256 ( 
.A1(n_75),
.A2(n_87),
.B1(n_107),
.B2(n_257),
.Y(n_256)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_80),
.A2(n_136),
.B1(n_137),
.B2(n_139),
.Y(n_135)
);

INVx4_ASAP7_75t_L g456 ( 
.A(n_80),
.Y(n_456)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_81),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_81),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_84),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_SL g313 ( 
.A(n_85),
.Y(n_313)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_85),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_86),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_86),
.Y(n_263)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_86),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_87),
.A2(n_107),
.B1(n_257),
.B2(n_309),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_87),
.A2(n_107),
.B1(n_309),
.B2(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_87),
.Y(n_389)
);

OAI22xp33_ASAP7_75t_SL g430 ( 
.A1(n_87),
.A2(n_98),
.B1(n_107),
.B2(n_431),
.Y(n_430)
);

OAI22x1_ASAP7_75t_L g512 ( 
.A1(n_87),
.A2(n_107),
.B1(n_513),
.B2(n_514),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_SL g538 ( 
.A(n_87),
.B(n_452),
.Y(n_538)
);

AO21x1_ASAP7_75t_L g604 ( 
.A1(n_87),
.A2(n_107),
.B(n_382),
.Y(n_604)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

AO21x2_ASAP7_75t_L g107 ( 
.A1(n_89),
.A2(n_108),
.B(n_114),
.Y(n_107)
);

INVxp67_ASAP7_75t_SL g379 ( 
.A(n_89),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_90),
.A2(n_92),
.B1(n_95),
.B2(n_96),
.Y(n_89)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_90),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_91),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_91),
.Y(n_190)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_91),
.Y(n_206)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_91),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_91),
.Y(n_501)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_91),
.Y(n_505)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_94),
.Y(n_493)
);

BUFx12f_ASAP7_75t_L g250 ( 
.A(n_95),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

INVx2_ASAP7_75t_SL g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_105),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_105),
.Y(n_438)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_105),
.Y(n_450)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_108),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_112),
.Y(n_108)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_113),
.Y(n_385)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_114),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_117),
.Y(n_114)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_119),
.A2(n_140),
.B1(n_145),
.B2(n_148),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g557 ( 
.A1(n_119),
.A2(n_147),
.B1(n_222),
.B2(n_558),
.Y(n_557)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_120),
.A2(n_146),
.B1(n_316),
.B2(n_318),
.Y(n_315)
);

INVx2_ASAP7_75t_SL g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_121),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_121),
.A2(n_145),
.B1(n_148),
.B2(n_270),
.Y(n_269)
);

OAI22x1_ASAP7_75t_L g360 ( 
.A1(n_121),
.A2(n_145),
.B1(n_270),
.B2(n_319),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g605 ( 
.A1(n_121),
.A2(n_145),
.B1(n_606),
.B2(n_607),
.Y(n_605)
);

AO21x2_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_128),
.B(n_135),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_125),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g141 ( 
.A(n_123),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_124),
.Y(n_181)
);

INVx8_ASAP7_75t_L g229 ( 
.A(n_124),
.Y(n_229)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_127),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_132),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_134),
.Y(n_143)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_135),
.Y(n_147)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_136),
.Y(n_139)
);

HB1xp67_ASAP7_75t_L g310 ( 
.A(n_137),
.Y(n_310)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_140),
.A2(n_145),
.B1(n_220),
.B2(n_222),
.Y(n_219)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_146),
.A2(n_221),
.B1(n_316),
.B2(n_372),
.Y(n_371)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_SL g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_SL g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_155),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_156),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g612 ( 
.A(n_156),
.Y(n_612)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_158),
.B(n_218),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_183),
.B1(n_211),
.B2(n_217),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_159),
.B(n_217),
.Y(n_291)
);

OAI32xp33_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_164),
.A3(n_169),
.B1(n_174),
.B2(n_182),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

OAI32xp33_ASAP7_75t_L g212 ( 
.A1(n_164),
.A2(n_169),
.A3(n_174),
.B1(n_182),
.B2(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx4_ASAP7_75t_L g275 ( 
.A(n_173),
.Y(n_275)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_173),
.Y(n_374)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_173),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_175),
.B(n_179),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_183),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_191),
.B1(n_201),
.B2(n_203),
.Y(n_183)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_184),
.Y(n_298)
);

OA21x2_ASAP7_75t_L g353 ( 
.A1(n_184),
.A2(n_354),
.B(n_356),
.Y(n_353)
);

AO22x1_ASAP7_75t_L g457 ( 
.A1(n_184),
.A2(n_201),
.B1(n_236),
.B2(n_458),
.Y(n_457)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_185),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_185),
.A2(n_204),
.B1(n_248),
.B2(n_252),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g532 ( 
.A1(n_185),
.A2(n_522),
.B1(n_533),
.B2(n_536),
.Y(n_532)
);

OR2x2_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_190),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_189),
.Y(n_302)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_190),
.Y(n_195)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_190),
.Y(n_237)
);

AO22x1_ASAP7_75t_SL g230 ( 
.A1(n_191),
.A2(n_231),
.B1(n_235),
.B2(n_236),
.Y(n_230)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_199),
.Y(n_239)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_199),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx6_ASAP7_75t_L g486 ( 
.A(n_200),
.Y(n_486)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_200),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g548 ( 
.A(n_200),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx4_ASAP7_75t_L g306 ( 
.A(n_206),
.Y(n_306)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx2_ASAP7_75t_SL g213 ( 
.A(n_214),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_230),
.C(n_240),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_219),
.B(n_428),
.Y(n_427)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx5_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx5_ASAP7_75t_L g317 ( 
.A(n_229),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_230),
.B(n_241),
.Y(n_428)
);

INVx3_ASAP7_75t_SL g231 ( 
.A(n_232),
.Y(n_231)
);

INVx8_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_234),
.Y(n_508)
);

HB1xp67_ASAP7_75t_L g537 ( 
.A(n_234),
.Y(n_537)
);

BUFx3_ASAP7_75t_L g545 ( 
.A(n_234),
.Y(n_545)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_235),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_SL g520 ( 
.A1(n_235),
.A2(n_253),
.B1(n_521),
.B2(n_528),
.Y(n_520)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_266),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_246),
.B1(n_264),
.B2(n_265),
.Y(n_244)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_245),
.Y(n_264)
);

INVxp33_ASAP7_75t_L g417 ( 
.A(n_245),
.Y(n_417)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_246),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_256),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_247),
.B(n_256),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_248),
.A2(n_298),
.B1(n_299),
.B2(n_303),
.Y(n_297)
);

INVx2_ASAP7_75t_SL g304 ( 
.A(n_250),
.Y(n_304)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx5_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx8_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx8_ASAP7_75t_L g355 ( 
.A(n_255),
.Y(n_355)
);

INVx4_ASAP7_75t_SL g541 ( 
.A(n_255),
.Y(n_541)
);

BUFx4f_ASAP7_75t_SL g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_261),
.Y(n_435)
);

INVx4_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

BUFx3_ASAP7_75t_L g349 ( 
.A(n_263),
.Y(n_349)
);

INVx4_ASAP7_75t_L g388 ( 
.A(n_263),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_265),
.B(n_267),
.C(n_417),
.Y(n_416)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_291),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_278),
.B1(n_289),
.B2(n_290),
.Y(n_268)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_269),
.Y(n_289)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx4_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_278),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g410 ( 
.A(n_278),
.Y(n_410)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_286),
.Y(n_395)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_289),
.Y(n_411)
);

INVxp33_ASAP7_75t_L g409 ( 
.A(n_291),
.Y(n_409)
);

A2O1A1O1Ixp25_ASAP7_75t_L g579 ( 
.A1(n_292),
.A2(n_402),
.B(n_580),
.C(n_582),
.D(n_583),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_364),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_293),
.B(n_364),
.Y(n_583)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_344),
.C(n_357),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_295),
.B(n_414),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_SL g295 ( 
.A(n_296),
.B(n_314),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_296),
.B(n_343),
.C(n_366),
.Y(n_365)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_308),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_297),
.B(n_308),
.Y(n_412)
);

INVx4_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx4_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx2_ASAP7_75t_SL g301 ( 
.A(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_303),
.Y(n_356)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g311 ( 
.A(n_312),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

OAI22xp33_ASAP7_75t_L g314 ( 
.A1(n_315),
.A2(n_327),
.B1(n_342),
.B2(n_343),
.Y(n_314)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_315),
.Y(n_343)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_327),
.Y(n_342)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_327),
.Y(n_366)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_345),
.B(n_358),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_SL g345 ( 
.A(n_346),
.B(n_353),
.Y(n_345)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_346),
.B(n_353),
.Y(n_392)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_347),
.Y(n_380)
);

INVx2_ASAP7_75t_SL g348 ( 
.A(n_349),
.Y(n_348)
);

BUFx6f_ASAP7_75t_SL g350 ( 
.A(n_351),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_353),
.Y(n_401)
);

AOI21xp5_ASAP7_75t_L g619 ( 
.A1(n_353),
.A2(n_620),
.B(n_621),
.Y(n_619)
);

INVx4_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

MAJx2_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_361),
.C(n_363),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_359),
.A2(n_360),
.B1(n_362),
.B2(n_407),
.Y(n_406)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVxp67_ASAP7_75t_SL g361 ( 
.A(n_362),
.Y(n_361)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_362),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_363),
.B(n_406),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_367),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g587 ( 
.A(n_365),
.B(n_588),
.C(n_589),
.Y(n_587)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_391),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g589 ( 
.A(n_369),
.Y(n_589)
);

NOR2xp67_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_390),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_375),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_371),
.B(n_375),
.Y(n_390)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_372),
.Y(n_606)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_376),
.A2(n_380),
.B1(n_381),
.B2(n_389),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_376),
.A2(n_474),
.B1(n_479),
.B2(n_480),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g567 ( 
.A1(n_376),
.A2(n_389),
.B1(n_432),
.B2(n_568),
.Y(n_567)
);

OA21x2_ASAP7_75t_SL g376 ( 
.A1(n_377),
.A2(n_378),
.B(n_379),
.Y(n_376)
);

AOI21xp33_ASAP7_75t_L g483 ( 
.A1(n_378),
.A2(n_484),
.B(n_487),
.Y(n_483)
);

INVxp67_ASAP7_75t_L g479 ( 
.A(n_379),
.Y(n_479)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx2_ASAP7_75t_SL g386 ( 
.A(n_387),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g592 ( 
.A1(n_390),
.A2(n_593),
.B1(n_594),
.B2(n_595),
.Y(n_592)
);

INVx1_ASAP7_75t_SL g593 ( 
.A(n_390),
.Y(n_593)
);

INVxp33_ASAP7_75t_L g588 ( 
.A(n_391),
.Y(n_588)
);

XNOR2x1_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_393),
.Y(n_391)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_392),
.Y(n_620)
);

XNOR2x1_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_401),
.Y(n_393)
);

INVxp33_ASAP7_75t_L g621 ( 
.A(n_394),
.Y(n_621)
);

OAI21x1_ASAP7_75t_L g394 ( 
.A1(n_395),
.A2(n_396),
.B(n_400),
.Y(n_394)
);

OA21x2_ASAP7_75t_L g595 ( 
.A1(n_395),
.A2(n_596),
.B(n_601),
.Y(n_595)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_413),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_403),
.B(n_413),
.Y(n_582)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_408),
.C(n_412),
.Y(n_403)
);

HB1xp67_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_405),
.B(n_421),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_410),
.C(n_411),
.Y(n_408)
);

MAJx2_ASAP7_75t_L g419 ( 
.A(n_409),
.B(n_410),
.C(n_411),
.Y(n_419)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_412),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_418),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g580 ( 
.A(n_416),
.B(n_418),
.C(n_581),
.Y(n_580)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_420),
.Y(n_418)
);

AOI21x1_ASAP7_75t_L g422 ( 
.A1(n_423),
.A2(n_467),
.B(n_578),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_424),
.B(n_426),
.Y(n_423)
);

NOR2xp67_ASAP7_75t_SL g578 ( 
.A(n_424),
.B(n_426),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_429),
.C(n_439),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_SL g573 ( 
.A(n_427),
.B(n_574),
.Y(n_573)
);

AOI21xp5_ASAP7_75t_L g574 ( 
.A1(n_429),
.A2(n_440),
.B(n_575),
.Y(n_574)
);

HB1xp67_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_SL g575 ( 
.A(n_430),
.B(n_440),
.Y(n_575)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx4_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVx5_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_438),
.Y(n_476)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_457),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_SL g555 ( 
.A(n_441),
.B(n_457),
.Y(n_555)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

BUFx3_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

INVx3_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

INVxp67_ASAP7_75t_SL g478 ( 
.A(n_448),
.Y(n_478)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

BUFx3_ASAP7_75t_L g481 ( 
.A(n_449),
.Y(n_481)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_453),
.Y(n_451)
);

OAI21xp33_ASAP7_75t_SL g474 ( 
.A1(n_452),
.A2(n_475),
.B(n_477),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_452),
.B(n_478),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_452),
.B(n_544),
.Y(n_543)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

INVx3_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

INVxp67_ASAP7_75t_L g509 ( 
.A(n_458),
.Y(n_509)
);

INVx3_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

INVx5_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

INVx4_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx4_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_466),
.Y(n_490)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_466),
.Y(n_534)
);

OAI21xp5_ASAP7_75t_L g467 ( 
.A1(n_468),
.A2(n_572),
.B(n_577),
.Y(n_467)
);

AOI21x1_ASAP7_75t_L g468 ( 
.A1(n_469),
.A2(n_552),
.B(n_571),
.Y(n_468)
);

OAI21x1_ASAP7_75t_L g469 ( 
.A1(n_470),
.A2(n_518),
.B(n_551),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_471),
.B(n_494),
.Y(n_470)
);

OR2x2_ASAP7_75t_L g551 ( 
.A(n_471),
.B(n_494),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_472),
.B(n_482),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g529 ( 
.A1(n_472),
.A2(n_473),
.B1(n_482),
.B2(n_483),
.Y(n_529)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

AOI21xp5_ASAP7_75t_L g487 ( 
.A1(n_477),
.A2(n_488),
.B(n_491),
.Y(n_487)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_480),
.Y(n_513)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

BUFx2_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

BUFx2_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

INVx1_ASAP7_75t_SL g488 ( 
.A(n_489),
.Y(n_488)
);

BUFx2_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

BUFx2_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_495),
.B(n_510),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_495),
.B(n_512),
.C(n_516),
.Y(n_553)
);

OAI22xp5_ASAP7_75t_L g495 ( 
.A1(n_496),
.A2(n_497),
.B1(n_506),
.B2(n_509),
.Y(n_495)
);

INVxp67_ASAP7_75t_L g528 ( 
.A(n_497),
.Y(n_528)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_499),
.Y(n_498)
);

BUFx3_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_500),
.Y(n_523)
);

INVx6_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

BUFx3_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

INVx4_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

BUFx2_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_L g510 ( 
.A1(n_511),
.A2(n_512),
.B1(n_516),
.B2(n_517),
.Y(n_510)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_511),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_512),
.Y(n_517)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_514),
.Y(n_568)
);

AOI21xp5_ASAP7_75t_L g518 ( 
.A1(n_519),
.A2(n_530),
.B(n_550),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_520),
.B(n_529),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_520),
.B(n_529),
.Y(n_550)
);

INVxp67_ASAP7_75t_L g521 ( 
.A(n_522),
.Y(n_521)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_523),
.Y(n_535)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_525),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_526),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_527),
.Y(n_526)
);

OAI21xp5_ASAP7_75t_SL g530 ( 
.A1(n_531),
.A2(n_539),
.B(n_549),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_532),
.B(n_538),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_532),
.B(n_538),
.Y(n_549)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_537),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_540),
.B(n_542),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_R g542 ( 
.A(n_543),
.B(n_546),
.Y(n_542)
);

INVx3_ASAP7_75t_L g544 ( 
.A(n_545),
.Y(n_544)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_547),
.Y(n_546)
);

HB1xp67_ASAP7_75t_L g547 ( 
.A(n_548),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_553),
.B(n_554),
.Y(n_552)
);

NOR2x1_ASAP7_75t_SL g571 ( 
.A(n_553),
.B(n_554),
.Y(n_571)
);

XNOR2xp5_ASAP7_75t_L g554 ( 
.A(n_555),
.B(n_556),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_555),
.B(n_567),
.C(n_570),
.Y(n_576)
);

AOI22xp5_ASAP7_75t_L g556 ( 
.A1(n_557),
.A2(n_567),
.B1(n_569),
.B2(n_570),
.Y(n_556)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_557),
.Y(n_570)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_560),
.Y(n_559)
);

INVx3_ASAP7_75t_L g560 ( 
.A(n_561),
.Y(n_560)
);

BUFx3_ASAP7_75t_L g561 ( 
.A(n_562),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_563),
.Y(n_562)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_565),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_566),
.Y(n_565)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_567),
.Y(n_569)
);

NOR2x1_ASAP7_75t_SL g572 ( 
.A(n_573),
.B(n_576),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_573),
.B(n_576),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_585),
.B(n_622),
.Y(n_584)
);

INVxp33_ASAP7_75t_SL g585 ( 
.A(n_586),
.Y(n_585)
);

NOR2xp67_ASAP7_75t_SL g586 ( 
.A(n_587),
.B(n_590),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_587),
.B(n_590),
.Y(n_623)
);

XNOR2xp5_ASAP7_75t_L g590 ( 
.A(n_591),
.B(n_619),
.Y(n_590)
);

OAI22xp5_ASAP7_75t_L g591 ( 
.A1(n_592),
.A2(n_602),
.B1(n_603),
.B2(n_618),
.Y(n_591)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_592),
.Y(n_618)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_595),
.Y(n_594)
);

INVxp67_ASAP7_75t_L g596 ( 
.A(n_597),
.Y(n_596)
);

INVx11_ASAP7_75t_L g598 ( 
.A(n_599),
.Y(n_598)
);

BUFx12f_ASAP7_75t_L g599 ( 
.A(n_600),
.Y(n_599)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_603),
.Y(n_602)
);

AOI22xp33_ASAP7_75t_SL g603 ( 
.A1(n_604),
.A2(n_605),
.B1(n_616),
.B2(n_617),
.Y(n_603)
);

INVx1_ASAP7_75t_SL g616 ( 
.A(n_604),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_605),
.Y(n_617)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_609),
.Y(n_608)
);

INVxp67_ASAP7_75t_L g609 ( 
.A(n_610),
.Y(n_609)
);

INVx3_ASAP7_75t_L g610 ( 
.A(n_611),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_612),
.Y(n_611)
);

INVx3_ASAP7_75t_L g613 ( 
.A(n_614),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_615),
.Y(n_614)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_623),
.Y(n_622)
);


endmodule