module fake_jpeg_56_n_167 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_167);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_167;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_SL g12 ( 
.A(n_8),
.B(n_10),
.Y(n_12)
);

INVx13_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

INVx6_ASAP7_75t_SL g16 ( 
.A(n_8),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_12),
.B(n_9),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_28),
.B(n_43),
.Y(n_60)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_29),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_31),
.Y(n_75)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_32),
.Y(n_66)
);

INVx4_ASAP7_75t_SL g33 ( 
.A(n_16),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_35),
.Y(n_79)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx4_ASAP7_75t_SL g37 ( 
.A(n_13),
.Y(n_37)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_37),
.Y(n_77)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_38),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_41),
.Y(n_87)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_12),
.B(n_0),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_45),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_22),
.B(n_6),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_46),
.B(n_47),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_48),
.B(n_51),
.Y(n_70)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_49),
.A2(n_55),
.B1(n_36),
.B2(n_40),
.Y(n_86)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_54),
.Y(n_59)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_52),
.B(n_53),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_26),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_29),
.A2(n_26),
.B1(n_14),
.B2(n_21),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_63),
.B(n_53),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_64),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_33),
.B(n_23),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_65),
.B(n_67),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_35),
.B(n_23),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_30),
.A2(n_14),
.B1(n_21),
.B2(n_15),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_69),
.B(n_71),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_39),
.A2(n_15),
.B1(n_2),
.B2(n_3),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_35),
.B(n_1),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_83),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_42),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_56),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_31),
.B(n_2),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_37),
.B(n_4),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_85),
.B(n_50),
.Y(n_91)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_66),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_91),
.B(n_100),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

AND2x2_ASAP7_75t_SL g94 ( 
.A(n_61),
.B(n_41),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_SL g121 ( 
.A(n_94),
.B(n_101),
.Y(n_121)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_103),
.Y(n_116)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_87),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_96),
.B(n_97),
.Y(n_112)
);

A2O1A1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_70),
.A2(n_52),
.B(n_47),
.C(n_54),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_98),
.A2(n_72),
.B1(n_87),
.B2(n_57),
.Y(n_118)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_66),
.Y(n_99)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_99),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_60),
.B(n_78),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_82),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_78),
.B(n_82),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_59),
.B(n_63),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_106),
.B(n_107),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_72),
.B(n_80),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_96),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_109),
.B(n_111),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_107),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_118),
.A2(n_114),
.B1(n_110),
.B2(n_99),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_106),
.A2(n_86),
.B1(n_79),
.B2(n_57),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_119),
.A2(n_104),
.B1(n_105),
.B2(n_79),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_102),
.B(n_75),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_120),
.B(n_75),
.Y(n_125)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_90),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_122),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_112),
.A2(n_98),
.B1(n_93),
.B2(n_94),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_124),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_125),
.B(n_108),
.Y(n_139)
);

OA22x2_ASAP7_75t_L g126 ( 
.A1(n_110),
.A2(n_104),
.B1(n_97),
.B2(n_92),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_126),
.B(n_129),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_94),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_128),
.B(n_114),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_111),
.B(n_101),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_113),
.A2(n_92),
.B(n_102),
.Y(n_130)
);

NOR3xp33_ASAP7_75t_L g134 ( 
.A(n_130),
.B(n_132),
.C(n_117),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_131),
.B(n_118),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_121),
.B(n_88),
.Y(n_132)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_133),
.Y(n_138)
);

OAI21x1_ASAP7_75t_SL g149 ( 
.A1(n_134),
.A2(n_143),
.B(n_126),
.Y(n_149)
);

NOR3xp33_ASAP7_75t_L g135 ( 
.A(n_130),
.B(n_117),
.C(n_89),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_135),
.B(n_139),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_137),
.A2(n_138),
.B1(n_127),
.B2(n_142),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_140),
.B(n_132),
.Y(n_147)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_123),
.Y(n_141)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_141),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_116),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_142),
.A2(n_124),
.B1(n_129),
.B2(n_128),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_145),
.A2(n_146),
.B1(n_150),
.B2(n_109),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_147),
.B(n_149),
.C(n_126),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_136),
.A2(n_126),
.B1(n_127),
.B2(n_108),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_148),
.B(n_140),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_151),
.B(n_153),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_152),
.B(n_154),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_147),
.B(n_115),
.C(n_122),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_152),
.B(n_147),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_156),
.B(n_150),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_158),
.B(n_159),
.Y(n_161)
);

NAND3xp33_ASAP7_75t_L g159 ( 
.A(n_157),
.B(n_144),
.C(n_145),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_155),
.B(n_115),
.Y(n_160)
);

AOI21x1_ASAP7_75t_SL g162 ( 
.A1(n_160),
.A2(n_156),
.B(n_68),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_162),
.B(n_58),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_161),
.A2(n_58),
.B(n_68),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_163),
.B(n_164),
.Y(n_165)
);

NAND3xp33_ASAP7_75t_SL g166 ( 
.A(n_165),
.B(n_62),
.C(n_74),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_62),
.Y(n_167)
);


endmodule