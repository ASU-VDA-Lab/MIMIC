module fake_netlist_6_1271_n_1121 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_1121);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1121;

wire n_992;
wire n_591;
wire n_435;
wire n_1115;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_881;
wire n_875;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_1008;
wire n_1027;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_1079;
wire n_362;
wire n_341;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_1033;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_1103;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_1061;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_994;
wire n_1072;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_396;
wire n_495;
wire n_1065;
wire n_815;
wire n_350;
wire n_1100;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_1042;
wire n_1071;
wire n_628;
wire n_1067;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_1074;
wire n_1032;
wire n_845;
wire n_255;
wire n_807;
wire n_1036;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_955;
wire n_865;
wire n_893;
wire n_214;
wire n_925;
wire n_485;
wire n_1099;
wire n_1026;
wire n_443;
wire n_1101;
wire n_246;
wire n_892;
wire n_768;
wire n_1097;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_1095;
wire n_573;
wire n_769;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_1120;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_447;
wire n_872;
wire n_300;
wire n_222;
wire n_718;
wire n_248;
wire n_517;
wire n_1018;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_1105;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_1078;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_1015;
wire n_836;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1057;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_235;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_1108;
wire n_387;
wire n_452;
wire n_658;
wire n_616;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_1119;
wire n_581;
wire n_428;
wire n_785;
wire n_761;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_631;
wire n_516;
wire n_720;
wire n_758;
wire n_525;
wire n_842;
wire n_1116;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_772;
wire n_656;
wire n_843;
wire n_989;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_1035;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_343;
wire n_844;
wire n_448;
wire n_953;
wire n_1017;
wire n_1004;
wire n_886;
wire n_1094;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_1083;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_1112;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_910;
wire n_901;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_236;
wire n_653;
wire n_887;
wire n_1117;
wire n_1087;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_1043;
wire n_1011;
wire n_224;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_1088;
wire n_708;
wire n_919;
wire n_1081;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_779;
wire n_800;
wire n_929;
wire n_460;
wire n_1084;
wire n_1104;
wire n_907;
wire n_854;
wire n_1058;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_1109;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_1054;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_1070;
wire n_1085;
wire n_232;
wire n_650;
wire n_998;
wire n_1046;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_1102;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1073;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_1041;
wire n_252;
wire n_757;
wire n_228;
wire n_594;
wire n_565;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_1062;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_1090;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_1068;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_964;
wire n_982;
wire n_831;
wire n_802;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_1075;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_237;
wire n_584;
wire n_1110;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_707;
wire n_322;
wire n_993;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_1064;
wire n_403;
wire n_1080;
wire n_723;
wire n_253;
wire n_634;
wire n_1051;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_249;
wire n_386;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_1086;
wire n_1066;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_970;
wire n_849;
wire n_1107;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_569;
wire n_1092;
wire n_441;
wire n_221;
wire n_811;
wire n_882;
wire n_1060;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_1111;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_1053;
wire n_530;
wire n_277;
wire n_520;
wire n_1029;
wire n_418;
wire n_1093;
wire n_618;
wire n_1055;
wire n_790;
wire n_1106;
wire n_582;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_1069;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_1052;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_285;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_920;
wire n_257;
wire n_903;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_286;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_1089;
wire n_401;
wire n_324;
wire n_766;
wire n_743;
wire n_816;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_205;
wire n_604;
wire n_848;
wire n_251;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_1096;
wire n_1063;
wire n_729;
wire n_1091;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_983;
wire n_288;
wire n_427;
wire n_1059;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_1077;
wire n_961;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_1082;
wire n_259;
wire n_1113;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_1098;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_956;
wire n_960;
wire n_841;
wire n_531;
wire n_827;
wire n_1001;
wire n_508;
wire n_361;
wire n_663;
wire n_856;
wire n_1050;
wire n_379;
wire n_778;
wire n_1025;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_664;
wire n_949;
wire n_678;
wire n_1007;
wire n_649;
wire n_283;

INVx1_ASAP7_75t_L g205 ( 
.A(n_96),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_90),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_132),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_190),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_25),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_36),
.Y(n_210)
);

BUFx8_ASAP7_75t_SL g211 ( 
.A(n_50),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_74),
.Y(n_212)
);

BUFx5_ASAP7_75t_L g213 ( 
.A(n_147),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_180),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_80),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_116),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_140),
.Y(n_217)
);

INVx2_ASAP7_75t_SL g218 ( 
.A(n_56),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_29),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_199),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_43),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_11),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_7),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_47),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_204),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_122),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_197),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_150),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_177),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_77),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_148),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_168),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_5),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_24),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_193),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_88),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_195),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_33),
.Y(n_238)
);

BUFx10_ASAP7_75t_L g239 ( 
.A(n_89),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_83),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_18),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_173),
.Y(n_242)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_163),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_188),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_178),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_181),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_153),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_106),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_81),
.Y(n_249)
);

BUFx2_ASAP7_75t_L g250 ( 
.A(n_5),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_57),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_176),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_154),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_137),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_189),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_6),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_87),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_84),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_14),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_182),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_174),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_198),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_28),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_45),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_0),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_145),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_107),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_175),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_112),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_27),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_65),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_15),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_16),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_233),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_233),
.Y(n_275)
);

INVxp67_ASAP7_75t_SL g276 ( 
.A(n_226),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_209),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_217),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_265),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_259),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_241),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_223),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_273),
.Y(n_283)
);

INVxp67_ASAP7_75t_SL g284 ( 
.A(n_235),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_219),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_219),
.Y(n_286)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_235),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_222),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_222),
.Y(n_289)
);

BUFx3_ASAP7_75t_L g290 ( 
.A(n_239),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_213),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_205),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_242),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_206),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_207),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_212),
.Y(n_296)
);

INVxp67_ASAP7_75t_SL g297 ( 
.A(n_243),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_216),
.Y(n_298)
);

INVxp67_ASAP7_75t_SL g299 ( 
.A(n_243),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_229),
.Y(n_300)
);

INVxp67_ASAP7_75t_SL g301 ( 
.A(n_231),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_213),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_234),
.Y(n_303)
);

INVxp33_ASAP7_75t_SL g304 ( 
.A(n_250),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_256),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_236),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_211),
.Y(n_307)
);

BUFx2_ASAP7_75t_L g308 ( 
.A(n_263),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_237),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_246),
.Y(n_310)
);

INVxp67_ASAP7_75t_SL g311 ( 
.A(n_252),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_264),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_268),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_211),
.Y(n_314)
);

INVxp67_ASAP7_75t_SL g315 ( 
.A(n_269),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_270),
.Y(n_316)
);

BUFx2_ASAP7_75t_SL g317 ( 
.A(n_255),
.Y(n_317)
);

BUFx10_ASAP7_75t_L g318 ( 
.A(n_272),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_270),
.Y(n_319)
);

INVxp67_ASAP7_75t_SL g320 ( 
.A(n_218),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_213),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_213),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_213),
.Y(n_323)
);

AND2x4_ASAP7_75t_L g324 ( 
.A(n_297),
.B(n_299),
.Y(n_324)
);

AND2x4_ASAP7_75t_L g325 ( 
.A(n_301),
.B(n_217),
.Y(n_325)
);

AND2x4_ASAP7_75t_L g326 ( 
.A(n_311),
.B(n_315),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_292),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_294),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_284),
.B(n_239),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_274),
.B(n_275),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_278),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_295),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_320),
.B(n_208),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_282),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_278),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_317),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_296),
.Y(n_337)
);

OA21x2_ASAP7_75t_L g338 ( 
.A1(n_321),
.A2(n_214),
.B(n_210),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_278),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_298),
.Y(n_340)
);

AND2x4_ASAP7_75t_L g341 ( 
.A(n_287),
.B(n_217),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_300),
.Y(n_342)
);

AND2x4_ASAP7_75t_L g343 ( 
.A(n_287),
.B(n_217),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_278),
.Y(n_344)
);

OA21x2_ASAP7_75t_L g345 ( 
.A1(n_321),
.A2(n_220),
.B(n_215),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_306),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_280),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_278),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_309),
.Y(n_349)
);

CKINVDCx11_ASAP7_75t_R g350 ( 
.A(n_307),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_304),
.A2(n_260),
.B1(n_224),
.B2(n_225),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_304),
.A2(n_248),
.B1(n_267),
.B2(n_266),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g353 ( 
.A(n_282),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_291),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_310),
.Y(n_355)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_291),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_285),
.Y(n_357)
);

AND2x2_ASAP7_75t_SL g358 ( 
.A(n_293),
.B(n_251),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_302),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_308),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_312),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_302),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_280),
.A2(n_247),
.B1(n_262),
.B2(n_261),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_285),
.Y(n_364)
);

BUFx8_ASAP7_75t_L g365 ( 
.A(n_308),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_290),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_307),
.A2(n_244),
.B1(n_258),
.B2(n_257),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_287),
.B(n_221),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_276),
.B(n_313),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_286),
.Y(n_370)
);

NAND2x1p5_ASAP7_75t_L g371 ( 
.A(n_322),
.B(n_251),
.Y(n_371)
);

AOI22x1_ASAP7_75t_SL g372 ( 
.A1(n_314),
.A2(n_227),
.B1(n_228),
.B2(n_230),
.Y(n_372)
);

OAI21x1_ASAP7_75t_L g373 ( 
.A1(n_323),
.A2(n_213),
.B(n_251),
.Y(n_373)
);

BUFx3_ASAP7_75t_L g374 ( 
.A(n_277),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_322),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_281),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_317),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_286),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_324),
.B(n_288),
.Y(n_379)
);

NAND2xp33_ASAP7_75t_SL g380 ( 
.A(n_351),
.B(n_303),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_336),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_375),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_336),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_354),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_358),
.B(n_303),
.Y(n_385)
);

INVx2_ASAP7_75t_SL g386 ( 
.A(n_329),
.Y(n_386)
);

BUFx3_ASAP7_75t_L g387 ( 
.A(n_324),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_354),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_329),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_359),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_359),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_375),
.Y(n_392)
);

INVx8_ASAP7_75t_L g393 ( 
.A(n_324),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_358),
.B(n_305),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_377),
.Y(n_395)
);

OAI22xp33_ASAP7_75t_L g396 ( 
.A1(n_352),
.A2(n_279),
.B1(n_305),
.B2(n_290),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_362),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_326),
.B(n_323),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_362),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_326),
.B(n_232),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_356),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_356),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_356),
.Y(n_403)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_331),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_364),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_364),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_331),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_364),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_333),
.B(n_318),
.Y(n_409)
);

INVx3_ASAP7_75t_L g410 ( 
.A(n_331),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_326),
.B(n_318),
.Y(n_411)
);

NOR2x1p5_ASAP7_75t_L g412 ( 
.A(n_377),
.B(n_283),
.Y(n_412)
);

NOR2x1p5_ASAP7_75t_L g413 ( 
.A(n_369),
.B(n_238),
.Y(n_413)
);

NOR2x1p5_ASAP7_75t_L g414 ( 
.A(n_374),
.B(n_240),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_331),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_364),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_364),
.Y(n_417)
);

INVx2_ASAP7_75t_SL g418 ( 
.A(n_341),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_360),
.B(n_318),
.Y(n_419)
);

INVx5_ASAP7_75t_L g420 ( 
.A(n_339),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_330),
.B(n_288),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_327),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_378),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_378),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_378),
.Y(n_425)
);

INVx2_ASAP7_75t_SL g426 ( 
.A(n_341),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_366),
.B(n_245),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_328),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_339),
.Y(n_429)
);

AND2x2_ASAP7_75t_SL g430 ( 
.A(n_338),
.B(n_251),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_378),
.Y(n_431)
);

INVx2_ASAP7_75t_SL g432 ( 
.A(n_341),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_378),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_363),
.B(n_325),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_332),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_357),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_330),
.B(n_319),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_337),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_340),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_367),
.A2(n_314),
.B1(n_249),
.B2(n_253),
.Y(n_440)
);

INVx4_ASAP7_75t_L g441 ( 
.A(n_339),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_357),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_357),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g444 ( 
.A(n_325),
.B(n_289),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_357),
.Y(n_445)
);

OR2x6_ASAP7_75t_L g446 ( 
.A(n_368),
.B(n_271),
.Y(n_446)
);

INVxp33_ASAP7_75t_SL g447 ( 
.A(n_334),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_342),
.Y(n_448)
);

INVx3_ASAP7_75t_L g449 ( 
.A(n_339),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_370),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_370),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_346),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_370),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_325),
.B(n_374),
.Y(n_454)
);

CKINVDCx16_ASAP7_75t_R g455 ( 
.A(n_380),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_387),
.B(n_338),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_418),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_386),
.B(n_353),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_418),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_426),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_426),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_401),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_386),
.B(n_365),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_432),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_389),
.B(n_349),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_381),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_432),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_454),
.B(n_355),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_381),
.B(n_347),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_387),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_383),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_383),
.B(n_347),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_393),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_395),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_454),
.B(n_361),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_387),
.B(n_376),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_395),
.B(n_372),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_393),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_421),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_447),
.Y(n_480)
);

INVxp67_ASAP7_75t_L g481 ( 
.A(n_444),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_421),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_437),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_437),
.Y(n_484)
);

CKINVDCx16_ASAP7_75t_R g485 ( 
.A(n_440),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_422),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_385),
.B(n_365),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_379),
.B(n_338),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_440),
.B(n_350),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_422),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_428),
.Y(n_491)
);

NAND2x1p5_ASAP7_75t_L g492 ( 
.A(n_379),
.B(n_343),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g493 ( 
.A(n_400),
.Y(n_493)
);

OR2x2_ASAP7_75t_L g494 ( 
.A(n_394),
.B(n_345),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_428),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_435),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_438),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_438),
.Y(n_498)
);

OAI21xp5_ASAP7_75t_L g499 ( 
.A1(n_430),
.A2(n_345),
.B(n_373),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_409),
.B(n_365),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_411),
.B(n_345),
.Y(n_501)
);

INVxp67_ASAP7_75t_L g502 ( 
.A(n_444),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_439),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_447),
.B(n_350),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_448),
.Y(n_505)
);

INVx2_ASAP7_75t_SL g506 ( 
.A(n_414),
.Y(n_506)
);

INVxp33_ASAP7_75t_L g507 ( 
.A(n_419),
.Y(n_507)
);

XOR2x2_ASAP7_75t_L g508 ( 
.A(n_434),
.B(n_0),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_396),
.B(n_427),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_448),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_398),
.B(n_343),
.Y(n_511)
);

CKINVDCx16_ASAP7_75t_R g512 ( 
.A(n_452),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_393),
.B(n_343),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_452),
.Y(n_514)
);

NAND2x1p5_ASAP7_75t_L g515 ( 
.A(n_436),
.B(n_373),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_SL g516 ( 
.A(n_393),
.B(n_430),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g517 ( 
.A(n_430),
.B(n_254),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_393),
.B(n_370),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_382),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_453),
.B(n_271),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_412),
.B(n_316),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_453),
.B(n_271),
.Y(n_522)
);

NOR2xp67_ASAP7_75t_L g523 ( 
.A(n_436),
.B(n_34),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_382),
.Y(n_524)
);

AND2x4_ASAP7_75t_L g525 ( 
.A(n_414),
.B(n_289),
.Y(n_525)
);

INVxp33_ASAP7_75t_L g526 ( 
.A(n_413),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_392),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_451),
.B(n_271),
.Y(n_528)
);

INVxp33_ASAP7_75t_L g529 ( 
.A(n_413),
.Y(n_529)
);

AND2x4_ASAP7_75t_L g530 ( 
.A(n_412),
.B(n_442),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_392),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_399),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_399),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_384),
.Y(n_534)
);

INVxp67_ASAP7_75t_L g535 ( 
.A(n_446),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_384),
.Y(n_536)
);

AND2x4_ASAP7_75t_L g537 ( 
.A(n_442),
.B(n_319),
.Y(n_537)
);

AOI22xp33_ASAP7_75t_L g538 ( 
.A1(n_508),
.A2(n_488),
.B1(n_509),
.B2(n_479),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_493),
.B(n_443),
.Y(n_539)
);

AOI22xp33_ASAP7_75t_L g540 ( 
.A1(n_482),
.A2(n_388),
.B1(n_391),
.B2(n_390),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_537),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_481),
.B(n_502),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_481),
.B(n_443),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_537),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_512),
.B(n_445),
.Y(n_545)
);

BUFx3_ASAP7_75t_L g546 ( 
.A(n_466),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_502),
.B(n_451),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_507),
.B(n_445),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_486),
.B(n_450),
.Y(n_549)
);

AND2x6_ASAP7_75t_SL g550 ( 
.A(n_500),
.B(n_446),
.Y(n_550)
);

AOI22xp5_ASAP7_75t_L g551 ( 
.A1(n_501),
.A2(n_446),
.B1(n_450),
.B2(n_406),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_490),
.B(n_388),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_516),
.B(n_405),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_470),
.Y(n_554)
);

NAND2xp33_ASAP7_75t_L g555 ( 
.A(n_473),
.B(n_405),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_462),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_491),
.B(n_390),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_458),
.B(n_446),
.Y(n_558)
);

NAND3xp33_ASAP7_75t_L g559 ( 
.A(n_474),
.B(n_446),
.C(n_408),
.Y(n_559)
);

HB1xp67_ASAP7_75t_L g560 ( 
.A(n_492),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_495),
.B(n_391),
.Y(n_561)
);

INVx6_ASAP7_75t_L g562 ( 
.A(n_530),
.Y(n_562)
);

AOI22xp33_ASAP7_75t_L g563 ( 
.A1(n_483),
.A2(n_397),
.B1(n_403),
.B2(n_402),
.Y(n_563)
);

OR2x6_ASAP7_75t_L g564 ( 
.A(n_506),
.B(n_406),
.Y(n_564)
);

AOI22x1_ASAP7_75t_L g565 ( 
.A1(n_494),
.A2(n_515),
.B1(n_517),
.B2(n_499),
.Y(n_565)
);

AND2x2_ASAP7_75t_SL g566 ( 
.A(n_516),
.B(n_408),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_473),
.B(n_416),
.Y(n_567)
);

INVxp67_ASAP7_75t_L g568 ( 
.A(n_521),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_465),
.B(n_402),
.Y(n_569)
);

AOI22xp5_ASAP7_75t_L g570 ( 
.A1(n_530),
.A2(n_476),
.B1(n_484),
.B2(n_459),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_496),
.B(n_403),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_532),
.Y(n_572)
);

HB1xp67_ASAP7_75t_L g573 ( 
.A(n_492),
.Y(n_573)
);

AND2x4_ASAP7_75t_L g574 ( 
.A(n_468),
.B(n_416),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_497),
.B(n_417),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_533),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_534),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_536),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_526),
.B(n_417),
.Y(n_579)
);

AOI22xp5_ASAP7_75t_L g580 ( 
.A1(n_457),
.A2(n_424),
.B1(n_423),
.B2(n_433),
.Y(n_580)
);

INVx2_ASAP7_75t_SL g581 ( 
.A(n_525),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_498),
.B(n_423),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_529),
.B(n_424),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_471),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_480),
.B(n_404),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_503),
.B(n_425),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_519),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_524),
.Y(n_588)
);

BUFx3_ASAP7_75t_L g589 ( 
.A(n_525),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_505),
.B(n_431),
.Y(n_590)
);

AOI21xp5_ASAP7_75t_L g591 ( 
.A1(n_513),
.A2(n_441),
.B(n_433),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_473),
.B(n_431),
.Y(n_592)
);

OAI22xp5_ASAP7_75t_L g593 ( 
.A1(n_511),
.A2(n_456),
.B1(n_535),
.B2(n_513),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_527),
.Y(n_594)
);

INVx2_ASAP7_75t_SL g595 ( 
.A(n_475),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_531),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_510),
.B(n_449),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_514),
.B(n_449),
.Y(n_598)
);

AOI22xp5_ASAP7_75t_L g599 ( 
.A1(n_460),
.A2(n_404),
.B1(n_410),
.B2(n_449),
.Y(n_599)
);

OAI22xp33_ASAP7_75t_L g600 ( 
.A1(n_485),
.A2(n_371),
.B1(n_449),
.B2(n_404),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_478),
.B(n_407),
.Y(n_601)
);

INVx2_ASAP7_75t_SL g602 ( 
.A(n_469),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_461),
.Y(n_603)
);

INVxp67_ASAP7_75t_SL g604 ( 
.A(n_574),
.Y(n_604)
);

INVx3_ASAP7_75t_L g605 ( 
.A(n_574),
.Y(n_605)
);

BUFx2_ASAP7_75t_L g606 ( 
.A(n_584),
.Y(n_606)
);

HB1xp67_ASAP7_75t_L g607 ( 
.A(n_595),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_572),
.Y(n_608)
);

INVx4_ASAP7_75t_L g609 ( 
.A(n_562),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_569),
.B(n_511),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_R g611 ( 
.A(n_602),
.B(n_455),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_576),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_542),
.B(n_464),
.Y(n_613)
);

AND2x4_ASAP7_75t_L g614 ( 
.A(n_589),
.B(n_467),
.Y(n_614)
);

OR2x6_ASAP7_75t_L g615 ( 
.A(n_546),
.B(n_463),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_550),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_577),
.Y(n_617)
);

NAND3xp33_ASAP7_75t_SL g618 ( 
.A(n_538),
.B(n_487),
.C(n_472),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_578),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_568),
.B(n_478),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_568),
.B(n_535),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_548),
.B(n_587),
.Y(n_622)
);

BUFx2_ASAP7_75t_L g623 ( 
.A(n_564),
.Y(n_623)
);

AND2x4_ASAP7_75t_L g624 ( 
.A(n_581),
.B(n_478),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_548),
.B(n_456),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_556),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_588),
.Y(n_627)
);

OR2x6_ASAP7_75t_L g628 ( 
.A(n_562),
.B(n_515),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_538),
.B(n_477),
.Y(n_629)
);

BUFx3_ASAP7_75t_L g630 ( 
.A(n_562),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_594),
.Y(n_631)
);

BUFx2_ASAP7_75t_L g632 ( 
.A(n_564),
.Y(n_632)
);

O2A1O1Ixp33_ASAP7_75t_L g633 ( 
.A1(n_600),
.A2(n_499),
.B(n_522),
.C(n_520),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_552),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_603),
.B(n_518),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_557),
.Y(n_636)
);

BUFx3_ASAP7_75t_L g637 ( 
.A(n_564),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_566),
.B(n_523),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_561),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_566),
.B(n_407),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_596),
.B(n_410),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_543),
.Y(n_642)
);

HB1xp67_ASAP7_75t_L g643 ( 
.A(n_541),
.Y(n_643)
);

INVxp67_ASAP7_75t_L g644 ( 
.A(n_545),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_547),
.B(n_410),
.Y(n_645)
);

BUFx6f_ASAP7_75t_L g646 ( 
.A(n_554),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_585),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_544),
.B(n_504),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_539),
.B(n_528),
.Y(n_649)
);

INVx2_ASAP7_75t_SL g650 ( 
.A(n_579),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_571),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_575),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_579),
.B(n_489),
.Y(n_653)
);

HB1xp67_ASAP7_75t_L g654 ( 
.A(n_560),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_582),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_586),
.Y(n_656)
);

BUFx6f_ASAP7_75t_L g657 ( 
.A(n_601),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_590),
.Y(n_658)
);

INVx6_ASAP7_75t_L g659 ( 
.A(n_583),
.Y(n_659)
);

NOR2x1_ASAP7_75t_R g660 ( 
.A(n_549),
.B(n_441),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_597),
.Y(n_661)
);

INVxp67_ASAP7_75t_L g662 ( 
.A(n_583),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_598),
.Y(n_663)
);

BUFx6f_ASAP7_75t_L g664 ( 
.A(n_567),
.Y(n_664)
);

INVxp67_ASAP7_75t_SL g665 ( 
.A(n_560),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_565),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_573),
.Y(n_667)
);

AOI21xp5_ASAP7_75t_L g668 ( 
.A1(n_610),
.A2(n_593),
.B(n_555),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_653),
.B(n_558),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_608),
.Y(n_670)
);

OAI21x1_ASAP7_75t_L g671 ( 
.A1(n_645),
.A2(n_591),
.B(n_553),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_662),
.B(n_570),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_662),
.B(n_558),
.Y(n_673)
);

OAI21x1_ASAP7_75t_L g674 ( 
.A1(n_633),
.A2(n_592),
.B(n_551),
.Y(n_674)
);

AOI21xp5_ASAP7_75t_L g675 ( 
.A1(n_638),
.A2(n_600),
.B(n_559),
.Y(n_675)
);

AO21x1_ASAP7_75t_L g676 ( 
.A1(n_638),
.A2(n_599),
.B(n_580),
.Y(n_676)
);

OAI21x1_ASAP7_75t_L g677 ( 
.A1(n_641),
.A2(n_640),
.B(n_625),
.Y(n_677)
);

OAI21xp5_ASAP7_75t_L g678 ( 
.A1(n_666),
.A2(n_563),
.B(n_540),
.Y(n_678)
);

OA22x2_ASAP7_75t_L g679 ( 
.A1(n_629),
.A2(n_573),
.B1(n_2),
.B2(n_3),
.Y(n_679)
);

O2A1O1Ixp5_ASAP7_75t_L g680 ( 
.A1(n_640),
.A2(n_441),
.B(n_348),
.C(n_344),
.Y(n_680)
);

OAI21xp5_ASAP7_75t_SL g681 ( 
.A1(n_618),
.A2(n_644),
.B(n_621),
.Y(n_681)
);

AOI21xp5_ASAP7_75t_L g682 ( 
.A1(n_649),
.A2(n_441),
.B(n_563),
.Y(n_682)
);

OAI21x1_ASAP7_75t_L g683 ( 
.A1(n_655),
.A2(n_540),
.B(n_344),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_650),
.B(n_371),
.Y(n_684)
);

INVx3_ASAP7_75t_L g685 ( 
.A(n_628),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_642),
.B(n_371),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_617),
.Y(n_687)
);

AOI21xp5_ASAP7_75t_L g688 ( 
.A1(n_635),
.A2(n_415),
.B(n_407),
.Y(n_688)
);

OAI21xp5_ASAP7_75t_L g689 ( 
.A1(n_661),
.A2(n_348),
.B(n_335),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_622),
.B(n_1),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_612),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_613),
.B(n_1),
.Y(n_692)
);

INVx2_ASAP7_75t_SL g693 ( 
.A(n_606),
.Y(n_693)
);

BUFx6f_ASAP7_75t_L g694 ( 
.A(n_630),
.Y(n_694)
);

AOI21xp5_ASAP7_75t_L g695 ( 
.A1(n_628),
.A2(n_415),
.B(n_407),
.Y(n_695)
);

AOI21x1_ASAP7_75t_L g696 ( 
.A1(n_663),
.A2(n_335),
.B(n_407),
.Y(n_696)
);

OA22x2_ASAP7_75t_L g697 ( 
.A1(n_647),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_634),
.B(n_415),
.Y(n_698)
);

AND2x2_ASAP7_75t_SL g699 ( 
.A(n_623),
.B(n_4),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_617),
.Y(n_700)
);

BUFx4_ASAP7_75t_SL g701 ( 
.A(n_615),
.Y(n_701)
);

OAI21xp5_ASAP7_75t_L g702 ( 
.A1(n_652),
.A2(n_420),
.B(n_415),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_627),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_631),
.Y(n_704)
);

AOI21xp33_ASAP7_75t_L g705 ( 
.A1(n_651),
.A2(n_6),
.B(n_7),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_619),
.Y(n_706)
);

OAI21x1_ASAP7_75t_L g707 ( 
.A1(n_655),
.A2(n_656),
.B(n_620),
.Y(n_707)
);

O2A1O1Ixp5_ASAP7_75t_L g708 ( 
.A1(n_621),
.A2(n_8),
.B(n_9),
.C(n_10),
.Y(n_708)
);

OAI21x1_ASAP7_75t_L g709 ( 
.A1(n_656),
.A2(n_619),
.B(n_626),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_644),
.B(n_643),
.Y(n_710)
);

OAI21x1_ASAP7_75t_L g711 ( 
.A1(n_626),
.A2(n_429),
.B(n_415),
.Y(n_711)
);

AOI21x1_ASAP7_75t_L g712 ( 
.A1(n_658),
.A2(n_429),
.B(n_420),
.Y(n_712)
);

OAI21xp5_ASAP7_75t_L g713 ( 
.A1(n_636),
.A2(n_420),
.B(n_429),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_659),
.B(n_8),
.Y(n_714)
);

BUFx3_ASAP7_75t_L g715 ( 
.A(n_607),
.Y(n_715)
);

INVx3_ASAP7_75t_L g716 ( 
.A(n_628),
.Y(n_716)
);

OAI22xp5_ASAP7_75t_L g717 ( 
.A1(n_604),
.A2(n_429),
.B1(n_10),
.B2(n_11),
.Y(n_717)
);

AOI21x1_ASAP7_75t_SL g718 ( 
.A1(n_624),
.A2(n_9),
.B(n_12),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_639),
.B(n_12),
.Y(n_719)
);

AOI21xp5_ASAP7_75t_SL g720 ( 
.A1(n_604),
.A2(n_660),
.B(n_624),
.Y(n_720)
);

AOI21xp5_ASAP7_75t_L g721 ( 
.A1(n_665),
.A2(n_37),
.B(n_35),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_643),
.Y(n_722)
);

AOI21xp5_ASAP7_75t_L g723 ( 
.A1(n_665),
.A2(n_39),
.B(n_38),
.Y(n_723)
);

AOI21xp33_ASAP7_75t_L g724 ( 
.A1(n_615),
.A2(n_13),
.B(n_14),
.Y(n_724)
);

BUFx10_ASAP7_75t_L g725 ( 
.A(n_614),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_659),
.B(n_13),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_611),
.B(n_15),
.Y(n_727)
);

INVx2_ASAP7_75t_SL g728 ( 
.A(n_715),
.Y(n_728)
);

AOI21xp5_ASAP7_75t_L g729 ( 
.A1(n_668),
.A2(n_605),
.B(n_646),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_669),
.B(n_667),
.Y(n_730)
);

OAI21x1_ASAP7_75t_L g731 ( 
.A1(n_671),
.A2(n_605),
.B(n_654),
.Y(n_731)
);

AOI21x1_ASAP7_75t_L g732 ( 
.A1(n_696),
.A2(n_632),
.B(n_654),
.Y(n_732)
);

AOI221xp5_ASAP7_75t_L g733 ( 
.A1(n_724),
.A2(n_705),
.B1(n_717),
.B2(n_681),
.C(n_708),
.Y(n_733)
);

BUFx5_ASAP7_75t_L g734 ( 
.A(n_706),
.Y(n_734)
);

AOI21xp5_ASAP7_75t_L g735 ( 
.A1(n_678),
.A2(n_646),
.B(n_657),
.Y(n_735)
);

OAI21x1_ASAP7_75t_SL g736 ( 
.A1(n_676),
.A2(n_609),
.B(n_659),
.Y(n_736)
);

AO21x1_ASAP7_75t_L g737 ( 
.A1(n_717),
.A2(n_614),
.B(n_609),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_670),
.Y(n_738)
);

AND2x2_ASAP7_75t_L g739 ( 
.A(n_710),
.B(n_648),
.Y(n_739)
);

AO31x2_ASAP7_75t_L g740 ( 
.A1(n_688),
.A2(n_657),
.A3(n_664),
.B(n_646),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_701),
.Y(n_741)
);

HB1xp67_ASAP7_75t_L g742 ( 
.A(n_722),
.Y(n_742)
);

OA21x2_ASAP7_75t_L g743 ( 
.A1(n_674),
.A2(n_607),
.B(n_616),
.Y(n_743)
);

A2O1A1Ixp33_ASAP7_75t_L g744 ( 
.A1(n_675),
.A2(n_681),
.B(n_678),
.C(n_690),
.Y(n_744)
);

NAND3xp33_ASAP7_75t_L g745 ( 
.A(n_724),
.B(n_615),
.C(n_646),
.Y(n_745)
);

AOI21xp5_ASAP7_75t_L g746 ( 
.A1(n_682),
.A2(n_657),
.B(n_664),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_673),
.B(n_672),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_687),
.Y(n_748)
);

OAI21x1_ASAP7_75t_SL g749 ( 
.A1(n_702),
.A2(n_657),
.B(n_637),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_714),
.B(n_611),
.Y(n_750)
);

AOI22xp33_ASAP7_75t_L g751 ( 
.A1(n_679),
.A2(n_637),
.B1(n_664),
.B2(n_630),
.Y(n_751)
);

AOI21xp5_ASAP7_75t_L g752 ( 
.A1(n_702),
.A2(n_664),
.B(n_41),
.Y(n_752)
);

NOR4xp25_ASAP7_75t_L g753 ( 
.A(n_705),
.B(n_16),
.C(n_17),
.D(n_18),
.Y(n_753)
);

AO21x2_ASAP7_75t_L g754 ( 
.A1(n_713),
.A2(n_42),
.B(n_40),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_692),
.B(n_17),
.Y(n_755)
);

A2O1A1Ixp33_ASAP7_75t_L g756 ( 
.A1(n_726),
.A2(n_19),
.B(n_20),
.C(n_21),
.Y(n_756)
);

O2A1O1Ixp33_ASAP7_75t_SL g757 ( 
.A1(n_719),
.A2(n_686),
.B(n_698),
.C(n_727),
.Y(n_757)
);

OR2x6_ASAP7_75t_L g758 ( 
.A(n_720),
.B(n_44),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_719),
.B(n_19),
.Y(n_759)
);

AOI21xp5_ASAP7_75t_L g760 ( 
.A1(n_713),
.A2(n_203),
.B(n_48),
.Y(n_760)
);

AOI221x1_ASAP7_75t_L g761 ( 
.A1(n_721),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.C(n_23),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_691),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_703),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_699),
.B(n_22),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_709),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_704),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_700),
.Y(n_767)
);

AO21x1_ASAP7_75t_L g768 ( 
.A1(n_723),
.A2(n_23),
.B(n_24),
.Y(n_768)
);

AND2x2_ASAP7_75t_L g769 ( 
.A(n_679),
.B(n_25),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_707),
.Y(n_770)
);

AOI21xp5_ASAP7_75t_L g771 ( 
.A1(n_689),
.A2(n_202),
.B(n_121),
.Y(n_771)
);

BUFx4f_ASAP7_75t_L g772 ( 
.A(n_694),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_685),
.Y(n_773)
);

AO31x2_ASAP7_75t_L g774 ( 
.A1(n_695),
.A2(n_26),
.A3(n_27),
.B(n_28),
.Y(n_774)
);

NAND3xp33_ASAP7_75t_L g775 ( 
.A(n_693),
.B(n_26),
.C(n_29),
.Y(n_775)
);

A2O1A1Ixp33_ASAP7_75t_L g776 ( 
.A1(n_685),
.A2(n_30),
.B(n_31),
.C(n_32),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_716),
.Y(n_777)
);

OAI21x1_ASAP7_75t_L g778 ( 
.A1(n_711),
.A2(n_124),
.B(n_200),
.Y(n_778)
);

BUFx6f_ASAP7_75t_L g779 ( 
.A(n_694),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_684),
.B(n_30),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_694),
.B(n_46),
.Y(n_781)
);

AND2x2_ASAP7_75t_L g782 ( 
.A(n_697),
.B(n_725),
.Y(n_782)
);

INVx5_ASAP7_75t_L g783 ( 
.A(n_725),
.Y(n_783)
);

AOI221x1_ASAP7_75t_L g784 ( 
.A1(n_689),
.A2(n_31),
.B1(n_32),
.B2(n_49),
.C(n_51),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_697),
.B(n_52),
.Y(n_785)
);

OA21x2_ASAP7_75t_L g786 ( 
.A1(n_677),
.A2(n_53),
.B(n_54),
.Y(n_786)
);

AOI21xp5_ASAP7_75t_L g787 ( 
.A1(n_698),
.A2(n_55),
.B(n_58),
.Y(n_787)
);

BUFx2_ASAP7_75t_L g788 ( 
.A(n_716),
.Y(n_788)
);

BUFx10_ASAP7_75t_L g789 ( 
.A(n_718),
.Y(n_789)
);

A2O1A1Ixp33_ASAP7_75t_L g790 ( 
.A1(n_680),
.A2(n_59),
.B(n_60),
.C(n_61),
.Y(n_790)
);

AO31x2_ASAP7_75t_L g791 ( 
.A1(n_712),
.A2(n_201),
.A3(n_63),
.B(n_64),
.Y(n_791)
);

OAI21x1_ASAP7_75t_L g792 ( 
.A1(n_683),
.A2(n_62),
.B(n_66),
.Y(n_792)
);

NOR2x1_ASAP7_75t_SL g793 ( 
.A(n_712),
.B(n_67),
.Y(n_793)
);

NOR2x1_ASAP7_75t_L g794 ( 
.A(n_720),
.B(n_68),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_669),
.B(n_69),
.Y(n_795)
);

AOI22xp33_ASAP7_75t_SL g796 ( 
.A1(n_764),
.A2(n_70),
.B1(n_71),
.B2(n_72),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_748),
.Y(n_797)
);

CKINVDCx6p67_ASAP7_75t_R g798 ( 
.A(n_783),
.Y(n_798)
);

NAND2x1p5_ASAP7_75t_L g799 ( 
.A(n_794),
.B(n_73),
.Y(n_799)
);

INVx3_ASAP7_75t_L g800 ( 
.A(n_779),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_747),
.B(n_75),
.Y(n_801)
);

OAI22xp5_ASAP7_75t_L g802 ( 
.A1(n_751),
.A2(n_76),
.B1(n_78),
.B2(n_79),
.Y(n_802)
);

INVx1_ASAP7_75t_SL g803 ( 
.A(n_742),
.Y(n_803)
);

INVx8_ASAP7_75t_L g804 ( 
.A(n_758),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_767),
.Y(n_805)
);

AOI22xp33_ASAP7_75t_L g806 ( 
.A1(n_733),
.A2(n_82),
.B1(n_85),
.B2(n_86),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_741),
.Y(n_807)
);

INVx1_ASAP7_75t_SL g808 ( 
.A(n_788),
.Y(n_808)
);

CKINVDCx20_ASAP7_75t_R g809 ( 
.A(n_750),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_738),
.Y(n_810)
);

AOI22xp33_ASAP7_75t_SL g811 ( 
.A1(n_785),
.A2(n_91),
.B1(n_92),
.B2(n_93),
.Y(n_811)
);

OAI22xp5_ASAP7_75t_L g812 ( 
.A1(n_744),
.A2(n_94),
.B1(n_95),
.B2(n_97),
.Y(n_812)
);

NAND2x1p5_ASAP7_75t_L g813 ( 
.A(n_731),
.B(n_98),
.Y(n_813)
);

CKINVDCx6p67_ASAP7_75t_R g814 ( 
.A(n_783),
.Y(n_814)
);

INVxp67_ASAP7_75t_SL g815 ( 
.A(n_730),
.Y(n_815)
);

AOI22xp5_ASAP7_75t_L g816 ( 
.A1(n_795),
.A2(n_99),
.B1(n_100),
.B2(n_101),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_762),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_763),
.Y(n_818)
);

BUFx12f_ASAP7_75t_L g819 ( 
.A(n_779),
.Y(n_819)
);

AND2x2_ASAP7_75t_L g820 ( 
.A(n_739),
.B(n_102),
.Y(n_820)
);

AOI22xp33_ASAP7_75t_SL g821 ( 
.A1(n_769),
.A2(n_103),
.B1(n_104),
.B2(n_105),
.Y(n_821)
);

OAI22xp5_ASAP7_75t_L g822 ( 
.A1(n_745),
.A2(n_782),
.B1(n_755),
.B2(n_759),
.Y(n_822)
);

OAI22xp5_ASAP7_75t_L g823 ( 
.A1(n_728),
.A2(n_108),
.B1(n_109),
.B2(n_110),
.Y(n_823)
);

AOI22xp33_ASAP7_75t_L g824 ( 
.A1(n_768),
.A2(n_111),
.B1(n_113),
.B2(n_114),
.Y(n_824)
);

OAI21xp5_ASAP7_75t_L g825 ( 
.A1(n_752),
.A2(n_115),
.B(n_117),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_779),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_766),
.Y(n_827)
);

BUFx10_ASAP7_75t_L g828 ( 
.A(n_781),
.Y(n_828)
);

OAI21xp5_ASAP7_75t_L g829 ( 
.A1(n_771),
.A2(n_118),
.B(n_119),
.Y(n_829)
);

OAI22x1_ASAP7_75t_L g830 ( 
.A1(n_775),
.A2(n_120),
.B1(n_123),
.B2(n_125),
.Y(n_830)
);

INVx2_ASAP7_75t_SL g831 ( 
.A(n_772),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_773),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_774),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_774),
.Y(n_834)
);

AOI22xp33_ASAP7_75t_L g835 ( 
.A1(n_737),
.A2(n_126),
.B1(n_127),
.B2(n_128),
.Y(n_835)
);

AOI22xp33_ASAP7_75t_L g836 ( 
.A1(n_758),
.A2(n_129),
.B1(n_130),
.B2(n_131),
.Y(n_836)
);

OAI22xp33_ASAP7_75t_L g837 ( 
.A1(n_761),
.A2(n_133),
.B1(n_134),
.B2(n_135),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_734),
.Y(n_838)
);

INVx5_ASAP7_75t_L g839 ( 
.A(n_789),
.Y(n_839)
);

INVx3_ASAP7_75t_L g840 ( 
.A(n_777),
.Y(n_840)
);

AOI22xp33_ASAP7_75t_L g841 ( 
.A1(n_789),
.A2(n_136),
.B1(n_138),
.B2(n_139),
.Y(n_841)
);

HB1xp67_ASAP7_75t_L g842 ( 
.A(n_735),
.Y(n_842)
);

INVxp67_ASAP7_75t_SL g843 ( 
.A(n_734),
.Y(n_843)
);

CKINVDCx11_ASAP7_75t_R g844 ( 
.A(n_734),
.Y(n_844)
);

HB1xp67_ASAP7_75t_SL g845 ( 
.A(n_772),
.Y(n_845)
);

NAND2x1p5_ASAP7_75t_L g846 ( 
.A(n_783),
.B(n_141),
.Y(n_846)
);

AOI22xp33_ASAP7_75t_L g847 ( 
.A1(n_736),
.A2(n_142),
.B1(n_143),
.B2(n_144),
.Y(n_847)
);

HB1xp67_ASAP7_75t_L g848 ( 
.A(n_740),
.Y(n_848)
);

AOI22xp33_ASAP7_75t_L g849 ( 
.A1(n_780),
.A2(n_146),
.B1(n_149),
.B2(n_151),
.Y(n_849)
);

AOI22xp33_ASAP7_75t_SL g850 ( 
.A1(n_760),
.A2(n_152),
.B1(n_155),
.B2(n_156),
.Y(n_850)
);

BUFx12f_ASAP7_75t_L g851 ( 
.A(n_756),
.Y(n_851)
);

OAI21xp5_ASAP7_75t_L g852 ( 
.A1(n_729),
.A2(n_157),
.B(n_158),
.Y(n_852)
);

CKINVDCx11_ASAP7_75t_R g853 ( 
.A(n_734),
.Y(n_853)
);

BUFx2_ASAP7_75t_SL g854 ( 
.A(n_743),
.Y(n_854)
);

BUFx2_ASAP7_75t_L g855 ( 
.A(n_740),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_810),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_817),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_818),
.Y(n_858)
);

AOI211xp5_ASAP7_75t_L g859 ( 
.A1(n_822),
.A2(n_753),
.B(n_776),
.C(n_757),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_827),
.Y(n_860)
);

HB1xp67_ASAP7_75t_L g861 ( 
.A(n_803),
.Y(n_861)
);

INVx2_ASAP7_75t_SL g862 ( 
.A(n_803),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_805),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_833),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_834),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_842),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_838),
.Y(n_867)
);

AOI221xp5_ASAP7_75t_L g868 ( 
.A1(n_837),
.A2(n_787),
.B1(n_749),
.B2(n_746),
.C(n_770),
.Y(n_868)
);

INVx3_ASAP7_75t_L g869 ( 
.A(n_844),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_848),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_797),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_855),
.Y(n_872)
);

OAI21x1_ASAP7_75t_L g873 ( 
.A1(n_813),
.A2(n_732),
.B(n_792),
.Y(n_873)
);

OAI222xp33_ASAP7_75t_L g874 ( 
.A1(n_811),
.A2(n_784),
.B1(n_765),
.B2(n_754),
.C1(n_743),
.C2(n_791),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_815),
.B(n_854),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_832),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_808),
.Y(n_877)
);

BUFx4f_ASAP7_75t_L g878 ( 
.A(n_804),
.Y(n_878)
);

HB1xp67_ASAP7_75t_L g879 ( 
.A(n_808),
.Y(n_879)
);

INVx2_ASAP7_75t_SL g880 ( 
.A(n_798),
.Y(n_880)
);

AND2x4_ASAP7_75t_L g881 ( 
.A(n_843),
.B(n_740),
.Y(n_881)
);

HB1xp67_ASAP7_75t_L g882 ( 
.A(n_840),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_840),
.Y(n_883)
);

INVx2_ASAP7_75t_SL g884 ( 
.A(n_814),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_839),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_839),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_839),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_839),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_853),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_800),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_800),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_846),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_846),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_851),
.B(n_786),
.Y(n_894)
);

INVx3_ASAP7_75t_L g895 ( 
.A(n_804),
.Y(n_895)
);

BUFx8_ASAP7_75t_L g896 ( 
.A(n_819),
.Y(n_896)
);

HB1xp67_ASAP7_75t_L g897 ( 
.A(n_826),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_799),
.Y(n_898)
);

AOI221xp5_ASAP7_75t_L g899 ( 
.A1(n_830),
.A2(n_790),
.B1(n_791),
.B2(n_786),
.C(n_162),
.Y(n_899)
);

AOI222xp33_ASAP7_75t_L g900 ( 
.A1(n_829),
.A2(n_793),
.B1(n_778),
.B2(n_161),
.C1(n_164),
.C2(n_165),
.Y(n_900)
);

HB1xp67_ASAP7_75t_L g901 ( 
.A(n_870),
.Y(n_901)
);

OR2x2_ASAP7_75t_L g902 ( 
.A(n_861),
.B(n_791),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_856),
.Y(n_903)
);

AO21x2_ASAP7_75t_L g904 ( 
.A1(n_864),
.A2(n_825),
.B(n_852),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_865),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_866),
.B(n_828),
.Y(n_906)
);

BUFx2_ASAP7_75t_L g907 ( 
.A(n_875),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_856),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_857),
.Y(n_909)
);

OAI21x1_ASAP7_75t_SL g910 ( 
.A1(n_889),
.A2(n_862),
.B(n_825),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_867),
.B(n_828),
.Y(n_911)
);

BUFx3_ASAP7_75t_L g912 ( 
.A(n_878),
.Y(n_912)
);

INVx2_ASAP7_75t_SL g913 ( 
.A(n_885),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_858),
.Y(n_914)
);

OR2x2_ASAP7_75t_L g915 ( 
.A(n_872),
.B(n_804),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_881),
.B(n_820),
.Y(n_916)
);

AO21x2_ASAP7_75t_L g917 ( 
.A1(n_870),
.A2(n_793),
.B(n_812),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_881),
.B(n_835),
.Y(n_918)
);

OAI21xp5_ASAP7_75t_L g919 ( 
.A1(n_859),
.A2(n_824),
.B(n_806),
.Y(n_919)
);

OA21x2_ASAP7_75t_L g920 ( 
.A1(n_873),
.A2(n_847),
.B(n_801),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_860),
.Y(n_921)
);

BUFx3_ASAP7_75t_L g922 ( 
.A(n_878),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_881),
.B(n_821),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_863),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_871),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_876),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_862),
.B(n_877),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_872),
.Y(n_928)
);

BUFx3_ASAP7_75t_L g929 ( 
.A(n_878),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_909),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_909),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_909),
.Y(n_932)
);

OR2x6_ASAP7_75t_L g933 ( 
.A(n_910),
.B(n_912),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_905),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_907),
.B(n_913),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_907),
.B(n_875),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_913),
.B(n_879),
.Y(n_937)
);

AND2x4_ASAP7_75t_L g938 ( 
.A(n_913),
.B(n_869),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_906),
.B(n_882),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_916),
.B(n_889),
.Y(n_940)
);

AND2x2_ASAP7_75t_L g941 ( 
.A(n_916),
.B(n_911),
.Y(n_941)
);

OR2x6_ASAP7_75t_L g942 ( 
.A(n_910),
.B(n_869),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_914),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_905),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_916),
.B(n_869),
.Y(n_945)
);

INVx5_ASAP7_75t_L g946 ( 
.A(n_912),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_911),
.B(n_897),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_914),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_914),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_921),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_936),
.B(n_911),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_930),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_934),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_936),
.B(n_923),
.Y(n_954)
);

INVx1_ASAP7_75t_SL g955 ( 
.A(n_947),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_931),
.Y(n_956)
);

NOR2xp67_ASAP7_75t_L g957 ( 
.A(n_946),
.B(n_880),
.Y(n_957)
);

OR2x2_ASAP7_75t_L g958 ( 
.A(n_934),
.B(n_927),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_944),
.Y(n_959)
);

HB1xp67_ASAP7_75t_L g960 ( 
.A(n_937),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_935),
.B(n_923),
.Y(n_961)
);

AND2x4_ASAP7_75t_L g962 ( 
.A(n_946),
.B(n_928),
.Y(n_962)
);

AND2x2_ASAP7_75t_L g963 ( 
.A(n_935),
.B(n_923),
.Y(n_963)
);

INVx2_ASAP7_75t_SL g964 ( 
.A(n_938),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_945),
.B(n_906),
.Y(n_965)
);

OR2x2_ASAP7_75t_L g966 ( 
.A(n_960),
.B(n_939),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_952),
.Y(n_967)
);

INVx3_ASAP7_75t_L g968 ( 
.A(n_962),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_965),
.B(n_937),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_953),
.Y(n_970)
);

AND2x2_ASAP7_75t_L g971 ( 
.A(n_964),
.B(n_938),
.Y(n_971)
);

INVx2_ASAP7_75t_SL g972 ( 
.A(n_962),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_952),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_965),
.B(n_940),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_954),
.B(n_940),
.Y(n_975)
);

INVx3_ASAP7_75t_L g976 ( 
.A(n_962),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_956),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_953),
.Y(n_978)
);

AND2x2_ASAP7_75t_L g979 ( 
.A(n_964),
.B(n_938),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_970),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_967),
.B(n_954),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_973),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_971),
.B(n_961),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_968),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_977),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_970),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_978),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_983),
.B(n_957),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_982),
.B(n_961),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_985),
.B(n_963),
.Y(n_990)
);

NOR2x1_ASAP7_75t_L g991 ( 
.A(n_984),
.B(n_968),
.Y(n_991)
);

INVx3_ASAP7_75t_L g992 ( 
.A(n_980),
.Y(n_992)
);

AO221x2_ASAP7_75t_L g993 ( 
.A1(n_981),
.A2(n_919),
.B1(n_975),
.B2(n_969),
.C(n_974),
.Y(n_993)
);

INVx4_ASAP7_75t_L g994 ( 
.A(n_980),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_992),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_989),
.Y(n_996)
);

INVx1_ASAP7_75t_SL g997 ( 
.A(n_991),
.Y(n_997)
);

OAI21xp33_ASAP7_75t_L g998 ( 
.A1(n_990),
.A2(n_981),
.B(n_986),
.Y(n_998)
);

AND2x4_ASAP7_75t_L g999 ( 
.A(n_994),
.B(n_972),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_993),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_988),
.Y(n_1001)
);

OR2x2_ASAP7_75t_L g1002 ( 
.A(n_989),
.B(n_966),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_992),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_993),
.B(n_972),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_995),
.Y(n_1005)
);

AOI22xp5_ASAP7_75t_L g1006 ( 
.A1(n_1000),
.A2(n_968),
.B1(n_976),
.B2(n_987),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_1003),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_999),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_999),
.Y(n_1009)
);

AND2x2_ASAP7_75t_L g1010 ( 
.A(n_1001),
.B(n_971),
.Y(n_1010)
);

OAI22xp5_ASAP7_75t_L g1011 ( 
.A1(n_997),
.A2(n_976),
.B1(n_942),
.B2(n_955),
.Y(n_1011)
);

O2A1O1Ixp33_ASAP7_75t_L g1012 ( 
.A1(n_1004),
.A2(n_919),
.B(n_976),
.C(n_884),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_998),
.A2(n_807),
.B(n_978),
.Y(n_1013)
);

INVx1_ASAP7_75t_SL g1014 ( 
.A(n_1008),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_1009),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_1005),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_1007),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_1010),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_1006),
.Y(n_1019)
);

AOI21xp33_ASAP7_75t_L g1020 ( 
.A1(n_1012),
.A2(n_996),
.B(n_1002),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_1013),
.B(n_979),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_1011),
.B(n_979),
.Y(n_1022)
);

OAI21xp33_ASAP7_75t_L g1023 ( 
.A1(n_1022),
.A2(n_880),
.B(n_884),
.Y(n_1023)
);

AOI322xp5_ASAP7_75t_L g1024 ( 
.A1(n_1019),
.A2(n_963),
.A3(n_894),
.B1(n_947),
.B2(n_951),
.C1(n_809),
.C2(n_918),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_1018),
.Y(n_1025)
);

AOI221x1_ASAP7_75t_L g1026 ( 
.A1(n_1016),
.A2(n_823),
.B1(n_956),
.B2(n_927),
.C(n_959),
.Y(n_1026)
);

NAND3xp33_ASAP7_75t_SL g1027 ( 
.A(n_1014),
.B(n_900),
.C(n_796),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_1014),
.Y(n_1028)
);

AOI21xp33_ASAP7_75t_L g1029 ( 
.A1(n_1015),
.A2(n_942),
.B(n_933),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_1028),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_1025),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_1023),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_1027),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_1024),
.B(n_1017),
.Y(n_1034)
);

AND2x2_ASAP7_75t_L g1035 ( 
.A(n_1029),
.B(n_1021),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_1026),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_1028),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_1028),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_1028),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_1028),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_1030),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_1036),
.B(n_1020),
.Y(n_1042)
);

NOR3xp33_ASAP7_75t_L g1043 ( 
.A(n_1038),
.B(n_1040),
.C(n_1039),
.Y(n_1043)
);

INVx2_ASAP7_75t_SL g1044 ( 
.A(n_1037),
.Y(n_1044)
);

NOR3xp33_ASAP7_75t_L g1045 ( 
.A(n_1034),
.B(n_895),
.C(n_831),
.Y(n_1045)
);

AOI211xp5_ASAP7_75t_L g1046 ( 
.A1(n_1034),
.A2(n_802),
.B(n_912),
.C(n_922),
.Y(n_1046)
);

NOR3xp33_ASAP7_75t_L g1047 ( 
.A(n_1035),
.B(n_895),
.C(n_850),
.Y(n_1047)
);

NOR2xp33_ASAP7_75t_L g1048 ( 
.A(n_1033),
.B(n_896),
.Y(n_1048)
);

NOR3xp33_ASAP7_75t_L g1049 ( 
.A(n_1032),
.B(n_895),
.C(n_816),
.Y(n_1049)
);

NOR2x1_ASAP7_75t_L g1050 ( 
.A(n_1031),
.B(n_942),
.Y(n_1050)
);

NOR3xp33_ASAP7_75t_L g1051 ( 
.A(n_1030),
.B(n_922),
.C(n_929),
.Y(n_1051)
);

NAND3xp33_ASAP7_75t_SL g1052 ( 
.A(n_1043),
.B(n_1045),
.C(n_1042),
.Y(n_1052)
);

AOI211xp5_ASAP7_75t_L g1053 ( 
.A1(n_1048),
.A2(n_922),
.B(n_929),
.C(n_896),
.Y(n_1053)
);

NAND4xp25_ASAP7_75t_L g1054 ( 
.A(n_1051),
.B(n_929),
.C(n_836),
.D(n_896),
.Y(n_1054)
);

NOR3xp33_ASAP7_75t_L g1055 ( 
.A(n_1044),
.B(n_892),
.C(n_893),
.Y(n_1055)
);

NAND3xp33_ASAP7_75t_L g1056 ( 
.A(n_1041),
.B(n_841),
.C(n_946),
.Y(n_1056)
);

INVx1_ASAP7_75t_SL g1057 ( 
.A(n_1050),
.Y(n_1057)
);

INVx3_ASAP7_75t_L g1058 ( 
.A(n_1049),
.Y(n_1058)
);

O2A1O1Ixp33_ASAP7_75t_L g1059 ( 
.A1(n_1046),
.A2(n_799),
.B(n_942),
.C(n_933),
.Y(n_1059)
);

NOR3xp33_ASAP7_75t_L g1060 ( 
.A(n_1052),
.B(n_1047),
.C(n_892),
.Y(n_1060)
);

NAND3xp33_ASAP7_75t_L g1061 ( 
.A(n_1053),
.B(n_849),
.C(n_946),
.Y(n_1061)
);

OAI221xp5_ASAP7_75t_L g1062 ( 
.A1(n_1057),
.A2(n_933),
.B1(n_893),
.B2(n_894),
.C(n_899),
.Y(n_1062)
);

AND2x2_ASAP7_75t_L g1063 ( 
.A(n_1058),
.B(n_951),
.Y(n_1063)
);

OAI211xp5_ASAP7_75t_L g1064 ( 
.A1(n_1054),
.A2(n_845),
.B(n_888),
.C(n_887),
.Y(n_1064)
);

AOI221x1_ASAP7_75t_L g1065 ( 
.A1(n_1056),
.A2(n_959),
.B1(n_886),
.B2(n_945),
.C(n_890),
.Y(n_1065)
);

NAND4xp25_ASAP7_75t_SL g1066 ( 
.A(n_1059),
.B(n_915),
.C(n_958),
.D(n_898),
.Y(n_1066)
);

NAND3xp33_ASAP7_75t_SL g1067 ( 
.A(n_1055),
.B(n_915),
.C(n_898),
.Y(n_1067)
);

NAND5xp2_ASAP7_75t_L g1068 ( 
.A(n_1053),
.B(n_918),
.C(n_868),
.D(n_941),
.E(n_891),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_1063),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_1060),
.Y(n_1070)
);

NAND2x1p5_ASAP7_75t_L g1071 ( 
.A(n_1064),
.B(n_915),
.Y(n_1071)
);

NOR2x1_ASAP7_75t_L g1072 ( 
.A(n_1061),
.B(n_933),
.Y(n_1072)
);

NOR3xp33_ASAP7_75t_L g1073 ( 
.A(n_1066),
.B(n_874),
.C(n_902),
.Y(n_1073)
);

NOR3xp33_ASAP7_75t_L g1074 ( 
.A(n_1068),
.B(n_1062),
.C(n_1067),
.Y(n_1074)
);

AOI22xp5_ASAP7_75t_L g1075 ( 
.A1(n_1065),
.A2(n_958),
.B1(n_904),
.B2(n_928),
.Y(n_1075)
);

NOR3xp33_ASAP7_75t_L g1076 ( 
.A(n_1064),
.B(n_902),
.C(n_924),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_1063),
.Y(n_1077)
);

INVx1_ASAP7_75t_SL g1078 ( 
.A(n_1069),
.Y(n_1078)
);

AND2x2_ASAP7_75t_SL g1079 ( 
.A(n_1077),
.B(n_920),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_1072),
.Y(n_1080)
);

INVx3_ASAP7_75t_L g1081 ( 
.A(n_1071),
.Y(n_1081)
);

AND3x1_ASAP7_75t_L g1082 ( 
.A(n_1070),
.B(n_918),
.C(n_944),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_1074),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_1076),
.B(n_924),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_1075),
.Y(n_1085)
);

NAND3x1_ASAP7_75t_L g1086 ( 
.A(n_1073),
.B(n_932),
.C(n_949),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_1069),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_1069),
.Y(n_1088)
);

OR3x2_ASAP7_75t_L g1089 ( 
.A(n_1077),
.B(n_159),
.C(n_160),
.Y(n_1089)
);

NAND4xp25_ASAP7_75t_L g1090 ( 
.A(n_1077),
.B(n_883),
.C(n_926),
.D(n_925),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_1081),
.Y(n_1091)
);

CKINVDCx20_ASAP7_75t_R g1092 ( 
.A(n_1078),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1087),
.Y(n_1093)
);

OAI221xp5_ASAP7_75t_L g1094 ( 
.A1(n_1080),
.A2(n_950),
.B1(n_948),
.B2(n_943),
.C(n_901),
.Y(n_1094)
);

OAI311xp33_ASAP7_75t_L g1095 ( 
.A1(n_1083),
.A2(n_908),
.A3(n_903),
.B1(n_169),
.C1(n_170),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_1083),
.A2(n_904),
.B(n_920),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_1088),
.B(n_926),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_1085),
.A2(n_904),
.B(n_920),
.Y(n_1098)
);

XNOR2x1_ASAP7_75t_L g1099 ( 
.A(n_1082),
.B(n_166),
.Y(n_1099)
);

OAI22xp5_ASAP7_75t_L g1100 ( 
.A1(n_1092),
.A2(n_1089),
.B1(n_1086),
.B2(n_1084),
.Y(n_1100)
);

INVx2_ASAP7_75t_SL g1101 ( 
.A(n_1091),
.Y(n_1101)
);

OAI22xp5_ASAP7_75t_SL g1102 ( 
.A1(n_1093),
.A2(n_1097),
.B1(n_1099),
.B2(n_1094),
.Y(n_1102)
);

AO22x2_ASAP7_75t_L g1103 ( 
.A1(n_1095),
.A2(n_1090),
.B1(n_1079),
.B2(n_921),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_1096),
.Y(n_1104)
);

AO22x2_ASAP7_75t_L g1105 ( 
.A1(n_1098),
.A2(n_921),
.B1(n_925),
.B2(n_926),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1103),
.Y(n_1106)
);

INVx3_ASAP7_75t_L g1107 ( 
.A(n_1101),
.Y(n_1107)
);

XNOR2xp5_ASAP7_75t_L g1108 ( 
.A(n_1100),
.B(n_167),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_1107),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_1109),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_1110),
.A2(n_1102),
.B(n_1106),
.Y(n_1111)
);

OAI22xp5_ASAP7_75t_L g1112 ( 
.A1(n_1111),
.A2(n_1108),
.B1(n_1104),
.B2(n_1105),
.Y(n_1112)
);

AOI22xp33_ASAP7_75t_L g1113 ( 
.A1(n_1111),
.A2(n_901),
.B1(n_925),
.B2(n_920),
.Y(n_1113)
);

AOI22xp5_ASAP7_75t_L g1114 ( 
.A1(n_1111),
.A2(n_917),
.B1(n_904),
.B2(n_920),
.Y(n_1114)
);

AO21x2_ASAP7_75t_L g1115 ( 
.A1(n_1112),
.A2(n_171),
.B(n_172),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_SL g1116 ( 
.A(n_1113),
.B(n_1114),
.Y(n_1116)
);

AO21x2_ASAP7_75t_L g1117 ( 
.A1(n_1112),
.A2(n_179),
.B(n_183),
.Y(n_1117)
);

AO221x2_ASAP7_75t_L g1118 ( 
.A1(n_1115),
.A2(n_184),
.B1(n_185),
.B2(n_186),
.C(n_187),
.Y(n_1118)
);

AOI22xp33_ASAP7_75t_L g1119 ( 
.A1(n_1117),
.A2(n_903),
.B1(n_908),
.B2(n_917),
.Y(n_1119)
);

AOI31xp33_ASAP7_75t_L g1120 ( 
.A1(n_1118),
.A2(n_1116),
.A3(n_191),
.B(n_192),
.Y(n_1120)
);

AOI211xp5_ASAP7_75t_L g1121 ( 
.A1(n_1120),
.A2(n_1119),
.B(n_194),
.C(n_196),
.Y(n_1121)
);


endmodule