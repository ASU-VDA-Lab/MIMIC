module fake_jpeg_27958_n_270 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_270);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_270;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_16),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx2_ASAP7_75t_SL g35 ( 
.A(n_20),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_35),
.B(n_37),
.Y(n_63)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_22),
.B(n_17),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_18),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_31),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_22),
.B(n_1),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_39),
.B(n_19),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_37),
.B(n_19),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_45),
.B(n_47),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_39),
.B(n_19),
.Y(n_47)
);

OAI21xp33_ASAP7_75t_L g72 ( 
.A1(n_49),
.A2(n_64),
.B(n_26),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_50),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_25),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_51),
.B(n_62),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_36),
.A2(n_20),
.B1(n_24),
.B2(n_32),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_55),
.A2(n_35),
.B1(n_44),
.B2(n_20),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_36),
.B(n_33),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_56),
.B(n_59),
.Y(n_89)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_43),
.B(n_33),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_32),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_61),
.B(n_17),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_28),
.Y(n_62)
);

HAxp5_ASAP7_75t_SL g64 ( 
.A(n_35),
.B(n_25),
.CON(n_64),
.SN(n_64)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_61),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_66),
.B(n_67),
.Y(n_98)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_69),
.Y(n_108)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_57),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_70),
.B(n_79),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_71),
.B(n_72),
.Y(n_112)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_73),
.B(n_74),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_75),
.Y(n_118)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_77),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_78),
.A2(n_80),
.B1(n_92),
.B2(n_86),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_56),
.B(n_40),
.C(n_42),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_53),
.A2(n_44),
.B1(n_29),
.B2(n_26),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_82),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

AND2x2_ASAP7_75t_SL g86 ( 
.A(n_46),
.B(n_21),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_91),
.Y(n_97)
);

NOR2x1_ASAP7_75t_L g87 ( 
.A(n_47),
.B(n_29),
.Y(n_87)
);

NAND3xp33_ASAP7_75t_L g96 ( 
.A(n_87),
.B(n_94),
.C(n_67),
.Y(n_96)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_90),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_49),
.B(n_28),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_46),
.B(n_23),
.C(n_26),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_53),
.A2(n_33),
.B1(n_21),
.B2(n_34),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_57),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_71),
.A2(n_58),
.B1(n_54),
.B2(n_60),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_95),
.A2(n_119),
.B1(n_69),
.B2(n_81),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_96),
.B(n_104),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_74),
.A2(n_54),
.B1(n_60),
.B2(n_21),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_99),
.A2(n_94),
.B1(n_70),
.B2(n_18),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_107),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_54),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_113),
.Y(n_124)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_77),
.Y(n_104)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_77),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_111),
.Y(n_125)
);

AND2x4_ASAP7_75t_L g107 ( 
.A(n_86),
.B(n_48),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_84),
.B(n_30),
.Y(n_110)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_76),
.B(n_66),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_73),
.B(n_48),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_87),
.B(n_34),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_115),
.B(n_116),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_82),
.B(n_41),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_79),
.B(n_41),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_117),
.B(n_120),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_67),
.A2(n_68),
.B1(n_88),
.B2(n_75),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_68),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_91),
.B(n_2),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_2),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_100),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_122),
.B(n_127),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_105),
.A2(n_117),
.B(n_97),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_123),
.A2(n_128),
.B(n_126),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_105),
.B(n_83),
.C(n_85),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_126),
.B(n_31),
.C(n_27),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_95),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_99),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_131),
.B(n_132),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_97),
.A2(n_107),
.B1(n_114),
.B2(n_101),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_134),
.A2(n_136),
.B1(n_138),
.B2(n_147),
.Y(n_154)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_113),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_135),
.B(n_146),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_107),
.A2(n_118),
.B1(n_108),
.B2(n_85),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_98),
.B(n_23),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_137),
.B(n_121),
.Y(n_157)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_109),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_139),
.B(n_141),
.Y(n_161)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_118),
.Y(n_140)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_140),
.Y(n_173)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_119),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_116),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_142),
.B(n_144),
.Y(n_175)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_108),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_103),
.Y(n_145)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_145),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_111),
.A2(n_31),
.B1(n_27),
.B2(n_93),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_120),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_148),
.B(n_130),
.Y(n_171)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_107),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_149),
.B(n_105),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_151),
.B(n_152),
.Y(n_200)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_124),
.Y(n_152)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_124),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_156),
.B(n_158),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_157),
.B(n_168),
.Y(n_188)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_143),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_135),
.B(n_112),
.Y(n_159)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_159),
.Y(n_199)
);

OA21x2_ASAP7_75t_L g160 ( 
.A1(n_149),
.A2(n_106),
.B(n_104),
.Y(n_160)
);

OA22x2_ASAP7_75t_L g193 ( 
.A1(n_160),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_125),
.B(n_115),
.Y(n_162)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_162),
.Y(n_181)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_143),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_163),
.B(n_169),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_134),
.B(n_102),
.Y(n_164)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_164),
.Y(n_182)
);

INVx2_ASAP7_75t_SL g165 ( 
.A(n_140),
.Y(n_165)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_165),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_128),
.A2(n_102),
.B(n_93),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_166),
.A2(n_174),
.B(n_2),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_123),
.B(n_93),
.Y(n_167)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_167),
.Y(n_197)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_132),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_171),
.B(n_144),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_172),
.B(n_176),
.C(n_177),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_128),
.A2(n_27),
.B(n_30),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_137),
.B(n_30),
.C(n_15),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_130),
.B(n_133),
.C(n_146),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_154),
.A2(n_122),
.B1(n_129),
.B2(n_138),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_178),
.A2(n_151),
.B1(n_172),
.B2(n_177),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_180),
.B(n_184),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_166),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_175),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_185),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_186),
.B(n_193),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_162),
.B(n_15),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_187),
.B(n_192),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_153),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_190),
.A2(n_195),
.B1(n_198),
.B2(n_170),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_161),
.B(n_14),
.Y(n_191)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_191),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_155),
.Y(n_192)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_193),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_169),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_167),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_196),
.A2(n_164),
.B1(n_158),
.B2(n_163),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_174),
.Y(n_198)
);

AOI21x1_ASAP7_75t_L g201 ( 
.A1(n_186),
.A2(n_168),
.B(n_160),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_201),
.B(n_211),
.Y(n_233)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_202),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_193),
.B(n_159),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_204),
.A2(n_182),
.B(n_199),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_205),
.B(n_207),
.Y(n_220)
);

NOR2x1_ASAP7_75t_L g206 ( 
.A(n_178),
.B(n_160),
.Y(n_206)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_206),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_188),
.B(n_156),
.C(n_152),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_208),
.B(n_214),
.C(n_216),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_188),
.B(n_157),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_209),
.B(n_212),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_181),
.A2(n_189),
.B1(n_182),
.B2(n_199),
.Y(n_210)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_210),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_194),
.B(n_150),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_194),
.B(n_150),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_213),
.B(n_197),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_200),
.B(n_176),
.C(n_173),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_200),
.B(n_173),
.C(n_165),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_218),
.B(n_179),
.Y(n_225)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_225),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_203),
.B(n_181),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_226),
.B(n_227),
.Y(n_244)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_216),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_228),
.A2(n_183),
.B(n_212),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_230),
.B(n_209),
.C(n_215),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_204),
.B(n_197),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_231),
.B(n_165),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_217),
.A2(n_184),
.B1(n_198),
.B2(n_183),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_232),
.A2(n_214),
.B1(n_208),
.B2(n_193),
.Y(n_237)
);

O2A1O1Ixp33_ASAP7_75t_L g234 ( 
.A1(n_231),
.A2(n_219),
.B(n_206),
.C(n_211),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_234),
.A2(n_229),
.B1(n_222),
.B2(n_8),
.Y(n_251)
);

BUFx4f_ASAP7_75t_SL g236 ( 
.A(n_228),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_236),
.A2(n_223),
.B1(n_232),
.B2(n_233),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_237),
.B(n_238),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_229),
.B(n_213),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_239),
.B(n_240),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_241),
.B(n_233),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_221),
.B(n_13),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_242),
.B(n_243),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_224),
.B(n_13),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_245),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_249),
.B(n_251),
.Y(n_254)
);

OAI21x1_ASAP7_75t_L g250 ( 
.A1(n_244),
.A2(n_220),
.B(n_230),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_250),
.B(n_234),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_240),
.B(n_222),
.C(n_7),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_252),
.B(n_253),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_235),
.A2(n_6),
.B(n_8),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_255),
.A2(n_246),
.B(n_248),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_247),
.B(n_236),
.C(n_8),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_257),
.B(n_6),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_246),
.B(n_236),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_258),
.B(n_251),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_260),
.B(n_259),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_261),
.B(n_263),
.Y(n_265)
);

OAI21x1_ASAP7_75t_SL g262 ( 
.A1(n_258),
.A2(n_252),
.B(n_9),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_262),
.A2(n_254),
.B(n_256),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_264),
.B(n_266),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_265),
.B(n_10),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_268),
.B(n_267),
.C(n_10),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_269),
.B(n_10),
.Y(n_270)
);


endmodule