module fake_jpeg_30882_n_476 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_476);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_476;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_16),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx6f_ASAP7_75t_SL g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_6),
.B(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_12),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_8),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_13),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_50),
.Y(n_109)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_51),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_20),
.B(n_15),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_52),
.B(n_61),
.Y(n_103)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_54),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_26),
.B(n_15),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_55),
.B(n_88),
.Y(n_142)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_56),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_57),
.Y(n_140)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_58),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_59),
.Y(n_99)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_60),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_20),
.B(n_12),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_62),
.Y(n_138)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_17),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g150 ( 
.A(n_63),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_47),
.B(n_0),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_64),
.B(n_69),
.Y(n_117)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_65),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_66),
.Y(n_101)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_67),
.Y(n_133)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_68),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_24),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_24),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_70),
.B(n_75),
.Y(n_123)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_71),
.Y(n_104)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_72),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

INVx4_ASAP7_75t_SL g148 ( 
.A(n_73),
.Y(n_148)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_74),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_38),
.Y(n_75)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g135 ( 
.A(n_76),
.Y(n_135)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_21),
.Y(n_77)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_77),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_34),
.Y(n_78)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_78),
.Y(n_134)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_79),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_38),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_80),
.B(n_82),
.Y(n_128)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_81),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_47),
.B(n_26),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_21),
.Y(n_83)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_83),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_84),
.Y(n_129)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g120 ( 
.A(n_85),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_34),
.Y(n_86)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_86),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_41),
.B(n_0),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_87),
.B(n_91),
.Y(n_146)
);

INVx6_ASAP7_75t_SL g88 ( 
.A(n_32),
.Y(n_88)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_34),
.Y(n_89)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_89),
.Y(n_127)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_22),
.Y(n_90)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_90),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_92),
.A2(n_95),
.B1(n_96),
.B2(n_45),
.Y(n_98)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_31),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_93),
.B(n_94),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_41),
.B(n_31),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_22),
.Y(n_95)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_48),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_42),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_97),
.B(n_28),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_98),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_58),
.A2(n_33),
.B1(n_32),
.B2(n_48),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_100),
.A2(n_110),
.B1(n_115),
.B2(n_141),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_108),
.B(n_2),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_72),
.A2(n_33),
.B1(n_32),
.B2(n_43),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_88),
.A2(n_33),
.B1(n_49),
.B2(n_32),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_111),
.A2(n_113),
.B1(n_116),
.B2(n_119),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_67),
.A2(n_49),
.B1(n_45),
.B2(n_43),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_79),
.A2(n_18),
.B1(n_43),
.B2(n_49),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_56),
.A2(n_49),
.B1(n_45),
.B2(n_18),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_97),
.A2(n_44),
.B1(n_42),
.B2(n_18),
.Y(n_119)
);

AOI21xp33_ASAP7_75t_SL g126 ( 
.A1(n_50),
.A2(n_73),
.B(n_62),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_126),
.B(n_130),
.C(n_71),
.Y(n_183)
);

AND2x2_ASAP7_75t_SL g130 ( 
.A(n_59),
.B(n_1),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_60),
.A2(n_44),
.B1(n_37),
.B2(n_19),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_132),
.A2(n_27),
.B1(n_76),
.B2(n_95),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_54),
.A2(n_46),
.B1(n_29),
.B2(n_28),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_137),
.A2(n_92),
.B1(n_91),
.B2(n_84),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_57),
.A2(n_46),
.B1(n_23),
.B2(n_29),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_63),
.B(n_37),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_143),
.B(n_151),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_65),
.A2(n_23),
.B1(n_19),
.B2(n_39),
.Y(n_144)
);

OR2x2_ASAP7_75t_L g176 ( 
.A(n_144),
.B(n_36),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_68),
.B(n_39),
.Y(n_151)
);

OAI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_81),
.A2(n_39),
.B1(n_27),
.B2(n_17),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_152),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g153 ( 
.A(n_143),
.B(n_108),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_153),
.B(n_130),
.Y(n_226)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_145),
.Y(n_154)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_154),
.Y(n_219)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_109),
.Y(n_155)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_155),
.Y(n_242)
);

OAI21xp33_ASAP7_75t_L g156 ( 
.A1(n_126),
.A2(n_73),
.B(n_62),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_156),
.Y(n_218)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_105),
.Y(n_158)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_158),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_123),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_159),
.B(n_170),
.Y(n_204)
);

A2O1A1Ixp33_ASAP7_75t_L g161 ( 
.A1(n_151),
.A2(n_17),
.B(n_27),
.C(n_50),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_161),
.B(n_194),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_162),
.Y(n_220)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_145),
.Y(n_163)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_163),
.Y(n_247)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_147),
.Y(n_164)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_164),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_106),
.A2(n_74),
.B1(n_96),
.B2(n_89),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_165),
.A2(n_179),
.B1(n_148),
.B2(n_135),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_166),
.A2(n_192),
.B1(n_203),
.B2(n_144),
.Y(n_207)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_147),
.Y(n_167)
);

INVx5_ASAP7_75t_L g215 ( 
.A(n_167),
.Y(n_215)
);

INVx13_ASAP7_75t_L g168 ( 
.A(n_109),
.Y(n_168)
);

BUFx12f_ASAP7_75t_L g211 ( 
.A(n_168),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_99),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_169),
.Y(n_210)
);

INVx8_ASAP7_75t_L g170 ( 
.A(n_138),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_125),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_171),
.Y(n_225)
);

BUFx12f_ASAP7_75t_L g172 ( 
.A(n_99),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_172),
.Y(n_208)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_133),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_173),
.B(n_183),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_103),
.B(n_85),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_175),
.B(n_177),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_176),
.A2(n_134),
.B(n_104),
.Y(n_237)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_114),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_125),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_178),
.B(n_180),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_150),
.A2(n_86),
.B1(n_78),
.B2(n_66),
.Y(n_179)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_138),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_124),
.B(n_90),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_181),
.B(n_182),
.Y(n_217)
);

OR2x2_ASAP7_75t_L g182 ( 
.A(n_124),
.B(n_1),
.Y(n_182)
);

OAI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_121),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_184),
.A2(n_174),
.B1(n_157),
.B2(n_191),
.Y(n_229)
);

INVx8_ASAP7_75t_L g185 ( 
.A(n_129),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_185),
.B(n_186),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_128),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_117),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_187),
.B(n_188),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_142),
.B(n_146),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_150),
.B(n_2),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_189),
.B(n_5),
.Y(n_221)
);

BUFx12_ASAP7_75t_L g190 ( 
.A(n_104),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_190),
.B(n_191),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_112),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_192)
);

OA22x2_ASAP7_75t_SL g193 ( 
.A1(n_130),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_193)
);

O2A1O1Ixp33_ASAP7_75t_L g228 ( 
.A1(n_193),
.A2(n_149),
.B(n_7),
.C(n_8),
.Y(n_228)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_133),
.Y(n_194)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_120),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_196),
.B(n_197),
.Y(n_216)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_131),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_102),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_198),
.B(n_199),
.Y(n_205)
);

INVx2_ASAP7_75t_SL g199 ( 
.A(n_134),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_107),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_200),
.B(n_201),
.Y(n_223)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_149),
.Y(n_201)
);

INVx6_ASAP7_75t_L g202 ( 
.A(n_129),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_202),
.B(n_140),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_207),
.A2(n_224),
.B1(n_202),
.B2(n_185),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_176),
.A2(n_115),
.B1(n_112),
.B2(n_139),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_212),
.A2(n_233),
.B1(n_238),
.B2(n_199),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_221),
.B(n_170),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_226),
.B(n_240),
.C(n_244),
.Y(n_259)
);

AND2x2_ASAP7_75t_SL g227 ( 
.A(n_160),
.B(n_148),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g272 ( 
.A(n_227),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_228),
.B(n_248),
.Y(n_256)
);

CKINVDCx14_ASAP7_75t_R g261 ( 
.A(n_229),
.Y(n_261)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_230),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_174),
.A2(n_195),
.B1(n_191),
.B2(n_160),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_232),
.A2(n_154),
.B1(n_164),
.B2(n_167),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_195),
.A2(n_101),
.B1(n_139),
.B2(n_140),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_153),
.B(n_127),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_234),
.B(n_236),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_182),
.B(n_183),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_237),
.A2(n_169),
.B(n_172),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_203),
.A2(n_101),
.B1(n_122),
.B2(n_100),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_158),
.B(n_161),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_239),
.B(n_246),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_173),
.B(n_194),
.C(n_196),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_198),
.B(n_118),
.C(n_136),
.Y(n_244)
);

O2A1O1Ixp33_ASAP7_75t_L g245 ( 
.A1(n_193),
.A2(n_135),
.B(n_136),
.C(n_118),
.Y(n_245)
);

OA21x2_ASAP7_75t_L g249 ( 
.A1(n_245),
.A2(n_199),
.B(n_193),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_197),
.B(n_122),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_200),
.B(n_6),
.C(n_8),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_249),
.A2(n_270),
.B(n_285),
.Y(n_313)
);

NAND3xp33_ASAP7_75t_L g311 ( 
.A(n_250),
.B(n_263),
.C(n_271),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_213),
.Y(n_251)
);

INVx13_ASAP7_75t_L g308 ( 
.A(n_251),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_204),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_253),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_206),
.B(n_180),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_254),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_243),
.B(n_155),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_255),
.Y(n_289)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_246),
.Y(n_257)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_257),
.Y(n_291)
);

BUFx8_ASAP7_75t_L g260 ( 
.A(n_211),
.Y(n_260)
);

BUFx2_ASAP7_75t_L g314 ( 
.A(n_260),
.Y(n_314)
);

BUFx3_ASAP7_75t_L g262 ( 
.A(n_208),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_262),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_231),
.B(n_168),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_265),
.A2(n_275),
.B1(n_230),
.B2(n_244),
.Y(n_290)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_222),
.Y(n_266)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_266),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_223),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_267),
.B(n_273),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_239),
.A2(n_171),
.B(n_178),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_268),
.A2(n_279),
.B(n_216),
.Y(n_298)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_222),
.Y(n_269)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_269),
.Y(n_295)
);

NOR2xp67_ASAP7_75t_L g271 ( 
.A(n_227),
.B(n_172),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_217),
.B(n_201),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_205),
.Y(n_274)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_274),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_214),
.B(n_163),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_276),
.B(n_278),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_277),
.A2(n_287),
.B1(n_233),
.B2(n_272),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_214),
.B(n_8),
.Y(n_278)
);

A2O1A1Ixp33_ASAP7_75t_L g279 ( 
.A1(n_218),
.A2(n_9),
.B(n_10),
.C(n_190),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_234),
.B(n_190),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_280),
.B(n_283),
.Y(n_303)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_219),
.Y(n_281)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_281),
.Y(n_302)
);

OAI32xp33_ASAP7_75t_L g282 ( 
.A1(n_236),
.A2(n_232),
.A3(n_238),
.B1(n_229),
.B2(n_218),
.Y(n_282)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_282),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_227),
.B(n_226),
.Y(n_283)
);

CKINVDCx14_ASAP7_75t_R g284 ( 
.A(n_208),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_L g312 ( 
.A1(n_284),
.A2(n_211),
.B1(n_210),
.B2(n_242),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_228),
.A2(n_237),
.B(n_220),
.Y(n_285)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_211),
.Y(n_286)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_286),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_220),
.A2(n_207),
.B1(n_212),
.B2(n_209),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_205),
.Y(n_288)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_288),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_290),
.B(n_293),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_261),
.A2(n_209),
.B1(n_245),
.B2(n_240),
.Y(n_293)
);

AO21x1_ASAP7_75t_L g355 ( 
.A1(n_298),
.A2(n_300),
.B(n_249),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_299),
.A2(n_251),
.B1(n_282),
.B2(n_277),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_256),
.A2(n_224),
.B(n_209),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_SL g304 ( 
.A(n_283),
.B(n_241),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_SL g328 ( 
.A(n_304),
.B(n_264),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_259),
.B(n_241),
.C(n_223),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_306),
.B(n_307),
.C(n_318),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_259),
.B(n_241),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_265),
.A2(n_216),
.B1(n_248),
.B2(n_225),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_310),
.B(n_321),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_312),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_272),
.B(n_210),
.C(n_247),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_258),
.B(n_247),
.C(n_225),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_319),
.B(n_322),
.C(n_323),
.Y(n_348)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_266),
.Y(n_320)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_320),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_275),
.A2(n_219),
.B1(n_235),
.B2(n_215),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_258),
.B(n_242),
.C(n_235),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_280),
.B(n_221),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_269),
.Y(n_324)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_324),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_301),
.B(n_253),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_325),
.B(n_330),
.Y(n_367)
);

CKINVDCx16_ASAP7_75t_R g327 ( 
.A(n_294),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_327),
.B(n_331),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_SL g369 ( 
.A(n_328),
.B(n_293),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_294),
.B(n_264),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_309),
.B(n_278),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_313),
.A2(n_256),
.B(n_271),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_333),
.A2(n_342),
.B(n_355),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_297),
.B(n_267),
.Y(n_334)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_334),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_313),
.A2(n_270),
.B(n_285),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g364 ( 
.A1(n_335),
.A2(n_341),
.B(n_353),
.Y(n_364)
);

CKINVDCx16_ASAP7_75t_R g336 ( 
.A(n_292),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_336),
.B(n_339),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_296),
.B(n_257),
.Y(n_337)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_337),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_315),
.A2(n_252),
.B1(n_288),
.B2(n_274),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_338),
.A2(n_349),
.B1(n_290),
.B2(n_310),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_314),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_300),
.A2(n_262),
.B(n_287),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_315),
.A2(n_279),
.B(n_276),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_292),
.Y(n_343)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_343),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_305),
.B(n_252),
.Y(n_345)
);

OAI21xp33_ASAP7_75t_L g376 ( 
.A1(n_345),
.A2(n_347),
.B(n_352),
.Y(n_376)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_295),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_346),
.A2(n_351),
.B1(n_354),
.B2(n_356),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_314),
.Y(n_347)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_295),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_297),
.B(n_268),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_L g353 ( 
.A1(n_311),
.A2(n_249),
.B(n_260),
.Y(n_353)
);

INVx13_ASAP7_75t_L g354 ( 
.A(n_316),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_320),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_356),
.A2(n_324),
.B(n_316),
.Y(n_374)
);

XOR2x1_ASAP7_75t_L g357 ( 
.A(n_335),
.B(n_355),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_357),
.B(n_341),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_329),
.A2(n_299),
.B1(n_296),
.B2(n_317),
.Y(n_358)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_358),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_344),
.B(n_307),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_359),
.B(n_361),
.C(n_362),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_344),
.B(n_306),
.C(n_304),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_344),
.B(n_318),
.C(n_303),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_348),
.B(n_303),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_363),
.B(n_368),
.C(n_372),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_366),
.A2(n_349),
.B1(n_337),
.B2(n_353),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_348),
.B(n_319),
.C(n_322),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_369),
.B(n_379),
.Y(n_400)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_370),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_348),
.B(n_323),
.C(n_317),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_326),
.B(n_291),
.C(n_289),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_373),
.B(n_377),
.C(n_382),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_374),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_329),
.A2(n_291),
.B1(n_289),
.B2(n_321),
.Y(n_375)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_375),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_326),
.B(n_298),
.C(n_302),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_333),
.B(n_308),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_352),
.A2(n_334),
.B1(n_330),
.B2(n_327),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_381),
.B(n_338),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_335),
.B(n_308),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_L g414 ( 
.A1(n_384),
.A2(n_389),
.B(n_394),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_386),
.A2(n_404),
.B1(n_406),
.B2(n_375),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_387),
.B(n_397),
.Y(n_424)
);

AOI22xp33_ASAP7_75t_L g388 ( 
.A1(n_360),
.A2(n_353),
.B1(n_339),
.B2(n_347),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_388),
.A2(n_405),
.B1(n_368),
.B2(n_362),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g389 ( 
.A1(n_364),
.A2(n_341),
.B(n_355),
.Y(n_389)
);

BUFx2_ASAP7_75t_L g393 ( 
.A(n_380),
.Y(n_393)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_393),
.Y(n_417)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_364),
.A2(n_355),
.B(n_342),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_365),
.A2(n_325),
.B(n_338),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_395),
.B(n_399),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_367),
.B(n_345),
.Y(n_397)
);

INVx13_ASAP7_75t_L g399 ( 
.A(n_376),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_383),
.B(n_331),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_401),
.B(n_402),
.Y(n_422)
);

BUFx12_ASAP7_75t_L g402 ( 
.A(n_357),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_366),
.A2(n_371),
.B1(n_377),
.B2(n_373),
.Y(n_404)
);

INVx1_ASAP7_75t_SL g405 ( 
.A(n_379),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_358),
.A2(n_350),
.B1(n_336),
.B2(n_351),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_407),
.B(n_411),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_391),
.B(n_359),
.C(n_361),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_408),
.B(n_413),
.C(n_415),
.Y(n_434)
);

NOR2xp67_ASAP7_75t_L g409 ( 
.A(n_395),
.B(n_365),
.Y(n_409)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_409),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_398),
.B(n_363),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_410),
.B(n_416),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_398),
.B(n_390),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_390),
.B(n_372),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_412),
.B(n_423),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_400),
.B(n_382),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_400),
.B(n_404),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_391),
.B(n_369),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_SL g418 ( 
.A(n_386),
.B(n_394),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_418),
.B(n_420),
.C(n_421),
.Y(n_435)
);

XNOR2x1_ASAP7_75t_L g420 ( 
.A(n_387),
.B(n_381),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_405),
.B(n_328),
.C(n_374),
.Y(n_421)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_417),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_427),
.B(n_436),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_422),
.A2(n_392),
.B1(n_396),
.B2(n_385),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_428),
.A2(n_396),
.B1(n_385),
.B2(n_406),
.Y(n_444)
);

BUFx24_ASAP7_75t_SL g430 ( 
.A(n_411),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_SL g442 ( 
.A(n_430),
.B(n_416),
.Y(n_442)
);

CKINVDCx16_ASAP7_75t_R g431 ( 
.A(n_424),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_431),
.B(n_433),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_419),
.B(n_378),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_410),
.B(n_397),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g437 ( 
.A1(n_414),
.A2(n_389),
.B(n_403),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_437),
.B(n_420),
.Y(n_440)
);

A2O1A1Ixp33_ASAP7_75t_SL g438 ( 
.A1(n_418),
.A2(n_402),
.B(n_403),
.C(n_399),
.Y(n_438)
);

NOR3xp33_ASAP7_75t_L g446 ( 
.A(n_438),
.B(n_402),
.C(n_332),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_SL g439 ( 
.A1(n_408),
.A2(n_402),
.B(n_392),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_439),
.B(n_328),
.Y(n_449)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_440),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_442),
.B(n_445),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_426),
.B(n_421),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_443),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_444),
.A2(n_438),
.B1(n_428),
.B2(n_432),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_SL g445 ( 
.A(n_437),
.B(n_415),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_446),
.B(n_449),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_432),
.B(n_413),
.C(n_332),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_447),
.B(n_451),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_435),
.B(n_346),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_450),
.B(n_435),
.C(n_434),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_434),
.B(n_343),
.Y(n_451)
);

OR2x2_ASAP7_75t_L g452 ( 
.A(n_438),
.B(n_340),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_452),
.B(n_393),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_453),
.B(n_457),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_460),
.B(n_461),
.Y(n_468)
);

FAx1_ASAP7_75t_SL g461 ( 
.A(n_440),
.B(n_438),
.CI(n_429),
.CON(n_461),
.SN(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_441),
.B(n_425),
.Y(n_462)
);

OAI21xp33_ASAP7_75t_L g469 ( 
.A1(n_462),
.A2(n_463),
.B(n_454),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_SL g463 ( 
.A(n_448),
.B(n_340),
.Y(n_463)
);

AOI22xp33_ASAP7_75t_SL g464 ( 
.A1(n_459),
.A2(n_446),
.B1(n_452),
.B2(n_443),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_L g470 ( 
.A1(n_464),
.A2(n_469),
.B1(n_456),
.B2(n_455),
.Y(n_470)
);

NOR3xp33_ASAP7_75t_SL g466 ( 
.A(n_458),
.B(n_450),
.C(n_354),
.Y(n_466)
);

FAx1_ASAP7_75t_SL g472 ( 
.A(n_466),
.B(n_461),
.CI(n_260),
.CON(n_472),
.SN(n_472)
);

MAJx2_ASAP7_75t_L g467 ( 
.A(n_457),
.B(n_302),
.C(n_354),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_467),
.B(n_456),
.C(n_461),
.Y(n_471)
);

AOI21xp5_ASAP7_75t_L g473 ( 
.A1(n_470),
.A2(n_472),
.B(n_468),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_L g474 ( 
.A1(n_471),
.A2(n_211),
.B(n_465),
.Y(n_474)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_473),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_475),
.B(n_474),
.Y(n_476)
);


endmodule