module fake_jpeg_16124_n_94 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_8, n_15, n_7, n_94);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_94;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_24),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_9),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx2_ASAP7_75t_R g40 ( 
.A(n_15),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_41),
.Y(n_42)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

BUFx24_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_40),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_44),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_49)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_46),
.Y(n_56)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_37),
.B(n_0),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_6),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_1),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_48),
.B(n_3),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_52),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_44),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_55),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_34),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_57),
.Y(n_72)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_41),
.C(n_38),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_46),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_58)
);

AOI22x1_ASAP7_75t_L g75 ( 
.A1(n_58),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_59),
.B(n_10),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_42),
.A2(n_36),
.B1(n_33),
.B2(n_32),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_60),
.A2(n_12),
.B1(n_13),
.B2(n_16),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_57),
.B(n_7),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_61),
.B(n_71),
.Y(n_82)
);

AND2x2_ASAP7_75t_SL g62 ( 
.A(n_51),
.B(n_35),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_63),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_60),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_67),
.Y(n_81)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g78 ( 
.A(n_69),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_70),
.A2(n_73),
.B1(n_74),
.B2(n_75),
.Y(n_80)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_52),
.B(n_17),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_60),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_64),
.A2(n_22),
.B1(n_23),
.B2(n_26),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_76),
.B(n_75),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_61),
.C(n_72),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_83),
.B(n_84),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_79),
.Y(n_84)
);

AOI322xp5_ASAP7_75t_SL g87 ( 
.A1(n_85),
.A2(n_80),
.A3(n_76),
.B1(n_77),
.B2(n_72),
.C1(n_66),
.C2(n_62),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_87),
.A2(n_66),
.B(n_82),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_88),
.A2(n_86),
.B(n_81),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_89),
.B(n_86),
.Y(n_90)
);

OAI21xp33_ASAP7_75t_L g91 ( 
.A1(n_90),
.A2(n_28),
.B(n_29),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_91),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_92),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_78),
.C(n_30),
.Y(n_94)
);


endmodule