module fake_jpeg_10752_n_110 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_110);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_110;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

INVx6_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

BUFx16f_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_20),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_35),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_14),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_45),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_51),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_L g49 ( 
.A1(n_44),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_49)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_19),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_36),
.A2(n_21),
.B1(n_33),
.B2(n_32),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_52),
.B(n_55),
.C(n_42),
.Y(n_63)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_46),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_55),
.B(n_37),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_47),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_59),
.Y(n_80)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_42),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_63),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_52),
.B(n_41),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_37),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_67),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_57),
.A2(n_54),
.B1(n_43),
.B2(n_40),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_68),
.A2(n_70),
.B1(n_74),
.B2(n_75),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_L g70 ( 
.A1(n_66),
.A2(n_39),
.B1(n_38),
.B2(n_43),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_59),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_62),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_73),
.B(n_76),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_56),
.A2(n_40),
.B1(n_37),
.B2(n_7),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_58),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_56),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_65),
.A2(n_8),
.B1(n_9),
.B2(n_34),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_77),
.A2(n_11),
.B(n_12),
.Y(n_88)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_79),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_71),
.B(n_67),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_81),
.B(n_82),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_80),
.B(n_62),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_84),
.A2(n_88),
.B(n_93),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_13),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_89),
.B(n_90),
.C(n_91),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_77),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_69),
.B(n_16),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_17),
.Y(n_92)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_92),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_69),
.B(n_18),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_84),
.B(n_22),
.C(n_23),
.Y(n_94)
);

AND2x2_ASAP7_75t_SL g103 ( 
.A(n_94),
.B(n_28),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_83),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_99),
.A2(n_87),
.B1(n_86),
.B2(n_91),
.Y(n_102)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_98),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_101),
.B(n_102),
.C(n_103),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_103),
.A2(n_96),
.B(n_95),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_100),
.Y(n_106)
);

NOR4xp25_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_104),
.C(n_85),
.D(n_94),
.Y(n_107)
);

AO21x1_ASAP7_75t_L g108 ( 
.A1(n_107),
.A2(n_97),
.B(n_29),
.Y(n_108)
);

BUFx24_ASAP7_75t_SL g109 ( 
.A(n_108),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_30),
.Y(n_110)
);


endmodule