module fake_jpeg_4249_n_279 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_279);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_279;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_21;
wire n_57;
wire n_187;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx24_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_32),
.B(n_35),
.Y(n_51)
);

INVx4_ASAP7_75t_SL g33 ( 
.A(n_22),
.Y(n_33)
);

INVx3_ASAP7_75t_SL g56 ( 
.A(n_33),
.Y(n_56)
);

BUFx24_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_22),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_15),
.B(n_26),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_37),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_27),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_42),
.B(n_49),
.Y(n_77)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_39),
.A2(n_16),
.B1(n_24),
.B2(n_28),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_46),
.A2(n_21),
.B1(n_28),
.B2(n_17),
.Y(n_87)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_48),
.Y(n_88)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx6_ASAP7_75t_SL g50 ( 
.A(n_34),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_53),
.B(n_58),
.Y(n_78)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_37),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_61),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_32),
.A2(n_16),
.B1(n_24),
.B2(n_23),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_62),
.A2(n_23),
.B1(n_29),
.B2(n_35),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_32),
.B(n_26),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_18),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_65),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_52),
.A2(n_39),
.B1(n_41),
.B2(n_24),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_67),
.A2(n_71),
.B1(n_81),
.B2(n_62),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_SL g103 ( 
.A(n_68),
.B(n_31),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_69),
.A2(n_73),
.B(n_50),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_52),
.A2(n_29),
.B1(n_35),
.B2(n_23),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_70),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_L g71 ( 
.A1(n_63),
.A2(n_39),
.B1(n_40),
.B2(n_29),
.Y(n_71)
);

AND2x4_ASAP7_75t_SL g73 ( 
.A(n_56),
.B(n_34),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_42),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_75),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_61),
.A2(n_35),
.B1(n_28),
.B2(n_21),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_79),
.A2(n_87),
.B1(n_15),
.B2(n_18),
.Y(n_100)
);

OA22x2_ASAP7_75t_L g81 ( 
.A1(n_56),
.A2(n_34),
.B1(n_22),
.B2(n_30),
.Y(n_81)
);

OAI32xp33_ASAP7_75t_L g85 ( 
.A1(n_56),
.A2(n_15),
.A3(n_18),
.B1(n_26),
.B2(n_31),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_44),
.Y(n_98)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_89),
.B(n_92),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_90),
.A2(n_91),
.B1(n_97),
.B2(n_108),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_75),
.A2(n_65),
.B1(n_53),
.B2(n_48),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_93),
.B(n_96),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_84),
.B(n_51),
.Y(n_94)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_94),
.Y(n_129)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_66),
.A2(n_49),
.B1(n_45),
.B2(n_43),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_98),
.B(n_73),
.Y(n_121)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_74),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_99),
.A2(n_109),
.B1(n_112),
.B2(n_80),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_100),
.A2(n_102),
.B(n_73),
.Y(n_119)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_101),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_103),
.B(n_78),
.Y(n_127)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_104),
.B(n_105),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_20),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_66),
.B(n_30),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_106),
.B(n_76),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_81),
.A2(n_57),
.B1(n_21),
.B2(n_17),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_81),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_84),
.B(n_19),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_110),
.Y(n_114)
);

BUFx8_ASAP7_75t_L g111 ( 
.A(n_73),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_111),
.Y(n_124)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_78),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_113),
.B(n_128),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_107),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_115),
.Y(n_153)
);

AOI322xp5_ASAP7_75t_L g116 ( 
.A1(n_104),
.A2(n_98),
.A3(n_111),
.B1(n_102),
.B2(n_96),
.C1(n_93),
.C2(n_89),
.Y(n_116)
);

BUFx24_ASAP7_75t_SL g154 ( 
.A(n_116),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_119),
.A2(n_123),
.B1(n_136),
.B2(n_31),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_121),
.A2(n_126),
.B1(n_133),
.B2(n_88),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_111),
.A2(n_81),
.B(n_85),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_125),
.A2(n_124),
.B(n_136),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_109),
.A2(n_81),
.B1(n_82),
.B2(n_76),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_134),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_106),
.B(n_82),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_112),
.B(n_103),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_131),
.B(n_47),
.Y(n_156)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_92),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_132),
.B(n_135),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_95),
.A2(n_72),
.B1(n_80),
.B2(n_83),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_90),
.B(n_86),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_97),
.Y(n_135)
);

AO21x2_ASAP7_75t_L g136 ( 
.A1(n_108),
.A2(n_88),
.B(n_34),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_117),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_137),
.B(n_138),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_115),
.B(n_99),
.Y(n_138)
);

INVx13_ASAP7_75t_L g139 ( 
.A(n_129),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_139),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_131),
.B(n_91),
.C(n_72),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_140),
.B(n_149),
.C(n_158),
.Y(n_162)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_113),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_141),
.B(n_145),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_143),
.A2(n_47),
.B(n_27),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_124),
.A2(n_95),
.B1(n_17),
.B2(n_83),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_144),
.A2(n_151),
.B1(n_152),
.B2(n_153),
.Y(n_163)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_118),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_119),
.A2(n_88),
.B(n_22),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_146),
.A2(n_27),
.B(n_25),
.Y(n_178)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_117),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_147),
.A2(n_150),
.B1(n_159),
.B2(n_137),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_127),
.B(n_134),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_122),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_136),
.A2(n_135),
.B1(n_121),
.B2(n_125),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_152),
.A2(n_130),
.B1(n_114),
.B2(n_129),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_156),
.B(n_126),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_130),
.A2(n_121),
.B1(n_136),
.B2(n_120),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_157),
.A2(n_160),
.B1(n_57),
.B2(n_30),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_128),
.B(n_30),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_133),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_136),
.Y(n_161)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_161),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_163),
.B(n_60),
.Y(n_202)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_165),
.Y(n_187)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_166),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_143),
.A2(n_114),
.B1(n_132),
.B2(n_101),
.Y(n_167)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_167),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_155),
.B(n_30),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_168),
.B(n_174),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_169),
.B(n_171),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_148),
.B(n_47),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_172),
.B(n_181),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_155),
.B(n_30),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_175),
.A2(n_19),
.B(n_25),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_149),
.B(n_148),
.C(n_156),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_176),
.B(n_177),
.C(n_179),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_140),
.B(n_31),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_178),
.A2(n_145),
.B(n_147),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_158),
.B(n_54),
.C(n_60),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_141),
.B(n_31),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_180),
.B(n_182),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_157),
.B(n_27),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_142),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_151),
.A2(n_19),
.B1(n_25),
.B2(n_11),
.Y(n_184)
);

A2O1A1Ixp33_ASAP7_75t_SL g203 ( 
.A1(n_184),
.A2(n_0),
.B(n_2),
.C(n_3),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_176),
.B(n_146),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_185),
.B(n_194),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_173),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_188),
.B(n_199),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_190),
.A2(n_191),
.B(n_192),
.Y(n_214)
);

AO22x1_ASAP7_75t_L g191 ( 
.A1(n_175),
.A2(n_161),
.B1(n_144),
.B2(n_139),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_172),
.B(n_162),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_162),
.B(n_177),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_196),
.B(n_198),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_170),
.A2(n_154),
.B1(n_25),
.B2(n_19),
.Y(n_197)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_197),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_181),
.B(n_60),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_183),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_163),
.B(n_64),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_201),
.B(n_179),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_202),
.A2(n_164),
.B1(n_184),
.B2(n_180),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_203),
.A2(n_178),
.B1(n_170),
.B2(n_191),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_206),
.B(n_217),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_207),
.A2(n_203),
.B1(n_2),
.B2(n_3),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_194),
.B(n_174),
.C(n_168),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_209),
.B(n_210),
.C(n_197),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_195),
.B(n_165),
.C(n_169),
.Y(n_210)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_213),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_185),
.B(n_164),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_215),
.B(n_222),
.Y(n_226)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_205),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_188),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_218),
.B(n_219),
.Y(n_232)
);

FAx1_ASAP7_75t_SL g219 ( 
.A(n_189),
.B(n_9),
.CI(n_14),
.CON(n_219),
.SN(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_186),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_220),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_200),
.A2(n_9),
.B(n_14),
.Y(n_221)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_221),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_189),
.B(n_54),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_215),
.B(n_195),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_223),
.B(n_211),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_214),
.A2(n_193),
.B1(n_187),
.B2(n_202),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_225),
.A2(n_227),
.B1(n_228),
.B2(n_231),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_218),
.A2(n_204),
.B1(n_203),
.B2(n_198),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_208),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_229),
.B(n_236),
.Y(n_246)
);

OR2x2_ASAP7_75t_L g231 ( 
.A(n_214),
.B(n_203),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_231),
.B(n_219),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_234),
.B(n_216),
.C(n_206),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_211),
.B(n_54),
.C(n_59),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_235),
.B(n_210),
.C(n_216),
.Y(n_240)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_209),
.Y(n_236)
);

AO21x1_ASAP7_75t_L g259 ( 
.A1(n_238),
.A2(n_249),
.B(n_5),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_239),
.B(n_243),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_240),
.B(n_244),
.Y(n_254)
);

BUFx24_ASAP7_75t_SL g241 ( 
.A(n_233),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_241),
.B(n_247),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_242),
.A2(n_6),
.B(n_11),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_223),
.B(n_222),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_235),
.B(n_212),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_245),
.B(n_237),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_226),
.B(n_8),
.C(n_14),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_226),
.B(n_234),
.C(n_224),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_248),
.B(n_239),
.Y(n_258)
);

A2O1A1O1Ixp25_ASAP7_75t_L g249 ( 
.A1(n_232),
.A2(n_7),
.B(n_13),
.C(n_12),
.D(n_11),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_246),
.A2(n_230),
.B1(n_227),
.B2(n_225),
.Y(n_250)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_250),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_249),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_251),
.A2(n_256),
.B(n_257),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_255),
.B(n_259),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_240),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_258),
.B(n_5),
.C(n_10),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_256),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_259),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_253),
.B(n_5),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_263),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_264),
.B(n_265),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_253),
.B(n_6),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_261),
.B(n_255),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_267),
.B(n_269),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_262),
.A2(n_254),
.B(n_252),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_271),
.A2(n_266),
.B(n_265),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_272),
.A2(n_274),
.B(n_8),
.Y(n_276)
);

MAJx2_ASAP7_75t_L g274 ( 
.A(n_268),
.B(n_264),
.C(n_58),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_273),
.A2(n_270),
.B(n_6),
.Y(n_275)
);

AOI322xp5_ASAP7_75t_L g277 ( 
.A1(n_275),
.A2(n_276),
.A3(n_10),
.B1(n_2),
.B2(n_3),
.C1(n_4),
.C2(n_0),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_277),
.A2(n_0),
.B(n_4),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_278),
.B(n_0),
.Y(n_279)
);


endmodule