module real_jpeg_7942_n_7 (n_5, n_4, n_36, n_0, n_39, n_37, n_40, n_1, n_41, n_2, n_38, n_6, n_3, n_7);

input n_5;
input n_4;
input n_36;
input n_0;
input n_39;
input n_37;
input n_40;
input n_1;
input n_41;
input n_2;
input n_38;
input n_6;
input n_3;

output n_7;

wire n_17;
wire n_8;
wire n_21;
wire n_33;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_22;
wire n_18;
wire n_26;
wire n_32;
wire n_20;
wire n_27;
wire n_19;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

OAI22xp5_ASAP7_75t_L g8 ( 
.A1(n_0),
.A2(n_9),
.B1(n_10),
.B2(n_14),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_0),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_1),
.B(n_20),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_2),
.B(n_18),
.C(n_26),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_4),
.B(n_16),
.C(n_32),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_5),
.B(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_5),
.B(n_25),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_5),
.B(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_5),
.B(n_31),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

XOR2xp5_ASAP7_75t_L g7 ( 
.A(n_8),
.B(n_15),
.Y(n_7)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_12),
.Y(n_10)
);

BUFx3_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_28),
.C(n_29),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_22),
.C(n_23),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_34),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_36),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_37),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_38),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_39),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_40),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_41),
.Y(n_33)
);


endmodule