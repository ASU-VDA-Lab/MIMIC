module fake_netlist_6_2800_n_787 (n_52, n_16, n_1, n_91, n_119, n_46, n_18, n_21, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_127, n_125, n_77, n_106, n_92, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_787);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_127;
input n_125;
input n_77;
input n_106;
input n_92;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_787;

wire n_591;
wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_148;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_144;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_783;
wire n_725;
wire n_358;
wire n_160;
wire n_751;
wire n_449;
wire n_749;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_255;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_781;
wire n_424;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_222;
wire n_179;
wire n_248;
wire n_300;
wire n_517;
wire n_718;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_147;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_693;
wire n_167;
wire n_631;
wire n_174;
wire n_516;
wire n_720;
wire n_153;
wire n_758;
wire n_525;
wire n_611;
wire n_156;
wire n_491;
wire n_145;
wire n_656;
wire n_772;
wire n_666;
wire n_371;
wire n_770;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_155;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_777;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_163;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_154;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_152;
wire n_623;
wire n_599;
wire n_513;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_325;
wire n_767;
wire n_329;
wire n_464;
wire n_600;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_159;
wire n_157;
wire n_162;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_146;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_193;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_149;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_728;
wire n_681;
wire n_729;
wire n_151;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_722;
wire n_688;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_170;
wire n_778;
wire n_332;
wire n_336;
wire n_410;
wire n_398;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_105),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_103),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_70),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_114),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_82),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_117),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_125),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_90),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g152 ( 
.A(n_36),
.B(n_25),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_12),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_121),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_137),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_88),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_86),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_31),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_53),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_40),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_122),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_89),
.B(n_133),
.Y(n_162)
);

INVx2_ASAP7_75t_SL g163 ( 
.A(n_84),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_12),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_61),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_96),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_47),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_1),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_13),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_85),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_46),
.Y(n_171)
);

INVx2_ASAP7_75t_SL g172 ( 
.A(n_11),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_104),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_59),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_129),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_115),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_116),
.Y(n_177)
);

BUFx2_ASAP7_75t_SL g178 ( 
.A(n_136),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_128),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_34),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_30),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_60),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_23),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_135),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_13),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_41),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_130),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_52),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_99),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_58),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_108),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_75),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_67),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_42),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_141),
.Y(n_195)
);

BUFx5_ASAP7_75t_L g196 ( 
.A(n_134),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_62),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_81),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_24),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_196),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_168),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_181),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_181),
.Y(n_203)
);

BUFx12f_ASAP7_75t_L g204 ( 
.A(n_185),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_164),
.Y(n_205)
);

BUFx12f_ASAP7_75t_L g206 ( 
.A(n_172),
.Y(n_206)
);

OAI22x1_ASAP7_75t_SL g207 ( 
.A1(n_153),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_145),
.Y(n_208)
);

OAI22x1_ASAP7_75t_R g209 ( 
.A1(n_171),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_209)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_164),
.Y(n_210)
);

AND2x4_ASAP7_75t_L g211 ( 
.A(n_163),
.B(n_18),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_166),
.B(n_3),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_196),
.B(n_4),
.Y(n_213)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_196),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_196),
.Y(n_215)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_144),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_196),
.Y(n_217)
);

INVx5_ASAP7_75t_L g218 ( 
.A(n_196),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_169),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_146),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_161),
.B(n_4),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_147),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_148),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_150),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_171),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_154),
.B(n_5),
.Y(n_226)
);

INVx2_ASAP7_75t_SL g227 ( 
.A(n_156),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_160),
.Y(n_228)
);

INVx5_ASAP7_75t_L g229 ( 
.A(n_178),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_165),
.Y(n_230)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_177),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_182),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_180),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_183),
.B(n_5),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_184),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_186),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_189),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_190),
.Y(n_238)
);

AND2x4_ASAP7_75t_L g239 ( 
.A(n_199),
.B(n_152),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_180),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_149),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_151),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_241),
.Y(n_243)
);

BUFx2_ASAP7_75t_L g244 ( 
.A(n_241),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_225),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_225),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_202),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_233),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_233),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_204),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_204),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_242),
.B(n_155),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_240),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_216),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_216),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_202),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_216),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_222),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_202),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_206),
.Y(n_260)
);

NOR2xp67_ASAP7_75t_L g261 ( 
.A(n_229),
.B(n_162),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_206),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_201),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_R g264 ( 
.A(n_212),
.B(n_167),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_202),
.Y(n_265)
);

BUFx2_ASAP7_75t_L g266 ( 
.A(n_219),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_202),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_203),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_203),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_203),
.Y(n_270)
);

NAND2xp33_ASAP7_75t_SL g271 ( 
.A(n_226),
.B(n_213),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_222),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_203),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_203),
.Y(n_274)
);

INVxp67_ASAP7_75t_SL g275 ( 
.A(n_235),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_229),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_229),
.Y(n_277)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_224),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_229),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_209),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_229),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_208),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_208),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_R g284 ( 
.A(n_231),
.B(n_197),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_230),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_223),
.Y(n_286)
);

NAND2x1p5_ASAP7_75t_L g287 ( 
.A(n_211),
.B(n_226),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_223),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_228),
.Y(n_289)
);

BUFx3_ASAP7_75t_L g290 ( 
.A(n_230),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_239),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_265),
.B(n_239),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_284),
.B(n_211),
.Y(n_293)
);

BUFx6f_ASAP7_75t_SL g294 ( 
.A(n_290),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_266),
.B(n_239),
.Y(n_295)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_247),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_247),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_282),
.B(n_283),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_268),
.B(n_211),
.Y(n_299)
);

INVx2_ASAP7_75t_SL g300 ( 
.A(n_285),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_290),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_278),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_269),
.B(n_220),
.Y(n_303)
);

AO221x1_ASAP7_75t_L g304 ( 
.A1(n_271),
.A2(n_231),
.B1(n_224),
.B2(n_237),
.C(n_220),
.Y(n_304)
);

INVx2_ASAP7_75t_SL g305 ( 
.A(n_252),
.Y(n_305)
);

BUFx6f_ASAP7_75t_SL g306 ( 
.A(n_286),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_291),
.B(n_254),
.Y(n_307)
);

INVx2_ASAP7_75t_SL g308 ( 
.A(n_253),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_255),
.B(n_221),
.Y(n_309)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_278),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_257),
.B(n_234),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_256),
.Y(n_312)
);

CKINVDCx14_ASAP7_75t_R g313 ( 
.A(n_264),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_278),
.Y(n_314)
);

INVx4_ASAP7_75t_L g315 ( 
.A(n_273),
.Y(n_315)
);

INVx2_ASAP7_75t_SL g316 ( 
.A(n_244),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_259),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_274),
.B(n_232),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_287),
.B(n_232),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_267),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_275),
.B(n_238),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_287),
.B(n_238),
.Y(n_322)
);

NAND3xp33_ASAP7_75t_L g323 ( 
.A(n_271),
.B(n_236),
.C(n_228),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_276),
.B(n_231),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_243),
.B(n_157),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_277),
.B(n_236),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_279),
.B(n_224),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_281),
.B(n_260),
.Y(n_328)
);

INVx1_ASAP7_75t_SL g329 ( 
.A(n_248),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_288),
.B(n_227),
.Y(n_330)
);

BUFx5_ASAP7_75t_L g331 ( 
.A(n_270),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_289),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_258),
.B(n_227),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_258),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_246),
.Y(n_335)
);

NAND2xp33_ASAP7_75t_L g336 ( 
.A(n_272),
.B(n_158),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_272),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_262),
.Y(n_338)
);

BUFx5_ASAP7_75t_L g339 ( 
.A(n_261),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_263),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_249),
.B(n_224),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_250),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_251),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_245),
.B(n_224),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_245),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_280),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_280),
.B(n_237),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_247),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_247),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_247),
.Y(n_350)
);

OAI221xp5_ASAP7_75t_L g351 ( 
.A1(n_271),
.A2(n_205),
.B1(n_210),
.B2(n_162),
.C(n_237),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_265),
.B(n_237),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_284),
.B(n_159),
.Y(n_353)
);

AND2x4_ASAP7_75t_L g354 ( 
.A(n_290),
.B(n_205),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_291),
.B(n_237),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_247),
.Y(n_356)
);

BUFx2_ASAP7_75t_L g357 ( 
.A(n_347),
.Y(n_357)
);

BUFx2_ASAP7_75t_L g358 ( 
.A(n_316),
.Y(n_358)
);

OR2x6_ASAP7_75t_L g359 ( 
.A(n_308),
.B(n_209),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_313),
.Y(n_360)
);

INVx2_ASAP7_75t_SL g361 ( 
.A(n_295),
.Y(n_361)
);

NAND2x1p5_ASAP7_75t_L g362 ( 
.A(n_301),
.B(n_210),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_354),
.Y(n_363)
);

AND2x4_ASAP7_75t_L g364 ( 
.A(n_354),
.B(n_301),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_305),
.B(n_170),
.Y(n_365)
);

NAND3xp33_ASAP7_75t_SL g366 ( 
.A(n_293),
.B(n_173),
.C(n_174),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_311),
.B(n_175),
.Y(n_367)
);

INVx4_ASAP7_75t_L g368 ( 
.A(n_301),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_334),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_315),
.B(n_176),
.Y(n_370)
);

BUFx3_ASAP7_75t_L g371 ( 
.A(n_338),
.Y(n_371)
);

AND2x4_ASAP7_75t_L g372 ( 
.A(n_323),
.B(n_210),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_319),
.B(n_200),
.Y(n_373)
);

INVx8_ASAP7_75t_L g374 ( 
.A(n_294),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_322),
.B(n_200),
.Y(n_375)
);

OAI22xp33_ASAP7_75t_L g376 ( 
.A1(n_292),
.A2(n_194),
.B1(n_187),
.B2(n_188),
.Y(n_376)
);

OR2x2_ASAP7_75t_L g377 ( 
.A(n_340),
.B(n_6),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_321),
.B(n_179),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_299),
.B(n_215),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_337),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_315),
.B(n_191),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_341),
.B(n_192),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_300),
.B(n_193),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_303),
.B(n_215),
.Y(n_384)
);

INVx2_ASAP7_75t_SL g385 ( 
.A(n_318),
.Y(n_385)
);

INVx3_ASAP7_75t_L g386 ( 
.A(n_349),
.Y(n_386)
);

INVx3_ASAP7_75t_L g387 ( 
.A(n_349),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_332),
.Y(n_388)
);

INVx3_ASAP7_75t_L g389 ( 
.A(n_349),
.Y(n_389)
);

AND2x4_ASAP7_75t_L g390 ( 
.A(n_297),
.B(n_195),
.Y(n_390)
);

BUFx12f_ASAP7_75t_SL g391 ( 
.A(n_338),
.Y(n_391)
);

AND2x6_ASAP7_75t_SL g392 ( 
.A(n_346),
.B(n_344),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_348),
.Y(n_393)
);

INVx6_ASAP7_75t_L g394 ( 
.A(n_338),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_310),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_355),
.B(n_217),
.Y(n_396)
);

INVx5_ASAP7_75t_L g397 ( 
.A(n_356),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_307),
.B(n_198),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_350),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_309),
.B(n_217),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_310),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_312),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_317),
.Y(n_403)
);

INVx5_ASAP7_75t_L g404 ( 
.A(n_356),
.Y(n_404)
);

INVx2_ASAP7_75t_SL g405 ( 
.A(n_324),
.Y(n_405)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_356),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_352),
.B(n_214),
.Y(n_407)
);

AOI22xp33_ASAP7_75t_L g408 ( 
.A1(n_304),
.A2(n_351),
.B1(n_314),
.B2(n_302),
.Y(n_408)
);

NOR3xp33_ASAP7_75t_SL g409 ( 
.A(n_346),
.B(n_207),
.C(n_7),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_331),
.B(n_214),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_335),
.A2(n_218),
.B1(n_214),
.B2(n_8),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_333),
.A2(n_214),
.B1(n_218),
.B2(n_8),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_296),
.Y(n_413)
);

AOI22xp33_ASAP7_75t_SL g414 ( 
.A1(n_306),
.A2(n_218),
.B1(n_214),
.B2(n_9),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_296),
.Y(n_415)
);

NOR2x1p5_ASAP7_75t_L g416 ( 
.A(n_343),
.B(n_6),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_325),
.B(n_7),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_330),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_320),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_320),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_320),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_336),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_327),
.Y(n_423)
);

BUFx12f_ASAP7_75t_SL g424 ( 
.A(n_294),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_326),
.Y(n_425)
);

AO22x1_ASAP7_75t_L g426 ( 
.A1(n_417),
.A2(n_345),
.B1(n_329),
.B2(n_342),
.Y(n_426)
);

OR2x6_ASAP7_75t_L g427 ( 
.A(n_374),
.B(n_298),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_R g428 ( 
.A(n_391),
.B(n_360),
.Y(n_428)
);

OR2x6_ASAP7_75t_L g429 ( 
.A(n_374),
.B(n_328),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_369),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_402),
.Y(n_431)
);

AOI21x1_ASAP7_75t_L g432 ( 
.A1(n_410),
.A2(n_353),
.B(n_331),
.Y(n_432)
);

O2A1O1Ixp33_ASAP7_75t_L g433 ( 
.A1(n_411),
.A2(n_306),
.B(n_10),
.C(n_11),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_425),
.A2(n_218),
.B1(n_339),
.B2(n_331),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_L g435 ( 
.A1(n_423),
.A2(n_218),
.B1(n_339),
.B2(n_331),
.Y(n_435)
);

OR2x6_ASAP7_75t_L g436 ( 
.A(n_374),
.B(n_9),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g437 ( 
.A1(n_373),
.A2(n_339),
.B(n_331),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_380),
.Y(n_438)
);

O2A1O1Ixp33_ASAP7_75t_SL g439 ( 
.A1(n_422),
.A2(n_367),
.B(n_379),
.C(n_375),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_L g440 ( 
.A1(n_373),
.A2(n_339),
.B(n_87),
.Y(n_440)
);

OA21x2_ASAP7_75t_L g441 ( 
.A1(n_375),
.A2(n_339),
.B(n_91),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_385),
.B(n_10),
.Y(n_442)
);

O2A1O1Ixp33_ASAP7_75t_SL g443 ( 
.A1(n_379),
.A2(n_14),
.B(n_15),
.C(n_16),
.Y(n_443)
);

OR2x6_ASAP7_75t_L g444 ( 
.A(n_394),
.B(n_14),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_403),
.Y(n_445)
);

INVx3_ASAP7_75t_L g446 ( 
.A(n_413),
.Y(n_446)
);

INVx3_ASAP7_75t_L g447 ( 
.A(n_394),
.Y(n_447)
);

AOI21xp5_ASAP7_75t_L g448 ( 
.A1(n_396),
.A2(n_92),
.B(n_142),
.Y(n_448)
);

NOR2x1_ASAP7_75t_SL g449 ( 
.A(n_366),
.B(n_397),
.Y(n_449)
);

INVx6_ASAP7_75t_L g450 ( 
.A(n_371),
.Y(n_450)
);

NOR2xp67_ASAP7_75t_L g451 ( 
.A(n_361),
.B(n_19),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_424),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_357),
.A2(n_83),
.B1(n_140),
.B2(n_139),
.Y(n_453)
);

A2O1A1Ixp33_ASAP7_75t_L g454 ( 
.A1(n_384),
.A2(n_405),
.B(n_378),
.C(n_372),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_L g455 ( 
.A1(n_418),
.A2(n_408),
.B1(n_396),
.B2(n_384),
.Y(n_455)
);

AOI21xp5_ASAP7_75t_L g456 ( 
.A1(n_407),
.A2(n_410),
.B(n_400),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_372),
.B(n_15),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_388),
.A2(n_80),
.B1(n_138),
.B2(n_20),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_364),
.B(n_21),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_358),
.B(n_16),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_415),
.B(n_17),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_SL g462 ( 
.A(n_359),
.B(n_22),
.Y(n_462)
);

O2A1O1Ixp33_ASAP7_75t_L g463 ( 
.A1(n_411),
.A2(n_376),
.B(n_377),
.C(n_363),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_393),
.B(n_17),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_L g465 ( 
.A1(n_407),
.A2(n_26),
.B(n_27),
.Y(n_465)
);

AND2x4_ASAP7_75t_L g466 ( 
.A(n_364),
.B(n_28),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_399),
.Y(n_467)
);

INVx1_ASAP7_75t_SL g468 ( 
.A(n_390),
.Y(n_468)
);

NOR2x1_ASAP7_75t_R g469 ( 
.A(n_368),
.B(n_29),
.Y(n_469)
);

BUFx12f_ASAP7_75t_L g470 ( 
.A(n_392),
.Y(n_470)
);

AOI21xp5_ASAP7_75t_L g471 ( 
.A1(n_395),
.A2(n_32),
.B(n_33),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_401),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_386),
.B(n_35),
.Y(n_473)
);

AND2x4_ASAP7_75t_L g474 ( 
.A(n_368),
.B(n_390),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_419),
.Y(n_475)
);

INVxp67_ASAP7_75t_SL g476 ( 
.A(n_386),
.Y(n_476)
);

CKINVDCx6p67_ASAP7_75t_R g477 ( 
.A(n_359),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_420),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_359),
.B(n_37),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_382),
.A2(n_38),
.B1(n_39),
.B2(n_43),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_398),
.B(n_44),
.Y(n_481)
);

AOI21x1_ASAP7_75t_L g482 ( 
.A1(n_421),
.A2(n_365),
.B(n_370),
.Y(n_482)
);

AOI21xp5_ASAP7_75t_L g483 ( 
.A1(n_397),
.A2(n_45),
.B(n_48),
.Y(n_483)
);

OR2x6_ASAP7_75t_L g484 ( 
.A(n_450),
.B(n_444),
.Y(n_484)
);

CKINVDCx11_ASAP7_75t_R g485 ( 
.A(n_470),
.Y(n_485)
);

BUFx2_ASAP7_75t_L g486 ( 
.A(n_450),
.Y(n_486)
);

NOR2xp67_ASAP7_75t_L g487 ( 
.A(n_452),
.B(n_383),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_431),
.Y(n_488)
);

INVx6_ASAP7_75t_L g489 ( 
.A(n_474),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_L g490 ( 
.A1(n_455),
.A2(n_412),
.B(n_381),
.Y(n_490)
);

BUFx12f_ASAP7_75t_L g491 ( 
.A(n_436),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_466),
.Y(n_492)
);

BUFx2_ASAP7_75t_L g493 ( 
.A(n_428),
.Y(n_493)
);

BUFx3_ASAP7_75t_L g494 ( 
.A(n_447),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_466),
.Y(n_495)
);

BUFx3_ASAP7_75t_L g496 ( 
.A(n_474),
.Y(n_496)
);

OAI21x1_ASAP7_75t_L g497 ( 
.A1(n_456),
.A2(n_406),
.B(n_387),
.Y(n_497)
);

INVx2_ASAP7_75t_SL g498 ( 
.A(n_460),
.Y(n_498)
);

AOI21xp33_ASAP7_75t_L g499 ( 
.A1(n_463),
.A2(n_468),
.B(n_481),
.Y(n_499)
);

OAI21xp5_ASAP7_75t_L g500 ( 
.A1(n_454),
.A2(n_437),
.B(n_440),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_445),
.B(n_387),
.Y(n_501)
);

INVx1_ASAP7_75t_SL g502 ( 
.A(n_444),
.Y(n_502)
);

HB1xp67_ASAP7_75t_L g503 ( 
.A(n_457),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_430),
.Y(n_504)
);

OAI21xp5_ASAP7_75t_L g505 ( 
.A1(n_439),
.A2(n_412),
.B(n_389),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_467),
.Y(n_506)
);

INVx1_ASAP7_75t_SL g507 ( 
.A(n_479),
.Y(n_507)
);

INVxp33_ASAP7_75t_L g508 ( 
.A(n_442),
.Y(n_508)
);

BUFx2_ASAP7_75t_R g509 ( 
.A(n_459),
.Y(n_509)
);

OAI21x1_ASAP7_75t_L g510 ( 
.A1(n_432),
.A2(n_406),
.B(n_389),
.Y(n_510)
);

BUFx2_ASAP7_75t_SL g511 ( 
.A(n_451),
.Y(n_511)
);

INVx2_ASAP7_75t_SL g512 ( 
.A(n_464),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_438),
.Y(n_513)
);

OAI21x1_ASAP7_75t_L g514 ( 
.A1(n_473),
.A2(n_362),
.B(n_416),
.Y(n_514)
);

AO21x2_ASAP7_75t_L g515 ( 
.A1(n_434),
.A2(n_435),
.B(n_465),
.Y(n_515)
);

INVx1_ASAP7_75t_SL g516 ( 
.A(n_477),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_482),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_475),
.B(n_392),
.Y(n_518)
);

AND2x4_ASAP7_75t_L g519 ( 
.A(n_472),
.B(n_397),
.Y(n_519)
);

INVx1_ASAP7_75t_SL g520 ( 
.A(n_426),
.Y(n_520)
);

OAI21x1_ASAP7_75t_L g521 ( 
.A1(n_448),
.A2(n_404),
.B(n_50),
.Y(n_521)
);

NAND2x1p5_ASAP7_75t_L g522 ( 
.A(n_446),
.B(n_404),
.Y(n_522)
);

AO21x2_ASAP7_75t_L g523 ( 
.A1(n_449),
.A2(n_409),
.B(n_404),
.Y(n_523)
);

AOI22x1_ASAP7_75t_L g524 ( 
.A1(n_478),
.A2(n_446),
.B1(n_476),
.B2(n_471),
.Y(n_524)
);

AO21x2_ASAP7_75t_L g525 ( 
.A1(n_461),
.A2(n_414),
.B(n_51),
.Y(n_525)
);

OR2x6_ASAP7_75t_L g526 ( 
.A(n_427),
.B(n_49),
.Y(n_526)
);

OAI21x1_ASAP7_75t_L g527 ( 
.A1(n_441),
.A2(n_54),
.B(n_55),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_427),
.B(n_56),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_443),
.Y(n_529)
);

OAI21x1_ASAP7_75t_L g530 ( 
.A1(n_441),
.A2(n_57),
.B(n_63),
.Y(n_530)
);

INVx3_ASAP7_75t_L g531 ( 
.A(n_429),
.Y(n_531)
);

INVx2_ASAP7_75t_SL g532 ( 
.A(n_436),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_504),
.Y(n_533)
);

NAND2x1p5_ASAP7_75t_L g534 ( 
.A(n_517),
.B(n_453),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_503),
.B(n_462),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_488),
.Y(n_536)
);

OAI21x1_ASAP7_75t_L g537 ( 
.A1(n_510),
.A2(n_483),
.B(n_480),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_504),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_503),
.B(n_433),
.Y(n_539)
);

BUFx4f_ASAP7_75t_SL g540 ( 
.A(n_486),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_485),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_506),
.Y(n_542)
);

BUFx12f_ASAP7_75t_L g543 ( 
.A(n_485),
.Y(n_543)
);

AOI22xp33_ASAP7_75t_SL g544 ( 
.A1(n_520),
.A2(n_429),
.B1(n_469),
.B2(n_458),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_529),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_513),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_501),
.Y(n_547)
);

BUFx3_ASAP7_75t_L g548 ( 
.A(n_493),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_512),
.B(n_64),
.Y(n_549)
);

CKINVDCx6p67_ASAP7_75t_R g550 ( 
.A(n_484),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_522),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_510),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_517),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_490),
.B(n_65),
.Y(n_554)
);

BUFx2_ASAP7_75t_L g555 ( 
.A(n_484),
.Y(n_555)
);

AOI22xp33_ASAP7_75t_SL g556 ( 
.A1(n_518),
.A2(n_66),
.B1(n_68),
.B2(n_69),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_517),
.Y(n_557)
);

AOI22xp33_ASAP7_75t_SL g558 ( 
.A1(n_518),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_558)
);

AOI21x1_ASAP7_75t_L g559 ( 
.A1(n_500),
.A2(n_74),
.B(n_76),
.Y(n_559)
);

OAI22xp33_ASAP7_75t_L g560 ( 
.A1(n_508),
.A2(n_77),
.B1(n_78),
.B2(n_79),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_517),
.Y(n_561)
);

BUFx8_ASAP7_75t_L g562 ( 
.A(n_491),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_497),
.Y(n_563)
);

BUFx2_ASAP7_75t_L g564 ( 
.A(n_484),
.Y(n_564)
);

OAI22xp33_ASAP7_75t_L g565 ( 
.A1(n_508),
.A2(n_93),
.B1(n_94),
.B2(n_95),
.Y(n_565)
);

HB1xp67_ASAP7_75t_L g566 ( 
.A(n_498),
.Y(n_566)
);

AOI22xp33_ASAP7_75t_L g567 ( 
.A1(n_499),
.A2(n_97),
.B1(n_98),
.B2(n_100),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_505),
.Y(n_568)
);

AOI22xp33_ASAP7_75t_L g569 ( 
.A1(n_525),
.A2(n_101),
.B1(n_102),
.B2(n_106),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_492),
.B(n_107),
.Y(n_570)
);

HB1xp67_ASAP7_75t_L g571 ( 
.A(n_502),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_497),
.Y(n_572)
);

INVx2_ASAP7_75t_SL g573 ( 
.A(n_494),
.Y(n_573)
);

CKINVDCx11_ASAP7_75t_R g574 ( 
.A(n_491),
.Y(n_574)
);

AOI22xp5_ASAP7_75t_L g575 ( 
.A1(n_507),
.A2(n_109),
.B1(n_110),
.B2(n_111),
.Y(n_575)
);

BUFx3_ASAP7_75t_L g576 ( 
.A(n_540),
.Y(n_576)
);

AOI22xp33_ASAP7_75t_L g577 ( 
.A1(n_554),
.A2(n_525),
.B1(n_526),
.B2(n_492),
.Y(n_577)
);

NOR3xp33_ASAP7_75t_SL g578 ( 
.A(n_535),
.B(n_509),
.C(n_511),
.Y(n_578)
);

INVx2_ASAP7_75t_SL g579 ( 
.A(n_548),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_542),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_542),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_536),
.Y(n_582)
);

OR2x2_ASAP7_75t_L g583 ( 
.A(n_555),
.B(n_531),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_539),
.B(n_555),
.Y(n_584)
);

OR2x2_ASAP7_75t_L g585 ( 
.A(n_564),
.B(n_531),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_543),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_548),
.B(n_528),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_543),
.Y(n_588)
);

BUFx3_ASAP7_75t_L g589 ( 
.A(n_564),
.Y(n_589)
);

NOR3xp33_ASAP7_75t_SL g590 ( 
.A(n_549),
.B(n_487),
.C(n_526),
.Y(n_590)
);

AOI22xp33_ASAP7_75t_L g591 ( 
.A1(n_554),
.A2(n_526),
.B1(n_492),
.B2(n_495),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_539),
.B(n_492),
.Y(n_592)
);

CKINVDCx16_ASAP7_75t_R g593 ( 
.A(n_541),
.Y(n_593)
);

CKINVDCx16_ASAP7_75t_R g594 ( 
.A(n_541),
.Y(n_594)
);

NOR2x1_ASAP7_75t_L g595 ( 
.A(n_551),
.B(n_523),
.Y(n_595)
);

AOI22xp33_ASAP7_75t_L g596 ( 
.A1(n_544),
.A2(n_495),
.B1(n_523),
.B2(n_532),
.Y(n_596)
);

INVxp67_ASAP7_75t_L g597 ( 
.A(n_566),
.Y(n_597)
);

HB1xp67_ASAP7_75t_L g598 ( 
.A(n_571),
.Y(n_598)
);

NAND2xp33_ASAP7_75t_R g599 ( 
.A(n_570),
.B(n_519),
.Y(n_599)
);

NOR3xp33_ASAP7_75t_SL g600 ( 
.A(n_560),
.B(n_516),
.C(n_514),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_550),
.B(n_495),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_546),
.Y(n_602)
);

AND2x4_ASAP7_75t_L g603 ( 
.A(n_573),
.B(n_496),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_574),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_550),
.B(n_494),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_562),
.Y(n_606)
);

AND2x2_ASAP7_75t_SL g607 ( 
.A(n_569),
.B(n_495),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_570),
.B(n_496),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_546),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_533),
.Y(n_610)
);

OAI22xp5_ASAP7_75t_L g611 ( 
.A1(n_545),
.A2(n_489),
.B1(n_519),
.B2(n_522),
.Y(n_611)
);

INVx2_ASAP7_75t_SL g612 ( 
.A(n_573),
.Y(n_612)
);

OR2x6_ASAP7_75t_L g613 ( 
.A(n_534),
.B(n_514),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_547),
.B(n_515),
.Y(n_614)
);

CKINVDCx16_ASAP7_75t_R g615 ( 
.A(n_575),
.Y(n_615)
);

OAI222xp33_ASAP7_75t_L g616 ( 
.A1(n_556),
.A2(n_524),
.B1(n_519),
.B2(n_515),
.C1(n_527),
.C2(n_530),
.Y(n_616)
);

NOR3xp33_ASAP7_75t_SL g617 ( 
.A(n_565),
.B(n_489),
.C(n_521),
.Y(n_617)
);

INVx2_ASAP7_75t_SL g618 ( 
.A(n_562),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_547),
.B(n_521),
.Y(n_619)
);

NAND2xp33_ASAP7_75t_L g620 ( 
.A(n_534),
.B(n_489),
.Y(n_620)
);

CKINVDCx16_ASAP7_75t_R g621 ( 
.A(n_562),
.Y(n_621)
);

AND2x4_ASAP7_75t_L g622 ( 
.A(n_533),
.B(n_530),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_538),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_538),
.Y(n_624)
);

NAND2xp33_ASAP7_75t_SL g625 ( 
.A(n_567),
.B(n_527),
.Y(n_625)
);

AND2x4_ASAP7_75t_L g626 ( 
.A(n_561),
.B(n_112),
.Y(n_626)
);

AOI22xp33_ASAP7_75t_L g627 ( 
.A1(n_558),
.A2(n_568),
.B1(n_534),
.B2(n_545),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_614),
.Y(n_628)
);

BUFx2_ASAP7_75t_SL g629 ( 
.A(n_579),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_602),
.Y(n_630)
);

OR2x2_ASAP7_75t_L g631 ( 
.A(n_614),
.B(n_568),
.Y(n_631)
);

OR2x2_ASAP7_75t_L g632 ( 
.A(n_584),
.B(n_572),
.Y(n_632)
);

BUFx2_ASAP7_75t_L g633 ( 
.A(n_613),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_592),
.B(n_561),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_580),
.B(n_557),
.Y(n_635)
);

OR2x2_ASAP7_75t_L g636 ( 
.A(n_619),
.B(n_572),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_609),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_582),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_581),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_610),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_623),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_624),
.Y(n_642)
);

OAI21x1_ASAP7_75t_L g643 ( 
.A1(n_619),
.A2(n_559),
.B(n_537),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_622),
.Y(n_644)
);

OR2x2_ASAP7_75t_L g645 ( 
.A(n_613),
.B(n_563),
.Y(n_645)
);

AND2x4_ASAP7_75t_L g646 ( 
.A(n_601),
.B(n_557),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_595),
.Y(n_647)
);

INVx4_ASAP7_75t_L g648 ( 
.A(n_603),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_598),
.B(n_553),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_583),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_622),
.Y(n_651)
);

BUFx2_ASAP7_75t_L g652 ( 
.A(n_613),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_585),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_597),
.B(n_608),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_627),
.B(n_553),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_626),
.B(n_589),
.Y(n_656)
);

AND2x4_ASAP7_75t_L g657 ( 
.A(n_626),
.B(n_552),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_612),
.Y(n_658)
);

BUFx3_ASAP7_75t_L g659 ( 
.A(n_576),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_620),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_577),
.B(n_563),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_600),
.B(n_552),
.Y(n_662)
);

AOI21x1_ASAP7_75t_L g663 ( 
.A1(n_611),
.A2(n_559),
.B(n_537),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_611),
.Y(n_664)
);

OR2x2_ASAP7_75t_L g665 ( 
.A(n_597),
.B(n_143),
.Y(n_665)
);

INVxp67_ASAP7_75t_L g666 ( 
.A(n_605),
.Y(n_666)
);

NAND2x1_ASAP7_75t_L g667 ( 
.A(n_617),
.B(n_113),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_628),
.B(n_600),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_637),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_628),
.B(n_607),
.Y(n_670)
);

AOI22xp33_ASAP7_75t_L g671 ( 
.A1(n_660),
.A2(n_615),
.B1(n_625),
.B2(n_596),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_650),
.B(n_587),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_653),
.B(n_590),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_630),
.Y(n_674)
);

AND2x4_ASAP7_75t_L g675 ( 
.A(n_633),
.B(n_603),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_649),
.B(n_591),
.Y(n_676)
);

NOR2x1_ASAP7_75t_L g677 ( 
.A(n_629),
.B(n_616),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_661),
.B(n_618),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_661),
.B(n_578),
.Y(n_679)
);

OR2x2_ASAP7_75t_L g680 ( 
.A(n_636),
.B(n_593),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_630),
.Y(n_681)
);

OR2x2_ASAP7_75t_L g682 ( 
.A(n_636),
.B(n_594),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_639),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_644),
.B(n_578),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_639),
.Y(n_685)
);

OR2x2_ASAP7_75t_L g686 ( 
.A(n_631),
.B(n_621),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_638),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_640),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_632),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_644),
.B(n_118),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_651),
.B(n_119),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_651),
.B(n_120),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_666),
.B(n_604),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_632),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_640),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_680),
.B(n_633),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_680),
.B(n_652),
.Y(n_697)
);

INVxp67_ASAP7_75t_L g698 ( 
.A(n_686),
.Y(n_698)
);

AND2x4_ASAP7_75t_L g699 ( 
.A(n_675),
.B(n_652),
.Y(n_699)
);

OR2x6_ASAP7_75t_L g700 ( 
.A(n_677),
.B(n_667),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_668),
.B(n_631),
.Y(n_701)
);

AND2x2_ASAP7_75t_L g702 ( 
.A(n_682),
.B(n_662),
.Y(n_702)
);

NOR3xp33_ASAP7_75t_SL g703 ( 
.A(n_673),
.B(n_586),
.C(n_588),
.Y(n_703)
);

OR2x2_ASAP7_75t_L g704 ( 
.A(n_682),
.B(n_645),
.Y(n_704)
);

AOI22xp5_ASAP7_75t_L g705 ( 
.A1(n_671),
.A2(n_599),
.B1(n_667),
.B2(n_656),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_674),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_678),
.B(n_662),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_687),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_674),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_686),
.B(n_654),
.Y(n_710)
);

OR2x2_ASAP7_75t_L g711 ( 
.A(n_689),
.B(n_645),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_683),
.Y(n_712)
);

OAI31xp33_ASAP7_75t_L g713 ( 
.A1(n_698),
.A2(n_679),
.A3(n_668),
.B(n_684),
.Y(n_713)
);

INVxp67_ASAP7_75t_L g714 ( 
.A(n_701),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_712),
.Y(n_715)
);

INVxp67_ASAP7_75t_SL g716 ( 
.A(n_701),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_706),
.Y(n_717)
);

AOI22xp5_ASAP7_75t_L g718 ( 
.A1(n_705),
.A2(n_679),
.B1(n_684),
.B2(n_678),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_704),
.Y(n_719)
);

OAI22xp33_ASAP7_75t_L g720 ( 
.A1(n_700),
.A2(n_676),
.B1(n_648),
.B2(n_664),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_708),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_709),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_717),
.Y(n_723)
);

XOR2x2_ASAP7_75t_L g724 ( 
.A(n_718),
.B(n_693),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_722),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_721),
.Y(n_726)
);

AOI21xp5_ASAP7_75t_L g727 ( 
.A1(n_720),
.A2(n_700),
.B(n_616),
.Y(n_727)
);

OR2x2_ASAP7_75t_L g728 ( 
.A(n_726),
.B(n_714),
.Y(n_728)
);

O2A1O1Ixp33_ASAP7_75t_L g729 ( 
.A1(n_727),
.A2(n_713),
.B(n_700),
.C(n_698),
.Y(n_729)
);

AOI21xp33_ASAP7_75t_SL g730 ( 
.A1(n_724),
.A2(n_606),
.B(n_710),
.Y(n_730)
);

INVx2_ASAP7_75t_SL g731 ( 
.A(n_723),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_725),
.B(n_714),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_730),
.B(n_659),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_732),
.Y(n_734)
);

AOI221xp5_ASAP7_75t_L g735 ( 
.A1(n_729),
.A2(n_727),
.B1(n_716),
.B2(n_710),
.C(n_702),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_728),
.B(n_659),
.Y(n_736)
);

XNOR2xp5_ASAP7_75t_L g737 ( 
.A(n_735),
.B(n_703),
.Y(n_737)
);

NOR2xp67_ASAP7_75t_L g738 ( 
.A(n_733),
.B(n_731),
.Y(n_738)
);

AOI22xp5_ASAP7_75t_L g739 ( 
.A1(n_737),
.A2(n_738),
.B1(n_734),
.B2(n_736),
.Y(n_739)
);

AOI22xp33_ASAP7_75t_L g740 ( 
.A1(n_737),
.A2(n_716),
.B1(n_697),
.B2(n_696),
.Y(n_740)
);

AOI222xp33_ASAP7_75t_L g741 ( 
.A1(n_737),
.A2(n_672),
.B1(n_658),
.B2(n_707),
.C1(n_670),
.C2(n_719),
.Y(n_741)
);

AOI22x1_ASAP7_75t_L g742 ( 
.A1(n_741),
.A2(n_629),
.B1(n_665),
.B2(n_703),
.Y(n_742)
);

AND2x4_ASAP7_75t_L g743 ( 
.A(n_739),
.B(n_699),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_740),
.Y(n_744)
);

OAI211xp5_ASAP7_75t_L g745 ( 
.A1(n_739),
.A2(n_665),
.B(n_692),
.C(n_691),
.Y(n_745)
);

NOR2x1_ASAP7_75t_L g746 ( 
.A(n_739),
.B(n_690),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_739),
.Y(n_747)
);

NOR2x1p5_ASAP7_75t_L g748 ( 
.A(n_747),
.B(n_648),
.Y(n_748)
);

NOR3xp33_ASAP7_75t_L g749 ( 
.A(n_744),
.B(n_690),
.C(n_691),
.Y(n_749)
);

OAI221xp5_ASAP7_75t_SL g750 ( 
.A1(n_745),
.A2(n_656),
.B1(n_670),
.B2(n_711),
.C(n_692),
.Y(n_750)
);

AOI22xp5_ASAP7_75t_L g751 ( 
.A1(n_743),
.A2(n_699),
.B1(n_675),
.B2(n_647),
.Y(n_751)
);

NOR3xp33_ASAP7_75t_L g752 ( 
.A(n_746),
.B(n_648),
.C(n_669),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_742),
.Y(n_753)
);

OAI211xp5_ASAP7_75t_L g754 ( 
.A1(n_747),
.A2(n_715),
.B(n_694),
.C(n_663),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_753),
.Y(n_755)
);

HB1xp67_ASAP7_75t_L g756 ( 
.A(n_748),
.Y(n_756)
);

BUFx4f_ASAP7_75t_SL g757 ( 
.A(n_749),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_752),
.Y(n_758)
);

OAI21xp5_ASAP7_75t_L g759 ( 
.A1(n_751),
.A2(n_642),
.B(n_655),
.Y(n_759)
);

INVx2_ASAP7_75t_SL g760 ( 
.A(n_750),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_R g761 ( 
.A(n_755),
.B(n_123),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_755),
.B(n_754),
.Y(n_762)
);

XNOR2x1_ASAP7_75t_L g763 ( 
.A(n_756),
.B(n_124),
.Y(n_763)
);

INVx3_ASAP7_75t_L g764 ( 
.A(n_757),
.Y(n_764)
);

OAI22xp5_ASAP7_75t_L g765 ( 
.A1(n_760),
.A2(n_758),
.B1(n_759),
.B2(n_675),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_755),
.Y(n_766)
);

XNOR2xp5_ASAP7_75t_L g767 ( 
.A(n_755),
.B(n_646),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_757),
.Y(n_768)
);

BUFx2_ASAP7_75t_L g769 ( 
.A(n_761),
.Y(n_769)
);

AND2x4_ASAP7_75t_L g770 ( 
.A(n_766),
.B(n_681),
.Y(n_770)
);

AOI22xp5_ASAP7_75t_L g771 ( 
.A1(n_768),
.A2(n_646),
.B1(n_655),
.B2(n_634),
.Y(n_771)
);

HB1xp67_ASAP7_75t_L g772 ( 
.A(n_763),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_764),
.Y(n_773)
);

AOI22xp5_ASAP7_75t_L g774 ( 
.A1(n_765),
.A2(n_646),
.B1(n_634),
.B2(n_664),
.Y(n_774)
);

AOI31xp33_ASAP7_75t_L g775 ( 
.A1(n_762),
.A2(n_635),
.A3(n_688),
.B(n_685),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_767),
.B(n_688),
.Y(n_776)
);

OAI22x1_ASAP7_75t_SL g777 ( 
.A1(n_773),
.A2(n_126),
.B1(n_127),
.B2(n_131),
.Y(n_777)
);

XOR2xp5_ASAP7_75t_L g778 ( 
.A(n_772),
.B(n_769),
.Y(n_778)
);

AOI22xp5_ASAP7_75t_L g779 ( 
.A1(n_774),
.A2(n_685),
.B1(n_683),
.B2(n_695),
.Y(n_779)
);

CKINVDCx20_ASAP7_75t_R g780 ( 
.A(n_771),
.Y(n_780)
);

INVxp67_ASAP7_75t_L g781 ( 
.A(n_770),
.Y(n_781)
);

AOI22xp5_ASAP7_75t_L g782 ( 
.A1(n_780),
.A2(n_776),
.B1(n_775),
.B2(n_695),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_778),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_783),
.B(n_781),
.Y(n_784)
);

AOI222xp33_ASAP7_75t_L g785 ( 
.A1(n_784),
.A2(n_777),
.B1(n_782),
.B2(n_779),
.C1(n_641),
.C2(n_635),
.Y(n_785)
);

OR2x6_ASAP7_75t_L g786 ( 
.A(n_785),
.B(n_132),
.Y(n_786)
);

AOI22xp33_ASAP7_75t_L g787 ( 
.A1(n_786),
.A2(n_641),
.B1(n_657),
.B2(n_643),
.Y(n_787)
);


endmodule