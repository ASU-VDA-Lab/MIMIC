module fake_jpeg_25146_n_201 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_201);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_201;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx6f_ASAP7_75t_SL g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_14),
.B(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_43),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_18),
.B(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_41),
.B(n_22),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_7),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_41),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_48),
.B(n_49),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_38),
.B(n_33),
.Y(n_49)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_31),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_58),
.Y(n_63)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_33),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_61),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_35),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_37),
.B(n_21),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_62),
.B(n_19),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_48),
.A2(n_24),
.B1(n_30),
.B2(n_21),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_64),
.B(n_25),
.Y(n_103)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_62),
.Y(n_65)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

NAND3xp33_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_9),
.C(n_15),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_66),
.B(n_29),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_44),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_67),
.B(n_75),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_69),
.B(n_73),
.Y(n_109)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_72),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_19),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_53),
.B(n_22),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_61),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_77),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_78),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_27),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_81),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_51),
.B(n_27),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_82),
.B(n_84),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_45),
.B(n_18),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_85),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_51),
.B(n_29),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_45),
.B(n_26),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_52),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_86),
.B(n_39),
.Y(n_93)
);

AO22x2_ASAP7_75t_L g87 ( 
.A1(n_67),
.A2(n_57),
.B1(n_35),
.B2(n_34),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_87),
.A2(n_72),
.B1(n_86),
.B2(n_71),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_91),
.B(n_100),
.Y(n_110)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_93),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_65),
.A2(n_57),
.B1(n_40),
.B2(n_47),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_95),
.A2(n_99),
.B1(n_79),
.B2(n_78),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_39),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_101),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_85),
.A2(n_30),
.B1(n_42),
.B2(n_52),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_68),
.B(n_32),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_77),
.B(n_39),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_59),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_81),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_103),
.A2(n_104),
.B(n_64),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_70),
.A2(n_0),
.B(n_2),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_74),
.B(n_32),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_108),
.B(n_17),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_98),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_111),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_112),
.A2(n_119),
.B1(n_120),
.B2(n_128),
.Y(n_148)
);

NOR2x1_ASAP7_75t_L g113 ( 
.A(n_103),
.B(n_63),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_113),
.B(n_125),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_114),
.B(n_118),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_115),
.A2(n_129),
.B1(n_119),
.B2(n_104),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_103),
.A2(n_78),
.B(n_71),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_117),
.A2(n_106),
.B(n_105),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_17),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_89),
.A2(n_34),
.B1(n_79),
.B2(n_76),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_101),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_122),
.B(n_123),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_88),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_124),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_109),
.B(n_23),
.Y(n_125)
);

A2O1A1O1Ixp25_ASAP7_75t_L g126 ( 
.A1(n_87),
.A2(n_90),
.B(n_89),
.C(n_97),
.D(n_102),
.Y(n_126)
);

XOR2x1_ASAP7_75t_L g138 ( 
.A(n_126),
.B(n_94),
.Y(n_138)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_107),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_127),
.B(n_107),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_87),
.A2(n_76),
.B1(n_23),
.B2(n_25),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_87),
.A2(n_23),
.B1(n_16),
.B2(n_5),
.Y(n_129)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_123),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_132),
.B(n_139),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_127),
.A2(n_87),
.B1(n_94),
.B2(n_106),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_133),
.A2(n_137),
.B1(n_129),
.B2(n_128),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_115),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_135),
.B(n_147),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_90),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_138),
.Y(n_159)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_120),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_116),
.B(n_108),
.C(n_96),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_140),
.B(n_142),
.C(n_3),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_122),
.B(n_111),
.Y(n_141)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_141),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_112),
.B(n_96),
.Y(n_142)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_144),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_145),
.A2(n_117),
.B(n_105),
.Y(n_149)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_126),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_149),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_150),
.A2(n_152),
.B1(n_154),
.B2(n_146),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_139),
.A2(n_121),
.B1(n_113),
.B2(n_91),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_141),
.A2(n_121),
.B(n_110),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_153),
.B(n_131),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_132),
.A2(n_16),
.B1(n_10),
.B2(n_11),
.Y(n_154)
);

NAND3xp33_ASAP7_75t_L g155 ( 
.A(n_138),
.B(n_12),
.C(n_14),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_155),
.B(n_161),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_156),
.B(n_163),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_147),
.B(n_3),
.C(n_4),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_158),
.B(n_140),
.C(n_142),
.Y(n_167)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_130),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_145),
.A2(n_3),
.B(n_4),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_164),
.B(n_174),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_157),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_165),
.B(n_166),
.Y(n_178)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_157),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_167),
.B(n_171),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_168),
.B(n_137),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_159),
.B(n_130),
.C(n_136),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_159),
.B(n_143),
.C(n_148),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_173),
.B(n_156),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_152),
.B(n_134),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_169),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_175),
.B(n_176),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_170),
.Y(n_176)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_177),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_179),
.B(n_182),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_173),
.B(n_154),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_180),
.B(n_171),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_183),
.B(n_184),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_175),
.B(n_167),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_178),
.A2(n_151),
.B1(n_172),
.B2(n_149),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_185),
.A2(n_160),
.B(n_153),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_177),
.A2(n_162),
.B(n_163),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_188),
.A2(n_169),
.B(n_5),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_190),
.A2(n_191),
.B(n_185),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_186),
.A2(n_181),
.B(n_160),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_187),
.B(n_158),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_192),
.B(n_189),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_193),
.A2(n_5),
.B(n_6),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_195),
.B(n_196),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_197),
.B(n_184),
.C(n_194),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_198),
.B(n_6),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_200),
.B(n_199),
.Y(n_201)
);


endmodule