module fake_netlist_6_4281_n_935 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_235, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_223, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_226, n_228, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_227, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_233, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_234, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_236, n_38, n_110, n_151, n_61, n_112, n_172, n_237, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_238, n_239, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_231, n_65, n_230, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_229, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_232, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_935);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_235;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_223;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_226;
input n_228;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_227;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_233;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_234;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_236;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_237;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_238;
input n_239;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_231;
input n_65;
input n_230;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_229;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_232;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_935;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_909;
wire n_580;
wire n_762;
wire n_881;
wire n_875;
wire n_465;
wire n_367;
wire n_760;
wire n_680;
wire n_741;
wire n_590;
wire n_625;
wire n_661;
wire n_278;
wire n_341;
wire n_362;
wire n_828;
wire n_462;
wire n_607;
wire n_726;
wire n_671;
wire n_316;
wire n_419;
wire n_304;
wire n_700;
wire n_694;
wire n_933;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_783;
wire n_725;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_628;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_698;
wire n_617;
wire n_898;
wire n_845;
wire n_255;
wire n_807;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_865;
wire n_893;
wire n_925;
wire n_485;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_573;
wire n_769;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_669;
wire n_447;
wire n_872;
wire n_248;
wire n_300;
wire n_517;
wire n_718;
wire n_747;
wire n_852;
wire n_667;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_901;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_822;
wire n_693;
wire n_758;
wire n_516;
wire n_720;
wire n_525;
wire n_631;
wire n_842;
wire n_611;
wire n_491;
wire n_878;
wire n_772;
wire n_656;
wire n_843;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_844;
wire n_343;
wire n_448;
wire n_886;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_454;
wire n_638;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_653;
wire n_887;
wire n_752;
wire n_908;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_803;
wire n_290;
wire n_809;
wire n_926;
wire n_927;
wire n_839;
wire n_734;
wire n_708;
wire n_919;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_800;
wire n_929;
wire n_460;
wire n_907;
wire n_854;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_650;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_594;
wire n_719;
wire n_565;
wire n_356;
wire n_577;
wire n_552;
wire n_619;
wire n_885;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_792;
wire n_880;
wire n_476;
wire n_714;
wire n_291;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_821;
wire n_325;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_523;
wire n_707;
wire n_322;
wire n_409;
wire n_345;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_787;
wire n_635;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_386;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_811;
wire n_882;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_299;
wire n_518;
wire n_679;
wire n_612;
wire n_453;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_247;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_257;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_286;
wire n_254;
wire n_834;
wire n_242;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_816;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_604;
wire n_848;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_385;
wire n_295;
wire n_701;
wire n_817;
wire n_629;
wire n_388;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_841;
wire n_531;
wire n_827;
wire n_508;
wire n_361;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_664;
wire n_678;
wire n_649;
wire n_283;

INVx1_ASAP7_75t_L g240 ( 
.A(n_228),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_115),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_105),
.Y(n_242)
);

BUFx10_ASAP7_75t_L g243 ( 
.A(n_76),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_95),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_17),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_141),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_102),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_203),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_123),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_109),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_100),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_171),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_164),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_218),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_25),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_79),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_7),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_219),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_129),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_88),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_126),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_157),
.Y(n_262)
);

CKINVDCx14_ASAP7_75t_R g263 ( 
.A(n_39),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_98),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_227),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_94),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_226),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_3),
.Y(n_268)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_208),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_222),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_7),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_49),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_212),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_131),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_207),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_195),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_31),
.Y(n_277)
);

BUFx2_ASAP7_75t_L g278 ( 
.A(n_18),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_35),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g280 ( 
.A(n_165),
.Y(n_280)
);

INVx2_ASAP7_75t_SL g281 ( 
.A(n_23),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_121),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_91),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_185),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_119),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_1),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_239),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_132),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_138),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_38),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_44),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_0),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_130),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_28),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_235),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_12),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_213),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_26),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_179),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_186),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_83),
.Y(n_301)
);

BUFx10_ASAP7_75t_L g302 ( 
.A(n_182),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_232),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_127),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_99),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_190),
.Y(n_306)
);

BUFx10_ASAP7_75t_L g307 ( 
.A(n_2),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_163),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_199),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_238),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_236),
.Y(n_311)
);

BUFx10_ASAP7_75t_L g312 ( 
.A(n_234),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_172),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_30),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_194),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_225),
.Y(n_316)
);

INVxp67_ASAP7_75t_SL g317 ( 
.A(n_191),
.Y(n_317)
);

BUFx3_ASAP7_75t_L g318 ( 
.A(n_54),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_224),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_167),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_70),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_215),
.Y(n_322)
);

BUFx2_ASAP7_75t_SL g323 ( 
.A(n_41),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_77),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_118),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_142),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_159),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_3),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_47),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_71),
.Y(n_330)
);

BUFx3_ASAP7_75t_L g331 ( 
.A(n_9),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_30),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_104),
.Y(n_333)
);

INVx2_ASAP7_75t_SL g334 ( 
.A(n_61),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_220),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_168),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_181),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_66),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_89),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_198),
.Y(n_340)
);

BUFx2_ASAP7_75t_SL g341 ( 
.A(n_52),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_122),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_107),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_128),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_97),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_92),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_184),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_192),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_86),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_16),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_188),
.Y(n_351)
);

BUFx5_ASAP7_75t_L g352 ( 
.A(n_158),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_174),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_149),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_152),
.Y(n_355)
);

BUFx3_ASAP7_75t_L g356 ( 
.A(n_180),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_139),
.Y(n_357)
);

INVx1_ASAP7_75t_SL g358 ( 
.A(n_231),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_90),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_93),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_144),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_153),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_117),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_205),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_229),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_230),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_73),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_58),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_106),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_223),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_25),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_56),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_151),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_210),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_84),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_18),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_50),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_196),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_8),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_96),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_237),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_43),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_176),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_75),
.Y(n_384)
);

CKINVDCx14_ASAP7_75t_R g385 ( 
.A(n_161),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_233),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_169),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_40),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_21),
.Y(n_389)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_148),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_11),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_202),
.Y(n_392)
);

INVx1_ASAP7_75t_SL g393 ( 
.A(n_24),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_124),
.Y(n_394)
);

BUFx3_ASAP7_75t_L g395 ( 
.A(n_19),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_67),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_57),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_120),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_217),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_204),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_278),
.B(n_1),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_273),
.B(n_2),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_267),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_296),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_296),
.B(n_4),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_296),
.B(n_4),
.Y(n_406)
);

BUFx2_ASAP7_75t_L g407 ( 
.A(n_331),
.Y(n_407)
);

HB1xp67_ASAP7_75t_L g408 ( 
.A(n_245),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_296),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_390),
.B(n_5),
.Y(n_410)
);

BUFx12f_ASAP7_75t_L g411 ( 
.A(n_307),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_352),
.Y(n_412)
);

AND2x4_ASAP7_75t_L g413 ( 
.A(n_318),
.B(n_6),
.Y(n_413)
);

INVx3_ASAP7_75t_L g414 ( 
.A(n_395),
.Y(n_414)
);

INVx5_ASAP7_75t_L g415 ( 
.A(n_267),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_267),
.Y(n_416)
);

BUFx3_ASAP7_75t_L g417 ( 
.A(n_243),
.Y(n_417)
);

INVx5_ASAP7_75t_L g418 ( 
.A(n_267),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_329),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_390),
.B(n_6),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_257),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_263),
.B(n_8),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_268),
.Y(n_423)
);

INVx5_ASAP7_75t_L g424 ( 
.A(n_329),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_352),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_263),
.B(n_10),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_317),
.B(n_10),
.Y(n_427)
);

BUFx3_ASAP7_75t_L g428 ( 
.A(n_302),
.Y(n_428)
);

INVx3_ASAP7_75t_L g429 ( 
.A(n_255),
.Y(n_429)
);

AND2x6_ASAP7_75t_L g430 ( 
.A(n_329),
.B(n_32),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g431 ( 
.A(n_385),
.B(n_11),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_334),
.B(n_12),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_352),
.Y(n_433)
);

BUFx2_ASAP7_75t_L g434 ( 
.A(n_286),
.Y(n_434)
);

INVx2_ASAP7_75t_SL g435 ( 
.A(n_307),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_352),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_385),
.B(n_13),
.Y(n_437)
);

AND2x4_ASAP7_75t_L g438 ( 
.A(n_318),
.B(n_13),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_281),
.B(n_14),
.Y(n_439)
);

XNOR2x1_ASAP7_75t_L g440 ( 
.A(n_292),
.B(n_14),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_256),
.B(n_15),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_246),
.B(n_15),
.Y(n_442)
);

BUFx12f_ASAP7_75t_L g443 ( 
.A(n_302),
.Y(n_443)
);

BUFx8_ASAP7_75t_SL g444 ( 
.A(n_391),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_269),
.B(n_16),
.Y(n_445)
);

BUFx3_ASAP7_75t_L g446 ( 
.A(n_312),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_249),
.B(n_17),
.Y(n_447)
);

INVx5_ASAP7_75t_L g448 ( 
.A(n_329),
.Y(n_448)
);

AND2x4_ASAP7_75t_L g449 ( 
.A(n_280),
.B(n_19),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_253),
.B(n_356),
.Y(n_450)
);

BUFx3_ASAP7_75t_L g451 ( 
.A(n_312),
.Y(n_451)
);

INVx5_ASAP7_75t_L g452 ( 
.A(n_352),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_240),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_358),
.B(n_20),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_271),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_241),
.Y(n_456)
);

BUFx3_ASAP7_75t_L g457 ( 
.A(n_242),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_277),
.Y(n_458)
);

AND2x4_ASAP7_75t_L g459 ( 
.A(n_244),
.B(n_248),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_332),
.B(n_20),
.Y(n_460)
);

HB1xp67_ASAP7_75t_L g461 ( 
.A(n_294),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_298),
.B(n_21),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_276),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_393),
.B(n_22),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_252),
.Y(n_465)
);

AND2x4_ASAP7_75t_L g466 ( 
.A(n_259),
.B(n_24),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_260),
.B(n_27),
.Y(n_467)
);

BUFx12f_ASAP7_75t_L g468 ( 
.A(n_376),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_314),
.Y(n_469)
);

AND2x4_ASAP7_75t_L g470 ( 
.A(n_261),
.B(n_27),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_SL g471 ( 
.A(n_379),
.B(n_328),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_350),
.B(n_28),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_371),
.Y(n_473)
);

INVx5_ASAP7_75t_L g474 ( 
.A(n_323),
.Y(n_474)
);

BUFx6f_ASAP7_75t_L g475 ( 
.A(n_262),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_389),
.B(n_29),
.Y(n_476)
);

AND2x4_ASAP7_75t_L g477 ( 
.A(n_264),
.B(n_265),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_295),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_303),
.B(n_31),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_304),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_310),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_313),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_316),
.B(n_319),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_321),
.B(n_33),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g485 ( 
.A(n_325),
.B(n_34),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_333),
.B(n_36),
.Y(n_486)
);

BUFx12f_ASAP7_75t_L g487 ( 
.A(n_247),
.Y(n_487)
);

INVx2_ASAP7_75t_SL g488 ( 
.A(n_250),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_336),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_434),
.B(n_251),
.Y(n_490)
);

OAI22xp33_ASAP7_75t_L g491 ( 
.A1(n_471),
.A2(n_284),
.B1(n_287),
.B2(n_279),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_471),
.A2(n_426),
.B1(n_431),
.B2(n_422),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_404),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_409),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_403),
.Y(n_495)
);

AND2x2_ASAP7_75t_SL g496 ( 
.A(n_437),
.B(n_464),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_407),
.B(n_254),
.Y(n_497)
);

AO22x2_ASAP7_75t_L g498 ( 
.A1(n_402),
.A2(n_341),
.B1(n_347),
.B2(n_339),
.Y(n_498)
);

OAI22xp33_ASAP7_75t_SL g499 ( 
.A1(n_402),
.A2(n_360),
.B1(n_363),
.B2(n_348),
.Y(n_499)
);

OA22x2_ASAP7_75t_L g500 ( 
.A1(n_480),
.A2(n_372),
.B1(n_380),
.B2(n_368),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_454),
.A2(n_326),
.B1(n_338),
.B2(n_306),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_403),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g503 ( 
.A(n_457),
.B(n_258),
.Y(n_503)
);

INVx2_ASAP7_75t_SL g504 ( 
.A(n_417),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_454),
.A2(n_361),
.B1(n_369),
.B2(n_344),
.Y(n_505)
);

AO22x2_ASAP7_75t_L g506 ( 
.A1(n_460),
.A2(n_392),
.B1(n_383),
.B2(n_386),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_488),
.B(n_266),
.Y(n_507)
);

AO22x2_ASAP7_75t_L g508 ( 
.A1(n_460),
.A2(n_394),
.B1(n_387),
.B2(n_388),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_428),
.B(n_270),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_401),
.A2(n_370),
.B1(n_399),
.B2(n_374),
.Y(n_510)
);

BUFx10_ASAP7_75t_L g511 ( 
.A(n_456),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_489),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_403),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_482),
.Y(n_514)
);

OAI22xp33_ASAP7_75t_SL g515 ( 
.A1(n_450),
.A2(n_381),
.B1(n_382),
.B2(n_384),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_427),
.A2(n_400),
.B1(n_398),
.B2(n_397),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_446),
.B(n_272),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_421),
.Y(n_518)
);

OAI22xp33_ASAP7_75t_L g519 ( 
.A1(n_410),
.A2(n_396),
.B1(n_378),
.B2(n_377),
.Y(n_519)
);

OR2x6_ASAP7_75t_L g520 ( 
.A(n_468),
.B(n_274),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_463),
.B(n_275),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_423),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_435),
.A2(n_322),
.B1(n_373),
.B2(n_367),
.Y(n_523)
);

OA22x2_ASAP7_75t_L g524 ( 
.A1(n_480),
.A2(n_375),
.B1(n_366),
.B2(n_365),
.Y(n_524)
);

OR2x2_ASAP7_75t_L g525 ( 
.A(n_414),
.B(n_282),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_L g526 ( 
.A1(n_410),
.A2(n_364),
.B1(n_362),
.B2(n_359),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_469),
.Y(n_527)
);

OAI22xp33_ASAP7_75t_L g528 ( 
.A1(n_420),
.A2(n_357),
.B1(n_355),
.B2(n_354),
.Y(n_528)
);

OAI22xp33_ASAP7_75t_L g529 ( 
.A1(n_420),
.A2(n_353),
.B1(n_351),
.B2(n_349),
.Y(n_529)
);

OAI22xp33_ASAP7_75t_L g530 ( 
.A1(n_447),
.A2(n_346),
.B1(n_345),
.B2(n_343),
.Y(n_530)
);

OR2x6_ASAP7_75t_L g531 ( 
.A(n_411),
.B(n_283),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_442),
.A2(n_342),
.B1(n_340),
.B2(n_337),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_450),
.B(n_285),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g534 ( 
.A(n_451),
.B(n_288),
.Y(n_534)
);

OAI22xp33_ASAP7_75t_L g535 ( 
.A1(n_447),
.A2(n_335),
.B1(n_330),
.B2(n_327),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_414),
.B(n_289),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_445),
.B(n_290),
.Y(n_537)
);

AOI22xp5_ASAP7_75t_L g538 ( 
.A1(n_443),
.A2(n_324),
.B1(n_320),
.B2(n_315),
.Y(n_538)
);

OAI22xp33_ASAP7_75t_SL g539 ( 
.A1(n_432),
.A2(n_311),
.B1(n_309),
.B2(n_308),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_473),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_432),
.B(n_291),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_459),
.B(n_293),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_416),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_416),
.Y(n_544)
);

OAI22xp5_ASAP7_75t_L g545 ( 
.A1(n_479),
.A2(n_305),
.B1(n_301),
.B2(n_300),
.Y(n_545)
);

AO22x2_ASAP7_75t_L g546 ( 
.A1(n_413),
.A2(n_299),
.B1(n_297),
.B2(n_45),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_487),
.Y(n_547)
);

AOI22xp5_ASAP7_75t_L g548 ( 
.A1(n_485),
.A2(n_37),
.B1(n_42),
.B2(n_46),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_477),
.B(n_48),
.Y(n_549)
);

INVx2_ASAP7_75t_SL g550 ( 
.A(n_408),
.Y(n_550)
);

AOI22xp5_ASAP7_75t_L g551 ( 
.A1(n_449),
.A2(n_51),
.B1(n_53),
.B2(n_55),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_419),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_419),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_518),
.Y(n_554)
);

BUFx2_ASAP7_75t_L g555 ( 
.A(n_497),
.Y(n_555)
);

NOR2xp67_ASAP7_75t_L g556 ( 
.A(n_541),
.B(n_415),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_550),
.B(n_477),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_495),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_533),
.B(n_474),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_502),
.Y(n_560)
);

CKINVDCx20_ASAP7_75t_R g561 ( 
.A(n_511),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_513),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_522),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_527),
.Y(n_564)
);

XNOR2xp5_ASAP7_75t_SL g565 ( 
.A(n_521),
.B(n_444),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g566 ( 
.A(n_536),
.B(n_408),
.Y(n_566)
);

OAI21xp5_ASAP7_75t_L g567 ( 
.A1(n_492),
.A2(n_483),
.B(n_484),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_540),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_516),
.B(n_474),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_514),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_553),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_553),
.Y(n_572)
);

XOR2x2_ASAP7_75t_L g573 ( 
.A(n_501),
.B(n_440),
.Y(n_573)
);

NOR2xp67_ASAP7_75t_L g574 ( 
.A(n_548),
.B(n_415),
.Y(n_574)
);

AND2x6_ASAP7_75t_L g575 ( 
.A(n_549),
.B(n_438),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_496),
.B(n_461),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_543),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_552),
.Y(n_578)
);

XNOR2x2_ASAP7_75t_L g579 ( 
.A(n_546),
.B(n_439),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_490),
.B(n_461),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_499),
.B(n_449),
.Y(n_581)
);

BUFx6f_ASAP7_75t_SL g582 ( 
.A(n_511),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_544),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_544),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_544),
.Y(n_585)
);

XNOR2xp5_ASAP7_75t_L g586 ( 
.A(n_491),
.B(n_505),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_525),
.B(n_483),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_493),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g589 ( 
.A(n_504),
.B(n_429),
.Y(n_589)
);

OR2x6_ASAP7_75t_L g590 ( 
.A(n_546),
.B(n_439),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_512),
.Y(n_591)
);

AND2x4_ASAP7_75t_L g592 ( 
.A(n_542),
.B(n_438),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_494),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_507),
.B(n_479),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_500),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_534),
.B(n_429),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_537),
.B(n_412),
.Y(n_597)
);

CKINVDCx20_ASAP7_75t_R g598 ( 
.A(n_510),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_503),
.Y(n_599)
);

OR2x2_ASAP7_75t_L g600 ( 
.A(n_532),
.B(n_509),
.Y(n_600)
);

INVxp33_ASAP7_75t_L g601 ( 
.A(n_524),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_551),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_506),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_528),
.B(n_529),
.Y(n_604)
);

OAI21xp5_ASAP7_75t_L g605 ( 
.A1(n_526),
.A2(n_484),
.B(n_466),
.Y(n_605)
);

CKINVDCx20_ASAP7_75t_R g606 ( 
.A(n_547),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_506),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_508),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_523),
.B(n_455),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_545),
.B(n_466),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_508),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_498),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_SL g613 ( 
.A(n_519),
.B(n_430),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_498),
.B(n_425),
.Y(n_614)
);

OR2x2_ASAP7_75t_L g615 ( 
.A(n_517),
.B(n_470),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_515),
.Y(n_616)
);

NAND2xp33_ASAP7_75t_R g617 ( 
.A(n_520),
.B(n_470),
.Y(n_617)
);

XNOR2x2_ASAP7_75t_L g618 ( 
.A(n_538),
.B(n_467),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_539),
.Y(n_619)
);

INVx2_ASAP7_75t_SL g620 ( 
.A(n_520),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_531),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_530),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_535),
.Y(n_623)
);

AND2x2_ASAP7_75t_SL g624 ( 
.A(n_613),
.B(n_486),
.Y(n_624)
);

HB1xp67_ASAP7_75t_L g625 ( 
.A(n_616),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_594),
.B(n_486),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_554),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_587),
.B(n_566),
.Y(n_628)
);

INVx1_ASAP7_75t_SL g629 ( 
.A(n_580),
.Y(n_629)
);

INVxp67_ASAP7_75t_SL g630 ( 
.A(n_563),
.Y(n_630)
);

OAI21x1_ASAP7_75t_L g631 ( 
.A1(n_597),
.A2(n_614),
.B(n_581),
.Y(n_631)
);

INVx3_ASAP7_75t_L g632 ( 
.A(n_558),
.Y(n_632)
);

BUFx3_ASAP7_75t_L g633 ( 
.A(n_564),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_567),
.B(n_458),
.Y(n_634)
);

HB1xp67_ASAP7_75t_L g635 ( 
.A(n_612),
.Y(n_635)
);

INVx2_ASAP7_75t_SL g636 ( 
.A(n_596),
.Y(n_636)
);

INVx2_ASAP7_75t_SL g637 ( 
.A(n_589),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_557),
.B(n_531),
.Y(n_638)
);

AND2x4_ASAP7_75t_L g639 ( 
.A(n_595),
.B(n_462),
.Y(n_639)
);

BUFx2_ASAP7_75t_L g640 ( 
.A(n_576),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_571),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_567),
.B(n_430),
.Y(n_642)
);

BUFx3_ASAP7_75t_L g643 ( 
.A(n_568),
.Y(n_643)
);

INVx4_ASAP7_75t_L g644 ( 
.A(n_575),
.Y(n_644)
);

BUFx3_ASAP7_75t_L g645 ( 
.A(n_570),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_597),
.B(n_430),
.Y(n_646)
);

OAI21xp5_ASAP7_75t_L g647 ( 
.A1(n_605),
.A2(n_441),
.B(n_467),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_572),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_592),
.B(n_405),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_559),
.B(n_453),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_610),
.B(n_465),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_592),
.B(n_405),
.Y(n_652)
);

INVxp67_ASAP7_75t_L g653 ( 
.A(n_555),
.Y(n_653)
);

INVx4_ASAP7_75t_L g654 ( 
.A(n_575),
.Y(n_654)
);

OAI21xp5_ASAP7_75t_L g655 ( 
.A1(n_605),
.A2(n_441),
.B(n_406),
.Y(n_655)
);

OR2x2_ASAP7_75t_L g656 ( 
.A(n_622),
.B(n_462),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_608),
.B(n_406),
.Y(n_657)
);

BUFx4_ASAP7_75t_SL g658 ( 
.A(n_561),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_623),
.B(n_472),
.Y(n_659)
);

INVx3_ASAP7_75t_L g660 ( 
.A(n_560),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_591),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_575),
.B(n_465),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_588),
.Y(n_663)
);

INVx3_ASAP7_75t_L g664 ( 
.A(n_562),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_599),
.B(n_472),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_614),
.B(n_476),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_593),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_603),
.B(n_433),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_601),
.B(n_475),
.Y(n_669)
);

HB1xp67_ASAP7_75t_L g670 ( 
.A(n_607),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_578),
.Y(n_671)
);

BUFx3_ASAP7_75t_L g672 ( 
.A(n_606),
.Y(n_672)
);

BUFx6f_ASAP7_75t_L g673 ( 
.A(n_584),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_611),
.B(n_436),
.Y(n_674)
);

INVx1_ASAP7_75t_SL g675 ( 
.A(n_609),
.Y(n_675)
);

BUFx8_ASAP7_75t_L g676 ( 
.A(n_582),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_577),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_575),
.B(n_475),
.Y(n_678)
);

BUFx6f_ASAP7_75t_L g679 ( 
.A(n_583),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_585),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_615),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_602),
.B(n_478),
.Y(n_682)
);

OAI21xp5_ASAP7_75t_L g683 ( 
.A1(n_604),
.A2(n_424),
.B(n_418),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_619),
.B(n_478),
.Y(n_684)
);

INVx3_ASAP7_75t_L g685 ( 
.A(n_600),
.Y(n_685)
);

OR2x2_ASAP7_75t_SL g686 ( 
.A(n_573),
.B(n_478),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_586),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_641),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_641),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_648),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_628),
.B(n_569),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_675),
.B(n_598),
.Y(n_692)
);

INVx5_ASAP7_75t_L g693 ( 
.A(n_685),
.Y(n_693)
);

INVx3_ASAP7_75t_L g694 ( 
.A(n_673),
.Y(n_694)
);

BUFx6f_ASAP7_75t_L g695 ( 
.A(n_633),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_628),
.B(n_618),
.Y(n_696)
);

NAND2x1_ASAP7_75t_SL g697 ( 
.A(n_638),
.B(n_574),
.Y(n_697)
);

INVx4_ASAP7_75t_L g698 ( 
.A(n_673),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_658),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_672),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_629),
.B(n_665),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_SL g702 ( 
.A(n_624),
.B(n_590),
.Y(n_702)
);

OR2x2_ASAP7_75t_L g703 ( 
.A(n_687),
.B(n_640),
.Y(n_703)
);

BUFx3_ASAP7_75t_L g704 ( 
.A(n_672),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_648),
.Y(n_705)
);

INVx4_ASAP7_75t_L g706 ( 
.A(n_673),
.Y(n_706)
);

AND2x4_ASAP7_75t_L g707 ( 
.A(n_636),
.B(n_621),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_SL g708 ( 
.A(n_624),
.B(n_590),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_627),
.Y(n_709)
);

AND2x2_ASAP7_75t_SL g710 ( 
.A(n_626),
.B(n_613),
.Y(n_710)
);

BUFx6f_ASAP7_75t_L g711 ( 
.A(n_633),
.Y(n_711)
);

BUFx2_ASAP7_75t_L g712 ( 
.A(n_653),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_663),
.Y(n_713)
);

NAND2x1p5_ASAP7_75t_L g714 ( 
.A(n_644),
.B(n_620),
.Y(n_714)
);

BUFx6f_ASAP7_75t_L g715 ( 
.A(n_643),
.Y(n_715)
);

INVx3_ASAP7_75t_L g716 ( 
.A(n_673),
.Y(n_716)
);

HB1xp67_ASAP7_75t_L g717 ( 
.A(n_670),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_685),
.B(n_681),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_666),
.B(n_590),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_663),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_666),
.B(n_556),
.Y(n_721)
);

BUFx2_ASAP7_75t_L g722 ( 
.A(n_685),
.Y(n_722)
);

BUFx2_ASAP7_75t_L g723 ( 
.A(n_686),
.Y(n_723)
);

NOR2xp67_ASAP7_75t_L g724 ( 
.A(n_644),
.B(n_556),
.Y(n_724)
);

BUFx6f_ASAP7_75t_L g725 ( 
.A(n_643),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_SL g726 ( 
.A(n_644),
.B(n_579),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_634),
.B(n_659),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_634),
.B(n_481),
.Y(n_728)
);

INVx3_ASAP7_75t_L g729 ( 
.A(n_679),
.Y(n_729)
);

AND2x4_ASAP7_75t_L g730 ( 
.A(n_645),
.B(n_59),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_688),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_727),
.B(n_659),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_689),
.Y(n_733)
);

BUFx6f_ASAP7_75t_L g734 ( 
.A(n_695),
.Y(n_734)
);

BUFx6f_ASAP7_75t_L g735 ( 
.A(n_695),
.Y(n_735)
);

HB1xp67_ASAP7_75t_L g736 ( 
.A(n_712),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_705),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_690),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_713),
.Y(n_739)
);

BUFx3_ASAP7_75t_L g740 ( 
.A(n_704),
.Y(n_740)
);

INVx3_ASAP7_75t_L g741 ( 
.A(n_698),
.Y(n_741)
);

INVx4_ASAP7_75t_L g742 ( 
.A(n_695),
.Y(n_742)
);

BUFx3_ASAP7_75t_L g743 ( 
.A(n_711),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_720),
.Y(n_744)
);

INVx4_ASAP7_75t_L g745 ( 
.A(n_711),
.Y(n_745)
);

BUFx6f_ASAP7_75t_L g746 ( 
.A(n_711),
.Y(n_746)
);

AND2x4_ASAP7_75t_L g747 ( 
.A(n_730),
.B(n_645),
.Y(n_747)
);

NOR2x1_ASAP7_75t_SL g748 ( 
.A(n_693),
.B(n_654),
.Y(n_748)
);

BUFx3_ASAP7_75t_L g749 ( 
.A(n_715),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_709),
.Y(n_750)
);

INVx3_ASAP7_75t_L g751 ( 
.A(n_698),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_728),
.Y(n_752)
);

INVx2_ASAP7_75t_SL g753 ( 
.A(n_717),
.Y(n_753)
);

NAND2x1p5_ASAP7_75t_L g754 ( 
.A(n_693),
.B(n_654),
.Y(n_754)
);

INVx5_ASAP7_75t_L g755 ( 
.A(n_729),
.Y(n_755)
);

INVx3_ASAP7_75t_L g756 ( 
.A(n_706),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_729),
.Y(n_757)
);

INVx2_ASAP7_75t_SL g758 ( 
.A(n_701),
.Y(n_758)
);

BUFx12f_ASAP7_75t_L g759 ( 
.A(n_699),
.Y(n_759)
);

BUFx3_ASAP7_75t_L g760 ( 
.A(n_715),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_727),
.B(n_682),
.Y(n_761)
);

OAI22xp33_ASAP7_75t_L g762 ( 
.A1(n_758),
.A2(n_708),
.B1(n_702),
.B2(n_726),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_759),
.Y(n_763)
);

BUFx6f_ASAP7_75t_SL g764 ( 
.A(n_740),
.Y(n_764)
);

AOI22xp33_ASAP7_75t_L g765 ( 
.A1(n_758),
.A2(n_696),
.B1(n_710),
.B2(n_647),
.Y(n_765)
);

INVx3_ASAP7_75t_L g766 ( 
.A(n_754),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_750),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_739),
.Y(n_768)
);

INVx3_ASAP7_75t_L g769 ( 
.A(n_754),
.Y(n_769)
);

AOI22xp33_ASAP7_75t_L g770 ( 
.A1(n_747),
.A2(n_708),
.B1(n_655),
.B2(n_723),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_732),
.B(n_691),
.Y(n_771)
);

CKINVDCx20_ASAP7_75t_R g772 ( 
.A(n_740),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_750),
.Y(n_773)
);

INVx2_ASAP7_75t_SL g774 ( 
.A(n_743),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_739),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_731),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_744),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_744),
.Y(n_778)
);

BUFx3_ASAP7_75t_L g779 ( 
.A(n_743),
.Y(n_779)
);

AOI22xp33_ASAP7_75t_SL g780 ( 
.A1(n_747),
.A2(n_692),
.B1(n_691),
.B2(n_700),
.Y(n_780)
);

AOI22xp33_ASAP7_75t_L g781 ( 
.A1(n_761),
.A2(n_625),
.B1(n_703),
.B2(n_719),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_731),
.Y(n_782)
);

AOI22xp33_ASAP7_75t_L g783 ( 
.A1(n_752),
.A2(n_707),
.B1(n_730),
.B2(n_722),
.Y(n_783)
);

BUFx3_ASAP7_75t_L g784 ( 
.A(n_749),
.Y(n_784)
);

INVx3_ASAP7_75t_L g785 ( 
.A(n_779),
.Y(n_785)
);

AOI22xp33_ASAP7_75t_SL g786 ( 
.A1(n_771),
.A2(n_676),
.B1(n_683),
.B2(n_651),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_773),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_765),
.B(n_718),
.Y(n_788)
);

AOI22xp33_ASAP7_75t_SL g789 ( 
.A1(n_772),
.A2(n_656),
.B1(n_565),
.B2(n_642),
.Y(n_789)
);

AOI22xp33_ASAP7_75t_L g790 ( 
.A1(n_780),
.A2(n_649),
.B1(n_652),
.B2(n_682),
.Y(n_790)
);

NAND3xp33_ASAP7_75t_L g791 ( 
.A(n_781),
.B(n_617),
.C(n_669),
.Y(n_791)
);

OAI21xp5_ASAP7_75t_SL g792 ( 
.A1(n_762),
.A2(n_669),
.B(n_684),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_770),
.B(n_736),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_773),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_768),
.Y(n_795)
);

OAI22xp5_ASAP7_75t_L g796 ( 
.A1(n_783),
.A2(n_725),
.B1(n_753),
.B2(n_721),
.Y(n_796)
);

AND2x4_ASAP7_75t_L g797 ( 
.A(n_784),
.B(n_749),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_767),
.Y(n_798)
);

AOI22xp33_ASAP7_75t_L g799 ( 
.A1(n_764),
.A2(n_657),
.B1(n_667),
.B2(n_661),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_776),
.Y(n_800)
);

BUFx4f_ASAP7_75t_SL g801 ( 
.A(n_784),
.Y(n_801)
);

INVx3_ASAP7_75t_SL g802 ( 
.A(n_763),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_782),
.Y(n_803)
);

INVx3_ASAP7_75t_L g804 ( 
.A(n_766),
.Y(n_804)
);

BUFx6f_ASAP7_75t_L g805 ( 
.A(n_774),
.Y(n_805)
);

HB1xp67_ASAP7_75t_L g806 ( 
.A(n_782),
.Y(n_806)
);

OAI22xp5_ASAP7_75t_L g807 ( 
.A1(n_774),
.A2(n_693),
.B1(n_630),
.B2(n_737),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_806),
.Y(n_808)
);

AOI22xp33_ASAP7_75t_L g809 ( 
.A1(n_791),
.A2(n_733),
.B1(n_737),
.B2(n_677),
.Y(n_809)
);

OAI222xp33_ASAP7_75t_L g810 ( 
.A1(n_786),
.A2(n_788),
.B1(n_790),
.B2(n_789),
.C1(n_799),
.C2(n_796),
.Y(n_810)
);

AOI22xp33_ASAP7_75t_L g811 ( 
.A1(n_789),
.A2(n_738),
.B1(n_631),
.B2(n_733),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_793),
.B(n_778),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_806),
.Y(n_813)
);

AOI22xp33_ASAP7_75t_L g814 ( 
.A1(n_798),
.A2(n_778),
.B1(n_777),
.B2(n_775),
.Y(n_814)
);

OAI22xp5_ASAP7_75t_L g815 ( 
.A1(n_792),
.A2(n_760),
.B1(n_714),
.B2(n_745),
.Y(n_815)
);

AOI22xp33_ASAP7_75t_L g816 ( 
.A1(n_802),
.A2(n_680),
.B1(n_760),
.B2(n_679),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_795),
.B(n_777),
.Y(n_817)
);

AOI22xp33_ASAP7_75t_SL g818 ( 
.A1(n_801),
.A2(n_769),
.B1(n_766),
.B2(n_748),
.Y(n_818)
);

OAI22xp5_ASAP7_75t_L g819 ( 
.A1(n_785),
.A2(n_742),
.B1(n_745),
.B2(n_746),
.Y(n_819)
);

OAI22xp5_ASAP7_75t_L g820 ( 
.A1(n_785),
.A2(n_742),
.B1(n_745),
.B2(n_746),
.Y(n_820)
);

AOI22xp33_ASAP7_75t_SL g821 ( 
.A1(n_807),
.A2(n_748),
.B1(n_735),
.B2(n_746),
.Y(n_821)
);

AOI22xp33_ASAP7_75t_L g822 ( 
.A1(n_805),
.A2(n_679),
.B1(n_678),
.B2(n_662),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_797),
.Y(n_823)
);

AOI22xp33_ASAP7_75t_L g824 ( 
.A1(n_787),
.A2(n_635),
.B1(n_481),
.B2(n_668),
.Y(n_824)
);

AOI22xp33_ASAP7_75t_L g825 ( 
.A1(n_805),
.A2(n_746),
.B1(n_734),
.B2(n_735),
.Y(n_825)
);

AOI22xp5_ASAP7_75t_L g826 ( 
.A1(n_804),
.A2(n_637),
.B1(n_639),
.B2(n_668),
.Y(n_826)
);

NAND3xp33_ASAP7_75t_L g827 ( 
.A(n_805),
.B(n_650),
.C(n_481),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_794),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_800),
.B(n_734),
.Y(n_829)
);

AOI22xp33_ASAP7_75t_L g830 ( 
.A1(n_804),
.A2(n_735),
.B1(n_671),
.B2(n_637),
.Y(n_830)
);

AOI22xp33_ASAP7_75t_L g831 ( 
.A1(n_803),
.A2(n_671),
.B1(n_632),
.B2(n_660),
.Y(n_831)
);

AOI22xp33_ASAP7_75t_L g832 ( 
.A1(n_791),
.A2(n_632),
.B1(n_660),
.B2(n_664),
.Y(n_832)
);

AOI22xp33_ASAP7_75t_SL g833 ( 
.A1(n_791),
.A2(n_751),
.B1(n_756),
.B2(n_741),
.Y(n_833)
);

OAI22xp5_ASAP7_75t_L g834 ( 
.A1(n_789),
.A2(n_756),
.B1(n_751),
.B2(n_741),
.Y(n_834)
);

NAND3xp33_ASAP7_75t_L g835 ( 
.A(n_811),
.B(n_757),
.C(n_674),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_828),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_812),
.B(n_757),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_808),
.B(n_639),
.Y(n_838)
);

NAND3xp33_ASAP7_75t_L g839 ( 
.A(n_809),
.B(n_674),
.C(n_660),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_813),
.B(n_419),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_829),
.B(n_697),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_817),
.B(n_664),
.Y(n_842)
);

AND2x2_ASAP7_75t_L g843 ( 
.A(n_823),
.B(n_694),
.Y(n_843)
);

AOI221xp5_ASAP7_75t_L g844 ( 
.A1(n_810),
.A2(n_664),
.B1(n_452),
.B2(n_646),
.C(n_716),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_814),
.B(n_716),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_834),
.B(n_60),
.Y(n_846)
);

NAND3xp33_ASAP7_75t_L g847 ( 
.A(n_833),
.B(n_452),
.C(n_755),
.Y(n_847)
);

NOR3xp33_ASAP7_75t_L g848 ( 
.A(n_815),
.B(n_706),
.C(n_654),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_821),
.B(n_62),
.Y(n_849)
);

NAND3xp33_ASAP7_75t_L g850 ( 
.A(n_826),
.B(n_816),
.C(n_824),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_818),
.B(n_755),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_825),
.B(n_63),
.Y(n_852)
);

OAI21xp5_ASAP7_75t_SL g853 ( 
.A1(n_827),
.A2(n_64),
.B(n_65),
.Y(n_853)
);

AOI22xp33_ASAP7_75t_L g854 ( 
.A1(n_832),
.A2(n_452),
.B1(n_755),
.B2(n_724),
.Y(n_854)
);

OAI21xp5_ASAP7_75t_SL g855 ( 
.A1(n_830),
.A2(n_68),
.B(n_69),
.Y(n_855)
);

AOI22xp33_ASAP7_75t_L g856 ( 
.A1(n_831),
.A2(n_822),
.B1(n_820),
.B2(n_819),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_836),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_840),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_840),
.Y(n_859)
);

NOR3xp33_ASAP7_75t_L g860 ( 
.A(n_844),
.B(n_72),
.C(n_74),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_843),
.B(n_78),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_837),
.B(n_841),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_842),
.B(n_838),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_851),
.B(n_848),
.Y(n_864)
);

NAND4xp25_ASAP7_75t_L g865 ( 
.A(n_850),
.B(n_80),
.C(n_81),
.D(n_82),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_849),
.B(n_85),
.Y(n_866)
);

NAND2x1_ASAP7_75t_L g867 ( 
.A(n_847),
.B(n_755),
.Y(n_867)
);

HB1xp67_ASAP7_75t_L g868 ( 
.A(n_845),
.Y(n_868)
);

AOI22xp33_ASAP7_75t_L g869 ( 
.A1(n_846),
.A2(n_448),
.B1(n_424),
.B2(n_418),
.Y(n_869)
);

AOI22xp5_ASAP7_75t_L g870 ( 
.A1(n_855),
.A2(n_839),
.B1(n_853),
.B2(n_835),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_852),
.B(n_87),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_857),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_857),
.Y(n_873)
);

INVxp67_ASAP7_75t_SL g874 ( 
.A(n_868),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_859),
.Y(n_875)
);

AOI22xp5_ASAP7_75t_L g876 ( 
.A1(n_870),
.A2(n_856),
.B1(n_854),
.B2(n_448),
.Y(n_876)
);

INVx5_ASAP7_75t_L g877 ( 
.A(n_861),
.Y(n_877)
);

OR2x2_ASAP7_75t_L g878 ( 
.A(n_868),
.B(n_101),
.Y(n_878)
);

BUFx2_ASAP7_75t_L g879 ( 
.A(n_858),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_862),
.Y(n_880)
);

AOI22xp5_ASAP7_75t_L g881 ( 
.A1(n_865),
.A2(n_103),
.B1(n_108),
.B2(n_110),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_863),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_864),
.Y(n_883)
);

AOI22xp5_ASAP7_75t_L g884 ( 
.A1(n_883),
.A2(n_860),
.B1(n_869),
.B2(n_871),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_872),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_872),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_873),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_874),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_879),
.Y(n_889)
);

XNOR2xp5_ASAP7_75t_L g890 ( 
.A(n_876),
.B(n_866),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_875),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_882),
.Y(n_892)
);

OR2x2_ASAP7_75t_L g893 ( 
.A(n_880),
.B(n_867),
.Y(n_893)
);

OAI22x1_ASAP7_75t_L g894 ( 
.A1(n_877),
.A2(n_111),
.B1(n_112),
.B2(n_113),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_878),
.Y(n_895)
);

AND2x4_ASAP7_75t_L g896 ( 
.A(n_877),
.B(n_114),
.Y(n_896)
);

XOR2x2_ASAP7_75t_L g897 ( 
.A(n_881),
.B(n_116),
.Y(n_897)
);

INVx2_ASAP7_75t_SL g898 ( 
.A(n_893),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_887),
.Y(n_899)
);

OA22x2_ASAP7_75t_L g900 ( 
.A1(n_884),
.A2(n_125),
.B1(n_133),
.B2(n_134),
.Y(n_900)
);

AOI22xp5_ASAP7_75t_L g901 ( 
.A1(n_897),
.A2(n_135),
.B1(n_136),
.B2(n_137),
.Y(n_901)
);

AOI22xp5_ASAP7_75t_L g902 ( 
.A1(n_896),
.A2(n_140),
.B1(n_143),
.B2(n_145),
.Y(n_902)
);

AOI22x1_ASAP7_75t_L g903 ( 
.A1(n_894),
.A2(n_896),
.B1(n_890),
.B2(n_892),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_885),
.Y(n_904)
);

OA22x2_ASAP7_75t_L g905 ( 
.A1(n_889),
.A2(n_146),
.B1(n_147),
.B2(n_150),
.Y(n_905)
);

XNOR2xp5_ASAP7_75t_L g906 ( 
.A(n_895),
.B(n_888),
.Y(n_906)
);

INVx2_ASAP7_75t_SL g907 ( 
.A(n_892),
.Y(n_907)
);

AOI22xp5_ASAP7_75t_L g908 ( 
.A1(n_891),
.A2(n_154),
.B1(n_155),
.B2(n_156),
.Y(n_908)
);

OA22x2_ASAP7_75t_L g909 ( 
.A1(n_891),
.A2(n_160),
.B1(n_162),
.B2(n_166),
.Y(n_909)
);

AOI22xp5_ASAP7_75t_L g910 ( 
.A1(n_886),
.A2(n_170),
.B1(n_173),
.B2(n_175),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_904),
.Y(n_911)
);

INVxp67_ASAP7_75t_L g912 ( 
.A(n_903),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_899),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_907),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_911),
.Y(n_915)
);

AOI22xp5_ASAP7_75t_L g916 ( 
.A1(n_912),
.A2(n_900),
.B1(n_898),
.B2(n_901),
.Y(n_916)
);

AOI22xp5_ASAP7_75t_L g917 ( 
.A1(n_914),
.A2(n_906),
.B1(n_905),
.B2(n_909),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_913),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_915),
.Y(n_919)
);

OAI22xp5_ASAP7_75t_L g920 ( 
.A1(n_917),
.A2(n_908),
.B1(n_910),
.B2(n_902),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_918),
.Y(n_921)
);

INVx2_ASAP7_75t_SL g922 ( 
.A(n_921),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_919),
.Y(n_923)
);

AOI22xp5_ASAP7_75t_L g924 ( 
.A1(n_920),
.A2(n_916),
.B1(n_177),
.B2(n_178),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_922),
.Y(n_925)
);

OR3x2_ASAP7_75t_L g926 ( 
.A(n_925),
.B(n_923),
.C(n_924),
.Y(n_926)
);

BUFx2_ASAP7_75t_L g927 ( 
.A(n_926),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_927),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_928),
.Y(n_929)
);

AOI22xp5_ASAP7_75t_L g930 ( 
.A1(n_929),
.A2(n_183),
.B1(n_187),
.B2(n_189),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_930),
.Y(n_931)
);

AO22x2_ASAP7_75t_L g932 ( 
.A1(n_931),
.A2(n_193),
.B1(n_197),
.B2(n_200),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_932),
.Y(n_933)
);

AOI221xp5_ASAP7_75t_L g934 ( 
.A1(n_933),
.A2(n_201),
.B1(n_206),
.B2(n_209),
.C(n_211),
.Y(n_934)
);

AOI211xp5_ASAP7_75t_L g935 ( 
.A1(n_934),
.A2(n_214),
.B(n_216),
.C(n_221),
.Y(n_935)
);


endmodule