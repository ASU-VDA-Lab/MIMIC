module fake_jpeg_14886_n_84 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_84);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_84;

wire n_10;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_8;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx1_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

BUFx5_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_3),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_6),
.Y(n_11)
);

INVx6_ASAP7_75t_SL g12 ( 
.A(n_7),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_4),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_17),
.B(n_18),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_16),
.B(n_4),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_16),
.B(n_15),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_19),
.B(n_21),
.Y(n_23)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_8),
.B(n_0),
.Y(n_22)
);

NAND3xp33_ASAP7_75t_L g26 ( 
.A(n_22),
.B(n_10),
.C(n_11),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_19),
.B(n_9),
.C(n_15),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_26),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_20),
.A2(n_12),
.B1(n_14),
.B2(n_8),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_28),
.A2(n_14),
.B1(n_8),
.B2(n_20),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_29),
.A2(n_12),
.B1(n_10),
.B2(n_11),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_18),
.Y(n_30)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_19),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_32),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_23),
.A2(n_17),
.B1(n_21),
.B2(n_20),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_32),
.A2(n_21),
.B1(n_17),
.B2(n_14),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_13),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_34),
.B(n_10),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_27),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_36),
.Y(n_40)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_38),
.B(n_42),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_44),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_36),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_13),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_22),
.Y(n_45)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_0),
.Y(n_46)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

NOR3xp33_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_48),
.C(n_29),
.Y(n_51)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_51),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_9),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_53),
.C(n_39),
.Y(n_62)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_9),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_41),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_54),
.B(n_33),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_57),
.Y(n_61)
);

AOI322xp5_ASAP7_75t_SL g59 ( 
.A1(n_50),
.A2(n_45),
.A3(n_38),
.B1(n_2),
.B2(n_3),
.C1(n_7),
.C2(n_6),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_62),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_58),
.B(n_46),
.Y(n_60)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_64),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_56),
.B(n_33),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_65),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_63),
.A2(n_55),
.B1(n_50),
.B2(n_56),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_70),
.B(n_68),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_67),
.A2(n_61),
.B1(n_53),
.B2(n_62),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_71),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_69),
.A2(n_60),
.B(n_58),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_72),
.A2(n_73),
.B(n_74),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_70),
.A2(n_52),
.B(n_1),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_74),
.B(n_66),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_77),
.B(n_1),
.Y(n_80)
);

MAJx2_ASAP7_75t_L g78 ( 
.A(n_76),
.B(n_66),
.C(n_57),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_78),
.A2(n_79),
.B1(n_80),
.B2(n_12),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_75),
.B(n_54),
.C(n_49),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_81),
.B(n_2),
.Y(n_82)
);

OAI221xp5_ASAP7_75t_L g83 ( 
.A1(n_82),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.C(n_0),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_83),
.B(n_5),
.Y(n_84)
);


endmodule