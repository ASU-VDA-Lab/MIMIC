module fake_jpeg_23288_n_347 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_347);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_347;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_6),
.B(n_10),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_38),
.Y(n_74)
);

INVx11_ASAP7_75t_SL g39 ( 
.A(n_17),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_44),
.A2(n_32),
.B1(n_30),
.B2(n_24),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_17),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_46),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_20),
.B(n_16),
.Y(n_46)
);

BUFx6f_ASAP7_75t_SL g47 ( 
.A(n_22),
.Y(n_47)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_50),
.Y(n_69)
);

BUFx12_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_28),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_52),
.B(n_60),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_44),
.A2(n_27),
.B1(n_21),
.B2(n_25),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_55),
.A2(n_58),
.B1(n_70),
.B2(n_24),
.Y(n_118)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_57),
.B(n_29),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_49),
.A2(n_27),
.B1(n_21),
.B2(n_25),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_24),
.Y(n_60)
);

AND2x2_ASAP7_75t_SL g61 ( 
.A(n_40),
.B(n_33),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_63),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_28),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_34),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_71),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_66),
.A2(n_32),
.B1(n_30),
.B2(n_22),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_38),
.A2(n_27),
.B1(n_21),
.B2(n_30),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_42),
.B(n_34),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_42),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_72),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_43),
.B(n_34),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_23),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_35),
.Y(n_75)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_75),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_76),
.Y(n_122)
);

INVx2_ASAP7_75t_SL g79 ( 
.A(n_56),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_79),
.B(n_83),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_62),
.B(n_20),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_80),
.B(n_103),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_35),
.Y(n_81)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_81),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_82),
.B(n_96),
.Y(n_133)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_67),
.B(n_35),
.Y(n_84)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_84),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_52),
.B(n_35),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_86),
.B(n_90),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_66),
.A2(n_30),
.B1(n_24),
.B2(n_32),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_87),
.A2(n_54),
.B1(n_18),
.B2(n_74),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g123 ( 
.A(n_88),
.Y(n_123)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_89),
.A2(n_91),
.B1(n_95),
.B2(n_99),
.Y(n_147)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_71),
.Y(n_90)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_55),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_92),
.B(n_93),
.Y(n_145)
);

INVx4_ASAP7_75t_SL g93 ( 
.A(n_60),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g129 ( 
.A(n_94),
.Y(n_129)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_51),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_69),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_72),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_97),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

BUFx24_ASAP7_75t_SL g135 ( 
.A(n_98),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_61),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_53),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_106),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_101),
.A2(n_54),
.B1(n_57),
.B2(n_36),
.Y(n_134)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_65),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_102),
.A2(n_104),
.B(n_108),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_73),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_63),
.B(n_35),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_105),
.B(n_109),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_61),
.B(n_43),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_59),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_107),
.B(n_112),
.Y(n_130)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_59),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_62),
.B(n_26),
.Y(n_109)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_68),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_111),
.A2(n_114),
.B1(n_118),
.B2(n_93),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_60),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_113),
.A2(n_31),
.B(n_19),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_60),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_59),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_116),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_61),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_68),
.B(n_31),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_117),
.B(n_23),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_121),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_58),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_124),
.B(n_126),
.C(n_136),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_99),
.B(n_58),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_99),
.A2(n_33),
.B(n_36),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_127),
.A2(n_147),
.B(n_120),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_92),
.A2(n_68),
.B1(n_17),
.B2(n_70),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_128),
.A2(n_138),
.B1(n_141),
.B2(n_76),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_134),
.A2(n_142),
.B1(n_93),
.B2(n_87),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_77),
.B(n_48),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_139),
.B(n_50),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_116),
.A2(n_74),
.B1(n_18),
.B2(n_23),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_118),
.A2(n_18),
.B1(n_23),
.B2(n_26),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_149),
.B(n_19),
.Y(n_168)
);

BUFx2_ASAP7_75t_L g150 ( 
.A(n_123),
.Y(n_150)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_150),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_152),
.A2(n_158),
.B1(n_160),
.B2(n_165),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_136),
.B(n_78),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_153),
.B(n_157),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_140),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_154),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_124),
.B(n_106),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_155),
.A2(n_167),
.B(n_173),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_129),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_156),
.B(n_178),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_133),
.B(n_78),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_145),
.A2(n_112),
.B1(n_77),
.B2(n_103),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_140),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_159),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_145),
.A2(n_83),
.B1(n_90),
.B2(n_82),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_133),
.B(n_110),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_161),
.B(n_162),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_126),
.B(n_110),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_125),
.A2(n_101),
.B1(n_110),
.B2(n_96),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_163),
.A2(n_169),
.B1(n_175),
.B2(n_151),
.Y(n_212)
);

A2O1A1O1Ixp25_ASAP7_75t_L g164 ( 
.A1(n_127),
.A2(n_104),
.B(n_98),
.C(n_88),
.D(n_97),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_164),
.B(n_143),
.C(n_134),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_119),
.A2(n_111),
.B1(n_91),
.B2(n_79),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_135),
.Y(n_166)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_166),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_168),
.B(n_176),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_125),
.A2(n_85),
.B1(n_115),
.B2(n_107),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_146),
.B(n_85),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_170),
.A2(n_174),
.B(n_149),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g171 ( 
.A(n_122),
.Y(n_171)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_171),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_137),
.A2(n_89),
.B1(n_79),
.B2(n_100),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_172),
.A2(n_141),
.B1(n_130),
.B2(n_177),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_119),
.A2(n_95),
.B1(n_108),
.B2(n_102),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_146),
.B(n_94),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_120),
.A2(n_50),
.B(n_1),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_177),
.A2(n_139),
.B(n_142),
.Y(n_195)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_131),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_137),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_180),
.B(n_131),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_179),
.B(n_144),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_182),
.B(n_185),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_179),
.B(n_144),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_186),
.A2(n_204),
.B1(n_198),
.B2(n_175),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_161),
.A2(n_130),
.B(n_143),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_187),
.A2(n_188),
.B(n_195),
.Y(n_240)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_191),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_154),
.B(n_148),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_194),
.B(n_11),
.Y(n_239)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_169),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_197),
.B(n_201),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_162),
.B(n_153),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_200),
.B(n_211),
.Y(n_230)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_150),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_202),
.B(n_209),
.Y(n_229)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_150),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_203),
.B(n_205),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_152),
.A2(n_138),
.B1(n_148),
.B2(n_132),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_171),
.Y(n_205)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_172),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_207),
.B(n_210),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_163),
.B(n_132),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_208),
.B(n_164),
.C(n_167),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_157),
.B(n_0),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_174),
.Y(n_210)
);

MAJx2_ASAP7_75t_L g211 ( 
.A(n_155),
.B(n_158),
.C(n_164),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_212),
.B(n_213),
.Y(n_238)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_170),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_214),
.B(n_208),
.C(n_206),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_190),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_216),
.B(n_223),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_217),
.A2(n_221),
.B1(n_225),
.B2(n_11),
.Y(n_256)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_186),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_219),
.B(n_227),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_207),
.A2(n_197),
.B1(n_188),
.B2(n_204),
.Y(n_221)
);

A2O1A1Ixp33_ASAP7_75t_L g223 ( 
.A1(n_211),
.A2(n_160),
.B(n_159),
.C(n_155),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_189),
.A2(n_178),
.B1(n_168),
.B2(n_156),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_212),
.A2(n_176),
.B1(n_122),
.B2(n_50),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_226),
.A2(n_192),
.B1(n_181),
.B2(n_206),
.Y(n_252)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_183),
.Y(n_227)
);

BUFx2_ASAP7_75t_L g228 ( 
.A(n_205),
.Y(n_228)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_228),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_189),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_231),
.A2(n_233),
.B1(n_236),
.B2(n_12),
.Y(n_265)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_183),
.Y(n_232)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_232),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_195),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_233)
);

NOR2x1_ASAP7_75t_L g234 ( 
.A(n_213),
.B(n_4),
.Y(n_234)
);

NOR3xp33_ASAP7_75t_SL g264 ( 
.A(n_234),
.B(n_9),
.C(n_14),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_209),
.B(n_187),
.Y(n_235)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_235),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_193),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_202),
.Y(n_237)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_237),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_239),
.B(n_242),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_209),
.B(n_4),
.Y(n_241)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_241),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_199),
.B(n_11),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_228),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_244),
.B(n_215),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_230),
.B(n_221),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_245),
.B(n_246),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_222),
.B(n_182),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_222),
.B(n_185),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_247),
.B(n_255),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_SL g273 ( 
.A(n_248),
.B(n_256),
.C(n_264),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_252),
.A2(n_265),
.B1(n_235),
.B2(n_217),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_230),
.B(n_200),
.C(n_196),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_253),
.B(n_261),
.C(n_262),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_219),
.A2(n_184),
.B1(n_5),
.B2(n_7),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_254),
.A2(n_264),
.B1(n_233),
.B2(n_236),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_214),
.B(n_184),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_240),
.B(n_10),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_258),
.B(n_241),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_220),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_259),
.B(n_228),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_240),
.B(n_16),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_229),
.B(n_10),
.Y(n_262)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_268),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_260),
.A2(n_238),
.B(n_237),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_269),
.B(n_281),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_270),
.B(n_285),
.Y(n_301)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_251),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_271),
.B(n_272),
.Y(n_303)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_243),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_274),
.Y(n_294)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_250),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_276),
.B(n_278),
.Y(n_288)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_252),
.Y(n_278)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_279),
.Y(n_290)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_259),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_280),
.B(n_283),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_248),
.B(n_245),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_254),
.A2(n_225),
.B1(n_218),
.B2(n_224),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_282),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_249),
.B(n_215),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_266),
.B(n_232),
.Y(n_284)
);

BUFx24_ASAP7_75t_SL g295 ( 
.A(n_284),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_263),
.A2(n_223),
.B1(n_234),
.B2(n_229),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_262),
.B(n_227),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_286),
.B(n_253),
.C(n_261),
.Y(n_291)
);

FAx1_ASAP7_75t_SL g298 ( 
.A(n_287),
.B(n_226),
.CI(n_231),
.CON(n_298),
.SN(n_298)
);

XNOR2xp5_ASAP7_75t_SL g289 ( 
.A(n_275),
.B(n_247),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_289),
.B(n_302),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_291),
.B(n_299),
.C(n_13),
.Y(n_317)
);

MAJx2_ASAP7_75t_L g292 ( 
.A(n_275),
.B(n_246),
.C(n_255),
.Y(n_292)
);

MAJx2_ASAP7_75t_L g316 ( 
.A(n_292),
.B(n_12),
.C(n_13),
.Y(n_316)
);

BUFx12_ASAP7_75t_L g297 ( 
.A(n_273),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_297),
.B(n_303),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_298),
.B(n_270),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_277),
.B(n_258),
.C(n_239),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_267),
.B(n_257),
.Y(n_302)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_305),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_300),
.A2(n_269),
.B(n_268),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_SL g327 ( 
.A(n_306),
.B(n_307),
.C(n_310),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_297),
.B(n_287),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_309),
.B(n_312),
.Y(n_319)
);

XOR2x2_ASAP7_75t_SL g310 ( 
.A(n_297),
.B(n_273),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_296),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_311),
.B(n_313),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_304),
.A2(n_286),
.B1(n_277),
.B2(n_272),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_295),
.B(n_267),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_293),
.B(n_281),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_314),
.B(n_316),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_290),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_315),
.A2(n_294),
.B1(n_288),
.B2(n_298),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_317),
.B(n_318),
.Y(n_321)
);

OA21x2_ASAP7_75t_SL g318 ( 
.A1(n_301),
.A2(n_14),
.B(n_15),
.Y(n_318)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_323),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_306),
.B(n_293),
.C(n_289),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_324),
.A2(n_325),
.B(n_316),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_308),
.B(n_291),
.C(n_292),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_314),
.B(n_302),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_328),
.B(n_320),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_322),
.B(n_315),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_329),
.B(n_331),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_330),
.B(n_324),
.Y(n_337)
);

OR2x2_ASAP7_75t_L g331 ( 
.A(n_327),
.B(n_310),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_319),
.B(n_317),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_332),
.A2(n_333),
.B(n_325),
.Y(n_340)
);

OR2x2_ASAP7_75t_L g334 ( 
.A(n_320),
.B(n_299),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_334),
.B(n_328),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_336),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_337),
.A2(n_338),
.B(n_340),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_332),
.B(n_326),
.Y(n_338)
);

OAI321xp33_ASAP7_75t_L g343 ( 
.A1(n_341),
.A2(n_339),
.A3(n_335),
.B1(n_321),
.B2(n_308),
.C(n_15),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_343),
.A2(n_342),
.B1(n_14),
.B2(n_8),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_SL g345 ( 
.A1(n_344),
.A2(n_7),
.B(n_8),
.Y(n_345)
);

BUFx24_ASAP7_75t_SL g346 ( 
.A(n_345),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_346),
.B(n_8),
.Y(n_347)
);


endmodule