module fake_jpeg_17600_n_333 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_333);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_333;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx4f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx3_ASAP7_75t_SL g67 ( 
.A(n_35),
.Y(n_67)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_45),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_39),
.A2(n_20),
.B1(n_30),
.B2(n_23),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_48),
.A2(n_66),
.B1(n_27),
.B2(n_18),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_20),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_62),
.Y(n_72)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

OA22x2_ASAP7_75t_L g54 ( 
.A1(n_40),
.A2(n_25),
.B1(n_23),
.B2(n_36),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_54),
.A2(n_21),
.B1(n_42),
.B2(n_41),
.Y(n_77)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_34),
.A2(n_32),
.B1(n_29),
.B2(n_25),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_61),
.A2(n_21),
.B1(n_18),
.B2(n_28),
.Y(n_75)
);

INVx5_ASAP7_75t_SL g62 ( 
.A(n_34),
.Y(n_62)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_35),
.A2(n_32),
.B1(n_29),
.B2(n_25),
.Y(n_66)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_32),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_70),
.B(n_81),
.Y(n_109)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_71),
.B(n_78),
.Y(n_111)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_73),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_75),
.A2(n_68),
.B1(n_55),
.B2(n_49),
.Y(n_108)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_76),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_77),
.A2(n_86),
.B1(n_57),
.B2(n_58),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_80),
.B(n_88),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_59),
.B(n_28),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_67),
.Y(n_83)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_84),
.A2(n_80),
.B1(n_91),
.B2(n_71),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_52),
.B(n_16),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_85),
.B(n_90),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_54),
.A2(n_27),
.B1(n_16),
.B2(n_22),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_87),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_46),
.A2(n_22),
.B1(n_19),
.B2(n_15),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_89),
.A2(n_49),
.B1(n_15),
.B2(n_33),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_54),
.B(n_44),
.Y(n_90)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_60),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_93),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_62),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_94),
.B(n_33),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_90),
.B(n_54),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_96),
.B(n_110),
.C(n_119),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_81),
.B(n_85),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_97),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_86),
.B(n_19),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_98),
.B(n_106),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_SL g130 ( 
.A(n_100),
.B(n_112),
.C(n_120),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_77),
.A2(n_46),
.B1(n_51),
.B2(n_57),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_101),
.Y(n_144)
);

O2A1O1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_70),
.A2(n_63),
.B(n_38),
.C(n_37),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_102),
.A2(n_103),
.B(n_104),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_94),
.A2(n_67),
.B1(n_65),
.B2(n_63),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_60),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_72),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_108),
.A2(n_122),
.B1(n_104),
.B2(n_83),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_72),
.B(n_38),
.C(n_37),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_113),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_79),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_115),
.A2(n_121),
.B1(n_83),
.B2(n_69),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_92),
.B(n_38),
.C(n_44),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_84),
.B(n_0),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_95),
.Y(n_121)
);

A2O1A1O1Ixp25_ASAP7_75t_L g124 ( 
.A1(n_96),
.A2(n_79),
.B(n_73),
.C(n_76),
.D(n_82),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_124),
.A2(n_138),
.B(n_141),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_99),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_125),
.B(n_134),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_109),
.B(n_82),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_126),
.B(n_135),
.Y(n_154)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_99),
.Y(n_127)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_127),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_128),
.A2(n_131),
.B1(n_145),
.B2(n_149),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_114),
.A2(n_69),
.B1(n_93),
.B2(n_95),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_129),
.A2(n_140),
.B1(n_104),
.B2(n_108),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_120),
.A2(n_114),
.B1(n_96),
.B2(n_100),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_118),
.Y(n_132)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_132),
.Y(n_172)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_118),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_133),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_116),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_110),
.B(n_91),
.C(n_74),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_104),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_136),
.B(n_148),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_110),
.B(n_71),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_139),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_98),
.A2(n_53),
.B1(n_42),
.B2(n_44),
.Y(n_140)
);

MAJx2_ASAP7_75t_L g141 ( 
.A(n_97),
.B(n_31),
.C(n_26),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_109),
.B(n_74),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_143),
.B(n_102),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_101),
.A2(n_42),
.B1(n_41),
.B2(n_74),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_116),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_120),
.A2(n_41),
.B1(n_1),
.B2(n_2),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_144),
.A2(n_101),
.B1(n_119),
.B2(n_103),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_150),
.A2(n_157),
.B1(n_169),
.B2(n_171),
.Y(n_180)
);

OR2x2_ASAP7_75t_L g202 ( 
.A(n_152),
.B(n_17),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_144),
.A2(n_120),
.B1(n_122),
.B2(n_112),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_153),
.A2(n_149),
.B(n_148),
.Y(n_182)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_156),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_138),
.A2(n_119),
.B1(n_113),
.B2(n_102),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_127),
.Y(n_158)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_158),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_132),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_160),
.B(n_168),
.Y(n_176)
);

A2O1A1Ixp33_ASAP7_75t_L g161 ( 
.A1(n_136),
.A2(n_124),
.B(n_146),
.C(n_131),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_161),
.B(n_174),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_143),
.B(n_121),
.Y(n_162)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_162),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_137),
.A2(n_103),
.B(n_111),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_165),
.A2(n_173),
.B(n_130),
.Y(n_183)
);

INVxp33_ASAP7_75t_L g168 ( 
.A(n_137),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_138),
.A2(n_107),
.B1(n_105),
.B2(n_117),
.Y(n_169)
);

AO22x1_ASAP7_75t_L g170 ( 
.A1(n_128),
.A2(n_145),
.B1(n_146),
.B2(n_129),
.Y(n_170)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_170),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_123),
.A2(n_115),
.B1(n_107),
.B2(n_117),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_123),
.A2(n_111),
.B(n_31),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_134),
.B(n_87),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_125),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_175),
.B(n_87),
.Y(n_194)
);

XNOR2x1_ASAP7_75t_L g181 ( 
.A(n_154),
.B(n_126),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_181),
.B(n_183),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_182),
.A2(n_1),
.B(n_2),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_154),
.B(n_135),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_184),
.B(n_186),
.C(n_201),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_164),
.B(n_130),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_153),
.A2(n_156),
.B1(n_165),
.B2(n_152),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_187),
.A2(n_196),
.B1(n_167),
.B2(n_165),
.Y(n_206)
);

OAI32xp33_ASAP7_75t_L g188 ( 
.A1(n_155),
.A2(n_147),
.A3(n_140),
.B1(n_141),
.B2(n_142),
.Y(n_188)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_188),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_158),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_189),
.B(n_190),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_158),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_164),
.B(n_133),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_191),
.B(n_173),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_163),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_193),
.B(n_160),
.Y(n_203)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_194),
.Y(n_218)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_163),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_195),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_153),
.A2(n_31),
.B1(n_26),
.B2(n_17),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_162),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_197),
.Y(n_224)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_159),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_198),
.B(n_199),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_159),
.B(n_166),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_172),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_200),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_173),
.B(n_26),
.C(n_17),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_202),
.Y(n_227)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_203),
.Y(n_231)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_206),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_198),
.B(n_166),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_208),
.B(n_195),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_210),
.B(n_219),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_192),
.A2(n_155),
.B1(n_161),
.B2(n_170),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_211),
.A2(n_213),
.B1(n_187),
.B2(n_188),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_192),
.A2(n_175),
.B1(n_169),
.B2(n_170),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_178),
.A2(n_161),
.B1(n_170),
.B2(n_157),
.Y(n_214)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_214),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_184),
.B(n_171),
.C(n_150),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_215),
.B(n_223),
.C(n_226),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_200),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_216),
.B(n_189),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_199),
.B(n_172),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_217),
.A2(n_176),
.B(n_185),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_186),
.B(n_174),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_178),
.A2(n_175),
.B1(n_151),
.B2(n_2),
.Y(n_222)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_222),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_191),
.B(n_0),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_225),
.A2(n_190),
.B(n_4),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_183),
.B(n_3),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_215),
.B(n_181),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_228),
.B(n_242),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_209),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_229),
.B(n_236),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_230),
.B(n_232),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_227),
.A2(n_185),
.B(n_182),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_221),
.B(n_179),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_233),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_220),
.A2(n_179),
.B1(n_197),
.B2(n_180),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_234),
.A2(n_240),
.B1(n_248),
.B2(n_224),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_221),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_237),
.B(n_243),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_227),
.A2(n_180),
.B1(n_202),
.B2(n_196),
.Y(n_242)
);

XOR2x1_ASAP7_75t_SL g252 ( 
.A(n_244),
.B(n_225),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_209),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_245),
.B(n_246),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_217),
.B(n_201),
.Y(n_246)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_217),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_219),
.B(n_177),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_249),
.B(n_206),
.C(n_211),
.Y(n_262)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_250),
.Y(n_270)
);

O2A1O1Ixp33_ASAP7_75t_L g277 ( 
.A1(n_252),
.A2(n_254),
.B(n_229),
.C(n_242),
.Y(n_277)
);

XNOR2x1_ASAP7_75t_L g254 ( 
.A(n_249),
.B(n_207),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_239),
.B(n_212),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_256),
.B(n_258),
.C(n_262),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_239),
.B(n_228),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_235),
.A2(n_204),
.B1(n_218),
.B2(n_212),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_259),
.A2(n_265),
.B1(n_238),
.B2(n_241),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_247),
.B(n_210),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_260),
.B(n_234),
.Y(n_275)
);

MAJx2_ASAP7_75t_L g261 ( 
.A(n_247),
.B(n_207),
.C(n_223),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_261),
.B(n_232),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_246),
.B(n_248),
.C(n_233),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_264),
.B(n_266),
.C(n_268),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_235),
.A2(n_205),
.B1(n_214),
.B2(n_222),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_230),
.B(n_226),
.C(n_177),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_238),
.B(n_3),
.C(n_4),
.Y(n_268)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_271),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_255),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_272),
.B(n_273),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_264),
.B(n_231),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_254),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_275),
.B(n_282),
.Y(n_285)
);

MAJx2_ASAP7_75t_L g289 ( 
.A(n_277),
.B(n_252),
.C(n_263),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_267),
.B(n_231),
.Y(n_278)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_278),
.Y(n_290)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_253),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_279),
.A2(n_281),
.B1(n_284),
.B2(n_261),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_256),
.B(n_244),
.C(n_241),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_280),
.B(n_283),
.C(n_4),
.Y(n_294)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_266),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_258),
.B(n_251),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_251),
.B(n_262),
.C(n_257),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_268),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_287),
.A2(n_8),
.B(n_9),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_289),
.A2(n_8),
.B(n_9),
.Y(n_307)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_291),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_283),
.B(n_3),
.Y(n_292)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_292),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_270),
.A2(n_280),
.B1(n_272),
.B2(n_276),
.Y(n_293)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_293),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_294),
.A2(n_298),
.B(n_292),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_269),
.B(n_276),
.C(n_274),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_295),
.B(n_296),
.C(n_7),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_269),
.B(n_4),
.C(n_5),
.Y(n_296)
);

OA21x2_ASAP7_75t_SL g297 ( 
.A1(n_277),
.A2(n_5),
.B(n_6),
.Y(n_297)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_297),
.Y(n_310)
);

OR2x2_ASAP7_75t_L g298 ( 
.A(n_279),
.B(n_5),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_298),
.B(n_8),
.Y(n_306)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_299),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_290),
.B(n_7),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_301),
.B(n_304),
.Y(n_316)
);

HB1xp67_ASAP7_75t_L g303 ( 
.A(n_286),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_303),
.B(n_306),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_288),
.B(n_7),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_305),
.B(n_294),
.C(n_295),
.Y(n_315)
);

OAI21xp33_ASAP7_75t_SL g317 ( 
.A1(n_307),
.A2(n_289),
.B(n_10),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_309),
.B(n_287),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_307),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_312),
.B(n_314),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_303),
.B(n_296),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_315),
.B(n_319),
.C(n_9),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_317),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_285),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_318),
.A2(n_302),
.B(n_305),
.Y(n_321)
);

OR2x2_ASAP7_75t_L g327 ( 
.A(n_321),
.B(n_323),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_313),
.A2(n_300),
.B(n_310),
.Y(n_323)
);

A2O1A1Ixp33_ASAP7_75t_L g326 ( 
.A1(n_324),
.A2(n_316),
.B(n_311),
.C(n_12),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_311),
.B(n_9),
.C(n_10),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_325),
.A2(n_10),
.B(n_11),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_326),
.A2(n_328),
.B(n_320),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_329),
.A2(n_322),
.B(n_327),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_330),
.A2(n_11),
.B(n_12),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_14),
.C(n_11),
.Y(n_332)
);

FAx1_ASAP7_75t_SL g333 ( 
.A(n_332),
.B(n_13),
.CI(n_14),
.CON(n_333),
.SN(n_333)
);


endmodule