module fake_jpeg_21894_n_25 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_25);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_25;

wire n_13;
wire n_21;
wire n_23;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_24;
wire n_17;
wire n_15;

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_10),
.B(n_5),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_6),
.B(n_9),
.Y(n_14)
);

BUFx10_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_SL g17 ( 
.A1(n_13),
.A2(n_0),
.B(n_2),
.Y(n_17)
);

AO22x1_ASAP7_75t_L g20 ( 
.A1(n_17),
.A2(n_14),
.B1(n_4),
.B2(n_7),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_14),
.B(n_3),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_18),
.B(n_19),
.Y(n_21)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_20),
.B(n_22),
.Y(n_23)
);

OA21x2_ASAP7_75t_L g22 ( 
.A1(n_17),
.A2(n_15),
.B(n_8),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_23),
.B(n_21),
.Y(n_24)
);

A2O1A1Ixp33_ASAP7_75t_L g25 ( 
.A1(n_24),
.A2(n_15),
.B(n_11),
.C(n_12),
.Y(n_25)
);


endmodule