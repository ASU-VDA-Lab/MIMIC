module fake_jpeg_5762_n_120 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_120);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_120;

wire n_117;
wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g10 ( 
.A(n_7),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_7),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

INVx2_ASAP7_75t_SL g14 ( 
.A(n_6),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx5_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_17),
.Y(n_18)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_20),
.B(n_21),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

HB1xp67_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_24),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_25),
.B(n_10),
.Y(n_28)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_28),
.Y(n_38)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_29),
.B(n_32),
.Y(n_45)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_21),
.B(n_14),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_14),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_37),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_23),
.C(n_21),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_35),
.A2(n_18),
.B1(n_23),
.B2(n_20),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_39),
.A2(n_48),
.B1(n_35),
.B2(n_18),
.Y(n_51)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_42),
.Y(n_53)
);

OA22x2_ASAP7_75t_L g41 ( 
.A1(n_33),
.A2(n_22),
.B1(n_24),
.B2(n_18),
.Y(n_41)
);

OA22x2_ASAP7_75t_L g59 ( 
.A1(n_41),
.A2(n_39),
.B1(n_36),
.B2(n_22),
.Y(n_59)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

CKINVDCx14_ASAP7_75t_R g43 ( 
.A(n_30),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_28),
.Y(n_44)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_46),
.A2(n_29),
.B1(n_32),
.B2(n_27),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_33),
.B(n_25),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_33),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_35),
.A2(n_18),
.B1(n_14),
.B2(n_20),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_49),
.B(n_55),
.Y(n_71)
);

HB1xp67_ASAP7_75t_SL g50 ( 
.A(n_41),
.Y(n_50)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_51),
.A2(n_59),
.B1(n_41),
.B2(n_36),
.Y(n_65)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_52),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_37),
.Y(n_66)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_56),
.B(n_58),
.Y(n_72)
);

AOI22x1_ASAP7_75t_SL g57 ( 
.A1(n_41),
.A2(n_33),
.B1(n_24),
.B2(n_29),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_57),
.A2(n_47),
.B1(n_43),
.B2(n_40),
.Y(n_67)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_61),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_66),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_65),
.A2(n_67),
.B1(n_68),
.B2(n_73),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_52),
.A2(n_44),
.B1(n_20),
.B2(n_46),
.Y(n_68)
);

CKINVDCx12_ASAP7_75t_R g69 ( 
.A(n_57),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_69),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_59),
.A2(n_20),
.B1(n_46),
.B2(n_42),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_72),
.A2(n_54),
.B(n_58),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_74),
.A2(n_73),
.B1(n_62),
.B2(n_30),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_66),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_76),
.B(n_77),
.C(n_81),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_63),
.A2(n_59),
.B(n_60),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_63),
.A2(n_59),
.B1(n_60),
.B2(n_55),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_78),
.A2(n_75),
.B1(n_81),
.B2(n_62),
.Y(n_90)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_65),
.C(n_70),
.Y(n_81)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_80),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_83),
.B(n_84),
.Y(n_96)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_77),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_82),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_86),
.A2(n_87),
.B(n_91),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_71),
.Y(n_87)
);

FAx1_ASAP7_75t_SL g94 ( 
.A(n_89),
.B(n_90),
.CI(n_32),
.CON(n_94),
.SN(n_94)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_24),
.Y(n_91)
);

XNOR2x1_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_76),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_88),
.B(n_25),
.C(n_21),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_93),
.B(n_94),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_26),
.Y(n_95)
);

MAJx2_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_21),
.C(n_26),
.Y(n_98)
);

A2O1A1Ixp33_ASAP7_75t_SL g99 ( 
.A1(n_89),
.A2(n_0),
.B(n_21),
.C(n_22),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_92),
.B(n_21),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_96),
.B(n_8),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_102),
.A2(n_99),
.B(n_98),
.Y(n_106)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_97),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_103),
.B(n_104),
.Y(n_109)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_99),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_95),
.B(n_24),
.Y(n_105)
);

MAJx2_ASAP7_75t_L g107 ( 
.A(n_105),
.B(n_16),
.C(n_13),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_106),
.B(n_108),
.Y(n_111)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_100),
.Y(n_108)
);

NOR2xp67_ASAP7_75t_L g110 ( 
.A(n_107),
.B(n_101),
.Y(n_110)
);

AOI21x1_ASAP7_75t_L g114 ( 
.A1(n_110),
.A2(n_5),
.B(n_1),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_109),
.B(n_0),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_112),
.B(n_0),
.Y(n_113)
);

AO21x2_ASAP7_75t_SL g117 ( 
.A1(n_114),
.A2(n_115),
.B(n_4),
.Y(n_117)
);

AOI21x1_ASAP7_75t_L g115 ( 
.A1(n_111),
.A2(n_5),
.B(n_1),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_113),
.A2(n_0),
.B(n_3),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_116),
.B(n_117),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_118),
.Y(n_119)
);

INVxp67_ASAP7_75t_SL g120 ( 
.A(n_119),
.Y(n_120)
);


endmodule