module fake_jpeg_23798_n_8 (n_3, n_2, n_1, n_0, n_4, n_8);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;

output n_8;

wire n_6;
wire n_5;
wire n_7;

MAJx2_ASAP7_75t_L g5 ( 
.A(n_0),
.B(n_2),
.C(n_1),
.Y(n_5)
);

INVx2_ASAP7_75t_L g6 ( 
.A(n_1),
.Y(n_6)
);

O2A1O1Ixp33_ASAP7_75t_SL g7 ( 
.A1(n_4),
.A2(n_2),
.B(n_0),
.C(n_3),
.Y(n_7)
);

AOI22xp5_ASAP7_75t_L g8 ( 
.A1(n_7),
.A2(n_3),
.B1(n_6),
.B2(n_5),
.Y(n_8)
);


endmodule