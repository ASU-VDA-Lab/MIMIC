module fake_jpeg_26033_n_322 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_322);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_322;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_46),
.Y(n_49)
);

AND2x4_ASAP7_75t_SL g43 ( 
.A(n_30),
.B(n_0),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_38),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_25),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_48),
.B(n_60),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_30),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_50),
.B(n_57),
.Y(n_76)
);

CKINVDCx9p33_ASAP7_75t_R g51 ( 
.A(n_43),
.Y(n_51)
);

INVxp33_ASAP7_75t_L g106 ( 
.A(n_51),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_41),
.A2(n_25),
.B1(n_35),
.B2(n_26),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_52),
.A2(n_55),
.B1(n_29),
.B2(n_20),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_47),
.A2(n_25),
.B1(n_30),
.B2(n_23),
.Y(n_55)
);

CKINVDCx5p33_ASAP7_75t_R g57 ( 
.A(n_39),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_43),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_63),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_38),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_29),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_39),
.A2(n_27),
.B1(n_35),
.B2(n_26),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_61),
.A2(n_66),
.B1(n_33),
.B2(n_22),
.Y(n_97)
);

AOI21xp33_ASAP7_75t_L g62 ( 
.A1(n_38),
.A2(n_31),
.B(n_32),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_62),
.B(n_29),
.C(n_17),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_27),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_38),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_65),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_46),
.A2(n_20),
.B1(n_32),
.B2(n_31),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_67),
.B(n_71),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_45),
.B(n_33),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_69),
.B(n_73),
.Y(n_108)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_37),
.Y(n_72)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_77),
.B(n_89),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_78),
.B(n_88),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_48),
.B(n_44),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_81),
.A2(n_86),
.B(n_96),
.Y(n_144)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_84),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_L g85 ( 
.A1(n_53),
.A2(n_17),
.B1(n_28),
.B2(n_37),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_85),
.A2(n_107),
.B1(n_75),
.B2(n_74),
.Y(n_118)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_87),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_58),
.A2(n_36),
.B1(n_34),
.B2(n_19),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_65),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_90),
.B(n_92),
.Y(n_134)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_64),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_93),
.B(n_94),
.Y(n_135)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

O2A1O1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_51),
.A2(n_44),
.B(n_40),
.C(n_37),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_95),
.A2(n_100),
.B1(n_56),
.B2(n_68),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_60),
.A2(n_19),
.B(n_33),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_97),
.A2(n_101),
.B1(n_102),
.B2(n_75),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_63),
.Y(n_98)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_54),
.Y(n_99)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_99),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_59),
.A2(n_22),
.B1(n_28),
.B2(n_17),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_54),
.A2(n_22),
.B1(n_18),
.B2(n_16),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_54),
.A2(n_75),
.B1(n_74),
.B2(n_53),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_50),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_103),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_70),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_104),
.Y(n_130)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_53),
.Y(n_105)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_105),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_62),
.A2(n_28),
.B1(n_18),
.B2(n_44),
.Y(n_107)
);

AOI21xp33_ASAP7_75t_L g110 ( 
.A1(n_59),
.A2(n_18),
.B(n_16),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_110),
.B(n_14),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_72),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_111),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_59),
.B(n_40),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_113),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_67),
.B(n_40),
.C(n_28),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_72),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_114),
.Y(n_141)
);

OA21x2_ASAP7_75t_L g117 ( 
.A1(n_112),
.A2(n_71),
.B(n_73),
.Y(n_117)
);

OA22x2_ASAP7_75t_L g158 ( 
.A1(n_117),
.A2(n_82),
.B1(n_89),
.B2(n_104),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_118),
.A2(n_120),
.B1(n_122),
.B2(n_128),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_106),
.A2(n_74),
.B1(n_57),
.B2(n_68),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_56),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_127),
.B(n_83),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_86),
.A2(n_56),
.B1(n_68),
.B2(n_2),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_109),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_129),
.B(n_132),
.Y(n_154)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_109),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_95),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_133),
.B(n_3),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_137),
.B(n_143),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_138),
.A2(n_142),
.B1(n_1),
.B2(n_3),
.Y(n_171)
);

A2O1A1Ixp33_ASAP7_75t_L g140 ( 
.A1(n_83),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_140)
);

A2O1A1Ixp33_ASAP7_75t_L g146 ( 
.A1(n_140),
.A2(n_80),
.B(n_90),
.C(n_81),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_108),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_81),
.A2(n_13),
.B1(n_12),
.B2(n_11),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_143),
.A2(n_77),
.B1(n_98),
.B2(n_93),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_145),
.B(n_156),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_146),
.A2(n_148),
.B(n_136),
.Y(n_181)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_134),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_147),
.B(n_151),
.Y(n_201)
);

A2O1A1Ixp33_ASAP7_75t_L g148 ( 
.A1(n_136),
.A2(n_78),
.B(n_80),
.C(n_103),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_119),
.B(n_78),
.C(n_113),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_149),
.B(n_136),
.C(n_128),
.Y(n_182)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_123),
.Y(n_150)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_150),
.Y(n_199)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_134),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_130),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_152),
.Y(n_184)
);

A2O1A1O1Ixp25_ASAP7_75t_L g153 ( 
.A1(n_144),
.A2(n_95),
.B(n_96),
.C(n_88),
.D(n_100),
.Y(n_153)
);

AOI21xp33_ASAP7_75t_L g191 ( 
.A1(n_153),
.A2(n_174),
.B(n_176),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_126),
.B(n_82),
.Y(n_155)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_155),
.Y(n_203)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_117),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_123),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_157),
.B(n_167),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_158),
.B(n_160),
.Y(n_205)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_117),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_159),
.B(n_161),
.Y(n_198)
);

OA22x2_ASAP7_75t_L g160 ( 
.A1(n_117),
.A2(n_133),
.B1(n_120),
.B2(n_138),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_127),
.B(n_94),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_162),
.A2(n_163),
.B1(n_165),
.B2(n_168),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_119),
.A2(n_84),
.B1(n_99),
.B2(n_105),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_125),
.A2(n_92),
.B1(n_79),
.B2(n_91),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_144),
.B(n_76),
.Y(n_166)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_166),
.Y(n_180)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_135),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_125),
.A2(n_79),
.B1(n_87),
.B2(n_76),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_126),
.B(n_114),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_169),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_129),
.B(n_111),
.Y(n_170)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_170),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_171),
.A2(n_11),
.B1(n_115),
.B2(n_5),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_122),
.Y(n_172)
);

INVx13_ASAP7_75t_L g179 ( 
.A(n_172),
.Y(n_179)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_135),
.Y(n_173)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_173),
.Y(n_188)
);

OR2x2_ASAP7_75t_SL g174 ( 
.A(n_132),
.B(n_12),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_136),
.B(n_10),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_175),
.B(n_142),
.Y(n_189)
);

AO21x1_ASAP7_75t_L g190 ( 
.A1(n_177),
.A2(n_140),
.B(n_137),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_166),
.B(n_116),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g218 ( 
.A(n_178),
.B(n_181),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_182),
.B(n_161),
.C(n_145),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_156),
.A2(n_118),
.B1(n_116),
.B2(n_141),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_183),
.A2(n_194),
.B1(n_196),
.B2(n_200),
.Y(n_209)
);

CKINVDCx10_ASAP7_75t_R g186 ( 
.A(n_150),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_186),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_189),
.B(n_206),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_190),
.B(n_3),
.Y(n_228)
);

OAI22x1_ASAP7_75t_L g192 ( 
.A1(n_164),
.A2(n_140),
.B1(n_141),
.B2(n_131),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_192),
.A2(n_207),
.B1(n_172),
.B2(n_151),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_159),
.A2(n_131),
.B1(n_130),
.B2(n_121),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_160),
.A2(n_121),
.B1(n_139),
.B2(n_124),
.Y(n_196)
);

INVx11_ASAP7_75t_L g197 ( 
.A(n_157),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_197),
.B(n_3),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_160),
.A2(n_139),
.B1(n_124),
.B2(n_115),
.Y(n_200)
);

BUFx2_ASAP7_75t_L g202 ( 
.A(n_152),
.Y(n_202)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_202),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_175),
.B(n_149),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_162),
.A2(n_163),
.B1(n_160),
.B2(n_168),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_208),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_181),
.A2(n_146),
.B(n_148),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_211),
.A2(n_212),
.B(n_222),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_214),
.B(n_216),
.C(n_223),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_193),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_215),
.B(n_201),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_206),
.B(n_170),
.C(n_147),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_203),
.B(n_173),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_217),
.B(n_228),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_200),
.A2(n_165),
.B1(n_158),
.B2(n_176),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_220),
.A2(n_231),
.B1(n_207),
.B2(n_195),
.Y(n_247)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_202),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_221),
.B(n_233),
.Y(n_236)
);

OA21x2_ASAP7_75t_L g222 ( 
.A1(n_192),
.A2(n_158),
.B(n_153),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_182),
.B(n_154),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_178),
.B(n_167),
.C(n_158),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_224),
.B(n_232),
.C(n_234),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_205),
.A2(n_174),
.B(n_4),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_225),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_205),
.A2(n_115),
.B(n_5),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_226),
.B(n_194),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_184),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_227),
.Y(n_241)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_229),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_187),
.B(n_185),
.Y(n_230)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_230),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_196),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_180),
.B(n_6),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_180),
.B(n_6),
.C(n_7),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_239),
.B(n_256),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_215),
.B(n_187),
.Y(n_242)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_242),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_227),
.B(n_204),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_245),
.B(n_246),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_220),
.B(n_188),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_247),
.A2(n_250),
.B1(n_251),
.B2(n_233),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_249),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_209),
.A2(n_208),
.B1(n_198),
.B2(n_195),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_209),
.A2(n_198),
.B1(n_185),
.B2(n_188),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_230),
.B(n_183),
.Y(n_252)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_252),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_218),
.B(n_189),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_253),
.B(n_219),
.Y(n_262)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_226),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_254),
.B(n_222),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_223),
.B(n_205),
.C(n_191),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_255),
.B(n_219),
.C(n_218),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_210),
.B(n_199),
.Y(n_256)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_258),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_252),
.A2(n_236),
.B1(n_240),
.B2(n_250),
.Y(n_259)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_259),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_260),
.A2(n_274),
.B1(n_235),
.B2(n_254),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_262),
.B(n_265),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_236),
.A2(n_224),
.B1(n_211),
.B2(n_222),
.Y(n_263)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_263),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_242),
.B(n_210),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_266),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_247),
.A2(n_221),
.B1(n_213),
.B2(n_231),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_267),
.A2(n_268),
.B1(n_240),
.B2(n_255),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_251),
.A2(n_214),
.B1(n_179),
.B2(n_216),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_238),
.B(n_232),
.C(n_234),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_269),
.B(n_271),
.C(n_244),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_238),
.B(n_225),
.C(n_199),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_248),
.A2(n_190),
.B(n_179),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_272),
.B(n_243),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_248),
.A2(n_186),
.B1(n_197),
.B2(n_9),
.Y(n_274)
);

OAI21xp33_ASAP7_75t_L g275 ( 
.A1(n_270),
.A2(n_249),
.B(n_243),
.Y(n_275)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_275),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_277),
.A2(n_283),
.B1(n_288),
.B2(n_261),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_266),
.B(n_241),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_279),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_280),
.B(n_264),
.C(n_267),
.Y(n_299)
);

INVxp33_ASAP7_75t_L g282 ( 
.A(n_257),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_282),
.B(n_274),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_271),
.B(n_244),
.C(n_237),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_285),
.B(n_287),
.C(n_269),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_268),
.B(n_237),
.C(n_241),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_289),
.B(n_295),
.C(n_297),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_280),
.B(n_263),
.C(n_265),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_290),
.B(n_292),
.Y(n_302)
);

AOI221xp5_ASAP7_75t_L g291 ( 
.A1(n_281),
.A2(n_258),
.B1(n_259),
.B2(n_264),
.C(n_272),
.Y(n_291)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_291),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_287),
.B(n_261),
.C(n_273),
.Y(n_292)
);

OR2x2_ASAP7_75t_L g306 ( 
.A(n_294),
.B(n_298),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_285),
.B(n_262),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_283),
.B(n_253),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_299),
.B(n_284),
.C(n_286),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_296),
.A2(n_281),
.B1(n_278),
.B2(n_276),
.Y(n_300)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_300),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_291),
.A2(n_276),
.B1(n_286),
.B2(n_278),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_304),
.A2(n_293),
.B1(n_260),
.B2(n_235),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_292),
.B(n_279),
.Y(n_305)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_305),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_307),
.B(n_290),
.C(n_284),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_308),
.B(n_309),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_302),
.B(n_289),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_312),
.A2(n_313),
.B(n_306),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_305),
.A2(n_7),
.B(n_8),
.Y(n_313)
);

AO21x1_ASAP7_75t_L g314 ( 
.A1(n_311),
.A2(n_301),
.B(n_304),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_314),
.A2(n_315),
.B(n_312),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_310),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_317),
.B(n_318),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_319),
.A2(n_303),
.B1(n_8),
.B2(n_9),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_8),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_9),
.Y(n_322)
);


endmodule