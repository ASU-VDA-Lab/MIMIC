module real_aes_3391_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_503;
wire n_357;
wire n_635;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_577;
wire n_580;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_560;
wire n_260;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_453;
wire n_374;
wire n_379;
wire n_235;
wire n_399;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_570;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_547;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_250;
wire n_85;
wire n_605;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_87;
wire n_171;
wire n_78;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_637;
wire n_526;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_601;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
INVx1_ASAP7_75t_L g267 ( .A(n_0), .Y(n_267) );
AOI22xp33_ASAP7_75t_L g163 ( .A1(n_1), .A2(n_24), .B1(n_164), .B2(n_165), .Y(n_163) );
HB1xp67_ASAP7_75t_L g80 ( .A(n_2), .Y(n_80) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_3), .B(n_282), .Y(n_400) );
NAND2xp5_ASAP7_75t_SL g401 ( .A(n_4), .B(n_402), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g345 ( .A1(n_5), .A2(n_28), .B1(n_281), .B2(n_346), .Y(n_345) );
AOI22xp5_ASAP7_75t_L g321 ( .A1(n_6), .A2(n_34), .B1(n_256), .B2(n_322), .Y(n_321) );
AOI22xp5_ASAP7_75t_L g246 ( .A1(n_7), .A2(n_47), .B1(n_230), .B2(n_233), .Y(n_246) );
INVx1_ASAP7_75t_L g262 ( .A(n_8), .Y(n_262) );
INVx1_ASAP7_75t_L g106 ( .A(n_9), .Y(n_106) );
INVxp67_ASAP7_75t_L g123 ( .A(n_9), .Y(n_123) );
NOR2xp33_ASAP7_75t_L g141 ( .A(n_9), .B(n_55), .Y(n_141) );
INVx1_ASAP7_75t_L g265 ( .A(n_10), .Y(n_265) );
OA21x2_ASAP7_75t_L g225 ( .A1(n_11), .A2(n_51), .B(n_226), .Y(n_225) );
OA21x2_ASAP7_75t_L g241 ( .A1(n_11), .A2(n_51), .B(n_226), .Y(n_241) );
NAND2xp5_ASAP7_75t_SL g102 ( .A(n_12), .B(n_91), .Y(n_102) );
AOI22xp5_ASAP7_75t_L g229 ( .A1(n_13), .A2(n_49), .B1(n_230), .B2(n_233), .Y(n_229) );
AOI22xp33_ASAP7_75t_L g115 ( .A1(n_14), .A2(n_73), .B1(n_116), .B2(n_125), .Y(n_115) );
AOI22xp33_ASAP7_75t_L g155 ( .A1(n_15), .A2(n_29), .B1(n_156), .B2(n_159), .Y(n_155) );
INVx1_ASAP7_75t_L g255 ( .A(n_16), .Y(n_255) );
BUFx3_ASAP7_75t_L g184 ( .A(n_17), .Y(n_184) );
BUFx6f_ASAP7_75t_L g91 ( .A(n_18), .Y(n_91) );
HB1xp67_ASAP7_75t_L g171 ( .A(n_19), .Y(n_171) );
AO22x1_ASAP7_75t_L g395 ( .A1(n_19), .A2(n_61), .B1(n_268), .B2(n_396), .Y(n_395) );
CKINVDCx5p33_ASAP7_75t_R g285 ( .A(n_20), .Y(n_285) );
AND2x2_ASAP7_75t_L g299 ( .A(n_21), .B(n_256), .Y(n_299) );
AOI22xp33_ASAP7_75t_L g160 ( .A1(n_22), .A2(n_56), .B1(n_161), .B2(n_162), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_23), .B(n_268), .Y(n_291) );
AOI22x1_ASAP7_75t_L g328 ( .A1(n_25), .A2(n_75), .B1(n_230), .B2(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g92 ( .A(n_26), .Y(n_92) );
NAND2xp5_ASAP7_75t_L g120 ( .A(n_26), .B(n_54), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_27), .B(n_331), .Y(n_347) );
HB1xp67_ASAP7_75t_L g177 ( .A(n_30), .Y(n_177) );
AOI22xp33_ASAP7_75t_L g109 ( .A1(n_31), .A2(n_60), .B1(n_110), .B2(n_114), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g174 ( .A(n_32), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g307 ( .A(n_33), .B(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_35), .B(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_36), .B(n_260), .Y(n_290) );
INVx1_ASAP7_75t_L g226 ( .A(n_37), .Y(n_226) );
HB1xp67_ASAP7_75t_L g176 ( .A(n_38), .Y(n_176) );
HB1xp67_ASAP7_75t_L g195 ( .A(n_39), .Y(n_195) );
AND2x4_ASAP7_75t_L g210 ( .A(n_39), .B(n_193), .Y(n_210) );
BUFx6f_ASAP7_75t_L g208 ( .A(n_40), .Y(n_208) );
INVx2_ASAP7_75t_L g237 ( .A(n_41), .Y(n_237) );
AOI22xp33_ASAP7_75t_L g342 ( .A1(n_42), .A2(n_57), .B1(n_281), .B2(n_329), .Y(n_342) );
CKINVDCx14_ASAP7_75t_R g404 ( .A(n_43), .Y(n_404) );
AND2x2_ASAP7_75t_L g305 ( .A(n_44), .B(n_268), .Y(n_305) );
OA22x2_ASAP7_75t_L g96 ( .A1(n_45), .A2(n_55), .B1(n_91), .B2(n_95), .Y(n_96) );
INVx1_ASAP7_75t_L g130 ( .A(n_45), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_46), .B(n_367), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_48), .B(n_358), .Y(n_357) );
HB1xp67_ASAP7_75t_L g631 ( .A(n_49), .Y(n_631) );
NAND2x1p5_ASAP7_75t_L g309 ( .A(n_50), .B(n_239), .Y(n_309) );
CKINVDCx14_ASAP7_75t_R g334 ( .A(n_52), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g84 ( .A(n_53), .B(n_85), .Y(n_84) );
INVx1_ASAP7_75t_L g108 ( .A(n_54), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_54), .B(n_128), .Y(n_144) );
HB1xp67_ASAP7_75t_L g187 ( .A(n_54), .Y(n_187) );
OAI21xp33_ASAP7_75t_L g131 ( .A1(n_55), .A2(n_62), .B(n_124), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_58), .B(n_282), .Y(n_362) );
AOI22xp33_ASAP7_75t_L g146 ( .A1(n_59), .A2(n_70), .B1(n_147), .B2(n_153), .Y(n_146) );
INVx1_ASAP7_75t_L g94 ( .A(n_62), .Y(n_94) );
NOR2xp33_ASAP7_75t_L g142 ( .A(n_62), .B(n_74), .Y(n_142) );
OAI22xp5_ASAP7_75t_L g636 ( .A1(n_63), .A2(n_81), .B1(n_82), .B2(n_637), .Y(n_636) );
CKINVDCx5p33_ASAP7_75t_R g637 ( .A(n_63), .Y(n_637) );
BUFx6f_ASAP7_75t_L g203 ( .A(n_64), .Y(n_203) );
BUFx5_ASAP7_75t_L g232 ( .A(n_64), .Y(n_232) );
INVx1_ASAP7_75t_L g325 ( .A(n_64), .Y(n_325) );
INVx2_ASAP7_75t_L g270 ( .A(n_65), .Y(n_270) );
INVx1_ASAP7_75t_L g135 ( .A(n_66), .Y(n_135) );
AOI21xp33_ASAP7_75t_L g132 ( .A1(n_67), .A2(n_133), .B(n_134), .Y(n_132) );
NAND2xp33_ASAP7_75t_L g301 ( .A(n_68), .B(n_302), .Y(n_301) );
INVx2_ASAP7_75t_SL g193 ( .A(n_69), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_71), .B(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_72), .B(n_308), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g100 ( .A(n_74), .B(n_101), .Y(n_100) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_76), .B(n_296), .Y(n_295) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_179), .B1(n_196), .B2(n_211), .C(n_629), .Y(n_77) );
XNOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_167), .Y(n_78) );
AOI22xp5_ASAP7_75t_L g79 ( .A1(n_80), .A2(n_81), .B1(n_82), .B2(n_166), .Y(n_79) );
CKINVDCx5p33_ASAP7_75t_R g166 ( .A(n_80), .Y(n_166) );
AOI22xp5_ASAP7_75t_SL g630 ( .A1(n_81), .A2(n_82), .B1(n_631), .B2(n_632), .Y(n_630) );
INVx1_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
OR2x2_ASAP7_75t_L g82 ( .A(n_83), .B(n_145), .Y(n_82) );
NAND4xp25_ASAP7_75t_L g83 ( .A(n_84), .B(n_109), .C(n_115), .D(n_132), .Y(n_83) );
INVx2_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
INVx2_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
AND2x2_ASAP7_75t_L g87 ( .A(n_88), .B(n_97), .Y(n_87) );
AND2x4_ASAP7_75t_L g114 ( .A(n_88), .B(n_113), .Y(n_114) );
AND2x4_ASAP7_75t_L g156 ( .A(n_88), .B(n_157), .Y(n_156) );
AND2x4_ASAP7_75t_L g159 ( .A(n_88), .B(n_154), .Y(n_159) );
AND2x2_ASAP7_75t_L g88 ( .A(n_89), .B(n_96), .Y(n_88) );
INVx1_ASAP7_75t_L g112 ( .A(n_89), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g89 ( .A(n_90), .B(n_93), .Y(n_89) );
NAND2xp33_ASAP7_75t_L g90 ( .A(n_91), .B(n_92), .Y(n_90) );
INVx2_ASAP7_75t_L g95 ( .A(n_91), .Y(n_95) );
INVx3_ASAP7_75t_L g101 ( .A(n_91), .Y(n_101) );
NAND2xp33_ASAP7_75t_L g107 ( .A(n_91), .B(n_108), .Y(n_107) );
HB1xp67_ASAP7_75t_L g119 ( .A(n_91), .Y(n_119) );
INVx1_ASAP7_75t_L g124 ( .A(n_91), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_92), .B(n_130), .Y(n_129) );
INVxp67_ASAP7_75t_L g188 ( .A(n_92), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g93 ( .A(n_94), .B(n_95), .Y(n_93) );
OAI21xp5_ASAP7_75t_L g122 ( .A1(n_94), .A2(n_123), .B(n_124), .Y(n_122) );
AND2x2_ASAP7_75t_L g111 ( .A(n_96), .B(n_112), .Y(n_111) );
AND2x2_ASAP7_75t_L g121 ( .A(n_96), .B(n_122), .Y(n_121) );
INVx1_ASAP7_75t_L g149 ( .A(n_96), .Y(n_149) );
AND2x4_ASAP7_75t_L g125 ( .A(n_97), .B(n_126), .Y(n_125) );
AND2x2_ASAP7_75t_L g133 ( .A(n_97), .B(n_111), .Y(n_133) );
AND2x4_ASAP7_75t_L g162 ( .A(n_97), .B(n_148), .Y(n_162) );
AND2x4_ASAP7_75t_L g97 ( .A(n_98), .B(n_103), .Y(n_97) );
INVx2_ASAP7_75t_L g98 ( .A(n_99), .Y(n_98) );
AND2x4_ASAP7_75t_L g113 ( .A(n_99), .B(n_103), .Y(n_113) );
AND2x2_ASAP7_75t_L g117 ( .A(n_99), .B(n_118), .Y(n_117) );
OR2x2_ASAP7_75t_L g151 ( .A(n_99), .B(n_152), .Y(n_151) );
AND2x4_ASAP7_75t_L g157 ( .A(n_99), .B(n_158), .Y(n_157) );
AND2x4_ASAP7_75t_L g99 ( .A(n_100), .B(n_102), .Y(n_99) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_101), .B(n_106), .Y(n_105) );
INVxp67_ASAP7_75t_L g128 ( .A(n_101), .Y(n_128) );
NAND3xp33_ASAP7_75t_L g143 ( .A(n_102), .B(n_127), .C(n_144), .Y(n_143) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_L g152 ( .A(n_104), .Y(n_152) );
AND2x2_ASAP7_75t_L g104 ( .A(n_105), .B(n_107), .Y(n_104) );
AND2x4_ASAP7_75t_L g110 ( .A(n_111), .B(n_113), .Y(n_110) );
AND2x4_ASAP7_75t_L g148 ( .A(n_112), .B(n_149), .Y(n_148) );
AND2x4_ASAP7_75t_L g161 ( .A(n_113), .B(n_148), .Y(n_161) );
AND2x2_ASAP7_75t_L g116 ( .A(n_117), .B(n_121), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_119), .B(n_120), .Y(n_118) );
INVx1_ASAP7_75t_L g139 ( .A(n_119), .Y(n_139) );
HB1xp67_ASAP7_75t_L g185 ( .A(n_120), .Y(n_185) );
AND2x4_ASAP7_75t_L g153 ( .A(n_126), .B(n_154), .Y(n_153) );
AND2x4_ASAP7_75t_L g165 ( .A(n_126), .B(n_157), .Y(n_165) );
AND2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_131), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_128), .B(n_129), .Y(n_127) );
HB1xp67_ASAP7_75t_L g189 ( .A(n_130), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g134 ( .A(n_135), .B(n_136), .Y(n_134) );
INVx4_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx3_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
AO21x2_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_140), .B(n_143), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_141), .B(n_142), .Y(n_140) );
NAND4xp25_ASAP7_75t_L g145 ( .A(n_146), .B(n_155), .C(n_160), .D(n_163), .Y(n_145) );
AND2x4_ASAP7_75t_L g147 ( .A(n_148), .B(n_150), .Y(n_147) );
AND2x4_ASAP7_75t_L g164 ( .A(n_148), .B(n_157), .Y(n_164) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g154 ( .A(n_151), .Y(n_154) );
INVx1_ASAP7_75t_L g158 ( .A(n_152), .Y(n_158) );
OAI22xp5_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_169), .B1(n_175), .B2(n_178), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
OAI22xp5_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_171), .B1(n_172), .B2(n_173), .Y(n_169) );
CKINVDCx5p33_ASAP7_75t_R g170 ( .A(n_171), .Y(n_170) );
INVx1_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
HB1xp67_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx1_ASAP7_75t_L g178 ( .A(n_175), .Y(n_178) );
XOR2xp5_ASAP7_75t_L g175 ( .A(n_176), .B(n_177), .Y(n_175) );
BUFx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
CKINVDCx5p33_ASAP7_75t_R g180 ( .A(n_181), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_182), .B(n_190), .Y(n_181) );
INVxp67_ASAP7_75t_SL g182 ( .A(n_183), .Y(n_182) );
AND2x2_ASAP7_75t_L g634 ( .A(n_183), .B(n_190), .Y(n_634) );
AOI211xp5_ASAP7_75t_L g183 ( .A1(n_184), .A2(n_185), .B(n_186), .C(n_189), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_187), .B(n_188), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g190 ( .A(n_191), .B(n_194), .Y(n_190) );
OR2x2_ASAP7_75t_L g639 ( .A(n_191), .B(n_195), .Y(n_639) );
INVx1_ASAP7_75t_L g642 ( .A(n_191), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_191), .B(n_194), .Y(n_643) );
HB1xp67_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
HB1xp67_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
INVx1_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
BUFx2_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
AND2x2_ASAP7_75t_L g197 ( .A(n_198), .B(n_209), .Y(n_197) );
OA21x2_ASAP7_75t_L g641 ( .A1(n_198), .A2(n_642), .B(n_643), .Y(n_641) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_199), .B(n_204), .Y(n_198) );
CKINVDCx16_ASAP7_75t_R g199 ( .A(n_200), .Y(n_199) );
HB1xp67_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx2_ASAP7_75t_L g260 ( .A(n_202), .Y(n_260) );
INVx2_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
INVx3_ASAP7_75t_L g235 ( .A(n_203), .Y(n_235) );
INVx6_ASAP7_75t_L g258 ( .A(n_203), .Y(n_258) );
INVx2_ASAP7_75t_L g288 ( .A(n_203), .Y(n_288) );
CKINVDCx20_ASAP7_75t_R g204 ( .A(n_205), .Y(n_204) );
HB1xp67_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_206), .B(n_284), .Y(n_283) );
OAI22x1_ASAP7_75t_L g320 ( .A1(n_206), .A2(n_321), .B1(n_326), .B2(n_328), .Y(n_320) );
INVx4_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
OAI22xp5_ASAP7_75t_L g280 ( .A1(n_207), .A2(n_281), .B1(n_283), .B2(n_286), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_207), .B(n_340), .Y(n_339) );
AOI21xp5_ASAP7_75t_L g360 ( .A1(n_207), .A2(n_361), .B(n_362), .Y(n_360) );
BUFx6f_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
INVx4_ASAP7_75t_L g223 ( .A(n_208), .Y(n_223) );
INVx3_ASAP7_75t_L g245 ( .A(n_208), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g254 ( .A(n_208), .B(n_255), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g261 ( .A(n_208), .B(n_262), .Y(n_261) );
BUFx6f_ASAP7_75t_L g293 ( .A(n_208), .Y(n_293) );
INVxp67_ASAP7_75t_L g303 ( .A(n_208), .Y(n_303) );
INVx1_ASAP7_75t_L g327 ( .A(n_208), .Y(n_327) );
OAI21x1_ASAP7_75t_L g279 ( .A1(n_209), .A2(n_280), .B(n_289), .Y(n_279) );
AO31x2_ASAP7_75t_L g319 ( .A1(n_209), .A2(n_320), .A3(n_330), .B(n_333), .Y(n_319) );
AO31x2_ASAP7_75t_L g374 ( .A1(n_209), .A2(n_320), .A3(n_330), .B(n_333), .Y(n_374) );
BUFx6f_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
INVx3_ASAP7_75t_L g228 ( .A(n_210), .Y(n_228) );
INVx1_ASAP7_75t_L g251 ( .A(n_210), .Y(n_251) );
INVx3_ASAP7_75t_L g341 ( .A(n_210), .Y(n_341) );
INVx1_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
HB1xp67_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
NAND2x1p5_ASAP7_75t_L g214 ( .A(n_215), .B(n_503), .Y(n_214) );
NOR4xp75_ASAP7_75t_L g215 ( .A(n_216), .B(n_416), .C(n_434), .D(n_460), .Y(n_215) );
AO21x1_ASAP7_75t_L g216 ( .A1(n_217), .A2(n_272), .B(n_380), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
HB1xp67_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_219), .B(n_413), .Y(n_412) );
AND2x2_ASAP7_75t_L g424 ( .A(n_219), .B(n_390), .Y(n_424) );
INVx2_ASAP7_75t_L g486 ( .A(n_219), .Y(n_486) );
AND2x2_ASAP7_75t_L g219 ( .A(n_220), .B(n_247), .Y(n_219) );
INVx1_ASAP7_75t_L g351 ( .A(n_220), .Y(n_351) );
INVx1_ASAP7_75t_L g379 ( .A(n_220), .Y(n_379) );
AND2x2_ASAP7_75t_L g406 ( .A(n_220), .B(n_248), .Y(n_406) );
INVx1_ASAP7_75t_L g437 ( .A(n_220), .Y(n_437) );
INVx2_ASAP7_75t_L g469 ( .A(n_220), .Y(n_469) );
NOR2x1_ASAP7_75t_L g511 ( .A(n_220), .B(n_512), .Y(n_511) );
HB1xp67_ASAP7_75t_L g526 ( .A(n_220), .Y(n_526) );
AND2x2_ASAP7_75t_L g575 ( .A(n_220), .B(n_355), .Y(n_575) );
OR2x6_ASAP7_75t_L g220 ( .A(n_221), .B(n_242), .Y(n_220) );
OAI21x1_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_229), .B(n_236), .Y(n_221) );
NAND3xp33_ASAP7_75t_SL g222 ( .A(n_223), .B(n_224), .C(n_227), .Y(n_222) );
NOR2xp33_ASAP7_75t_SL g264 ( .A(n_223), .B(n_265), .Y(n_264) );
NOR2xp33_ASAP7_75t_L g266 ( .A(n_223), .B(n_267), .Y(n_266) );
NAND3xp33_ASAP7_75t_L g243 ( .A(n_224), .B(n_227), .C(n_244), .Y(n_243) );
INVx1_ASAP7_75t_L g250 ( .A(n_224), .Y(n_250) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
INVx1_ASAP7_75t_L g332 ( .A(n_225), .Y(n_332) );
NOR2xp33_ASAP7_75t_L g340 ( .A(n_225), .B(n_341), .Y(n_340) );
AOI21xp33_ASAP7_75t_SL g312 ( .A1(n_227), .A2(n_313), .B(n_315), .Y(n_312) );
INVx2_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
NOR2x1_ASAP7_75t_L g369 ( .A(n_228), .B(n_358), .Y(n_369) );
INVx2_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx2_ASAP7_75t_L g268 ( .A(n_232), .Y(n_268) );
INVx2_ASAP7_75t_L g282 ( .A(n_232), .Y(n_282) );
INVx2_ASAP7_75t_L g367 ( .A(n_232), .Y(n_367) );
INVx1_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
INVx1_ASAP7_75t_L g346 ( .A(n_234), .Y(n_346) );
INVx2_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
INVx2_ASAP7_75t_L g365 ( .A(n_235), .Y(n_365) );
INVx1_ASAP7_75t_L g402 ( .A(n_235), .Y(n_402) );
OR2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_238), .Y(n_236) );
INVx1_ASAP7_75t_L g296 ( .A(n_238), .Y(n_296) );
INVx1_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
INVx3_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
INVx2_ASAP7_75t_L g314 ( .A(n_240), .Y(n_314) );
INVx4_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
INVx2_ASAP7_75t_L g271 ( .A(n_241), .Y(n_271) );
BUFx3_ASAP7_75t_L g294 ( .A(n_241), .Y(n_294) );
NOR2xp67_ASAP7_75t_L g242 ( .A(n_243), .B(n_246), .Y(n_242) );
INVx3_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
AND2x2_ASAP7_75t_L g468 ( .A(n_247), .B(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
OR2x2_ASAP7_75t_L g473 ( .A(n_248), .B(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g493 ( .A(n_248), .Y(n_493) );
INVx1_ASAP7_75t_L g512 ( .A(n_248), .Y(n_512) );
AND2x2_ASAP7_75t_L g574 ( .A(n_248), .B(n_439), .Y(n_574) );
INVxp67_ASAP7_75t_L g604 ( .A(n_248), .Y(n_604) );
AO21x2_ASAP7_75t_L g248 ( .A1(n_249), .A2(n_252), .B(n_269), .Y(n_248) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_250), .B(n_251), .Y(n_249) );
OR2x2_ASAP7_75t_L g392 ( .A(n_251), .B(n_296), .Y(n_392) );
NAND3xp33_ASAP7_75t_SL g252 ( .A(n_253), .B(n_259), .C(n_263), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_254), .B(n_256), .Y(n_253) );
INVx2_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
INVx1_ASAP7_75t_L g302 ( .A(n_258), .Y(n_302) );
INVx1_ASAP7_75t_L g308 ( .A(n_258), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_260), .B(n_261), .Y(n_259) );
AOI22xp5_ASAP7_75t_L g263 ( .A1(n_260), .A2(n_264), .B1(n_266), .B2(n_268), .Y(n_263) );
NOR2xp33_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
INVx3_ASAP7_75t_L g358 ( .A(n_271), .Y(n_358) );
OAI22xp5_ASAP7_75t_L g272 ( .A1(n_273), .A2(n_348), .B1(n_370), .B2(n_377), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AND2x4_ASAP7_75t_L g274 ( .A(n_275), .B(n_316), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVx1_ASAP7_75t_L g545 ( .A(n_276), .Y(n_545) );
OR2x2_ASAP7_75t_L g627 ( .A(n_276), .B(n_459), .Y(n_627) );
INVx2_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g458 ( .A(n_277), .B(n_459), .Y(n_458) );
AND2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_297), .Y(n_277) );
AND2x2_ASAP7_75t_L g371 ( .A(n_278), .B(n_372), .Y(n_371) );
NAND2x1_ASAP7_75t_L g420 ( .A(n_278), .B(n_318), .Y(n_420) );
AND2x2_ASAP7_75t_L g555 ( .A(n_278), .B(n_337), .Y(n_555) );
OA21x2_ASAP7_75t_L g278 ( .A1(n_279), .A2(n_294), .B(n_295), .Y(n_278) );
OA21x2_ASAP7_75t_L g386 ( .A1(n_279), .A2(n_294), .B(n_295), .Y(n_386) );
INVx2_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AOI21xp5_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_291), .B(n_292), .Y(n_289) );
INVxp67_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
INVx2_ASAP7_75t_SL g311 ( .A(n_293), .Y(n_311) );
INVx1_ASAP7_75t_L g368 ( .A(n_293), .Y(n_368) );
INVx1_ASAP7_75t_L g394 ( .A(n_293), .Y(n_394) );
INVx3_ASAP7_75t_L g335 ( .A(n_294), .Y(n_335) );
AND2x2_ASAP7_75t_L g381 ( .A(n_297), .B(n_374), .Y(n_381) );
AND2x4_ASAP7_75t_L g409 ( .A(n_297), .B(n_410), .Y(n_409) );
OR2x2_ASAP7_75t_L g528 ( .A(n_297), .B(n_374), .Y(n_528) );
AO21x2_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_304), .B(n_312), .Y(n_297) );
AO21x2_ASAP7_75t_L g376 ( .A1(n_298), .A2(n_304), .B(n_312), .Y(n_376) );
OAI21x1_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_300), .B(n_303), .Y(n_298) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx2_ASAP7_75t_L g329 ( .A(n_302), .Y(n_329) );
OAI21x1_ASAP7_75t_SL g304 ( .A1(n_305), .A2(n_306), .B(n_310), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_307), .B(n_309), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_309), .B(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g315 ( .A(n_309), .Y(n_315) );
AOI21x1_ASAP7_75t_L g399 ( .A1(n_311), .A2(n_400), .B(n_401), .Y(n_399) );
INVx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g316 ( .A(n_317), .B(n_336), .Y(n_316) );
INVx2_ASAP7_75t_L g411 ( .A(n_317), .Y(n_411) );
INVx1_ASAP7_75t_L g443 ( .A(n_317), .Y(n_443) );
INVx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g433 ( .A(n_318), .B(n_376), .Y(n_433) );
INVx1_ASAP7_75t_L g447 ( .A(n_318), .Y(n_447) );
AND2x2_ASAP7_75t_L g587 ( .A(n_318), .B(n_387), .Y(n_587) );
INVx3_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx3_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx2_ASAP7_75t_L g398 ( .A(n_325), .Y(n_398) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_327), .B(n_340), .Y(n_344) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
NOR2xp67_ASAP7_75t_SL g333 ( .A(n_334), .B(n_335), .Y(n_333) );
OR2x2_ASAP7_75t_L g403 ( .A(n_335), .B(n_404), .Y(n_403) );
INVx2_ASAP7_75t_L g459 ( .A(n_336), .Y(n_459) );
OR2x2_ASAP7_75t_L g571 ( .A(n_336), .B(n_420), .Y(n_571) );
INVx2_ASAP7_75t_L g579 ( .A(n_336), .Y(n_579) );
INVx2_ASAP7_75t_SL g336 ( .A(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g337 ( .A(n_338), .B(n_343), .Y(n_337) );
NAND2x1p5_ASAP7_75t_L g372 ( .A(n_338), .B(n_343), .Y(n_372) );
OR2x2_ASAP7_75t_L g338 ( .A(n_339), .B(n_342), .Y(n_338) );
OA21x2_ASAP7_75t_L g343 ( .A1(n_344), .A2(n_345), .B(n_347), .Y(n_343) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_350), .B(n_352), .Y(n_349) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g494 ( .A(n_351), .B(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g519 ( .A(n_353), .B(n_479), .Y(n_519) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
OR2x2_ASAP7_75t_L g453 ( .A(n_354), .B(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
AND2x2_ASAP7_75t_L g390 ( .A(n_355), .B(n_391), .Y(n_390) );
INVx3_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx2_ASAP7_75t_L g415 ( .A(n_356), .Y(n_415) );
AND2x2_ASAP7_75t_L g438 ( .A(n_356), .B(n_439), .Y(n_438) );
AND2x2_ASAP7_75t_L g450 ( .A(n_356), .B(n_391), .Y(n_450) );
AND2x4_ASAP7_75t_L g356 ( .A(n_357), .B(n_359), .Y(n_356) );
OAI21x1_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_363), .B(n_369), .Y(n_359) );
AOI21xp5_ASAP7_75t_L g363 ( .A1(n_364), .A2(n_366), .B(n_368), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_371), .B(n_373), .Y(n_370) );
AND2x2_ASAP7_75t_L g475 ( .A(n_371), .B(n_419), .Y(n_475) );
INVx1_ASAP7_75t_L g588 ( .A(n_371), .Y(n_588) );
AND2x2_ASAP7_75t_L g620 ( .A(n_371), .B(n_447), .Y(n_620) );
INVx2_ASAP7_75t_L g387 ( .A(n_372), .Y(n_387) );
AND2x2_ASAP7_75t_L g430 ( .A(n_372), .B(n_385), .Y(n_430) );
INVx1_ASAP7_75t_L g480 ( .A(n_372), .Y(n_480) );
INVx1_ASAP7_75t_L g532 ( .A(n_372), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_372), .B(n_499), .Y(n_540) );
BUFx3_ASAP7_75t_L g427 ( .A(n_373), .Y(n_427) );
NOR2xp67_ASAP7_75t_L g547 ( .A(n_373), .B(n_429), .Y(n_547) );
AND2x4_ASAP7_75t_L g373 ( .A(n_374), .B(n_375), .Y(n_373) );
INVx1_ASAP7_75t_L g457 ( .A(n_374), .Y(n_457) );
INVx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVxp67_ASAP7_75t_L g419 ( .A(n_376), .Y(n_419) );
INVx1_ASAP7_75t_L g499 ( .A(n_376), .Y(n_499) );
INVx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
AND2x2_ASAP7_75t_L g449 ( .A(n_378), .B(n_450), .Y(n_449) );
OR2x2_ASAP7_75t_L g452 ( .A(n_378), .B(n_453), .Y(n_452) );
HB1xp67_ASAP7_75t_L g481 ( .A(n_378), .Y(n_481) );
OR2x2_ASAP7_75t_L g608 ( .A(n_378), .B(n_485), .Y(n_608) );
INVx2_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
AND2x2_ASAP7_75t_L g471 ( .A(n_379), .B(n_472), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_379), .B(n_537), .Y(n_536) );
OAI32xp33_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_382), .A3(n_388), .B1(n_407), .B2(n_412), .Y(n_380) );
INVx2_ASAP7_75t_L g543 ( .A(n_381), .Y(n_543) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g570 ( .A(n_383), .Y(n_570) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVxp67_ASAP7_75t_L g490 ( .A(n_384), .Y(n_490) );
OR2x2_ASAP7_75t_L g497 ( .A(n_384), .B(n_498), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_385), .B(n_387), .Y(n_384) );
INVx1_ASAP7_75t_L g582 ( .A(n_385), .Y(n_582) );
INVx2_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx2_ASAP7_75t_L g410 ( .A(n_386), .Y(n_410) );
HB1xp67_ASAP7_75t_L g538 ( .A(n_386), .Y(n_538) );
INVx1_ASAP7_75t_L g432 ( .A(n_387), .Y(n_432) );
INVx2_ASAP7_75t_L g422 ( .A(n_388), .Y(n_422) );
OR2x2_ASAP7_75t_L g388 ( .A(n_389), .B(n_405), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
AND2x4_ASAP7_75t_L g510 ( .A(n_390), .B(n_511), .Y(n_510) );
AND2x2_ASAP7_75t_L g597 ( .A(n_390), .B(n_468), .Y(n_597) );
INVx2_ASAP7_75t_SL g439 ( .A(n_391), .Y(n_439) );
OAI21x1_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_393), .B(n_403), .Y(n_391) );
OAI21xp5_ASAP7_75t_L g474 ( .A1(n_392), .A2(n_393), .B(n_403), .Y(n_474) );
AOI21x1_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_395), .B(n_399), .Y(n_393) );
INVx2_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
AND2x2_ASAP7_75t_L g546 ( .A(n_406), .B(n_450), .Y(n_546) );
NAND2x1_ASAP7_75t_SL g568 ( .A(n_406), .B(n_438), .Y(n_568) );
AND2x2_ASAP7_75t_L g577 ( .A(n_406), .B(n_466), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_406), .B(n_619), .Y(n_618) );
INVx2_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
AND2x2_ASAP7_75t_L g621 ( .A(n_408), .B(n_479), .Y(n_621) );
AND2x2_ASAP7_75t_L g408 ( .A(n_409), .B(n_411), .Y(n_408) );
AND2x4_ASAP7_75t_SL g446 ( .A(n_409), .B(n_447), .Y(n_446) );
BUFx3_ASAP7_75t_L g522 ( .A(n_409), .Y(n_522) );
INVxp67_ASAP7_75t_SL g515 ( .A(n_410), .Y(n_515) );
INVx1_ASAP7_75t_L g548 ( .A(n_412), .Y(n_548) );
AOI211xp5_ASAP7_75t_SL g535 ( .A1(n_413), .A2(n_447), .B(n_536), .C(n_538), .Y(n_535) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
AND2x2_ASAP7_75t_L g492 ( .A(n_414), .B(n_493), .Y(n_492) );
OR2x2_ASAP7_75t_L g550 ( .A(n_414), .B(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g617 ( .A(n_414), .B(n_468), .Y(n_617) );
INVx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
AND2x2_ASAP7_75t_L g501 ( .A(n_415), .B(n_437), .Y(n_501) );
OR2x2_ASAP7_75t_L g516 ( .A(n_415), .B(n_473), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g603 ( .A(n_415), .B(n_604), .Y(n_603) );
OAI22xp5_ASAP7_75t_SL g416 ( .A1(n_417), .A2(n_421), .B1(n_423), .B2(n_425), .Y(n_416) );
OR2x2_ASAP7_75t_L g417 ( .A(n_418), .B(n_420), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
HB1xp67_ASAP7_75t_L g514 ( .A(n_419), .Y(n_514) );
AND3x2_ASAP7_75t_L g594 ( .A(n_419), .B(n_579), .C(n_582), .Y(n_594) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
OA21x2_ASAP7_75t_L g425 ( .A1(n_426), .A2(n_428), .B(n_431), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g613 ( .A(n_428), .Y(n_613) );
INVx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g444 ( .A(n_430), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_432), .B(n_433), .Y(n_431) );
BUFx3_ASAP7_75t_L g508 ( .A(n_433), .Y(n_508) );
AND2x2_ASAP7_75t_L g578 ( .A(n_433), .B(n_579), .Y(n_578) );
OAI21xp5_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_440), .B(n_448), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_437), .B(n_438), .Y(n_436) );
AND2x2_ASAP7_75t_L g558 ( .A(n_438), .B(n_468), .Y(n_558) );
INVx2_ASAP7_75t_L g566 ( .A(n_438), .Y(n_566) );
INVx1_ASAP7_75t_L g454 ( .A(n_439), .Y(n_454) );
INVx1_ASAP7_75t_L g483 ( .A(n_439), .Y(n_483) );
INVxp67_ASAP7_75t_SL g440 ( .A(n_441), .Y(n_440) );
NAND2xp5_ASAP7_75t_SL g441 ( .A(n_442), .B(n_445), .Y(n_441) );
OAI22xp5_ASAP7_75t_L g477 ( .A1(n_442), .A2(n_463), .B1(n_478), .B2(n_484), .Y(n_477) );
OR2x2_ASAP7_75t_L g442 ( .A(n_443), .B(n_444), .Y(n_442) );
OR2x2_ASAP7_75t_L g553 ( .A(n_443), .B(n_554), .Y(n_553) );
INVx2_ASAP7_75t_SL g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g463 ( .A(n_446), .Y(n_463) );
OAI21xp5_ASAP7_75t_L g448 ( .A1(n_449), .A2(n_451), .B(n_455), .Y(n_448) );
INVx2_ASAP7_75t_L g485 ( .A(n_450), .Y(n_485) );
AND2x2_ASAP7_75t_L g530 ( .A(n_450), .B(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
OAI22xp5_ASAP7_75t_L g580 ( .A1(n_452), .A2(n_553), .B1(n_581), .B2(n_583), .Y(n_580) );
INVxp67_ASAP7_75t_SL g466 ( .A(n_454), .Y(n_466) );
AND2x2_ASAP7_75t_L g455 ( .A(n_456), .B(n_458), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_456), .B(n_490), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_456), .B(n_570), .Y(n_569) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
NAND3x1_ASAP7_75t_L g460 ( .A(n_461), .B(n_476), .C(n_487), .Y(n_460) );
AOI21x1_ASAP7_75t_L g461 ( .A1(n_462), .A2(n_464), .B(n_470), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
OAI22xp5_ASAP7_75t_L g626 ( .A1(n_465), .A2(n_550), .B1(n_627), .B2(n_628), .Y(n_626) );
OR2x2_ASAP7_75t_L g465 ( .A(n_466), .B(n_467), .Y(n_465) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
AND2x2_ASAP7_75t_L g470 ( .A(n_471), .B(n_475), .Y(n_470) );
INVx1_ASAP7_75t_L g520 ( .A(n_472), .Y(n_520) );
AND2x2_ASAP7_75t_L g600 ( .A(n_472), .B(n_526), .Y(n_600) );
INVx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g502 ( .A(n_473), .Y(n_502) );
BUFx2_ASAP7_75t_L g495 ( .A(n_474), .Y(n_495) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
NAND3xp33_ASAP7_75t_L g478 ( .A(n_479), .B(n_481), .C(n_482), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
AND2x2_ASAP7_75t_L g534 ( .A(n_483), .B(n_493), .Y(n_534) );
OR2x2_ASAP7_75t_L g484 ( .A(n_485), .B(n_486), .Y(n_484) );
INVxp67_ASAP7_75t_L g524 ( .A(n_486), .Y(n_524) );
AOI22xp5_ASAP7_75t_L g487 ( .A1(n_488), .A2(n_491), .B1(n_496), .B2(n_500), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
NAND3xp33_ASAP7_75t_SL g542 ( .A(n_489), .B(n_543), .C(n_544), .Y(n_542) );
AND2x2_ASAP7_75t_L g491 ( .A(n_492), .B(n_494), .Y(n_491) );
AND2x2_ASAP7_75t_L g602 ( .A(n_494), .B(n_603), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_494), .B(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g537 ( .A(n_495), .Y(n_537) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_498), .B(n_532), .Y(n_628) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
AOI22xp5_ASAP7_75t_L g523 ( .A1(n_499), .A2(n_524), .B1(n_525), .B2(n_527), .Y(n_523) );
AND2x2_ASAP7_75t_L g500 ( .A(n_501), .B(n_502), .Y(n_500) );
NAND2x2_ASAP7_75t_L g611 ( .A(n_501), .B(n_612), .Y(n_611) );
NOR2x1_ASAP7_75t_L g503 ( .A(n_504), .B(n_589), .Y(n_503) );
NAND4xp25_ASAP7_75t_L g504 ( .A(n_505), .B(n_541), .C(n_556), .D(n_576), .Y(n_504) );
NOR2xp67_ASAP7_75t_L g505 ( .A(n_506), .B(n_517), .Y(n_505) );
OAI22xp5_ASAP7_75t_L g506 ( .A1(n_507), .A2(n_509), .B1(n_513), .B2(n_516), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
AOI21xp33_ASAP7_75t_L g598 ( .A1(n_509), .A2(n_521), .B(n_599), .Y(n_598) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx2_ASAP7_75t_L g551 ( .A(n_511), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_514), .B(n_515), .Y(n_513) );
OAI211xp5_ASAP7_75t_SL g533 ( .A1(n_515), .A2(n_534), .B(n_535), .C(n_539), .Y(n_533) );
INVx1_ASAP7_75t_L g560 ( .A(n_515), .Y(n_560) );
AOI21xp33_ASAP7_75t_L g585 ( .A1(n_516), .A2(n_586), .B(n_588), .Y(n_585) );
OAI321xp33_ASAP7_75t_L g517 ( .A1(n_518), .A2(n_520), .A3(n_521), .B1(n_523), .B2(n_529), .C(n_533), .Y(n_517) );
INVx2_ASAP7_75t_SL g518 ( .A(n_519), .Y(n_518) );
OR2x2_ASAP7_75t_L g583 ( .A(n_520), .B(n_584), .Y(n_583) );
INVx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_522), .B(n_563), .Y(n_562) );
NOR2x1_ASAP7_75t_R g605 ( .A(n_522), .B(n_586), .Y(n_605) );
HB1xp67_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
AND2x2_ASAP7_75t_L g606 ( .A(n_527), .B(n_555), .Y(n_606) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
OR2x2_ASAP7_75t_L g581 ( .A(n_528), .B(n_582), .Y(n_581) );
INVx2_ASAP7_75t_L g593 ( .A(n_528), .Y(n_593) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g563 ( .A(n_532), .Y(n_563) );
INVxp67_ASAP7_75t_L g619 ( .A(n_537), .Y(n_619) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
AOI222xp33_ASAP7_75t_L g541 ( .A1(n_542), .A2(n_546), .B1(n_547), .B2(n_548), .C1(n_549), .C2(n_552), .Y(n_541) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g610 ( .A(n_545), .Y(n_610) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
OR2x2_ASAP7_75t_L g565 ( .A(n_551), .B(n_566), .Y(n_565) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
AOI221x1_ASAP7_75t_L g556 ( .A1(n_557), .A2(n_559), .B1(n_561), .B2(n_564), .C(n_567), .Y(n_556) );
HB1xp67_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
OAI22xp33_ASAP7_75t_SL g567 ( .A1(n_568), .A2(n_569), .B1(n_571), .B2(n_572), .Y(n_567) );
INVx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
AND2x4_ASAP7_75t_L g573 ( .A(n_574), .B(n_575), .Y(n_573) );
BUFx3_ASAP7_75t_L g612 ( .A(n_574), .Y(n_612) );
INVx2_ASAP7_75t_L g584 ( .A(n_575), .Y(n_584) );
AOI211xp5_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_578), .B(n_580), .C(n_585), .Y(n_576) );
NAND2x1_ASAP7_75t_L g592 ( .A(n_579), .B(n_593), .Y(n_592) );
OAI22xp5_ASAP7_75t_SL g609 ( .A1(n_583), .A2(n_610), .B1(n_611), .B2(n_613), .Y(n_609) );
INVx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
NAND3xp33_ASAP7_75t_SL g589 ( .A(n_590), .B(n_601), .C(n_614), .Y(n_589) );
O2A1O1Ixp33_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_594), .B(n_595), .C(n_598), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVx2_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
AOI221xp5_ASAP7_75t_L g601 ( .A1(n_602), .A2(n_605), .B1(n_606), .B2(n_607), .C(n_609), .Y(n_601) );
HB1xp67_ASAP7_75t_L g625 ( .A(n_604), .Y(n_625) );
INVxp67_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
AOI221xp5_ASAP7_75t_L g614 ( .A1(n_615), .A2(n_620), .B1(n_621), .B2(n_622), .C(n_626), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_616), .B(n_618), .Y(n_615) );
INVx2_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVxp67_ASAP7_75t_SL g622 ( .A(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
OAI222xp33_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_632), .B1(n_633), .B2(n_635), .C1(n_638), .C2(n_640), .Y(n_629) );
CKINVDCx20_ASAP7_75t_R g632 ( .A(n_631), .Y(n_632) );
INVx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
HB1xp67_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
BUFx2_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
endmodule