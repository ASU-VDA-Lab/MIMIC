module real_jpeg_25690_n_26 (n_17, n_8, n_0, n_21, n_2, n_10, n_9, n_12, n_154, n_152, n_147, n_24, n_146, n_6, n_153, n_151, n_23, n_11, n_14, n_25, n_7, n_22, n_18, n_3, n_145, n_5, n_4, n_150, n_1, n_20, n_19, n_148, n_149, n_16, n_15, n_13, n_155, n_26);

input n_17;
input n_8;
input n_0;
input n_21;
input n_2;
input n_10;
input n_9;
input n_12;
input n_154;
input n_152;
input n_147;
input n_24;
input n_146;
input n_6;
input n_153;
input n_151;
input n_23;
input n_11;
input n_14;
input n_25;
input n_7;
input n_22;
input n_18;
input n_3;
input n_145;
input n_5;
input n_4;
input n_150;
input n_1;
input n_20;
input n_19;
input n_148;
input n_149;
input n_16;
input n_15;
input n_13;
input n_155;

output n_26;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_131;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_141;
wire n_139;
wire n_33;
wire n_65;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_118;
wire n_123;
wire n_116;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_30;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

BUFx10_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVx6_ASAP7_75t_SL g69 ( 
.A(n_0),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_1),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_2),
.B(n_30),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_2),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_3),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_4),
.B(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_4),
.B(n_126),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_5),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_6),
.B(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_6),
.B(n_58),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_7),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_8),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_9),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_10),
.B(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_10),
.B(n_78),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_11),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_12),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_13),
.B(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_13),
.B(n_40),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_14),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_15),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_16),
.B(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_16),
.B(n_96),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_17),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_18),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_19),
.B(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_19),
.B(n_107),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_20),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_21),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_22),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_23),
.B(n_45),
.C(n_123),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_24),
.B(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_24),
.B(n_112),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_25),
.B(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_25),
.B(n_47),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_139),
.Y(n_26)
);

AO21x1_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_38),
.B(n_136),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_30),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_32),
.Y(n_30)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_34),
.B(n_104),
.Y(n_103)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_36),
.B(n_119),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_36),
.B(n_132),
.Y(n_131)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_37),
.B(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g85 ( 
.A(n_37),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_37),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_37),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_42),
.B(n_135),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_129),
.B(n_134),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_125),
.B(n_128),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_51),
.B(n_122),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_49),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_49),
.B(n_124),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_49),
.B(n_142),
.Y(n_141)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_50),
.B(n_127),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_116),
.B(n_121),
.Y(n_51)
);

OAI321xp33_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_106),
.A3(n_111),
.B1(n_114),
.B2(n_115),
.C(n_145),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_100),
.B(n_105),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_95),
.B(n_99),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_89),
.B(n_94),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_61),
.B(n_88),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_59),
.B(n_60),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_81),
.B(n_87),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_77),
.B(n_80),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_71),
.B(n_76),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_66),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_65),
.B(n_66),
.Y(n_76)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_68),
.B(n_70),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_68),
.B(n_74),
.Y(n_73)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_72),
.B(n_75),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_83),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_82),
.B(n_83),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_86),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_91),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_90),
.B(n_91),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_93),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_97),
.B(n_98),
.Y(n_96)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_97),
.B(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_102),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_101),
.B(n_102),
.Y(n_105)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_108),
.B(n_110),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_117),
.B(n_120),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_117),
.B(n_120),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_133),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_130),
.B(n_133),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_138),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_137),
.A2(n_140),
.B(n_143),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_137),
.B(n_140),
.Y(n_143)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_146),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_147),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_148),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_149),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_150),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_151),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_152),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_153),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_154),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_155),
.Y(n_113)
);


endmodule