module real_jpeg_9942_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_43;
wire n_37;
wire n_21;
wire n_33;
wire n_38;
wire n_35;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_44;
wire n_28;
wire n_46;
wire n_23;
wire n_47;
wire n_14;
wire n_11;
wire n_45;
wire n_25;
wire n_42;
wire n_7;
wire n_22;
wire n_18;
wire n_39;
wire n_36;
wire n_40;
wire n_41;
wire n_26;
wire n_27;
wire n_20;
wire n_19;
wire n_48;
wire n_32;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_0),
.Y(n_11)
);

OR2x2_ASAP7_75t_SL g12 ( 
.A(n_1),
.B(n_3),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

OR2x2_ASAP7_75t_SL g40 ( 
.A(n_1),
.B(n_24),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_SL g13 ( 
.A1(n_2),
.A2(n_14),
.B1(n_15),
.B2(n_18),
.Y(n_13)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_2),
.B(n_4),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_2),
.B(n_17),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_2),
.B(n_17),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_3),
.B(n_23),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g15 ( 
.A1(n_4),
.A2(n_5),
.B1(n_16),
.B2(n_17),
.Y(n_15)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

OA21x2_ASAP7_75t_L g30 ( 
.A1(n_5),
.A2(n_31),
.B(n_33),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_SL g37 ( 
.A1(n_5),
.A2(n_38),
.B(n_39),
.Y(n_37)
);

NOR5xp2_ASAP7_75t_L g6 ( 
.A(n_7),
.B(n_19),
.C(n_26),
.D(n_36),
.E(n_44),
.Y(n_6)
);

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_8),
.B(n_13),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_9),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_10),
.B(n_12),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_10),
.B(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_10),
.B(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_10),
.B(n_22),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_10),
.B(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_10),
.B(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_11),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_11),
.B(n_18),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_11),
.B(n_37),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_17),
.B(n_18),
.Y(n_32)
);

O2A1O1Ixp33_ASAP7_75t_L g44 ( 
.A1(n_18),
.A2(n_45),
.B(n_46),
.C(n_48),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_25),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

OR2x2_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_24),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_29),
.B1(n_30),
.B2(n_34),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

O2A1O1Ixp33_ASAP7_75t_SL g36 ( 
.A1(n_37),
.A2(n_40),
.B(n_41),
.C(n_43),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_40),
.Y(n_42)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);


endmodule