module fake_jpeg_12963_n_415 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_415);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_415;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_378;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx2_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx4f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_4),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_14),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_38),
.Y(n_79)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_39),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_15),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_40),
.B(n_49),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_41),
.Y(n_103)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_42),
.Y(n_85)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_48),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_15),
.B(n_0),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_50),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_29),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_51),
.B(n_54),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_20),
.B(n_0),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_52),
.B(n_56),
.Y(n_104)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_29),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g78 ( 
.A(n_55),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_20),
.B(n_1),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_57),
.B(n_65),
.Y(n_80)
);

BUFx2_ASAP7_75t_R g58 ( 
.A(n_21),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_58),
.B(n_64),
.Y(n_109)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_59),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_61),
.Y(n_100)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_62),
.Y(n_102)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_16),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_63),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_21),
.B(n_1),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_28),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_16),
.Y(n_66)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_66),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_28),
.Y(n_67)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_22),
.B(n_37),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_37),
.Y(n_82)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_16),
.Y(n_69)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_18),
.Y(n_70)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_19),
.Y(n_71)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_71),
.Y(n_101)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_18),
.Y(n_72)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_72),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_55),
.A2(n_19),
.B1(n_18),
.B2(n_25),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_74),
.A2(n_86),
.B1(n_93),
.B2(n_98),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_82),
.B(n_112),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_64),
.A2(n_19),
.B1(n_18),
.B2(n_26),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_83),
.A2(n_97),
.B1(n_35),
.B2(n_33),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_41),
.A2(n_18),
.B1(n_26),
.B2(n_27),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_39),
.A2(n_18),
.B1(n_26),
.B2(n_27),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_62),
.A2(n_27),
.B1(n_23),
.B2(n_24),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_60),
.A2(n_25),
.B1(n_23),
.B2(n_24),
.Y(n_98)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_63),
.Y(n_106)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_106),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_61),
.A2(n_25),
.B1(n_23),
.B2(n_24),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_108),
.A2(n_17),
.B1(n_32),
.B2(n_34),
.Y(n_129)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_66),
.Y(n_110)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_110),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_47),
.B(n_36),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_47),
.B(n_36),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_113),
.B(n_50),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_69),
.A2(n_34),
.B1(n_32),
.B2(n_17),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_114),
.B(n_58),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_91),
.B(n_50),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_116),
.Y(n_160)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_75),
.Y(n_118)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_118),
.Y(n_174)
);

BUFx12f_ASAP7_75t_L g119 ( 
.A(n_85),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_119),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_109),
.B(n_45),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_120),
.B(n_123),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_109),
.B(n_43),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_121),
.B(n_127),
.Y(n_162)
);

INVx13_ASAP7_75t_L g122 ( 
.A(n_85),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_122),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_109),
.B(n_53),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g164 ( 
.A(n_124),
.B(n_73),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g125 ( 
.A(n_107),
.Y(n_125)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_125),
.Y(n_165)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_103),
.Y(n_126)
);

HB1xp67_ASAP7_75t_L g171 ( 
.A(n_126),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_83),
.B(n_35),
.Y(n_127)
);

AOI21xp33_ASAP7_75t_L g128 ( 
.A1(n_104),
.A2(n_22),
.B(n_33),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_128),
.B(n_132),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_129),
.A2(n_130),
.B1(n_150),
.B2(n_78),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_97),
.A2(n_34),
.B1(n_32),
.B2(n_17),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_114),
.A2(n_46),
.B1(n_44),
.B2(n_48),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_131),
.A2(n_146),
.B1(n_81),
.B2(n_94),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_76),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_75),
.Y(n_133)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_133),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_80),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_134),
.B(n_136),
.Y(n_184)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_84),
.Y(n_135)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_135),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_96),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_78),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_138),
.B(n_139),
.Y(n_190)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_103),
.Y(n_140)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_140),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_141),
.A2(n_88),
.B1(n_95),
.B2(n_94),
.Y(n_191)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_106),
.B(n_38),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_142),
.A2(n_111),
.B(n_101),
.Y(n_179)
);

INVx2_ASAP7_75t_SL g143 ( 
.A(n_92),
.Y(n_143)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_143),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_96),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_144),
.B(n_147),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_88),
.A2(n_71),
.B1(n_67),
.B2(n_70),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_87),
.B(n_84),
.Y(n_147)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_100),
.Y(n_148)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_148),
.Y(n_186)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_73),
.Y(n_149)
);

INVx3_ASAP7_75t_SL g173 ( 
.A(n_149),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g150 ( 
.A(n_107),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_96),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_151),
.B(n_79),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_90),
.B(n_72),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_152),
.B(n_154),
.Y(n_175)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_89),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_153),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_87),
.B(n_59),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_90),
.B(n_2),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_155),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_89),
.B(n_2),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_156),
.B(n_136),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_157),
.A2(n_159),
.B1(n_131),
.B2(n_146),
.Y(n_206)
);

OAI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_115),
.A2(n_81),
.B1(n_100),
.B2(n_101),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_120),
.B(n_110),
.C(n_105),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_161),
.B(n_166),
.Y(n_233)
);

OAI21xp33_ASAP7_75t_L g200 ( 
.A1(n_164),
.A2(n_122),
.B(n_117),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_121),
.B(n_105),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_168),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_123),
.B(n_111),
.C(n_78),
.Y(n_172)
);

MAJx2_ASAP7_75t_L g213 ( 
.A(n_172),
.B(n_185),
.C(n_150),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_179),
.A2(n_183),
.B(n_188),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_182),
.B(n_152),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_124),
.A2(n_127),
.B(n_142),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_147),
.B(n_102),
.C(n_77),
.Y(n_185)
);

OR2x2_ASAP7_75t_L g187 ( 
.A(n_141),
.B(n_99),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_187),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_142),
.A2(n_99),
.B(n_92),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_191),
.A2(n_138),
.B1(n_143),
.B2(n_151),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_154),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_192),
.B(n_162),
.Y(n_212)
);

INVx8_ASAP7_75t_L g193 ( 
.A(n_122),
.Y(n_193)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_193),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_156),
.B(n_102),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_194),
.B(n_144),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_195),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_196),
.A2(n_234),
.B1(n_189),
.B2(n_173),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_198),
.B(n_199),
.Y(n_245)
);

OA21x2_ASAP7_75t_L g260 ( 
.A1(n_200),
.A2(n_186),
.B(n_177),
.Y(n_260)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_195),
.Y(n_201)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_201),
.Y(n_240)
);

BUFx5_ASAP7_75t_L g203 ( 
.A(n_158),
.Y(n_203)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_203),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_180),
.B(n_134),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_204),
.B(n_207),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_192),
.B(n_139),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_205),
.B(n_212),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_206),
.A2(n_214),
.B1(n_218),
.B2(n_223),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_182),
.B(n_137),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_163),
.B(n_137),
.Y(n_208)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_208),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_160),
.A2(n_143),
.B1(n_140),
.B2(n_126),
.Y(n_209)
);

A2O1A1Ixp33_ASAP7_75t_SL g269 ( 
.A1(n_209),
.A2(n_5),
.B(n_6),
.C(n_7),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_180),
.B(n_132),
.Y(n_210)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_210),
.Y(n_259)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_181),
.Y(n_211)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_211),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_213),
.B(n_169),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_157),
.A2(n_77),
.B1(n_145),
.B2(n_117),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_181),
.Y(n_215)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_215),
.Y(n_262)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_158),
.Y(n_217)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_217),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_162),
.A2(n_77),
.B1(n_145),
.B2(n_95),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_194),
.B(n_119),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_219),
.B(n_222),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_175),
.B(n_119),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_175),
.A2(n_94),
.B1(n_153),
.B2(n_135),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_176),
.Y(n_224)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_224),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_187),
.A2(n_133),
.B1(n_118),
.B2(n_148),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_225),
.A2(n_228),
.B1(n_165),
.B2(n_179),
.Y(n_241)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_176),
.Y(n_226)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_226),
.Y(n_270)
);

AND2x2_ASAP7_75t_SL g227 ( 
.A(n_170),
.B(n_119),
.Y(n_227)
);

AND2x2_ASAP7_75t_SL g267 ( 
.A(n_227),
.B(n_42),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_187),
.A2(n_125),
.B1(n_79),
.B2(n_149),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_184),
.B(n_2),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_229),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_190),
.B(n_3),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_230),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_171),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_231),
.B(n_232),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_170),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_160),
.B(n_3),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_233),
.B(n_166),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_235),
.B(n_236),
.C(n_239),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_233),
.B(n_213),
.C(n_232),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_238),
.A2(n_241),
.B1(n_242),
.B2(n_251),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_213),
.B(n_161),
.C(n_169),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_220),
.A2(n_183),
.B1(n_191),
.B2(n_185),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_243),
.B(n_218),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_220),
.A2(n_164),
.B(n_188),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_244),
.A2(n_211),
.B(n_197),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_201),
.A2(n_172),
.B1(n_164),
.B2(n_189),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_202),
.A2(n_193),
.B1(n_178),
.B2(n_167),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_254),
.A2(n_255),
.B1(n_263),
.B2(n_5),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_202),
.A2(n_193),
.B1(n_178),
.B2(n_167),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_206),
.A2(n_165),
.B1(n_177),
.B2(n_186),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_256),
.A2(n_196),
.B1(n_225),
.B2(n_228),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_227),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_258),
.B(n_266),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_260),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_221),
.A2(n_174),
.B1(n_158),
.B2(n_173),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_207),
.B(n_174),
.C(n_173),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_264),
.B(n_231),
.C(n_215),
.Y(n_288)
);

OAI32xp33_ASAP7_75t_L g266 ( 
.A1(n_212),
.A2(n_42),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_266)
);

CKINVDCx14_ASAP7_75t_R g285 ( 
.A(n_267),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_269),
.A2(n_214),
.B(n_223),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_272),
.A2(n_279),
.B1(n_281),
.B2(n_238),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_242),
.A2(n_216),
.B1(n_205),
.B2(n_221),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_273),
.A2(n_283),
.B1(n_249),
.B2(n_266),
.Y(n_322)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_268),
.Y(n_275)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_275),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_239),
.B(n_199),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_276),
.B(n_277),
.C(n_288),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_236),
.B(n_222),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_247),
.A2(n_256),
.B1(n_240),
.B2(n_265),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_244),
.A2(n_227),
.B(n_216),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_280),
.A2(n_290),
.B(n_294),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_247),
.A2(n_227),
.B1(n_219),
.B2(n_198),
.Y(n_281)
);

FAx1_ASAP7_75t_SL g282 ( 
.A(n_246),
.B(n_208),
.CI(n_234),
.CON(n_282),
.SN(n_282)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_282),
.B(n_296),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_257),
.A2(n_246),
.B1(n_245),
.B2(n_265),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_SL g314 ( 
.A(n_284),
.B(n_241),
.Y(n_314)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_268),
.Y(n_286)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_286),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_287),
.B(n_297),
.Y(n_307)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_270),
.Y(n_289)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_289),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_235),
.B(n_226),
.C(n_224),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_291),
.B(n_292),
.C(n_293),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_243),
.B(n_197),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_245),
.B(n_217),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_267),
.A2(n_203),
.B(n_6),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_254),
.Y(n_296)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_270),
.Y(n_298)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_298),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_257),
.B(n_6),
.C(n_7),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_299),
.B(n_300),
.C(n_253),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_251),
.B(n_8),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_277),
.B(n_274),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_301),
.B(n_309),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_305),
.B(n_318),
.Y(n_341)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_293),
.Y(n_308)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_308),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_274),
.B(n_264),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_276),
.B(n_267),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_310),
.B(n_313),
.C(n_317),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_292),
.B(n_260),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_314),
.B(n_278),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_315),
.A2(n_325),
.B1(n_307),
.B2(n_273),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_295),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_316),
.A2(n_326),
.B(n_280),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_291),
.B(n_260),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_290),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_283),
.B(n_259),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_319),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_299),
.B(n_248),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_321),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_322),
.A2(n_323),
.B1(n_272),
.B2(n_282),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_279),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_281),
.Y(n_324)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_324),
.Y(n_334)
);

OA21x2_ASAP7_75t_L g325 ( 
.A1(n_295),
.A2(n_263),
.B(n_255),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_325),
.B(n_316),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_SL g362 ( 
.A(n_328),
.B(n_314),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g364 ( 
.A1(n_329),
.A2(n_269),
.B(n_9),
.Y(n_364)
);

AND2x2_ASAP7_75t_SL g352 ( 
.A(n_330),
.B(n_332),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_301),
.B(n_288),
.C(n_284),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_333),
.B(n_304),
.C(n_303),
.Y(n_356)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_302),
.Y(n_336)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_336),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_320),
.B(n_262),
.Y(n_337)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_337),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_307),
.A2(n_271),
.B1(n_285),
.B2(n_294),
.Y(n_338)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_338),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_326),
.A2(n_282),
.B(n_261),
.Y(n_340)
);

AO21x1_ASAP7_75t_L g353 ( 
.A1(n_340),
.A2(n_307),
.B(n_313),
.Y(n_353)
);

CKINVDCx14_ASAP7_75t_R g350 ( 
.A(n_342),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_304),
.B(n_300),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_344),
.B(n_348),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_322),
.A2(n_250),
.B1(n_237),
.B2(n_252),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_L g359 ( 
.A1(n_345),
.A2(n_346),
.B1(n_347),
.B2(n_237),
.Y(n_359)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_306),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_311),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_325),
.B(n_252),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_SL g349 ( 
.A(n_339),
.B(n_305),
.Y(n_349)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_349),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_353),
.A2(n_338),
.B1(n_329),
.B2(n_330),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_356),
.B(n_360),
.C(n_343),
.Y(n_366)
);

NOR3xp33_ASAP7_75t_L g358 ( 
.A(n_340),
.B(n_312),
.C(n_303),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_358),
.B(n_363),
.Y(n_373)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_359),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_343),
.B(n_333),
.C(n_309),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_344),
.B(n_317),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_361),
.B(n_362),
.Y(n_377)
);

NOR3xp33_ASAP7_75t_L g363 ( 
.A(n_337),
.B(n_310),
.C(n_269),
.Y(n_363)
);

A2O1A1Ixp33_ASAP7_75t_SL g369 ( 
.A1(n_364),
.A2(n_334),
.B(n_332),
.C(n_269),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_SL g365 ( 
.A(n_341),
.B(n_8),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_365),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_366),
.B(n_367),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_360),
.B(n_356),
.C(n_361),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_368),
.A2(n_369),
.B1(n_352),
.B2(n_328),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_357),
.A2(n_348),
.B1(n_334),
.B2(n_335),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_370),
.A2(n_374),
.B1(n_376),
.B2(n_379),
.Y(n_389)
);

INVx1_ASAP7_75t_SL g374 ( 
.A(n_352),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_374),
.B(n_378),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_SL g375 ( 
.A1(n_357),
.A2(n_327),
.B(n_331),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_375),
.A2(n_352),
.B(n_362),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_355),
.B(n_331),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_354),
.B(n_327),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_379),
.B(n_350),
.Y(n_380)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_380),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_371),
.A2(n_353),
.B1(n_364),
.B2(n_351),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_381),
.A2(n_369),
.B1(n_336),
.B2(n_11),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_372),
.B(n_355),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_SL g395 ( 
.A(n_383),
.B(n_386),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_384),
.A2(n_389),
.B1(n_369),
.B2(n_346),
.Y(n_396)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_375),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_385),
.B(n_388),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_367),
.B(n_347),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_SL g390 ( 
.A(n_373),
.B(n_366),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_390),
.A2(n_373),
.B(n_378),
.Y(n_391)
);

AOI21x1_ASAP7_75t_SL g405 ( 
.A1(n_391),
.A2(n_12),
.B(n_13),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_382),
.B(n_377),
.C(n_370),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_392),
.B(n_394),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_387),
.B(n_377),
.C(n_369),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_396),
.B(n_399),
.Y(n_400)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_398),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_387),
.B(n_9),
.C(n_10),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_SL g402 ( 
.A1(n_393),
.A2(n_388),
.B(n_384),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g408 ( 
.A1(n_402),
.A2(n_12),
.B(n_13),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_SL g403 ( 
.A1(n_393),
.A2(n_11),
.B(n_12),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_403),
.B(n_12),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_405),
.B(n_397),
.C(n_399),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_401),
.B(n_395),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_406),
.B(n_407),
.Y(n_411)
);

A2O1A1O1Ixp25_ASAP7_75t_L g410 ( 
.A1(n_408),
.A2(n_409),
.B(n_404),
.C(n_403),
.D(n_14),
.Y(n_410)
);

CKINVDCx16_ASAP7_75t_R g412 ( 
.A(n_410),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_412),
.B(n_411),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_413),
.B(n_400),
.C(n_13),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_414),
.B(n_13),
.C(n_14),
.Y(n_415)
);


endmodule