module fake_aes_11502_n_28 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_28);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_28;
wire n_20;
wire n_23;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_27;
INVx1_ASAP7_75t_SL g14 ( .A(n_11), .Y(n_14) );
NAND2xp5_ASAP7_75t_SL g15 ( .A(n_9), .B(n_3), .Y(n_15) );
INVx6_ASAP7_75t_L g16 ( .A(n_8), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_6), .Y(n_17) );
OA21x2_ASAP7_75t_L g18 ( .A1(n_0), .A2(n_2), .B(n_5), .Y(n_18) );
NAND2xp5_ASAP7_75t_L g19 ( .A(n_17), .B(n_0), .Y(n_19) );
AND2x4_ASAP7_75t_SL g20 ( .A(n_16), .B(n_4), .Y(n_20) );
INVx4_ASAP7_75t_L g21 ( .A(n_20), .Y(n_21) );
OAI33xp33_ASAP7_75t_L g22 ( .A1(n_21), .A2(n_19), .A3(n_15), .B1(n_18), .B2(n_16), .B3(n_14), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_22), .Y(n_23) );
NAND2xp5_ASAP7_75t_L g24 ( .A(n_23), .B(n_21), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_24), .Y(n_25) );
OR3x2_ASAP7_75t_L g26 ( .A(n_25), .B(n_1), .C(n_2), .Y(n_26) );
AND3x1_ASAP7_75t_L g27 ( .A(n_26), .B(n_1), .C(n_18), .Y(n_27) );
AOI222xp33_ASAP7_75t_L g28 ( .A1(n_27), .A2(n_14), .B1(n_10), .B2(n_12), .C1(n_13), .C2(n_7), .Y(n_28) );
endmodule