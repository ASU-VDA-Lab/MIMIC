module fake_jpeg_365_n_324 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_324);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_324;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx8_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx8_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx8_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_11),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_4),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_49),
.Y(n_120)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_50),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_51),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_52),
.Y(n_130)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_53),
.Y(n_111)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_54),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_55),
.Y(n_137)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVx3_ASAP7_75t_SL g149 ( 
.A(n_57),
.Y(n_149)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

BUFx10_ASAP7_75t_L g106 ( 
.A(n_58),
.Y(n_106)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_59),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVx8_ASAP7_75t_L g148 ( 
.A(n_60),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g127 ( 
.A(n_61),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_62),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_63),
.Y(n_104)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_64),
.Y(n_134)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_65),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_66),
.Y(n_140)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_67),
.Y(n_135)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_68),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_22),
.B(n_2),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_69),
.A2(n_72),
.B(n_90),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_70),
.Y(n_136)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_30),
.Y(n_71)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_71),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_22),
.B(n_3),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_30),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g138 ( 
.A(n_73),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_24),
.Y(n_74)
);

BUFx4f_ASAP7_75t_SL g124 ( 
.A(n_74),
.Y(n_124)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_34),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_75),
.Y(n_144)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_76),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_17),
.Y(n_77)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_77),
.Y(n_146)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_34),
.Y(n_78)
);

BUFx4f_ASAP7_75t_L g141 ( 
.A(n_78),
.Y(n_141)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_34),
.Y(n_79)
);

BUFx4f_ASAP7_75t_SL g126 ( 
.A(n_79),
.Y(n_126)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

INVx13_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_18),
.B(n_3),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_84),
.Y(n_102)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_82),
.B(n_86),
.Y(n_105)
);

CKINVDCx6p67_ASAP7_75t_R g83 ( 
.A(n_17),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_83),
.B(n_85),
.Y(n_123)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_38),
.Y(n_84)
);

HAxp5_ASAP7_75t_SL g85 ( 
.A(n_17),
.B(n_3),
.CON(n_85),
.SN(n_85)
);

BUFx12_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_20),
.B(n_4),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_87),
.B(n_99),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

AOI21xp33_ASAP7_75t_SL g108 ( 
.A1(n_88),
.A2(n_94),
.B(n_96),
.Y(n_108)
);

BUFx24_ASAP7_75t_L g89 ( 
.A(n_42),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_92),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_27),
.B(n_6),
.Y(n_90)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_91),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_40),
.B(n_6),
.Y(n_92)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_44),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_97),
.Y(n_113)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_44),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_45),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_95),
.Y(n_116)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_48),
.Y(n_96)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_48),
.Y(n_97)
);

BUFx24_ASAP7_75t_L g98 ( 
.A(n_48),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_100),
.Y(n_114)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_45),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_23),
.Y(n_100)
);

AND2x2_ASAP7_75t_SL g118 ( 
.A(n_87),
.B(n_31),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_118),
.B(n_23),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_83),
.A2(n_31),
.B1(n_43),
.B2(n_37),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_121),
.A2(n_129),
.B1(n_133),
.B2(n_139),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_90),
.B(n_35),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_122),
.B(n_131),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_85),
.A2(n_98),
.B1(n_89),
.B2(n_72),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_69),
.B(n_46),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_70),
.A2(n_43),
.B1(n_37),
.B2(n_32),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_61),
.A2(n_63),
.B1(n_52),
.B2(n_60),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_95),
.B(n_33),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_142),
.B(n_145),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_49),
.B(n_32),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_113),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_152),
.B(n_158),
.Y(n_197)
);

OAI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_123),
.A2(n_57),
.B1(n_55),
.B2(n_51),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_154),
.A2(n_166),
.B1(n_110),
.B2(n_146),
.Y(n_188)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_134),
.Y(n_155)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_155),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_156),
.B(n_175),
.Y(n_204)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_147),
.Y(n_157)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_157),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_126),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_105),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_159),
.B(n_162),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_115),
.B(n_6),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_160),
.B(n_171),
.Y(n_198)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_149),
.Y(n_161)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_161),
.Y(n_194)
);

A2O1A1Ixp33_ASAP7_75t_L g162 ( 
.A1(n_132),
.A2(n_8),
.B(n_11),
.C(n_12),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_149),
.Y(n_163)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_163),
.Y(n_206)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_109),
.Y(n_164)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_164),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_123),
.A2(n_41),
.B1(n_11),
.B2(n_12),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_134),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_167),
.B(n_174),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_108),
.A2(n_41),
.B1(n_13),
.B2(n_14),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_168),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_129),
.A2(n_86),
.B(n_8),
.Y(n_169)
);

O2A1O1Ixp33_ASAP7_75t_L g208 ( 
.A1(n_169),
.A2(n_138),
.B(n_106),
.C(n_124),
.Y(n_208)
);

BUFx2_ASAP7_75t_L g170 ( 
.A(n_148),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_170),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_102),
.B(n_118),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_117),
.Y(n_172)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_172),
.Y(n_189)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_127),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_173),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_127),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_114),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_150),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_176),
.B(n_179),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_133),
.A2(n_15),
.B1(n_116),
.B2(n_104),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_177),
.A2(n_178),
.B1(n_180),
.B2(n_181),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_104),
.A2(n_15),
.B1(n_137),
.B2(n_125),
.Y(n_178)
);

AND2x2_ASAP7_75t_SL g179 ( 
.A(n_143),
.B(n_119),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_120),
.A2(n_137),
.B1(n_125),
.B2(n_130),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_120),
.A2(n_130),
.B1(n_103),
.B2(n_136),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_136),
.A2(n_111),
.B1(n_135),
.B2(n_110),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_182),
.A2(n_141),
.B1(n_112),
.B2(n_140),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_128),
.B(n_107),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_183),
.B(n_101),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_121),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_184),
.B(n_138),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_170),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_185),
.B(n_191),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_186),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_188),
.A2(n_195),
.B1(n_165),
.B2(n_180),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_177),
.A2(n_148),
.B1(n_144),
.B2(n_140),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_184),
.A2(n_138),
.B1(n_112),
.B2(n_144),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_196),
.A2(n_208),
.B(n_174),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_159),
.B(n_124),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_203),
.B(n_210),
.Y(n_228)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_207),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_170),
.Y(n_210)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_211),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_191),
.B(n_171),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_212),
.B(n_223),
.C(n_197),
.Y(n_236)
);

INVx8_ASAP7_75t_L g213 ( 
.A(n_187),
.Y(n_213)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_213),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_190),
.A2(n_153),
.B1(n_160),
.B2(n_175),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_214),
.A2(n_215),
.B1(n_217),
.B2(n_225),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_188),
.A2(n_195),
.B1(n_198),
.B2(n_209),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_202),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_216),
.B(n_220),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_198),
.A2(n_153),
.B1(n_152),
.B2(n_169),
.Y(n_217)
);

NOR2xp67_ASAP7_75t_L g220 ( 
.A(n_204),
.B(n_156),
.Y(n_220)
);

AND2x2_ASAP7_75t_SL g221 ( 
.A(n_209),
.B(n_156),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_221),
.Y(n_234)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_206),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_222),
.B(n_226),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_204),
.B(n_183),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_224),
.A2(n_208),
.B(n_192),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_185),
.A2(n_157),
.B1(n_167),
.B2(n_176),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_206),
.Y(n_226)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_205),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_229),
.B(n_194),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_201),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_230),
.B(n_193),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_216),
.B(n_200),
.Y(n_233)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_233),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_236),
.B(n_215),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_237),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_238),
.A2(n_239),
.B(n_211),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_227),
.A2(n_192),
.B(n_162),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_223),
.B(n_217),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_242),
.B(n_244),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_218),
.A2(n_179),
.B1(n_205),
.B2(n_210),
.Y(n_243)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_243),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_214),
.B(n_166),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_218),
.A2(n_179),
.B1(n_155),
.B2(n_172),
.Y(n_245)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_245),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_212),
.B(n_164),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_246),
.B(n_221),
.C(n_228),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_219),
.B(n_199),
.Y(n_247)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_247),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_248),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_232),
.A2(n_227),
.B(n_224),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_249),
.B(n_263),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_236),
.B(n_220),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_251),
.C(n_253),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_246),
.B(n_234),
.C(n_232),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_234),
.B(n_247),
.C(n_221),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_257),
.B(n_258),
.C(n_261),
.Y(n_273)
);

XNOR2x1_ASAP7_75t_SL g261 ( 
.A(n_233),
.B(n_229),
.Y(n_261)
);

BUFx24_ASAP7_75t_SL g264 ( 
.A(n_259),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_264),
.B(n_267),
.Y(n_280)
);

INVx2_ASAP7_75t_SL g265 ( 
.A(n_262),
.Y(n_265)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_265),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_254),
.B(n_235),
.Y(n_266)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_266),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_249),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_260),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_269),
.A2(n_270),
.B1(n_272),
.B2(n_274),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_255),
.A2(n_241),
.B1(n_240),
.B2(n_238),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_261),
.Y(n_272)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_262),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_254),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_275),
.B(n_235),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_258),
.B(n_240),
.C(n_241),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_276),
.B(n_251),
.C(n_263),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_271),
.B(n_250),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_281),
.Y(n_290)
);

NOR3xp33_ASAP7_75t_SL g279 ( 
.A(n_268),
.B(n_242),
.C(n_239),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_279),
.B(n_286),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_271),
.B(n_253),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_282),
.B(n_285),
.C(n_270),
.Y(n_289)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_284),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_273),
.B(n_257),
.C(n_252),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_273),
.B(n_244),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_276),
.B(n_255),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_288),
.B(n_265),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_289),
.B(n_231),
.C(n_222),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_277),
.A2(n_265),
.B(n_274),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_291),
.A2(n_297),
.B(n_226),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_292),
.B(n_294),
.Y(n_298)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_283),
.Y(n_294)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_287),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_296),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_280),
.A2(n_266),
.B(n_256),
.Y(n_297)
);

AO221x1_ASAP7_75t_L g300 ( 
.A1(n_293),
.A2(n_279),
.B1(n_285),
.B2(n_282),
.C(n_281),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_300),
.A2(n_302),
.B1(n_290),
.B2(n_230),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_289),
.B(n_278),
.C(n_256),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_301),
.B(n_290),
.C(n_291),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_295),
.A2(n_248),
.B(n_231),
.Y(n_302)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_303),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_304),
.B(n_213),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_305),
.B(n_306),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_299),
.A2(n_151),
.B1(n_243),
.B2(n_245),
.Y(n_308)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_308),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_298),
.A2(n_193),
.B1(n_201),
.B2(n_207),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_309),
.A2(n_173),
.B(n_163),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_310),
.A2(n_301),
.B(n_189),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_311),
.B(n_314),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_307),
.A2(n_187),
.B1(n_189),
.B2(n_194),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_315),
.A2(n_199),
.B(n_161),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_312),
.A2(n_305),
.B1(n_309),
.B2(n_187),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_317),
.B(n_314),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_318),
.B(n_313),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_319),
.A2(n_320),
.B(n_316),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_321),
.A2(n_141),
.B1(n_126),
.B2(n_106),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_106),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_323),
.B(n_101),
.Y(n_324)
);


endmodule