module real_jpeg_12962_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_356, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_356;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx4f_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_3),
.B(n_27),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_3),
.B(n_62),
.Y(n_72)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_3),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_3),
.B(n_31),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_3),
.B(n_53),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_3),
.B(n_67),
.Y(n_259)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_5),
.B(n_62),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_5),
.B(n_45),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_5),
.B(n_27),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_5),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_5),
.B(n_31),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_6),
.B(n_31),
.Y(n_30)
);

AND2x2_ASAP7_75t_SL g52 ( 
.A(n_6),
.B(n_53),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_6),
.B(n_67),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_6),
.B(n_45),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_6),
.B(n_51),
.Y(n_102)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_6),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_6),
.B(n_27),
.Y(n_139)
);

AND2x2_ASAP7_75t_SL g286 ( 
.A(n_6),
.B(n_62),
.Y(n_286)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_8),
.B(n_35),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_8),
.B(n_51),
.Y(n_155)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_8),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_8),
.B(n_53),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_8),
.B(n_62),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_8),
.B(n_31),
.Y(n_285)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_9),
.B(n_31),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_9),
.B(n_67),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_9),
.B(n_51),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_9),
.B(n_62),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_9),
.B(n_45),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_10),
.B(n_45),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g49 ( 
.A(n_10),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_10),
.B(n_62),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_10),
.B(n_67),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_10),
.B(n_31),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_10),
.B(n_27),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_10),
.B(n_53),
.Y(n_184)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_11),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_13),
.B(n_27),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_13),
.B(n_62),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_13),
.B(n_67),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_13),
.B(n_51),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_13),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_13),
.B(n_45),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_13),
.B(n_31),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_13),
.B(n_35),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_14),
.B(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_14),
.B(n_51),
.Y(n_80)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_14),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_14),
.B(n_45),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_14),
.B(n_67),
.Y(n_302)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_15),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_146),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_145),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_120),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_20),
.B(n_120),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_82),
.C(n_106),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_21),
.B(n_345),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_64),
.C(n_76),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_22),
.A2(n_23),
.B1(n_339),
.B2(n_340),
.Y(n_338)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_39),
.B2(n_40),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_24),
.B(n_41),
.C(n_58),
.Y(n_108)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

XOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_29),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_26),
.B(n_30),
.C(n_33),
.Y(n_105)
);

INVx5_ASAP7_75t_SL g172 ( 
.A(n_27),
.Y(n_172)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_30),
.A2(n_32),
.B1(n_33),
.B2(n_38),
.Y(n_29)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_37),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_34),
.B(n_117),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_34),
.B(n_49),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_34),
.B(n_203),
.Y(n_274)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_37),
.B(n_162),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_37),
.B(n_172),
.Y(n_224)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_42),
.B1(n_57),
.B2(n_58),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_44),
.B1(n_47),
.B2(n_56),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_44),
.B(n_52),
.C(n_54),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_45),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_52),
.B1(n_54),
.B2(n_55),
.Y(n_47)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_48),
.A2(n_54),
.B1(n_139),
.B2(n_140),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_49),
.B(n_50),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_50),
.B(n_203),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_50),
.B(n_90),
.Y(n_292)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_52),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_66),
.C(n_70),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_52),
.A2(n_55),
.B1(n_66),
.B2(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_52),
.A2(n_55),
.B1(n_164),
.B2(n_165),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_52),
.B(n_164),
.Y(n_180)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_53),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_54),
.B(n_139),
.C(n_274),
.Y(n_295)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_60),
.C(n_61),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_59),
.A2(n_61),
.B1(n_136),
.B2(n_314),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_59),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_60),
.B(n_313),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_61),
.A2(n_136),
.B1(n_137),
.B2(n_138),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_61),
.Y(n_136)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_63),
.B(n_92),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_64),
.B(n_76),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_71),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_65),
.B(n_72),
.C(n_74),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_66),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_66),
.A2(n_79),
.B1(n_231),
.B2(n_232),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_66),
.B(n_231),
.Y(n_263)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_68),
.B(n_160),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_68),
.B(n_203),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_78),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_72),
.A2(n_73),
.B1(n_74),
.B2(n_75),
.Y(n_71)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_72),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_73),
.A2(n_74),
.B1(n_101),
.B2(n_102),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_73),
.A2(n_74),
.B1(n_115),
.B2(n_116),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_73),
.B(n_116),
.C(n_118),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_73),
.B(n_98),
.C(n_102),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_73),
.A2(n_74),
.B1(n_184),
.B2(n_185),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_74),
.B(n_184),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_80),
.C(n_81),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_77),
.B(n_323),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_80),
.A2(n_81),
.B1(n_324),
.B2(n_325),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_80),
.Y(n_325)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_81),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_82),
.B(n_106),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_84),
.B1(n_94),
.B2(n_95),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_83),
.B(n_96),
.C(n_105),
.Y(n_121)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_86),
.B1(n_87),
.B2(n_93),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_85),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_85),
.B(n_88),
.C(n_91),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_91),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_90),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_89),
.B(n_160),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_92),
.B(n_162),
.Y(n_270)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_97),
.B1(n_104),
.B2(n_105),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_99),
.B1(n_100),
.B2(n_103),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_98),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_98),
.A2(n_103),
.B1(n_283),
.B2(n_284),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_98),
.B(n_286),
.C(n_287),
.Y(n_316)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_101),
.A2(n_102),
.B1(n_139),
.B2(n_140),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_101),
.A2(n_102),
.B1(n_226),
.B2(n_227),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_102),
.B(n_224),
.C(n_226),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_108),
.B1(n_109),
.B2(n_110),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_107),
.B(n_111),
.C(n_119),
.Y(n_144)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_119),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_112),
.A2(n_113),
.B1(n_114),
.B2(n_118),
.Y(n_111)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_112),
.Y(n_118)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx24_ASAP7_75t_SL g352 ( 
.A(n_120),
.Y(n_352)
);

FAx1_ASAP7_75t_SL g120 ( 
.A(n_121),
.B(n_122),
.CI(n_144),
.CON(n_120),
.SN(n_120)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_134),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_125),
.B1(n_126),
.B2(n_127),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_129),
.B1(n_130),
.B2(n_133),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_130),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_131),
.B(n_132),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_SL g134 ( 
.A(n_135),
.B(n_141),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_139),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

AOI321xp33_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_332),
.A3(n_342),
.B1(n_346),
.B2(n_351),
.C(n_356),
.Y(n_146)
);

NOR3xp33_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_277),
.C(n_327),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_248),
.B(n_276),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_150),
.A2(n_218),
.B(n_247),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_187),
.B(n_217),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_166),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_152),
.B(n_166),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_157),
.C(n_163),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_153),
.A2(n_169),
.B1(n_170),
.B2(n_178),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_153),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_153),
.B(n_214),
.Y(n_213)
);

FAx1_ASAP7_75t_SL g153 ( 
.A(n_154),
.B(n_155),
.CI(n_156),
.CON(n_153),
.SN(n_153)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_157),
.A2(n_158),
.B1(n_163),
.B2(n_215),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_161),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_159),
.B(n_161),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_160),
.B(n_172),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_162),
.B(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_163),
.Y(n_215)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_179),
.B2(n_186),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_169),
.B(n_178),
.C(n_186),
.Y(n_219)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_170),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_173),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_171),
.B(n_174),
.C(n_177),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_175),
.B1(n_176),
.B2(n_177),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_176),
.Y(n_177)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_179),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_180),
.B(n_182),
.C(n_183),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_184),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_184),
.A2(n_185),
.B1(n_302),
.B2(n_303),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_184),
.B(n_300),
.C(n_303),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_211),
.B(n_216),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_200),
.B(n_210),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_195),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_190),
.B(n_195),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_191),
.B(n_193),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_191),
.A2(n_192),
.B1(n_193),
.B2(n_194),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_196),
.B(n_198),
.C(n_199),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_205),
.B(n_209),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_204),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_202),
.B(n_204),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_206),
.B(n_208),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_212),
.B(n_213),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_219),
.B(n_220),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_222),
.B1(n_233),
.B2(n_234),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_221),
.B(n_235),
.C(n_246),
.Y(n_249)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_228),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_223),
.B(n_229),
.C(n_230),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_236),
.B1(n_245),
.B2(n_246),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_238),
.B1(n_239),
.B2(n_244),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_237),
.B(n_241),
.C(n_243),
.Y(n_267)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_239),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_241),
.B1(n_242),
.B2(n_243),
.Y(n_239)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_240),
.Y(n_243)
);

CKINVDCx14_ASAP7_75t_R g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_249),
.B(n_250),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_266),
.B2(n_275),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_254),
.B1(n_255),
.B2(n_265),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_253),
.B(n_265),
.C(n_275),
.Y(n_328)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_255),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_257),
.B1(n_261),
.B2(n_262),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_256),
.B(n_263),
.C(n_264),
.Y(n_296)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

BUFx24_ASAP7_75t_SL g353 ( 
.A(n_257),
.Y(n_353)
);

FAx1_ASAP7_75t_SL g257 ( 
.A(n_258),
.B(n_259),
.CI(n_260),
.CON(n_257),
.SN(n_257)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_258),
.B(n_259),
.C(n_260),
.Y(n_305)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_266),
.Y(n_275)
);

BUFx24_ASAP7_75t_SL g355 ( 
.A(n_266),
.Y(n_355)
);

FAx1_ASAP7_75t_SL g266 ( 
.A(n_267),
.B(n_268),
.CI(n_272),
.CON(n_266),
.SN(n_266)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_267),
.B(n_268),
.C(n_272),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_270),
.B(n_271),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_269),
.B(n_270),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_271),
.A2(n_305),
.B1(n_306),
.B2(n_307),
.Y(n_304)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_271),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_SL g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

AOI21xp33_ASAP7_75t_L g347 ( 
.A1(n_278),
.A2(n_348),
.B(n_349),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_309),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_279),
.B(n_309),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_297),
.C(n_308),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_280),
.B(n_330),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_281),
.B(n_296),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_289),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_282),
.B(n_289),
.C(n_296),
.Y(n_326)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_286),
.B1(n_287),
.B2(n_288),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_285),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_286),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_295),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_291),
.A2(n_292),
.B1(n_293),
.B2(n_294),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_292),
.B(n_293),
.C(n_295),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_294),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_297),
.A2(n_298),
.B1(n_308),
.B2(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_SL g298 ( 
.A(n_299),
.B(n_304),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_299),
.B(n_305),
.C(n_307),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_300),
.B(n_301),
.Y(n_299)
);

CKINVDCx14_ASAP7_75t_R g303 ( 
.A(n_302),
.Y(n_303)
);

CKINVDCx14_ASAP7_75t_R g306 ( 
.A(n_305),
.Y(n_306)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_308),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_326),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_318),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_311),
.B(n_318),
.C(n_326),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_315),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_312),
.B(n_316),
.C(n_317),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_SL g318 ( 
.A(n_319),
.B(n_320),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_319),
.B(n_321),
.C(n_322),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_322),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_329),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_328),
.B(n_329),
.Y(n_348)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g346 ( 
.A1(n_333),
.A2(n_347),
.B(n_350),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_335),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_334),
.B(n_335),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_341),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_338),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_337),
.B(n_338),
.C(n_341),
.Y(n_343)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_344),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_343),
.B(n_344),
.Y(n_351)
);


endmodule