module real_jpeg_15527_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_0),
.A2(n_50),
.B1(n_55),
.B2(n_56),
.Y(n_49)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_0),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_0),
.A2(n_55),
.B1(n_161),
.B2(n_165),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_1),
.A2(n_15),
.B(n_425),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_1),
.B(n_426),
.Y(n_425)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_2),
.Y(n_87)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_2),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_2),
.Y(n_95)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_2),
.Y(n_99)
);

BUFx5_ASAP7_75t_L g170 ( 
.A(n_3),
.Y(n_170)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_3),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_3),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_3),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_4),
.A2(n_76),
.B1(n_79),
.B2(n_80),
.Y(n_75)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_4),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_4),
.A2(n_79),
.B1(n_138),
.B2(n_139),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_4),
.A2(n_79),
.B1(n_278),
.B2(n_300),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_L g335 ( 
.A1(n_4),
.A2(n_79),
.B1(n_336),
.B2(n_339),
.Y(n_335)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_5),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_5),
.Y(n_69)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_6),
.Y(n_426)
);

INVx2_ASAP7_75t_SL g25 ( 
.A(n_7),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_7),
.B(n_103),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_7),
.A2(n_25),
.B1(n_147),
.B2(n_150),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_7),
.A2(n_25),
.B1(n_202),
.B2(n_204),
.Y(n_201)
);

OAI32xp33_ASAP7_75t_L g310 ( 
.A1(n_7),
.A2(n_311),
.A3(n_314),
.B1(n_317),
.B2(n_321),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_7),
.B(n_93),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_7),
.B(n_356),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_7),
.B(n_168),
.Y(n_365)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_8),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_8),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_8),
.Y(n_164)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_8),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_8),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_8),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_8),
.Y(n_279)
);

BUFx5_ASAP7_75t_L g301 ( 
.A(n_8),
.Y(n_301)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_9),
.B(n_71),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_9),
.A2(n_111),
.B1(n_115),
.B2(n_116),
.Y(n_110)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_9),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_9),
.A2(n_115),
.B1(n_181),
.B2(n_182),
.Y(n_180)
);

OAI22xp33_ASAP7_75t_L g242 ( 
.A1(n_9),
.A2(n_45),
.B1(n_115),
.B2(n_243),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_10),
.Y(n_122)
);

BUFx5_ASAP7_75t_L g124 ( 
.A(n_10),
.Y(n_124)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_10),
.Y(n_131)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_10),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_12),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_12),
.Y(n_57)
);

BUFx4f_ASAP7_75t_L g72 ( 
.A(n_12),
.Y(n_72)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_12),
.Y(n_153)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_13),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_400),
.Y(n_15)
);

AOI21xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_262),
.B(n_396),
.Y(n_16)
);

INVxp33_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_246),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_19),
.B(n_399),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_227),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g397 ( 
.A(n_20),
.B(n_227),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_142),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_21),
.B(n_143),
.C(n_403),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_73),
.C(n_107),
.Y(n_21)
);

XOR2x1_ASAP7_75t_SL g229 ( 
.A(n_22),
.B(n_230),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_48),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_23),
.B(n_48),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_30),
.B1(n_40),
.B2(n_44),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_26),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_25),
.B(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_25),
.B(n_106),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_25),
.A2(n_40),
.B(n_238),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_R g256 ( 
.A(n_25),
.B(n_120),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_25),
.B(n_318),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OA22x2_ASAP7_75t_L g120 ( 
.A1(n_28),
.A2(n_121),
.B1(n_123),
.B2(n_124),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_29),
.Y(n_78)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_29),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_29),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_29),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_36),
.Y(n_30)
);

INVx2_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_35),
.Y(n_114)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_42),
.Y(n_136)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_46),
.A2(n_86),
.B1(n_88),
.B2(n_91),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_58),
.B(n_61),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_49),
.A2(n_63),
.B(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g316 ( 
.A(n_54),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_57),
.Y(n_171)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_57),
.Y(n_177)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_57),
.Y(n_338)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_59),
.Y(n_216)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_60),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_61),
.B(n_369),
.Y(n_368)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_62),
.A2(n_145),
.B(n_154),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_70),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_63),
.B(n_146),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_63),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_63),
.B(n_335),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_66),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_66),
.Y(n_333)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_69),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_70),
.A2(n_212),
.B(n_215),
.Y(n_211)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_72),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_73),
.A2(n_107),
.B1(n_108),
.B2(n_231),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_73),
.Y(n_231)
);

AND2x4_ASAP7_75t_SL g73 ( 
.A(n_74),
.B(n_100),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_74),
.B(n_255),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_84),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_75),
.B(n_93),
.Y(n_240)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_78),
.Y(n_123)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_SL g223 ( 
.A(n_84),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_84),
.B(n_242),
.Y(n_241)
);

NOR2x1_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_93),
.Y(n_84)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_89),
.Y(n_283)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_89),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_91),
.Y(n_274)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_92),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_93),
.B(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_93),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_93),
.B(n_242),
.Y(n_255)
);

AO22x2_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_96),
.B1(n_97),
.B2(n_98),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_96),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_101),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_105),
.Y(n_101)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_104),
.Y(n_244)
);

OAI32xp33_ASAP7_75t_L g270 ( 
.A1(n_105),
.A2(n_271),
.A3(n_275),
.B1(n_280),
.B2(n_284),
.Y(n_270)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_125),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_119),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_110),
.B(n_126),
.Y(n_220)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_112),
.A2(n_128),
.B1(n_132),
.B2(n_136),
.Y(n_127)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx2_ASAP7_75t_L g238 ( 
.A(n_113),
.Y(n_238)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_114),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_115),
.B(n_214),
.Y(n_213)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx3_ASAP7_75t_SL g138 ( 
.A(n_118),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_119),
.B(n_137),
.Y(n_219)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_120),
.B(n_127),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_120),
.A2(n_417),
.B1(n_418),
.B2(n_419),
.Y(n_416)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_126),
.B(n_137),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_126),
.B(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_126),
.Y(n_418)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_137),
.Y(n_417)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_197),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_158),
.Y(n_143)
);

AOI21x1_ASAP7_75t_SL g420 ( 
.A1(n_144),
.A2(n_159),
.B(n_178),
.Y(n_420)
);

OA21x2_ASAP7_75t_L g290 ( 
.A1(n_145),
.A2(n_291),
.B(n_293),
.Y(n_290)
);

AO21x1_ASAP7_75t_L g331 ( 
.A1(n_145),
.A2(n_332),
.B(n_334),
.Y(n_331)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_149),
.Y(n_320)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_151),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx3_ASAP7_75t_L g354 ( 
.A(n_152),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_153),
.Y(n_342)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx4_ASAP7_75t_SL g155 ( 
.A(n_156),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_156),
.Y(n_292)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_156),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_178),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_160),
.B(n_168),
.Y(n_159)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_160),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

BUFx2_ASAP7_75t_L g181 ( 
.A(n_162),
.Y(n_181)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_164),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_164),
.Y(n_189)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_168),
.B(n_180),
.Y(n_208)
);

OA21x2_ASAP7_75t_L g234 ( 
.A1(n_168),
.A2(n_186),
.B(n_201),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_168),
.B(n_201),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_168),
.B(n_299),
.Y(n_329)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

AND2x2_ASAP7_75t_SL g186 ( 
.A(n_169),
.B(n_187),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_171),
.B1(n_172),
.B2(n_176),
.Y(n_169)
);

OAI22xp33_ASAP7_75t_L g187 ( 
.A1(n_172),
.A2(n_188),
.B1(n_190),
.B2(n_193),
.Y(n_187)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_179),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_179),
.B(n_380),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_186),
.Y(n_179)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_186),
.B(n_201),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_186),
.B(n_299),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_186),
.Y(n_411)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx8_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_196),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_197),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_217),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_198),
.B(n_221),
.C(n_226),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_209),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_199),
.B(n_209),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_200),
.B(n_208),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_200),
.B(n_329),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

BUFx12f_ASAP7_75t_L g289 ( 
.A(n_207),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_208),
.B(n_298),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g409 ( 
.A1(n_208),
.A2(n_410),
.B(n_411),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_211),
.B(n_259),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g364 ( 
.A(n_211),
.B(n_334),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_221),
.B1(n_222),
.B2(n_226),
.Y(n_217)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_218),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_219),
.B(n_236),
.Y(n_235)
);

INVx2_ASAP7_75t_SL g221 ( 
.A(n_222),
.Y(n_221)
);

AOI21x1_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_224),
.B(n_225),
.Y(n_222)
);

NOR2x1_ASAP7_75t_L g384 ( 
.A(n_223),
.B(n_225),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_232),
.C(n_245),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_229),
.B(n_261),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_232),
.B(n_245),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_235),
.C(n_239),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_233),
.A2(n_234),
.B1(n_239),
.B2(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_235),
.B(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_237),
.Y(n_419)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_239),
.Y(n_250)
);

AND2x4_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_240),
.B(n_383),
.Y(n_382)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_260),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_247),
.B(n_260),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_251),
.C(n_252),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_248),
.B(n_303),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_251),
.A2(n_252),
.B1(n_253),
.B2(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_251),
.Y(n_304)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_256),
.C(n_257),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_254),
.B(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_255),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_256),
.A2(n_257),
.B1(n_258),
.B2(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_256),
.Y(n_268)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g358 ( 
.A(n_259),
.B(n_359),
.Y(n_358)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_305),
.B(n_395),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_302),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_265),
.B(n_302),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_269),
.C(n_294),
.Y(n_265)
);

XOR2x1_ASAP7_75t_L g390 ( 
.A(n_266),
.B(n_391),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_269),
.A2(n_294),
.B1(n_295),
.B2(n_392),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_269),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_290),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_270),
.A2(n_290),
.B1(n_386),
.B2(n_387),
.Y(n_385)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_270),
.Y(n_387)
);

INVx1_ASAP7_75t_SL g271 ( 
.A(n_272),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_278),
.Y(n_313)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_288),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_290),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_290),
.A2(n_386),
.B1(n_408),
.B2(n_409),
.Y(n_407)
);

BUFx3_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_298),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

AOI21x1_ASAP7_75t_SL g305 ( 
.A1(n_306),
.A2(n_389),
.B(n_394),
.Y(n_305)
);

OAI21x1_ASAP7_75t_L g306 ( 
.A1(n_307),
.A2(n_373),
.B(n_388),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_308),
.A2(n_348),
.B(n_372),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_330),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_309),
.B(n_330),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_328),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_310),
.B(n_328),
.Y(n_370)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

BUFx3_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

BUFx3_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_325),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx5_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

BUFx2_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_329),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_343),
.Y(n_330)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_331),
.Y(n_375)
);

BUFx2_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_335),
.B(n_360),
.Y(n_359)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_344),
.A2(n_345),
.B1(n_346),
.B2(n_347),
.Y(n_343)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_344),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_345),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_345),
.B(n_346),
.C(n_375),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_L g348 ( 
.A1(n_349),
.A2(n_367),
.B(n_371),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_350),
.A2(n_363),
.B(n_366),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_358),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_355),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_359),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_364),
.B(n_365),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_364),
.B(n_365),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_370),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_368),
.B(n_370),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_376),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_374),
.B(n_376),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_385),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_378),
.A2(n_379),
.B1(n_381),
.B2(n_382),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_378),
.B(n_382),
.C(n_385),
.Y(n_393)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

NOR2xp67_ASAP7_75t_SL g414 ( 
.A(n_384),
.B(n_415),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_390),
.B(n_393),
.Y(n_389)
);

NOR2xp67_ASAP7_75t_L g394 ( 
.A(n_390),
.B(n_393),
.Y(n_394)
);

NAND2xp33_ASAP7_75t_R g396 ( 
.A(n_397),
.B(n_398),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_423),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_404),
.Y(n_401)
);

OR2x2_ASAP7_75t_L g424 ( 
.A(n_402),
.B(n_404),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_406),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_407),
.A2(n_412),
.B1(n_421),
.B2(n_422),
.Y(n_406)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_407),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_412),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_413),
.B(n_420),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_416),
.Y(n_413)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);


endmodule