module fake_jpeg_24174_n_191 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_191);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_191;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_15),
.B(n_0),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_34),
.B(n_3),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_38),
.B(n_42),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_40),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_17),
.B(n_1),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_45),
.Y(n_46)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_28),
.Y(n_58)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_44),
.A2(n_30),
.B1(n_31),
.B2(n_4),
.Y(n_65)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_18),
.C(n_15),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_48),
.B(n_53),
.C(n_10),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_17),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_49),
.B(n_51),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_45),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_SL g53 ( 
.A1(n_38),
.A2(n_23),
.B(n_21),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_26),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_54),
.B(n_56),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_44),
.A2(n_21),
.B1(n_23),
.B2(n_22),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_55),
.A2(n_64),
.B1(n_66),
.B2(n_9),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_32),
.B(n_29),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_43),
.A2(n_22),
.B1(n_29),
.B2(n_24),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_57),
.A2(n_60),
.B1(n_62),
.B2(n_5),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_58),
.B(n_9),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_43),
.A2(n_24),
.B1(n_19),
.B2(n_25),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_32),
.A2(n_26),
.B1(n_25),
.B2(n_28),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_40),
.A2(n_16),
.B1(n_31),
.B2(n_30),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_40),
.A2(n_30),
.B1(n_3),
.B2(n_5),
.Y(n_66)
);

BUFx12_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_67),
.B(n_74),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_33),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_68),
.B(n_70),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_39),
.B(n_2),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_39),
.B(n_2),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_71),
.B(n_72),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_35),
.B(n_2),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_73),
.B(n_30),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_35),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_76),
.B(n_82),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_73),
.B(n_37),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_77),
.B(n_78),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_73),
.B(n_37),
.Y(n_78)
);

AND2x4_ASAP7_75t_L g79 ( 
.A(n_53),
.B(n_3),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_79),
.A2(n_95),
.B(n_52),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_81),
.A2(n_88),
.B1(n_62),
.B2(n_63),
.Y(n_110)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

A2O1A1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_46),
.A2(n_6),
.B(n_7),
.C(n_8),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_84),
.B(n_72),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_61),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_85),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_48),
.B(n_7),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_86),
.B(n_94),
.C(n_70),
.Y(n_113)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_93),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_89),
.B(n_99),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_51),
.B(n_10),
.Y(n_91)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_91),
.Y(n_112)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_57),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_58),
.B(n_10),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_54),
.B(n_11),
.Y(n_96)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_49),
.B(n_71),
.Y(n_97)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_47),
.B(n_46),
.Y(n_99)
);

INVxp33_ASAP7_75t_L g100 ( 
.A(n_50),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_100),
.B(n_63),
.Y(n_104)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_101),
.B(n_103),
.Y(n_126)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_104),
.B(n_105),
.Y(n_131)
);

NAND3xp33_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_47),
.C(n_59),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_75),
.B(n_69),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_106),
.B(n_122),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_93),
.A2(n_66),
.B1(n_64),
.B2(n_63),
.Y(n_107)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_107),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_79),
.B(n_74),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_108),
.B(n_89),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_110),
.B(n_88),
.Y(n_125)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_79),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_111),
.B(n_118),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_SL g128 ( 
.A(n_113),
.B(n_98),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_82),
.A2(n_68),
.B1(n_59),
.B2(n_61),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_120),
.B(n_83),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_121),
.A2(n_79),
.B(n_77),
.Y(n_124)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_75),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_116),
.B(n_99),
.C(n_95),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_123),
.B(n_113),
.C(n_119),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_124),
.B(n_128),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_125),
.A2(n_107),
.B1(n_103),
.B2(n_115),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_111),
.A2(n_80),
.B(n_78),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_127),
.A2(n_130),
.B(n_137),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_101),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_129),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_121),
.A2(n_80),
.B(n_92),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_115),
.A2(n_76),
.B(n_98),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_135),
.A2(n_139),
.B(n_140),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_102),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_136),
.B(n_138),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_108),
.A2(n_92),
.B(n_84),
.Y(n_137)
);

BUFx12_ASAP7_75t_L g138 ( 
.A(n_108),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_122),
.B(n_83),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_141),
.B(n_119),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_142),
.B(n_152),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_145),
.B(n_123),
.C(n_128),
.Y(n_161)
);

INVx2_ASAP7_75t_SL g148 ( 
.A(n_129),
.Y(n_148)
);

AO221x1_ASAP7_75t_L g165 ( 
.A1(n_148),
.A2(n_155),
.B1(n_89),
.B2(n_94),
.C(n_129),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_130),
.A2(n_127),
.B(n_137),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_149),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_132),
.A2(n_103),
.B1(n_81),
.B2(n_116),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_150),
.A2(n_125),
.B1(n_141),
.B2(n_139),
.Y(n_164)
);

NAND3xp33_ASAP7_75t_L g152 ( 
.A(n_140),
.B(n_117),
.C(n_112),
.Y(n_152)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_153),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_133),
.A2(n_120),
.B(n_109),
.Y(n_154)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_154),
.Y(n_159)
);

NAND4xp25_ASAP7_75t_L g155 ( 
.A(n_136),
.B(n_118),
.C(n_109),
.D(n_86),
.Y(n_155)
);

A2O1A1O1Ixp25_ASAP7_75t_L g157 ( 
.A1(n_151),
.A2(n_124),
.B(n_126),
.C(n_138),
.D(n_135),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g170 ( 
.A(n_157),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_161),
.B(n_162),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_145),
.B(n_138),
.C(n_132),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_147),
.B(n_138),
.C(n_131),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_163),
.B(n_143),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_164),
.A2(n_165),
.B1(n_153),
.B2(n_147),
.Y(n_167)
);

A2O1A1O1Ixp25_ASAP7_75t_L g166 ( 
.A1(n_151),
.A2(n_134),
.B(n_94),
.C(n_117),
.D(n_112),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g174 ( 
.A(n_166),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_167),
.A2(n_168),
.B(n_172),
.Y(n_177)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_164),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_159),
.B(n_146),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_169),
.B(n_162),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_158),
.B(n_143),
.Y(n_173)
);

OAI21xp33_ASAP7_75t_L g178 ( 
.A1(n_173),
.A2(n_175),
.B(n_174),
.Y(n_178)
);

A2O1A1Ixp33_ASAP7_75t_SL g175 ( 
.A1(n_160),
.A2(n_156),
.B(n_157),
.C(n_163),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_175),
.A2(n_166),
.B(n_161),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_176),
.B(n_181),
.Y(n_183)
);

OR2x2_ASAP7_75t_L g185 ( 
.A(n_178),
.B(n_180),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_179),
.B(n_170),
.C(n_171),
.Y(n_182)
);

NAND2xp33_ASAP7_75t_SL g180 ( 
.A(n_175),
.B(n_150),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_173),
.A2(n_134),
.B(n_114),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_182),
.A2(n_144),
.B(n_114),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_177),
.B(n_148),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_184),
.B(n_52),
.Y(n_188)
);

AO221x1_ASAP7_75t_L g186 ( 
.A1(n_185),
.A2(n_148),
.B1(n_144),
.B2(n_175),
.C(n_52),
.Y(n_186)
);

AOI31xp33_ASAP7_75t_L g189 ( 
.A1(n_186),
.A2(n_67),
.A3(n_183),
.B(n_165),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_187),
.B(n_188),
.C(n_67),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_189),
.B(n_190),
.Y(n_191)
);


endmodule