module fake_jpeg_281_n_517 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_517);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_517;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_331;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_SL g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_1),
.B(n_5),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_2),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_13),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_15),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_45),
.B(n_56),
.Y(n_115)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_46),
.Y(n_101)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_47),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_22),
.B(n_14),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_48),
.B(n_53),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_49),
.Y(n_154)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g145 ( 
.A(n_50),
.Y(n_145)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx11_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_52),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_22),
.B(n_0),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_54),
.Y(n_121)
);

BUFx12_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx6_ASAP7_75t_SL g114 ( 
.A(n_55),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_22),
.Y(n_56)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_57),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_58),
.Y(n_148)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_59),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_34),
.B(n_7),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_60),
.B(n_61),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_14),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_62),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_63),
.Y(n_116)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_64),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_16),
.B(n_7),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_65),
.B(n_71),
.Y(n_150)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_66),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_39),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_67),
.B(n_74),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_68),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_69),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_70),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_16),
.B(n_6),
.Y(n_71)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx11_ASAP7_75t_L g136 ( 
.A(n_72),
.Y(n_136)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_21),
.Y(n_73)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_73),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_42),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_42),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_75),
.B(n_85),
.Y(n_137)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_76),
.Y(n_127)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_77),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_78),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_17),
.B(n_6),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_79),
.B(n_82),
.Y(n_152)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_33),
.Y(n_80)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_80),
.Y(n_149)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_33),
.Y(n_81)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_81),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_44),
.B(n_0),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_40),
.Y(n_83)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_83),
.Y(n_155)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_18),
.Y(n_84)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_84),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_17),
.B(n_6),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_21),
.Y(n_86)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_86),
.Y(n_156)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_21),
.Y(n_87)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_18),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_88),
.B(n_92),
.Y(n_142)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_40),
.Y(n_89)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_89),
.Y(n_157)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_35),
.Y(n_90)
);

BUFx5_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_19),
.B(n_6),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_91),
.B(n_28),
.Y(n_112)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_18),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_32),
.Y(n_93)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

INVx3_ASAP7_75t_SL g94 ( 
.A(n_35),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g147 ( 
.A(n_94),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_19),
.B(n_8),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_95),
.B(n_98),
.Y(n_146)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_35),
.Y(n_96)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_96),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_35),
.Y(n_97)
);

BUFx2_ASAP7_75t_R g106 ( 
.A(n_97),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_35),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_53),
.B(n_36),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_100),
.B(n_135),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_112),
.B(n_117),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_95),
.B(n_30),
.Y(n_117)
);

A2O1A1Ixp33_ASAP7_75t_L g119 ( 
.A1(n_82),
.A2(n_30),
.B(n_28),
.C(n_37),
.Y(n_119)
);

AOI21xp33_ASAP7_75t_L g169 ( 
.A1(n_119),
.A2(n_41),
.B(n_20),
.Y(n_169)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_81),
.B(n_38),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_122),
.B(n_123),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_70),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_50),
.A2(n_38),
.B1(n_24),
.B2(n_27),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_126),
.A2(n_32),
.B1(n_29),
.B2(n_27),
.Y(n_165)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_93),
.Y(n_130)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_130),
.Y(n_164)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_62),
.Y(n_131)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_131),
.Y(n_168)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_52),
.B(n_38),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_133),
.B(n_143),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_89),
.B(n_25),
.Y(n_135)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_64),
.Y(n_138)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_138),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_46),
.A2(n_37),
.B1(n_25),
.B2(n_24),
.Y(n_140)
);

AO22x1_ASAP7_75t_SL g166 ( 
.A1(n_140),
.A2(n_29),
.B1(n_27),
.B2(n_68),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_78),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_76),
.B(n_35),
.C(n_29),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_144),
.B(n_41),
.Y(n_198)
);

CKINVDCx12_ASAP7_75t_R g158 ( 
.A(n_55),
.Y(n_158)
);

CKINVDCx12_ASAP7_75t_R g161 ( 
.A(n_158),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_94),
.B(n_24),
.Y(n_159)
);

OAI21xp33_ASAP7_75t_L g187 ( 
.A1(n_159),
.A2(n_0),
.B(n_1),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_100),
.B(n_32),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_160),
.B(n_188),
.Y(n_223)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_111),
.Y(n_162)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_162),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_122),
.B(n_50),
.Y(n_163)
);

NAND2x1_ASAP7_75t_L g221 ( 
.A(n_163),
.B(n_177),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_165),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_166),
.A2(n_178),
.B1(n_181),
.B2(n_145),
.Y(n_214)
);

AOI21xp33_ASAP7_75t_L g230 ( 
.A1(n_169),
.A2(n_176),
.B(n_187),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_140),
.A2(n_73),
.B1(n_86),
.B2(n_51),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_171),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_133),
.Y(n_174)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_174),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_142),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_175),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_115),
.B(n_137),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_135),
.B(n_96),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_152),
.A2(n_57),
.B1(n_66),
.B2(n_87),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_109),
.A2(n_69),
.B1(n_63),
.B2(n_58),
.Y(n_179)
);

OAI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_179),
.A2(n_195),
.B1(n_200),
.B2(n_202),
.Y(n_210)
);

INVx6_ASAP7_75t_L g180 ( 
.A(n_148),
.Y(n_180)
);

BUFx2_ASAP7_75t_L g219 ( 
.A(n_180),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_144),
.A2(n_49),
.B1(n_86),
.B2(n_83),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_127),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_182),
.Y(n_218)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_129),
.Y(n_183)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_183),
.Y(n_207)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_129),
.Y(n_184)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_184),
.Y(n_209)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_148),
.Y(n_185)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_185),
.Y(n_212)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_145),
.Y(n_186)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_186),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_113),
.B(n_1),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_119),
.B(n_90),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_189),
.B(n_193),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_150),
.B(n_77),
.Y(n_190)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_190),
.Y(n_208)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_99),
.Y(n_191)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_191),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_116),
.Y(n_192)
);

INVx6_ASAP7_75t_L g215 ( 
.A(n_192),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_118),
.B(n_97),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_146),
.A2(n_72),
.B1(n_90),
.B2(n_97),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_194),
.A2(n_199),
.B1(n_205),
.B2(n_114),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_110),
.A2(n_20),
.B1(n_41),
.B2(n_4),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_127),
.Y(n_196)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_196),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_125),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_197),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_198),
.B(n_154),
.C(n_156),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_121),
.B(n_139),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_153),
.A2(n_20),
.B1(n_3),
.B2(n_4),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_147),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_105),
.Y(n_203)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_203),
.Y(n_234)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_149),
.Y(n_204)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_204),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_114),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_128),
.Y(n_206)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_206),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_189),
.A2(n_124),
.B1(n_151),
.B2(n_102),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_213),
.A2(n_220),
.B1(n_226),
.B2(n_232),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_214),
.B(n_231),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_217),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_163),
.A2(n_157),
.B1(n_108),
.B2(n_120),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_163),
.A2(n_157),
.B1(n_108),
.B2(n_120),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_227),
.B(n_198),
.Y(n_244)
);

AND2x4_ASAP7_75t_L g231 ( 
.A(n_177),
.B(n_99),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_172),
.A2(n_170),
.B1(n_181),
.B2(n_177),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_178),
.A2(n_151),
.B1(n_102),
.B2(n_101),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_233),
.A2(n_240),
.B1(n_214),
.B2(n_126),
.Y(n_262)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_186),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_237),
.Y(n_261)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_183),
.Y(n_239)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_239),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_174),
.A2(n_101),
.B1(n_107),
.B2(n_132),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_244),
.B(n_269),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_241),
.B(n_175),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_245),
.B(n_249),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_218),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_247),
.B(n_253),
.Y(n_289)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_238),
.Y(n_248)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_248),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_223),
.B(n_188),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_238),
.Y(n_250)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_250),
.Y(n_286)
);

OAI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_225),
.A2(n_160),
.B1(n_166),
.B2(n_205),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_251),
.A2(n_263),
.B1(n_248),
.B2(n_250),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_223),
.B(n_201),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_252),
.B(n_259),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_225),
.Y(n_253)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_207),
.Y(n_255)
);

INVx2_ASAP7_75t_SL g279 ( 
.A(n_255),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_231),
.B(n_166),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_256),
.B(n_262),
.Y(n_300)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_222),
.Y(n_257)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_257),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_208),
.B(n_167),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_258),
.B(n_263),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_229),
.B(n_197),
.Y(n_259)
);

OR2x2_ASAP7_75t_L g260 ( 
.A(n_224),
.B(n_201),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_260),
.A2(n_164),
.B(n_235),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_213),
.B(n_167),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_236),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_264),
.B(n_267),
.Y(n_294)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_207),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_265),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_224),
.B(n_202),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_222),
.Y(n_268)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_268),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_227),
.B(n_166),
.Y(n_269)
);

AND2x6_ASAP7_75t_L g270 ( 
.A(n_230),
.B(n_204),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_270),
.Y(n_293)
);

OAI22xp33_ASAP7_75t_L g271 ( 
.A1(n_228),
.A2(n_185),
.B1(n_180),
.B2(n_132),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_271),
.A2(n_262),
.B1(n_219),
.B2(n_256),
.Y(n_281)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_234),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_272),
.Y(n_290)
);

MAJx2_ASAP7_75t_L g273 ( 
.A(n_244),
.B(n_221),
.C(n_231),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g303 ( 
.A(n_273),
.B(n_260),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_269),
.A2(n_233),
.B1(n_211),
.B2(n_228),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_274),
.A2(n_275),
.B1(n_277),
.B2(n_265),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_266),
.A2(n_211),
.B1(n_240),
.B2(n_210),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_266),
.A2(n_221),
.B1(n_231),
.B2(n_234),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_281),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_243),
.A2(n_221),
.B(n_242),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_284),
.B(n_260),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_244),
.B(n_161),
.C(n_162),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_285),
.B(n_291),
.C(n_297),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_266),
.A2(n_242),
.B1(n_219),
.B2(n_212),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_287),
.A2(n_288),
.B1(n_247),
.B2(n_268),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_266),
.A2(n_212),
.B1(n_192),
.B2(n_216),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_252),
.B(n_161),
.C(n_203),
.Y(n_291)
);

OAI22x1_ASAP7_75t_L g295 ( 
.A1(n_256),
.A2(n_270),
.B1(n_267),
.B2(n_259),
.Y(n_295)
);

OAI22x1_ASAP7_75t_L g328 ( 
.A1(n_295),
.A2(n_296),
.B1(n_287),
.B2(n_281),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_246),
.A2(n_235),
.B(n_216),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_249),
.B(n_206),
.Y(n_297)
);

OR2x2_ASAP7_75t_L g331 ( 
.A(n_299),
.B(n_302),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_303),
.B(n_321),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_304),
.B(n_329),
.Y(n_353)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_279),
.Y(n_305)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_305),
.Y(n_335)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_279),
.Y(n_306)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_306),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_283),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_307),
.B(n_314),
.Y(n_342)
);

INVx4_ASAP7_75t_L g309 ( 
.A(n_279),
.Y(n_309)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_309),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_282),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_310),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_298),
.B(n_258),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g349 ( 
.A(n_311),
.B(n_323),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_289),
.B(n_298),
.Y(n_312)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_312),
.Y(n_346)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_282),
.Y(n_313)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_313),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_294),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_283),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_315),
.B(n_320),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_316),
.A2(n_277),
.B(n_302),
.Y(n_345)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_286),
.Y(n_317)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_317),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_299),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_318),
.B(n_322),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_290),
.Y(n_320)
);

XOR2x2_ASAP7_75t_L g321 ( 
.A(n_278),
.B(n_270),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_286),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_280),
.B(n_245),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_278),
.B(n_272),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_324),
.B(n_330),
.C(n_301),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_SL g325 ( 
.A(n_280),
.B(n_257),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_325),
.B(n_301),
.Y(n_356)
);

INVx6_ASAP7_75t_SL g326 ( 
.A(n_295),
.Y(n_326)
);

CKINVDCx14_ASAP7_75t_R g364 ( 
.A(n_326),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_276),
.B(n_237),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g363 ( 
.A(n_327),
.B(n_261),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_328),
.A2(n_300),
.B(n_284),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_273),
.B(n_164),
.C(n_196),
.Y(n_330)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_292),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_332),
.B(n_333),
.Y(n_358)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_292),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_324),
.B(n_285),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_334),
.B(n_339),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_312),
.B(n_297),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_SL g368 ( 
.A(n_337),
.B(n_344),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_308),
.B(n_291),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g387 ( 
.A1(n_341),
.A2(n_355),
.B(n_261),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_325),
.B(n_293),
.Y(n_344)
);

AO21x1_ASAP7_75t_L g371 ( 
.A1(n_345),
.A2(n_347),
.B(n_362),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_331),
.A2(n_300),
.B(n_293),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_310),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_348),
.B(n_309),
.Y(n_372)
);

CKINVDCx16_ASAP7_75t_R g350 ( 
.A(n_331),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_350),
.B(n_363),
.Y(n_365)
);

AOI21xp5_ASAP7_75t_L g355 ( 
.A1(n_326),
.A2(n_328),
.B(n_300),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_SL g380 ( 
.A(n_356),
.B(n_305),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_357),
.B(n_360),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_321),
.B(n_274),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_329),
.A2(n_288),
.B1(n_290),
.B2(n_296),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_361),
.A2(n_261),
.B1(n_254),
.B2(n_236),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_318),
.A2(n_275),
.B(n_255),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_349),
.B(n_308),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_SL g395 ( 
.A(n_366),
.B(n_391),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_339),
.B(n_330),
.C(n_303),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_367),
.B(n_369),
.C(n_393),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_357),
.B(n_319),
.C(n_332),
.Y(n_369)
);

FAx1_ASAP7_75t_SL g370 ( 
.A(n_354),
.B(n_304),
.CI(n_322),
.CON(n_370),
.SN(n_370)
);

FAx1_ASAP7_75t_SL g419 ( 
.A(n_370),
.B(n_367),
.CI(n_393),
.CON(n_419),
.SN(n_419)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_372),
.B(n_385),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_358),
.B(n_333),
.Y(n_373)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_373),
.Y(n_397)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_336),
.Y(n_374)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_374),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_358),
.B(n_313),
.Y(n_375)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_375),
.Y(n_411)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_351),
.Y(n_376)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_376),
.Y(n_413)
);

CKINVDCx16_ASAP7_75t_R g377 ( 
.A(n_342),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_377),
.B(n_378),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_351),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_353),
.A2(n_319),
.B1(n_317),
.B2(n_306),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_379),
.A2(n_384),
.B1(n_389),
.B2(n_361),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_380),
.B(n_386),
.Y(n_407)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_352),
.Y(n_382)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_382),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_340),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_334),
.B(n_254),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_387),
.A2(n_392),
.B(n_362),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_340),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_388),
.B(n_348),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_353),
.A2(n_192),
.B1(n_209),
.B2(n_239),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_364),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_390),
.B(n_374),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_346),
.B(n_209),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_SL g392 ( 
.A1(n_341),
.A2(n_141),
.B(n_155),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_360),
.B(n_191),
.C(n_141),
.Y(n_393)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_396),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_372),
.Y(n_398)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_398),
.Y(n_422)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_399),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_L g400 ( 
.A1(n_371),
.A2(n_355),
.B(n_347),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_400),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_381),
.B(n_354),
.C(n_356),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_401),
.B(n_404),
.Y(n_426)
);

INVxp33_ASAP7_75t_L g428 ( 
.A(n_403),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_369),
.B(n_346),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_368),
.B(n_359),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_405),
.B(n_415),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_386),
.B(n_345),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_408),
.B(n_412),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_409),
.A2(n_378),
.B1(n_376),
.B2(n_365),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_381),
.B(n_353),
.Y(n_412)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_373),
.Y(n_415)
);

A2O1A1Ixp33_ASAP7_75t_SL g416 ( 
.A1(n_387),
.A2(n_343),
.B(n_338),
.C(n_359),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_L g440 ( 
.A1(n_416),
.A2(n_419),
.B(n_370),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_383),
.B(n_343),
.C(n_338),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_417),
.B(n_418),
.Y(n_424)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_375),
.Y(n_418)
);

CKINVDCx16_ASAP7_75t_R g421 ( 
.A(n_406),
.Y(n_421)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_421),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_423),
.A2(n_403),
.B1(n_416),
.B2(n_352),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_417),
.B(n_371),
.Y(n_425)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_425),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_410),
.A2(n_409),
.B1(n_397),
.B2(n_411),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_429),
.A2(n_430),
.B1(n_155),
.B2(n_107),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_413),
.A2(n_384),
.B1(n_389),
.B2(n_388),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_401),
.B(n_383),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_431),
.B(n_433),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_412),
.B(n_380),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_408),
.B(n_379),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_434),
.B(n_437),
.Y(n_455)
);

BUFx24_ASAP7_75t_SL g436 ( 
.A(n_395),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_SL g451 ( 
.A(n_436),
.B(n_442),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_407),
.B(n_392),
.Y(n_437)
);

AOI322xp5_ASAP7_75t_L g439 ( 
.A1(n_402),
.A2(n_398),
.A3(n_385),
.B1(n_400),
.B2(n_414),
.C1(n_382),
.C2(n_416),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_439),
.B(n_441),
.Y(n_446)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_440),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_407),
.B(n_370),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_402),
.Y(n_442)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_445),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_435),
.A2(n_416),
.B1(n_394),
.B2(n_419),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_447),
.A2(n_435),
.B1(n_441),
.B2(n_437),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_424),
.B(n_394),
.C(n_419),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_449),
.B(n_450),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_438),
.B(n_335),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_425),
.B(n_335),
.C(n_184),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_452),
.B(n_454),
.Y(n_467)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_453),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_434),
.B(n_156),
.C(n_168),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_427),
.A2(n_215),
.B1(n_185),
.B2(n_180),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_456),
.B(n_461),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_431),
.B(n_168),
.C(n_154),
.Y(n_457)
);

HB1xp67_ASAP7_75t_L g477 ( 
.A(n_457),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_420),
.B(n_215),
.Y(n_458)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_458),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_426),
.B(n_173),
.C(n_136),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_460),
.B(n_432),
.C(n_433),
.Y(n_462)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_422),
.Y(n_461)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_462),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_SL g463 ( 
.A1(n_446),
.A2(n_448),
.B(n_447),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_463),
.B(n_464),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_449),
.B(n_432),
.C(n_428),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_451),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_465),
.B(n_472),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_468),
.B(n_473),
.Y(n_487)
);

MAJx2_ASAP7_75t_L g469 ( 
.A(n_459),
.B(n_428),
.C(n_173),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_469),
.B(n_106),
.C(n_103),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_445),
.A2(n_134),
.B1(n_116),
.B2(n_136),
.Y(n_471)
);

INVxp67_ASAP7_75t_L g478 ( 
.A(n_471),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_455),
.B(n_134),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_455),
.B(n_103),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_SL g479 ( 
.A(n_476),
.B(n_444),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_479),
.B(n_482),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_464),
.B(n_474),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_SL g497 ( 
.A(n_480),
.B(n_486),
.Y(n_497)
);

NAND4xp25_ASAP7_75t_SL g482 ( 
.A(n_477),
.B(n_452),
.C(n_460),
.D(n_454),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_L g483 ( 
.A1(n_466),
.A2(n_457),
.B1(n_443),
.B2(n_104),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_483),
.B(n_488),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_475),
.B(n_443),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_470),
.B(n_462),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g500 ( 
.A(n_489),
.B(n_55),
.Y(n_500)
);

CKINVDCx16_ASAP7_75t_R g490 ( 
.A(n_467),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_490),
.A2(n_106),
.B1(n_3),
.B2(n_4),
.Y(n_495)
);

AOI21xp5_ASAP7_75t_L g492 ( 
.A1(n_481),
.A2(n_473),
.B(n_469),
.Y(n_492)
);

AOI21x1_ASAP7_75t_L g503 ( 
.A1(n_492),
.A2(n_499),
.B(n_478),
.Y(n_503)
);

A2O1A1Ixp33_ASAP7_75t_L g494 ( 
.A1(n_484),
.A2(n_472),
.B(n_471),
.C(n_104),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_494),
.B(n_500),
.Y(n_504)
);

OAI21xp5_ASAP7_75t_SL g506 ( 
.A1(n_495),
.A2(n_13),
.B(n_8),
.Y(n_506)
);

INVxp33_ASAP7_75t_SL g496 ( 
.A(n_485),
.Y(n_496)
);

AOI22xp33_ASAP7_75t_SL g505 ( 
.A1(n_496),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_505)
);

INVx6_ASAP7_75t_L g498 ( 
.A(n_482),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_498),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_487),
.A2(n_10),
.B(n_3),
.Y(n_499)
);

AOI21xp5_ASAP7_75t_SL g502 ( 
.A1(n_497),
.A2(n_487),
.B(n_478),
.Y(n_502)
);

AOI21xp5_ASAP7_75t_L g508 ( 
.A1(n_502),
.A2(n_505),
.B(n_506),
.Y(n_508)
);

INVxp67_ASAP7_75t_L g511 ( 
.A(n_503),
.Y(n_511)
);

INVxp67_ASAP7_75t_L g507 ( 
.A(n_497),
.Y(n_507)
);

AO22x1_ASAP7_75t_L g510 ( 
.A1(n_507),
.A2(n_9),
.B1(n_11),
.B2(n_13),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_501),
.B(n_491),
.C(n_493),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_509),
.B(n_510),
.Y(n_512)
);

INVxp67_ASAP7_75t_L g513 ( 
.A(n_511),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_513),
.B(n_504),
.C(n_508),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_514),
.Y(n_515)
);

AOI211xp5_ASAP7_75t_L g516 ( 
.A1(n_515),
.A2(n_2),
.B(n_512),
.C(n_501),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g517 ( 
.A(n_516),
.B(n_2),
.Y(n_517)
);


endmodule