module fake_jpeg_1934_n_129 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_129);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_129;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_122;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_10),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_10),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

INVx13_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx5_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_15),
.B(n_27),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_28),
.B(n_41),
.Y(n_55)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_30),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_33),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_20),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_34),
.B(n_35),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_39),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

HB1xp67_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_25),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_42),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_43),
.Y(n_60)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_44),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

BUFx24_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_48),
.A2(n_50),
.B1(n_52),
.B2(n_18),
.Y(n_64)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_51),
.Y(n_69)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

INVx3_ASAP7_75t_SL g51 ( 
.A(n_11),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_54),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_14),
.B(n_4),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

A2O1A1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_40),
.A2(n_22),
.B(n_18),
.C(n_4),
.Y(n_66)
);

A2O1A1O1Ixp25_ASAP7_75t_L g83 ( 
.A1(n_66),
.A2(n_37),
.B(n_47),
.C(n_39),
.D(n_50),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g67 ( 
.A1(n_42),
.A2(n_51),
.B(n_43),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_29),
.Y(n_79)
);

AO22x1_ASAP7_75t_SL g70 ( 
.A1(n_39),
.A2(n_22),
.B1(n_1),
.B2(n_3),
.Y(n_70)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_30),
.A2(n_1),
.B1(n_3),
.B2(n_45),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_74),
.A2(n_76),
.B1(n_47),
.B2(n_62),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_30),
.A2(n_3),
.B1(n_45),
.B2(n_46),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_69),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_77),
.B(n_81),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_79),
.A2(n_83),
.B(n_86),
.Y(n_100)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_71),
.B(n_52),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_52),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_82),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_66),
.B(n_31),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_90),
.Y(n_99)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_60),
.A2(n_67),
.B1(n_70),
.B2(n_72),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_88),
.A2(n_61),
.B1(n_63),
.B2(n_70),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_55),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_89),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_62),
.B(n_63),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_91),
.B(n_63),
.C(n_59),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_85),
.C(n_81),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_95),
.A2(n_97),
.B1(n_101),
.B2(n_90),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_78),
.A2(n_61),
.B1(n_56),
.B2(n_58),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_78),
.A2(n_88),
.B1(n_84),
.B2(n_79),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_102),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_103),
.Y(n_113)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_98),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_106),
.Y(n_112)
);

OA21x2_ASAP7_75t_L g115 ( 
.A1(n_105),
.A2(n_97),
.B(n_100),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_96),
.B(n_92),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_77),
.Y(n_107)
);

OAI321xp33_ASAP7_75t_L g111 ( 
.A1(n_107),
.A2(n_110),
.A3(n_101),
.B1(n_83),
.B2(n_100),
.C(n_95),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_108),
.B(n_109),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_82),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_99),
.B(n_80),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_111),
.B(n_94),
.Y(n_119)
);

OAI21xp33_ASAP7_75t_L g117 ( 
.A1(n_115),
.A2(n_105),
.B(n_110),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_114),
.B(n_108),
.C(n_109),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_116),
.B(n_114),
.C(n_113),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_117),
.B(n_119),
.Y(n_122)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_112),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_118),
.B(n_115),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_120),
.B(n_121),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_122),
.A2(n_117),
.B1(n_87),
.B2(n_65),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_124),
.A2(n_65),
.B1(n_75),
.B2(n_57),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_123),
.B(n_56),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_125),
.B(n_126),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_57),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_75),
.Y(n_129)
);


endmodule