module fake_jpeg_3578_n_121 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_121);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_121;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_25),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_28),
.Y(n_36)
);

INVx6_ASAP7_75t_SL g37 ( 
.A(n_4),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g41 ( 
.A1(n_24),
.A2(n_10),
.B(n_6),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

BUFx8_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_38),
.B(n_0),
.Y(n_48)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_41),
.Y(n_56)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_0),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_50),
.B(n_43),
.Y(n_55)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

AND2x2_ASAP7_75t_SL g57 ( 
.A(n_51),
.B(n_39),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_47),
.A2(n_41),
.B(n_44),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_55),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_57),
.Y(n_63)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_49),
.A2(n_37),
.B1(n_44),
.B2(n_34),
.Y(n_60)
);

BUFx24_ASAP7_75t_L g64 ( 
.A(n_60),
.Y(n_64)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_62),
.Y(n_84)
);

AO22x1_ASAP7_75t_SL g65 ( 
.A1(n_57),
.A2(n_51),
.B1(n_34),
.B2(n_42),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_67),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_61),
.B(n_33),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_66),
.B(n_1),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_61),
.A2(n_36),
.B1(n_2),
.B2(n_3),
.Y(n_67)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

AO22x1_ASAP7_75t_SL g69 ( 
.A1(n_60),
.A2(n_42),
.B1(n_13),
.B2(n_14),
.Y(n_69)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_73),
.B(n_12),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_79),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_70),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_SL g87 ( 
.A(n_75),
.B(n_76),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_70),
.B(n_54),
.C(n_42),
.Y(n_76)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_1),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_16),
.C(n_29),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_SL g92 ( 
.A(n_81),
.B(n_68),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_64),
.A2(n_2),
.B(n_4),
.Y(n_85)
);

OAI21xp33_ASAP7_75t_L g94 ( 
.A1(n_85),
.A2(n_5),
.B(n_6),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_89),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_71),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_69),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_90),
.A2(n_93),
.B(n_94),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_72),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_92),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_64),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_5),
.Y(n_95)
);

AOI322xp5_ASAP7_75t_SL g106 ( 
.A1(n_95),
.A2(n_8),
.A3(n_10),
.B1(n_11),
.B2(n_19),
.C1(n_22),
.C2(n_31),
.Y(n_106)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_97),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_7),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_98),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_93),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_100),
.A2(n_94),
.B1(n_101),
.B2(n_86),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_21),
.C(n_26),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_103),
.B(n_105),
.C(n_101),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_20),
.C(n_23),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_106),
.B(n_108),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_96),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_109),
.B(n_110),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_107),
.Y(n_112)
);

NOR2xp67_ASAP7_75t_SL g114 ( 
.A(n_112),
.B(n_113),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_102),
.B(n_99),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_115),
.A2(n_112),
.B(n_104),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_116),
.B(n_114),
.C(n_103),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_105),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_118),
.Y(n_119)
);

BUFx24_ASAP7_75t_SL g120 ( 
.A(n_119),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_111),
.Y(n_121)
);


endmodule