module fake_jpeg_21225_n_129 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_129);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_129;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_6),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g16 ( 
.A(n_5),
.B(n_9),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_2),
.B(n_5),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_12),
.B(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_30),
.B(n_37),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_34),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_16),
.B(n_1),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_36),
.Y(n_38)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_37),
.A2(n_23),
.B1(n_25),
.B2(n_24),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_39),
.A2(n_46),
.B1(n_50),
.B2(n_19),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_29),
.B(n_23),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_36),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_28),
.A2(n_25),
.B1(n_24),
.B2(n_20),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_30),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_15),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_35),
.A2(n_20),
.B1(n_15),
.B2(n_13),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_51),
.B(n_61),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_16),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_52),
.B(n_58),
.Y(n_73)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_55),
.B(n_57),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_56),
.B(n_62),
.Y(n_81)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_46),
.B(n_34),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_59),
.A2(n_36),
.B1(n_33),
.B2(n_32),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_13),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_60),
.B(n_67),
.Y(n_78)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_31),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_65),
.C(n_71),
.Y(n_82)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVxp33_ASAP7_75t_SL g75 ( 
.A(n_64),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_31),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_70),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_27),
.Y(n_67)
);

NOR2x1_ASAP7_75t_L g68 ( 
.A(n_38),
.B(n_26),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_68),
.B(n_69),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_21),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_38),
.B(n_17),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_41),
.B(n_31),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_26),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_72),
.A2(n_17),
.B(n_7),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_76),
.A2(n_72),
.B(n_68),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_SL g77 ( 
.A(n_56),
.B(n_17),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_63),
.C(n_62),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_33),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_65),
.C(n_61),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_85),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_87),
.Y(n_89)
);

AO221x1_ASAP7_75t_L g104 ( 
.A1(n_89),
.A2(n_80),
.B1(n_86),
.B2(n_82),
.C(n_10),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_63),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_90),
.B(n_96),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_71),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_94),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_92),
.A2(n_95),
.B(n_76),
.Y(n_102)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_84),
.Y(n_93)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_93),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_65),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_78),
.B(n_66),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_97),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_32),
.C(n_29),
.Y(n_98)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_98),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_88),
.A2(n_75),
.B1(n_86),
.B2(n_79),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_101),
.A2(n_88),
.B1(n_98),
.B2(n_74),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_102),
.B(n_55),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_104),
.B(n_4),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_103),
.B(n_95),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_107),
.B(n_112),
.C(n_113),
.Y(n_116)
);

XNOR2x1_ASAP7_75t_L g108 ( 
.A(n_99),
.B(n_96),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_108),
.A2(n_109),
.B(n_102),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_101),
.B(n_82),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_110),
.A2(n_111),
.B1(n_106),
.B2(n_100),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_103),
.B(n_83),
.C(n_54),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_114),
.Y(n_122)
);

BUFx5_ASAP7_75t_L g115 ( 
.A(n_108),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_115),
.B(n_118),
.Y(n_119)
);

AOI221xp5_ASAP7_75t_L g121 ( 
.A1(n_117),
.A2(n_74),
.B1(n_7),
.B2(n_8),
.C(n_11),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_107),
.B(n_105),
.C(n_100),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_116),
.B(n_109),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_120),
.B(n_121),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_119),
.B(n_4),
.Y(n_123)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_123),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_122),
.B(n_8),
.Y(n_124)
);

OAI21xp33_ASAP7_75t_L g127 ( 
.A1(n_124),
.A2(n_11),
.B(n_12),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_127),
.B(n_125),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_126),
.Y(n_129)
);


endmodule