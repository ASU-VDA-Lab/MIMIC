module fake_jpeg_10477_n_203 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_203);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_203;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx8_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx8_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_38),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_18),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_35),
.A2(n_22),
.B1(n_17),
.B2(n_29),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_20),
.B(n_27),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_28),
.Y(n_52)
);

BUFx8_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_41),
.Y(n_61)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_44),
.Y(n_55)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_0),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_35),
.A2(n_18),
.B1(n_27),
.B2(n_25),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_47),
.A2(n_29),
.B1(n_32),
.B2(n_24),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_1),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_49),
.B(n_64),
.Y(n_83)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_60),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_62),
.Y(n_67)
);

OA22x2_ASAP7_75t_L g53 ( 
.A1(n_41),
.A2(n_42),
.B1(n_28),
.B2(n_25),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_53),
.A2(n_57),
.B1(n_38),
.B2(n_31),
.Y(n_73)
);

O2A1O1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_54),
.A2(n_58),
.B(n_32),
.C(n_23),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_21),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_56),
.B(n_59),
.Y(n_91)
);

OA22x2_ASAP7_75t_L g57 ( 
.A1(n_42),
.A2(n_22),
.B1(n_32),
.B2(n_24),
.Y(n_57)
);

NAND2xp33_ASAP7_75t_SL g58 ( 
.A(n_34),
.B(n_2),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_21),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_31),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_37),
.B(n_33),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_37),
.B(n_17),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_55),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_47),
.A2(n_38),
.B1(n_34),
.B2(n_33),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_66),
.A2(n_76),
.B1(n_60),
.B2(n_4),
.Y(n_114)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_68),
.B(n_70),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_52),
.B(n_56),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_69),
.B(n_77),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_60),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_30),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_72),
.B(n_82),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_73),
.Y(n_94)
);

CKINVDCx10_ASAP7_75t_R g74 ( 
.A(n_60),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_74),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_75),
.A2(n_50),
.B1(n_45),
.B2(n_19),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_77),
.B(n_78),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_10),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_12),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_79),
.B(n_81),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_46),
.B(n_3),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_59),
.B(n_21),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_54),
.B(n_32),
.C(n_23),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_93),
.C(n_57),
.Y(n_97)
);

INVx13_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_85),
.B(n_86),
.Y(n_113)
);

INVx13_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_48),
.B(n_3),
.Y(n_87)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_53),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_90),
.B(n_92),
.Y(n_110)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_58),
.B(n_23),
.C(n_19),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_97),
.B(n_93),
.Y(n_122)
);

AND2x2_ASAP7_75t_SL g98 ( 
.A(n_91),
.B(n_49),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_98),
.B(n_100),
.C(n_83),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_91),
.B(n_57),
.C(n_48),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_71),
.Y(n_101)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_105),
.B(n_108),
.Y(n_129)
);

OA22x2_ASAP7_75t_L g106 ( 
.A1(n_92),
.A2(n_51),
.B1(n_45),
.B2(n_49),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_106),
.A2(n_76),
.B1(n_90),
.B2(n_89),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_74),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_107),
.B(n_85),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_69),
.B(n_63),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_67),
.B(n_63),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_SL g133 ( 
.A(n_109),
.B(n_81),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_111),
.A2(n_114),
.B1(n_88),
.B2(n_84),
.Y(n_125)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_96),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_116),
.B(n_119),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_117),
.A2(n_136),
.B(n_110),
.Y(n_143)
);

OAI221xp5_ASAP7_75t_L g118 ( 
.A1(n_105),
.A2(n_73),
.B1(n_83),
.B2(n_66),
.C(n_67),
.Y(n_118)
);

BUFx24_ASAP7_75t_SL g141 ( 
.A(n_118),
.Y(n_141)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_108),
.Y(n_119)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_109),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_121),
.B(n_123),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_122),
.B(n_130),
.C(n_132),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_68),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_124),
.B(n_126),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_125),
.B(n_127),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_95),
.B(n_78),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_113),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_99),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_128),
.B(n_131),
.Y(n_139)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_95),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_100),
.B(n_70),
.C(n_83),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_133),
.B(n_134),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_97),
.B(n_79),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_106),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_135),
.B(n_110),
.Y(n_142)
);

XNOR2x2_ASAP7_75t_L g136 ( 
.A(n_98),
.B(n_81),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_142),
.B(n_144),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_143),
.A2(n_154),
.B(n_3),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_125),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_136),
.A2(n_135),
.B(n_130),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_145),
.A2(n_103),
.B(n_106),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_119),
.B(n_98),
.Y(n_146)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_146),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_129),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_147),
.B(n_151),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_129),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_120),
.B(n_102),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_152),
.B(n_153),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_134),
.B(n_98),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_133),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_138),
.B(n_122),
.C(n_132),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_155),
.B(n_162),
.C(n_164),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_144),
.A2(n_94),
.B1(n_115),
.B2(n_104),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_157),
.A2(n_159),
.B1(n_163),
.B2(n_168),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_150),
.A2(n_94),
.B1(n_115),
.B2(n_104),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_138),
.B(n_117),
.C(n_114),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_148),
.A2(n_120),
.B1(n_106),
.B2(n_101),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_153),
.B(n_112),
.C(n_103),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_165),
.B(n_143),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_140),
.B(n_112),
.C(n_107),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_166),
.B(n_146),
.C(n_86),
.Y(n_177)
);

AO21x1_ASAP7_75t_L g179 ( 
.A1(n_167),
.A2(n_4),
.B(n_5),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_154),
.A2(n_80),
.B1(n_85),
.B2(n_86),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_169),
.B(n_170),
.C(n_172),
.Y(n_182)
);

MAJx2_ASAP7_75t_L g170 ( 
.A(n_156),
.B(n_145),
.C(n_140),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_166),
.B(n_141),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_160),
.B(n_137),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_173),
.B(n_177),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_159),
.B(n_139),
.Y(n_174)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_174),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_168),
.A2(n_149),
.B1(n_151),
.B2(n_147),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_175),
.A2(n_164),
.B(n_155),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_158),
.B(n_80),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_178),
.B(n_157),
.Y(n_181)
);

NOR3xp33_ASAP7_75t_L g187 ( 
.A(n_179),
.B(n_7),
.C(n_8),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_181),
.B(n_186),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_177),
.A2(n_161),
.B(n_162),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_183),
.A2(n_176),
.B(n_171),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_184),
.B(n_187),
.Y(n_191)
);

AOI31xp67_ASAP7_75t_L g186 ( 
.A1(n_179),
.A2(n_6),
.A3(n_7),
.B(n_8),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_182),
.B(n_176),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_189),
.B(n_190),
.C(n_180),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_185),
.B(n_169),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_192),
.B(n_193),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_187),
.B(n_14),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_194),
.B(n_195),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_189),
.B(n_170),
.Y(n_195)
);

BUFx4f_ASAP7_75t_SL g196 ( 
.A(n_191),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_196),
.A2(n_188),
.B(n_14),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_198),
.B(n_200),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_197),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_199),
.A2(n_197),
.B(n_7),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_202),
.A2(n_8),
.B(n_201),
.Y(n_203)
);


endmodule