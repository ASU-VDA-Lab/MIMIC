module fake_netlist_1_2213_n_888 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_204, n_221, n_185, n_22, n_203, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_9, n_161, n_10, n_177, n_130, n_189, n_103, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_181, n_101, n_62, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_16, n_13, n_198, n_169, n_193, n_152, n_113, n_95, n_124, n_156, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_197, n_201, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_191, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_205, n_12, n_86, n_143, n_213, n_182, n_166, n_162, n_186, n_75, n_163, n_105, n_159, n_174, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_92, n_11, n_223, n_25, n_30, n_59, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_66, n_134, n_222, n_1, n_164, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_224, n_96, n_225, n_39, n_888);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_204;
input n_221;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_181;
input n_101;
input n_62;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_152;
input n_113;
input n_95;
input n_124;
input n_156;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_197;
input n_201;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_191;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_182;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_105;
input n_159;
input n_174;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_92;
input n_11;
input n_223;
input n_25;
input n_30;
input n_59;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_222;
input n_1;
input n_164;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_224;
input n_96;
input n_225;
input n_39;
output n_888;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_838;
wire n_705;
wire n_603;
wire n_604;
wire n_858;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_848;
wire n_607;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_667;
wire n_496;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_878;
wire n_814;
wire n_637;
wire n_817;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_288;
wire n_383;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_787;
wire n_853;
wire n_296;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_462;
wire n_232;
wire n_316;
wire n_545;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_789;
wire n_330;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_434;
wire n_384;
wire n_227;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_752;
wire n_732;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_857;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_479;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_567;
wire n_809;
wire n_580;
wire n_502;
wire n_543;
wire n_854;
wire n_455;
wire n_312;
wire n_529;
wire n_880;
wire n_630;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_865;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_255;
wire n_426;
wire n_624;
wire n_769;
wire n_725;
wire n_818;
wire n_844;
wire n_230;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_506;
wire n_533;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_708;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_501;
wire n_248;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_876;
wire n_886;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_466;
wire n_302;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_788;
wire n_475;
wire n_578;
wire n_542;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_450;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_446;
wire n_420;
wire n_285;
wire n_423;
wire n_342;
wire n_621;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_874;
wire n_388;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_823;
wire n_822;
wire n_390;
wire n_682;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_881;
wire n_260;
wire n_806;
wire n_539;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_265;
wire n_522;
wire n_264;
wire n_883;
wire n_573;
wire n_673;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_861;
wire n_295;
wire n_654;
wire n_263;
wire n_495;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_577;
wire n_870;
wire n_790;
wire n_761;
wire n_615;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_835;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_267;
wire n_456;
wire n_782;
wire n_449;
wire n_300;
wire n_734;
wire n_524;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_240;
wire n_841;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_306;
wire n_242;
wire n_766;
wire n_602;
wire n_831;
wire n_859;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_837;
wire n_410;
wire n_774;
wire n_867;
wire n_377;
wire n_510;
wire n_343;
wire n_675;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_493;
wire n_418;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_266;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_845;
wire n_713;
wire n_457;
wire n_595;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_781;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g226 ( .A(n_30), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_95), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_56), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_24), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_221), .Y(n_230) );
CKINVDCx5p33_ASAP7_75t_R g231 ( .A(n_147), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_160), .Y(n_232) );
INVxp33_ASAP7_75t_SL g233 ( .A(n_222), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_2), .Y(n_234) );
CKINVDCx20_ASAP7_75t_R g235 ( .A(n_126), .Y(n_235) );
CKINVDCx14_ASAP7_75t_R g236 ( .A(n_58), .Y(n_236) );
BUFx6f_ASAP7_75t_L g237 ( .A(n_213), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_8), .Y(n_238) );
BUFx6f_ASAP7_75t_L g239 ( .A(n_71), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_191), .Y(n_240) );
CKINVDCx5p33_ASAP7_75t_R g241 ( .A(n_39), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_220), .Y(n_242) );
HB1xp67_ASAP7_75t_L g243 ( .A(n_125), .Y(n_243) );
INVxp67_ASAP7_75t_L g244 ( .A(n_67), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_73), .Y(n_245) );
INVxp33_ASAP7_75t_SL g246 ( .A(n_41), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_190), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_117), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_60), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_175), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_210), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_163), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_208), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_112), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_143), .Y(n_255) );
INVx3_ASAP7_75t_L g256 ( .A(n_128), .Y(n_256) );
CKINVDCx20_ASAP7_75t_R g257 ( .A(n_145), .Y(n_257) );
CKINVDCx16_ASAP7_75t_R g258 ( .A(n_9), .Y(n_258) );
INVx2_ASAP7_75t_L g259 ( .A(n_7), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_198), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_184), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_14), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_193), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_177), .Y(n_264) );
INVxp67_ASAP7_75t_L g265 ( .A(n_114), .Y(n_265) );
INVxp67_ASAP7_75t_SL g266 ( .A(n_94), .Y(n_266) );
CKINVDCx16_ASAP7_75t_R g267 ( .A(n_102), .Y(n_267) );
INVxp33_ASAP7_75t_SL g268 ( .A(n_148), .Y(n_268) );
INVxp67_ASAP7_75t_L g269 ( .A(n_155), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_121), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_224), .Y(n_271) );
INVxp33_ASAP7_75t_SL g272 ( .A(n_166), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_139), .Y(n_273) );
INVx1_ASAP7_75t_SL g274 ( .A(n_98), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_120), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_87), .Y(n_276) );
CKINVDCx5p33_ASAP7_75t_R g277 ( .A(n_153), .Y(n_277) );
CKINVDCx5p33_ASAP7_75t_R g278 ( .A(n_186), .Y(n_278) );
HB1xp67_ASAP7_75t_L g279 ( .A(n_129), .Y(n_279) );
BUFx6f_ASAP7_75t_L g280 ( .A(n_3), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_109), .Y(n_281) );
CKINVDCx5p33_ASAP7_75t_R g282 ( .A(n_169), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_176), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_131), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_212), .Y(n_285) );
CKINVDCx5p33_ASAP7_75t_R g286 ( .A(n_35), .Y(n_286) );
CKINVDCx5p33_ASAP7_75t_R g287 ( .A(n_56), .Y(n_287) );
CKINVDCx5p33_ASAP7_75t_R g288 ( .A(n_49), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_66), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_51), .Y(n_290) );
CKINVDCx5p33_ASAP7_75t_R g291 ( .A(n_12), .Y(n_291) );
INVxp33_ASAP7_75t_SL g292 ( .A(n_24), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_30), .Y(n_293) );
BUFx2_ASAP7_75t_L g294 ( .A(n_81), .Y(n_294) );
BUFx3_ASAP7_75t_L g295 ( .A(n_158), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_13), .Y(n_296) );
INVxp67_ASAP7_75t_SL g297 ( .A(n_188), .Y(n_297) );
HB1xp67_ASAP7_75t_L g298 ( .A(n_110), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_4), .Y(n_299) );
INVxp33_ASAP7_75t_L g300 ( .A(n_72), .Y(n_300) );
CKINVDCx14_ASAP7_75t_R g301 ( .A(n_200), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_54), .Y(n_302) );
BUFx3_ASAP7_75t_L g303 ( .A(n_182), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_93), .Y(n_304) );
CKINVDCx16_ASAP7_75t_R g305 ( .A(n_34), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_194), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_40), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_20), .Y(n_308) );
BUFx3_ASAP7_75t_L g309 ( .A(n_171), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_167), .Y(n_310) );
CKINVDCx5p33_ASAP7_75t_R g311 ( .A(n_204), .Y(n_311) );
INVxp67_ASAP7_75t_SL g312 ( .A(n_218), .Y(n_312) );
BUFx3_ASAP7_75t_L g313 ( .A(n_43), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_215), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_80), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_107), .Y(n_316) );
INVxp67_ASAP7_75t_L g317 ( .A(n_135), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_142), .Y(n_318) );
INVxp67_ASAP7_75t_SL g319 ( .A(n_165), .Y(n_319) );
CKINVDCx5p33_ASAP7_75t_R g320 ( .A(n_63), .Y(n_320) );
CKINVDCx16_ASAP7_75t_R g321 ( .A(n_4), .Y(n_321) );
BUFx3_ASAP7_75t_L g322 ( .A(n_170), .Y(n_322) );
BUFx6f_ASAP7_75t_SL g323 ( .A(n_219), .Y(n_323) );
CKINVDCx5p33_ASAP7_75t_R g324 ( .A(n_65), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_62), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_214), .B(n_130), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_211), .Y(n_327) );
BUFx3_ASAP7_75t_L g328 ( .A(n_150), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_82), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_67), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_185), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_50), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_123), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_59), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_55), .Y(n_335) );
INVxp67_ASAP7_75t_SL g336 ( .A(n_124), .Y(n_336) );
NOR2xp67_ASAP7_75t_L g337 ( .A(n_33), .B(n_183), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_25), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_181), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_19), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_206), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_179), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_225), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_240), .Y(n_344) );
AND2x4_ASAP7_75t_L g345 ( .A(n_256), .B(n_0), .Y(n_345) );
NAND2xp5_ASAP7_75t_SL g346 ( .A(n_256), .B(n_0), .Y(n_346) );
NOR2xp33_ASAP7_75t_L g347 ( .A(n_243), .B(n_1), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_294), .B(n_1), .Y(n_348) );
BUFx6f_ASAP7_75t_L g349 ( .A(n_237), .Y(n_349) );
BUFx6f_ASAP7_75t_L g350 ( .A(n_237), .Y(n_350) );
CKINVDCx16_ASAP7_75t_R g351 ( .A(n_267), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_237), .Y(n_352) );
BUFx6f_ASAP7_75t_L g353 ( .A(n_237), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_240), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_242), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_237), .Y(n_356) );
OAI22xp5_ASAP7_75t_SL g357 ( .A1(n_258), .A2(n_5), .B1(n_2), .B2(n_3), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_294), .B(n_5), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_242), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_256), .Y(n_360) );
INVxp67_ASAP7_75t_L g361 ( .A(n_279), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_247), .Y(n_362) );
INVx3_ASAP7_75t_L g363 ( .A(n_239), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_247), .Y(n_364) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_236), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_300), .B(n_6), .Y(n_366) );
INVx2_ASAP7_75t_L g367 ( .A(n_254), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_248), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_248), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_298), .B(n_6), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_238), .B(n_7), .Y(n_371) );
CKINVDCx5p33_ASAP7_75t_R g372 ( .A(n_301), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_250), .Y(n_373) );
BUFx6f_ASAP7_75t_L g374 ( .A(n_295), .Y(n_374) );
OAI21x1_ASAP7_75t_L g375 ( .A1(n_254), .A2(n_85), .B(n_84), .Y(n_375) );
BUFx6f_ASAP7_75t_L g376 ( .A(n_295), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_273), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_238), .B(n_8), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_245), .B(n_9), .Y(n_379) );
NAND2xp5_ASAP7_75t_SL g380 ( .A(n_345), .B(n_273), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_361), .B(n_313), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_360), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_360), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_359), .B(n_327), .Y(n_384) );
AOI22xp5_ASAP7_75t_L g385 ( .A1(n_358), .A2(n_292), .B1(n_246), .B2(n_305), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_360), .Y(n_386) );
BUFx10_ASAP7_75t_L g387 ( .A(n_345), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_349), .Y(n_388) );
AND2x6_ASAP7_75t_L g389 ( .A(n_345), .B(n_250), .Y(n_389) );
HB1xp67_ASAP7_75t_L g390 ( .A(n_365), .Y(n_390) );
BUFx6f_ASAP7_75t_L g391 ( .A(n_349), .Y(n_391) );
INVxp67_ASAP7_75t_SL g392 ( .A(n_348), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_345), .Y(n_393) );
OR2x2_ASAP7_75t_L g394 ( .A(n_365), .B(n_321), .Y(n_394) );
INVx1_ASAP7_75t_SL g395 ( .A(n_358), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_345), .Y(n_396) );
CKINVDCx5p33_ASAP7_75t_R g397 ( .A(n_351), .Y(n_397) );
NOR2xp33_ASAP7_75t_L g398 ( .A(n_361), .B(n_265), .Y(n_398) );
INVx3_ASAP7_75t_L g399 ( .A(n_367), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_359), .B(n_327), .Y(n_400) );
INVx3_ASAP7_75t_L g401 ( .A(n_367), .Y(n_401) );
NOR2xp33_ASAP7_75t_L g402 ( .A(n_344), .B(n_269), .Y(n_402) );
HB1xp67_ASAP7_75t_L g403 ( .A(n_366), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_367), .Y(n_404) );
AND2x6_ASAP7_75t_L g405 ( .A(n_358), .B(n_251), .Y(n_405) );
BUFx2_ASAP7_75t_L g406 ( .A(n_372), .Y(n_406) );
INVx5_ASAP7_75t_L g407 ( .A(n_349), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_366), .B(n_313), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_349), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_377), .Y(n_410) );
NOR2xp33_ASAP7_75t_L g411 ( .A(n_354), .B(n_317), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_349), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_366), .B(n_245), .Y(n_413) );
INVx4_ASAP7_75t_L g414 ( .A(n_374), .Y(n_414) );
NAND2xp5_ASAP7_75t_SL g415 ( .A(n_359), .B(n_343), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_377), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g417 ( .A1(n_354), .A2(n_262), .B1(n_330), .B2(n_249), .Y(n_417) );
BUFx6f_ASAP7_75t_L g418 ( .A(n_349), .Y(n_418) );
INVx1_ASAP7_75t_SL g419 ( .A(n_351), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_382), .Y(n_420) );
INVx2_ASAP7_75t_SL g421 ( .A(n_387), .Y(n_421) );
INVx2_ASAP7_75t_SL g422 ( .A(n_387), .Y(n_422) );
BUFx6f_ASAP7_75t_L g423 ( .A(n_387), .Y(n_423) );
INVx3_ASAP7_75t_L g424 ( .A(n_387), .Y(n_424) );
NOR2xp67_ASAP7_75t_L g425 ( .A(n_385), .B(n_372), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_382), .Y(n_426) );
NOR2xp33_ASAP7_75t_L g427 ( .A(n_392), .B(n_370), .Y(n_427) );
OR2x6_ASAP7_75t_L g428 ( .A(n_403), .B(n_357), .Y(n_428) );
NOR2xp33_ASAP7_75t_SL g429 ( .A(n_395), .B(n_235), .Y(n_429) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_392), .B(n_370), .Y(n_430) );
BUFx3_ASAP7_75t_L g431 ( .A(n_389), .Y(n_431) );
BUFx4f_ASAP7_75t_L g432 ( .A(n_405), .Y(n_432) );
INVx5_ASAP7_75t_L g433 ( .A(n_389), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_383), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_398), .B(n_355), .Y(n_435) );
AO22x1_ASAP7_75t_L g436 ( .A1(n_397), .A2(n_292), .B1(n_246), .B2(n_268), .Y(n_436) );
NOR2xp33_ASAP7_75t_L g437 ( .A(n_398), .B(n_362), .Y(n_437) );
NAND2xp5_ASAP7_75t_SL g438 ( .A(n_387), .B(n_362), .Y(n_438) );
OR2x2_ASAP7_75t_L g439 ( .A(n_394), .B(n_348), .Y(n_439) );
NOR2xp33_ASAP7_75t_L g440 ( .A(n_408), .B(n_364), .Y(n_440) );
HB1xp67_ASAP7_75t_L g441 ( .A(n_390), .Y(n_441) );
BUFx3_ASAP7_75t_L g442 ( .A(n_389), .Y(n_442) );
BUFx2_ASAP7_75t_L g443 ( .A(n_405), .Y(n_443) );
INVx5_ASAP7_75t_L g444 ( .A(n_389), .Y(n_444) );
AOI211xp5_ASAP7_75t_L g445 ( .A1(n_385), .A2(n_357), .B(n_347), .C(n_346), .Y(n_445) );
OAI22xp33_ASAP7_75t_L g446 ( .A1(n_395), .A2(n_235), .B1(n_257), .B2(n_241), .Y(n_446) );
AND3x1_ASAP7_75t_SL g447 ( .A(n_394), .B(n_229), .C(n_228), .Y(n_447) );
NOR2xp33_ASAP7_75t_L g448 ( .A(n_408), .B(n_381), .Y(n_448) );
INVx5_ASAP7_75t_L g449 ( .A(n_389), .Y(n_449) );
BUFx8_ASAP7_75t_L g450 ( .A(n_405), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_405), .A2(n_364), .B1(n_369), .B2(n_368), .Y(n_451) );
BUFx2_ASAP7_75t_L g452 ( .A(n_405), .Y(n_452) );
BUFx4f_ASAP7_75t_L g453 ( .A(n_405), .Y(n_453) );
NAND2xp33_ASAP7_75t_SL g454 ( .A(n_393), .B(n_257), .Y(n_454) );
INVx1_ASAP7_75t_SL g455 ( .A(n_419), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_386), .Y(n_456) );
INVx4_ASAP7_75t_L g457 ( .A(n_389), .Y(n_457) );
BUFx3_ASAP7_75t_L g458 ( .A(n_389), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_414), .Y(n_459) );
BUFx6f_ASAP7_75t_SL g460 ( .A(n_405), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_381), .B(n_368), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_414), .Y(n_462) );
BUFx3_ASAP7_75t_L g463 ( .A(n_389), .Y(n_463) );
AND2x4_ASAP7_75t_L g464 ( .A(n_413), .B(n_346), .Y(n_464) );
OR2x6_ASAP7_75t_L g465 ( .A(n_413), .B(n_371), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_404), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_413), .B(n_369), .Y(n_467) );
NAND2xp33_ASAP7_75t_SL g468 ( .A(n_393), .B(n_323), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_414), .Y(n_469) );
AND2x4_ASAP7_75t_L g470 ( .A(n_405), .B(n_347), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_402), .B(n_373), .Y(n_471) );
OAI22xp5_ASAP7_75t_SL g472 ( .A1(n_419), .A2(n_286), .B1(n_287), .B2(n_226), .Y(n_472) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_402), .B(n_373), .Y(n_473) );
OR2x6_ASAP7_75t_L g474 ( .A(n_406), .B(n_378), .Y(n_474) );
AND2x4_ASAP7_75t_SL g475 ( .A(n_396), .B(n_262), .Y(n_475) );
INVx5_ASAP7_75t_L g476 ( .A(n_389), .Y(n_476) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_405), .A2(n_379), .B1(n_268), .B2(n_272), .Y(n_477) );
HB1xp67_ASAP7_75t_L g478 ( .A(n_384), .Y(n_478) );
INVxp67_ASAP7_75t_SL g479 ( .A(n_396), .Y(n_479) );
NAND2xp5_ASAP7_75t_SL g480 ( .A(n_380), .B(n_227), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_410), .Y(n_481) );
HB1xp67_ASAP7_75t_L g482 ( .A(n_478), .Y(n_482) );
INVx2_ASAP7_75t_SL g483 ( .A(n_455), .Y(n_483) );
OAI22xp5_ASAP7_75t_L g484 ( .A1(n_465), .A2(n_380), .B1(n_417), .B2(n_411), .Y(n_484) );
AOI22xp5_ASAP7_75t_L g485 ( .A1(n_427), .A2(n_417), .B1(n_288), .B2(n_291), .Y(n_485) );
A2O1A1Ixp33_ASAP7_75t_L g486 ( .A1(n_473), .A2(n_416), .B(n_410), .C(n_384), .Y(n_486) );
BUFx6f_ASAP7_75t_L g487 ( .A(n_423), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_420), .Y(n_488) );
BUFx6f_ASAP7_75t_L g489 ( .A(n_423), .Y(n_489) );
OAI22xp5_ASAP7_75t_L g490 ( .A1(n_465), .A2(n_400), .B1(n_233), .B2(n_272), .Y(n_490) );
A2O1A1Ixp33_ASAP7_75t_L g491 ( .A1(n_473), .A2(n_416), .B(n_399), .C(n_401), .Y(n_491) );
NAND2xp5_ASAP7_75t_SL g492 ( .A(n_423), .B(n_414), .Y(n_492) );
BUFx6f_ASAP7_75t_L g493 ( .A(n_423), .Y(n_493) );
AOI22xp5_ASAP7_75t_L g494 ( .A1(n_430), .A2(n_288), .B1(n_291), .B2(n_287), .Y(n_494) );
OAI22xp5_ASAP7_75t_L g495 ( .A1(n_465), .A2(n_233), .B1(n_415), .B2(n_401), .Y(n_495) );
NOR2x1_ASAP7_75t_R g496 ( .A(n_429), .B(n_320), .Y(n_496) );
BUFx3_ASAP7_75t_L g497 ( .A(n_441), .Y(n_497) );
AOI22xp33_ASAP7_75t_L g498 ( .A1(n_464), .A2(n_399), .B1(n_401), .B2(n_415), .Y(n_498) );
NOR2x1_ASAP7_75t_L g499 ( .A(n_439), .B(n_474), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_420), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_426), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_426), .Y(n_502) );
BUFx2_ASAP7_75t_L g503 ( .A(n_450), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_434), .Y(n_504) );
BUFx2_ASAP7_75t_L g505 ( .A(n_450), .Y(n_505) );
NOR2xp33_ASAP7_75t_L g506 ( .A(n_448), .B(n_244), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_467), .Y(n_507) );
NOR2xp33_ASAP7_75t_L g508 ( .A(n_448), .B(n_320), .Y(n_508) );
OAI21x1_ASAP7_75t_L g509 ( .A1(n_424), .A2(n_375), .B(n_399), .Y(n_509) );
INVx5_ASAP7_75t_L g510 ( .A(n_457), .Y(n_510) );
BUFx2_ASAP7_75t_L g511 ( .A(n_450), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_464), .A2(n_399), .B1(n_401), .B2(n_377), .Y(n_512) );
INVx2_ASAP7_75t_SL g513 ( .A(n_474), .Y(n_513) );
A2O1A1Ixp33_ASAP7_75t_L g514 ( .A1(n_437), .A2(n_440), .B(n_430), .C(n_471), .Y(n_514) );
BUFx6f_ASAP7_75t_L g515 ( .A(n_431), .Y(n_515) );
OAI21x1_ASAP7_75t_L g516 ( .A1(n_424), .A2(n_375), .B(n_399), .Y(n_516) );
INVx3_ASAP7_75t_L g517 ( .A(n_424), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_475), .Y(n_518) );
INVx6_ASAP7_75t_L g519 ( .A(n_433), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_438), .A2(n_435), .B(n_479), .Y(n_520) );
BUFx8_ASAP7_75t_L g521 ( .A(n_460), .Y(n_521) );
BUFx2_ASAP7_75t_L g522 ( .A(n_474), .Y(n_522) );
INVx5_ASAP7_75t_L g523 ( .A(n_433), .Y(n_523) );
NAND3xp33_ASAP7_75t_L g524 ( .A(n_445), .B(n_324), .C(n_414), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_460), .A2(n_377), .B1(n_332), .B2(n_334), .Y(n_525) );
A2O1A1Ixp33_ASAP7_75t_L g526 ( .A1(n_437), .A2(n_375), .B(n_335), .C(n_338), .Y(n_526) );
AOI21xp33_ASAP7_75t_L g527 ( .A1(n_440), .A2(n_297), .B(n_266), .Y(n_527) );
BUFx2_ASAP7_75t_L g528 ( .A(n_454), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_459), .Y(n_529) );
BUFx12f_ASAP7_75t_L g530 ( .A(n_428), .Y(n_530) );
AOI22xp33_ASAP7_75t_SL g531 ( .A1(n_428), .A2(n_324), .B1(n_340), .B2(n_330), .Y(n_531) );
CKINVDCx11_ASAP7_75t_R g532 ( .A(n_442), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_438), .A2(n_326), .B(n_252), .Y(n_533) );
BUFx6f_ASAP7_75t_L g534 ( .A(n_442), .Y(n_534) );
BUFx6f_ASAP7_75t_L g535 ( .A(n_458), .Y(n_535) );
BUFx6f_ASAP7_75t_SL g536 ( .A(n_470), .Y(n_536) );
OR2x2_ASAP7_75t_L g537 ( .A(n_446), .B(n_340), .Y(n_537) );
AND2x4_ASAP7_75t_L g538 ( .A(n_444), .B(n_234), .Y(n_538) );
BUFx6f_ASAP7_75t_L g539 ( .A(n_458), .Y(n_539) );
OAI22xp5_ASAP7_75t_L g540 ( .A1(n_432), .A2(n_277), .B1(n_278), .B2(n_231), .Y(n_540) );
HB1xp67_ASAP7_75t_L g541 ( .A(n_463), .Y(n_541) );
AND2x6_ASAP7_75t_L g542 ( .A(n_463), .B(n_432), .Y(n_542) );
CKINVDCx5p33_ASAP7_75t_R g543 ( .A(n_472), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_462), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_461), .Y(n_545) );
INVx2_ASAP7_75t_L g546 ( .A(n_469), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_466), .Y(n_547) );
INVx3_ASAP7_75t_L g548 ( .A(n_453), .Y(n_548) );
INVx1_ASAP7_75t_SL g549 ( .A(n_454), .Y(n_549) );
BUFx4f_ASAP7_75t_L g550 ( .A(n_470), .Y(n_550) );
BUFx6f_ASAP7_75t_L g551 ( .A(n_444), .Y(n_551) );
AOI22xp5_ASAP7_75t_L g552 ( .A1(n_447), .A2(n_278), .B1(n_282), .B2(n_277), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_451), .B(n_289), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_477), .B(n_290), .Y(n_554) );
INVx5_ASAP7_75t_L g555 ( .A(n_449), .Y(n_555) );
AND2x6_ASAP7_75t_L g556 ( .A(n_453), .B(n_253), .Y(n_556) );
BUFx6f_ASAP7_75t_L g557 ( .A(n_449), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_481), .Y(n_558) );
AND2x4_ASAP7_75t_L g559 ( .A(n_449), .B(n_293), .Y(n_559) );
BUFx6f_ASAP7_75t_L g560 ( .A(n_476), .Y(n_560) );
AND2x4_ASAP7_75t_L g561 ( .A(n_482), .B(n_443), .Y(n_561) );
AOI22xp33_ASAP7_75t_SL g562 ( .A1(n_522), .A2(n_470), .B1(n_452), .B2(n_436), .Y(n_562) );
O2A1O1Ixp33_ASAP7_75t_L g563 ( .A1(n_514), .A2(n_480), .B(n_425), .C(n_456), .Y(n_563) );
BUFx6f_ASAP7_75t_L g564 ( .A(n_487), .Y(n_564) );
OAI22xp5_ASAP7_75t_L g565 ( .A1(n_514), .A2(n_476), .B1(n_299), .B2(n_302), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_483), .B(n_296), .Y(n_566) );
BUFx6f_ASAP7_75t_L g567 ( .A(n_487), .Y(n_567) );
OR2x6_ASAP7_75t_L g568 ( .A(n_530), .B(n_503), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_531), .A2(n_468), .B1(n_469), .B2(n_421), .Y(n_569) );
A2O1A1Ixp33_ASAP7_75t_L g570 ( .A1(n_520), .A2(n_421), .B(n_422), .C(n_337), .Y(n_570) );
OAI22xp5_ASAP7_75t_L g571 ( .A1(n_486), .A2(n_259), .B1(n_260), .B2(n_255), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_531), .A2(n_422), .B1(n_323), .B2(n_308), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_497), .B(n_307), .Y(n_573) );
OAI22xp5_ASAP7_75t_L g574 ( .A1(n_507), .A2(n_255), .B1(n_261), .B2(n_260), .Y(n_574) );
OAI22xp5_ASAP7_75t_L g575 ( .A1(n_545), .A2(n_261), .B1(n_264), .B2(n_263), .Y(n_575) );
NOR2xp67_ASAP7_75t_L g576 ( .A(n_543), .B(n_10), .Y(n_576) );
BUFx4f_ASAP7_75t_L g577 ( .A(n_505), .Y(n_577) );
AOI22xp5_ASAP7_75t_L g578 ( .A1(n_499), .A2(n_311), .B1(n_282), .B2(n_315), .Y(n_578) );
OAI22xp5_ASAP7_75t_L g579 ( .A1(n_500), .A2(n_263), .B1(n_270), .B2(n_264), .Y(n_579) );
INVx8_ASAP7_75t_L g580 ( .A(n_523), .Y(n_580) );
AND2x4_ASAP7_75t_L g581 ( .A(n_513), .B(n_325), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_536), .A2(n_329), .B1(n_280), .B2(n_239), .Y(n_582) );
CKINVDCx6p67_ASAP7_75t_R g583 ( .A(n_532), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_550), .A2(n_280), .B1(n_239), .B2(n_271), .Y(n_584) );
NAND2x1p5_ASAP7_75t_L g585 ( .A(n_510), .B(n_239), .Y(n_585) );
INVx1_ASAP7_75t_SL g586 ( .A(n_518), .Y(n_586) );
AOI22xp33_ASAP7_75t_SL g587 ( .A1(n_528), .A2(n_311), .B1(n_319), .B2(n_312), .Y(n_587) );
BUFx6f_ASAP7_75t_L g588 ( .A(n_487), .Y(n_588) );
INVx4_ASAP7_75t_L g589 ( .A(n_523), .Y(n_589) );
A2O1A1Ixp33_ASAP7_75t_L g590 ( .A1(n_520), .A2(n_271), .B(n_275), .C(n_270), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_547), .Y(n_591) );
AOI22xp5_ASAP7_75t_L g592 ( .A1(n_490), .A2(n_508), .B1(n_549), .B2(n_484), .Y(n_592) );
OAI22xp33_ASAP7_75t_L g593 ( .A1(n_485), .A2(n_280), .B1(n_239), .B2(n_275), .Y(n_593) );
OAI221xp5_ASAP7_75t_L g594 ( .A1(n_552), .A2(n_336), .B1(n_341), .B2(n_339), .C(n_342), .Y(n_594) );
OAI22xp5_ASAP7_75t_L g595 ( .A1(n_501), .A2(n_331), .B1(n_339), .B2(n_333), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_558), .Y(n_596) );
OAI22xp5_ASAP7_75t_L g597 ( .A1(n_504), .A2(n_333), .B1(n_342), .B2(n_341), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_550), .A2(n_280), .B1(n_230), .B2(n_232), .Y(n_598) );
OAI22xp5_ASAP7_75t_L g599 ( .A1(n_491), .A2(n_524), .B1(n_512), .B2(n_525), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_494), .B(n_10), .Y(n_600) );
NAND2xp5_ASAP7_75t_SL g601 ( .A(n_487), .B(n_274), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_553), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_553), .Y(n_603) );
INVx6_ASAP7_75t_L g604 ( .A(n_521), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_506), .B(n_276), .Y(n_605) );
OAI21xp5_ASAP7_75t_L g606 ( .A1(n_526), .A2(n_283), .B(n_281), .Y(n_606) );
INVx6_ASAP7_75t_L g607 ( .A(n_521), .Y(n_607) );
INVx2_ASAP7_75t_L g608 ( .A(n_488), .Y(n_608) );
AOI21xp33_ASAP7_75t_L g609 ( .A1(n_495), .A2(n_285), .B(n_284), .Y(n_609) );
CKINVDCx11_ASAP7_75t_R g610 ( .A(n_511), .Y(n_610) );
AOI22xp33_ASAP7_75t_SL g611 ( .A1(n_496), .A2(n_556), .B1(n_537), .B2(n_506), .Y(n_611) );
OAI22xp33_ASAP7_75t_L g612 ( .A1(n_554), .A2(n_309), .B1(n_322), .B2(n_303), .Y(n_612) );
O2A1O1Ixp33_ASAP7_75t_SL g613 ( .A1(n_491), .A2(n_526), .B(n_492), .C(n_502), .Y(n_613) );
INVxp67_ASAP7_75t_L g614 ( .A(n_540), .Y(n_614) );
OAI22xp33_ASAP7_75t_L g615 ( .A1(n_510), .A2(n_309), .B1(n_322), .B2(n_303), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_512), .Y(n_616) );
AOI22xp33_ASAP7_75t_L g617 ( .A1(n_527), .A2(n_306), .B1(n_310), .B2(n_304), .Y(n_617) );
OAI22xp5_ASAP7_75t_L g618 ( .A1(n_525), .A2(n_316), .B1(n_318), .B2(n_314), .Y(n_618) );
HB1xp67_ASAP7_75t_L g619 ( .A(n_541), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_538), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_538), .Y(n_621) );
AOI22xp33_ASAP7_75t_L g622 ( .A1(n_556), .A2(n_328), .B1(n_376), .B2(n_374), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_498), .B(n_11), .Y(n_623) );
AOI21xp33_ASAP7_75t_L g624 ( .A1(n_559), .A2(n_376), .B(n_374), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_533), .B(n_374), .Y(n_625) );
AOI221xp5_ASAP7_75t_L g626 ( .A1(n_559), .A2(n_374), .B1(n_376), .B2(n_363), .C(n_356), .Y(n_626) );
OAI22xp5_ASAP7_75t_SL g627 ( .A1(n_510), .A2(n_16), .B1(n_11), .B2(n_15), .Y(n_627) );
INVx2_ASAP7_75t_L g628 ( .A(n_529), .Y(n_628) );
AND2x4_ASAP7_75t_L g629 ( .A(n_510), .B(n_15), .Y(n_629) );
AND2x4_ASAP7_75t_L g630 ( .A(n_548), .B(n_16), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_517), .B(n_17), .Y(n_631) );
BUFx6f_ASAP7_75t_L g632 ( .A(n_489), .Y(n_632) );
OA21x2_ASAP7_75t_L g633 ( .A1(n_509), .A2(n_409), .B(n_388), .Y(n_633) );
INVx2_ASAP7_75t_L g634 ( .A(n_544), .Y(n_634) );
INVx2_ASAP7_75t_L g635 ( .A(n_546), .Y(n_635) );
OR2x2_ASAP7_75t_L g636 ( .A(n_517), .B(n_18), .Y(n_636) );
CKINVDCx5p33_ASAP7_75t_R g637 ( .A(n_523), .Y(n_637) );
AOI22xp5_ASAP7_75t_L g638 ( .A1(n_548), .A2(n_374), .B1(n_376), .B2(n_363), .Y(n_638) );
OAI22xp5_ASAP7_75t_L g639 ( .A1(n_489), .A2(n_376), .B1(n_374), .B2(n_356), .Y(n_639) );
AO21x2_ASAP7_75t_L g640 ( .A1(n_516), .A2(n_356), .B(n_352), .Y(n_640) );
BUFx6f_ASAP7_75t_L g641 ( .A(n_493), .Y(n_641) );
AOI22xp33_ASAP7_75t_L g642 ( .A1(n_611), .A2(n_493), .B1(n_376), .B2(n_374), .Y(n_642) );
OAI21xp33_ASAP7_75t_L g643 ( .A1(n_572), .A2(n_376), .B(n_363), .Y(n_643) );
AND2x2_ASAP7_75t_L g644 ( .A(n_573), .B(n_21), .Y(n_644) );
AOI22xp33_ASAP7_75t_L g645 ( .A1(n_616), .A2(n_542), .B1(n_515), .B2(n_535), .Y(n_645) );
AOI21xp5_ASAP7_75t_L g646 ( .A1(n_613), .A2(n_534), .B(n_515), .Y(n_646) );
AOI22xp33_ASAP7_75t_SL g647 ( .A1(n_627), .A2(n_539), .B1(n_519), .B2(n_560), .Y(n_647) );
AND2x2_ASAP7_75t_L g648 ( .A(n_566), .B(n_22), .Y(n_648) );
OAI22xp5_ASAP7_75t_L g649 ( .A1(n_592), .A2(n_555), .B1(n_519), .B2(n_551), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_591), .Y(n_650) );
AOI21xp33_ASAP7_75t_L g651 ( .A1(n_563), .A2(n_557), .B(n_551), .Y(n_651) );
AOI22xp33_ASAP7_75t_L g652 ( .A1(n_600), .A2(n_352), .B1(n_557), .B2(n_551), .Y(n_652) );
OAI22xp5_ASAP7_75t_L g653 ( .A1(n_569), .A2(n_555), .B1(n_557), .B2(n_560), .Y(n_653) );
AOI221xp5_ASAP7_75t_L g654 ( .A1(n_605), .A2(n_560), .B1(n_557), .B2(n_551), .C(n_349), .Y(n_654) );
AOI221xp5_ASAP7_75t_L g655 ( .A1(n_574), .A2(n_575), .B1(n_571), .B2(n_609), .C(n_594), .Y(n_655) );
NOR2xp33_ASAP7_75t_L g656 ( .A(n_586), .B(n_555), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_596), .Y(n_657) );
INVx2_ASAP7_75t_L g658 ( .A(n_608), .Y(n_658) );
INVxp67_ASAP7_75t_L g659 ( .A(n_630), .Y(n_659) );
OAI22xp5_ASAP7_75t_L g660 ( .A1(n_614), .A2(n_349), .B1(n_350), .B2(n_353), .Y(n_660) );
AND2x4_ASAP7_75t_L g661 ( .A(n_561), .B(n_23), .Y(n_661) );
AND2x2_ASAP7_75t_L g662 ( .A(n_577), .B(n_23), .Y(n_662) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_602), .A2(n_353), .B1(n_350), .B2(n_412), .Y(n_663) );
OAI21x1_ASAP7_75t_L g664 ( .A1(n_633), .A2(n_353), .B(n_350), .Y(n_664) );
BUFx4f_ASAP7_75t_L g665 ( .A(n_604), .Y(n_665) );
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_603), .A2(n_418), .B1(n_391), .B2(n_26), .Y(n_666) );
OAI211xp5_ASAP7_75t_L g667 ( .A1(n_576), .A2(n_587), .B(n_617), .C(n_562), .Y(n_667) );
AOI22xp33_ASAP7_75t_L g668 ( .A1(n_609), .A2(n_418), .B1(n_391), .B2(n_27), .Y(n_668) );
AOI221xp5_ASAP7_75t_L g669 ( .A1(n_574), .A2(n_418), .B1(n_391), .B2(n_29), .C(n_31), .Y(n_669) );
AO21x2_ASAP7_75t_L g670 ( .A1(n_606), .A2(n_418), .B(n_391), .Y(n_670) );
OAI21x1_ASAP7_75t_L g671 ( .A1(n_625), .A2(n_418), .B(n_391), .Y(n_671) );
AOI22xp33_ASAP7_75t_L g672 ( .A1(n_565), .A2(n_418), .B1(n_391), .B2(n_29), .Y(n_672) );
OA21x2_ASAP7_75t_L g673 ( .A1(n_606), .A2(n_88), .B(n_86), .Y(n_673) );
AOI22xp33_ASAP7_75t_L g674 ( .A1(n_599), .A2(n_25), .B1(n_28), .B2(n_31), .Y(n_674) );
AND2x4_ASAP7_75t_L g675 ( .A(n_589), .B(n_32), .Y(n_675) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_599), .A2(n_36), .B1(n_37), .B2(n_38), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_581), .Y(n_677) );
CKINVDCx5p33_ASAP7_75t_R g678 ( .A(n_583), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_636), .Y(n_679) );
AND2x2_ASAP7_75t_L g680 ( .A(n_619), .B(n_42), .Y(n_680) );
OAI21xp5_ASAP7_75t_L g681 ( .A1(n_590), .A2(n_407), .B(n_42), .Y(n_681) );
OAI21x1_ASAP7_75t_L g682 ( .A1(n_625), .A2(n_90), .B(n_89), .Y(n_682) );
INVx2_ASAP7_75t_L g683 ( .A(n_628), .Y(n_683) );
OAI22xp33_ASAP7_75t_L g684 ( .A1(n_579), .A2(n_44), .B1(n_45), .B2(n_46), .Y(n_684) );
CKINVDCx20_ASAP7_75t_R g685 ( .A(n_610), .Y(n_685) );
AOI22xp33_ASAP7_75t_L g686 ( .A1(n_623), .A2(n_45), .B1(n_46), .B2(n_47), .Y(n_686) );
AOI222xp33_ASAP7_75t_L g687 ( .A1(n_575), .A2(n_48), .B1(n_50), .B2(n_52), .C1(n_53), .C2(n_54), .Y(n_687) );
OR2x6_ASAP7_75t_L g688 ( .A(n_580), .B(n_52), .Y(n_688) );
NOR2xp33_ASAP7_75t_L g689 ( .A(n_578), .B(n_55), .Y(n_689) );
AND2x2_ASAP7_75t_L g690 ( .A(n_568), .B(n_57), .Y(n_690) );
INVx2_ASAP7_75t_L g691 ( .A(n_634), .Y(n_691) );
INVx2_ASAP7_75t_L g692 ( .A(n_635), .Y(n_692) );
INVx3_ASAP7_75t_L g693 ( .A(n_580), .Y(n_693) );
A2O1A1Ixp33_ASAP7_75t_L g694 ( .A1(n_570), .A2(n_407), .B(n_61), .C(n_62), .Y(n_694) );
AND2x2_ASAP7_75t_L g695 ( .A(n_568), .B(n_60), .Y(n_695) );
INVx5_ASAP7_75t_L g696 ( .A(n_580), .Y(n_696) );
AOI22xp33_ASAP7_75t_L g697 ( .A1(n_618), .A2(n_63), .B1(n_64), .B2(n_65), .Y(n_697) );
AOI22xp5_ASAP7_75t_L g698 ( .A1(n_620), .A2(n_68), .B1(n_69), .B2(n_70), .Y(n_698) );
NOR2xp33_ASAP7_75t_L g699 ( .A(n_568), .B(n_69), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_631), .Y(n_700) );
OAI22xp5_ASAP7_75t_L g701 ( .A1(n_595), .A2(n_74), .B1(n_75), .B2(n_76), .Y(n_701) );
INVx4_ASAP7_75t_L g702 ( .A(n_607), .Y(n_702) );
INVx3_ASAP7_75t_L g703 ( .A(n_589), .Y(n_703) );
OAI211xp5_ASAP7_75t_L g704 ( .A1(n_582), .A2(n_407), .B(n_75), .C(n_76), .Y(n_704) );
AOI21xp33_ASAP7_75t_L g705 ( .A1(n_593), .A2(n_74), .B(n_77), .Y(n_705) );
AOI22xp33_ASAP7_75t_L g706 ( .A1(n_597), .A2(n_78), .B1(n_79), .B2(n_80), .Y(n_706) );
AOI22xp33_ASAP7_75t_L g707 ( .A1(n_597), .A2(n_81), .B1(n_83), .B2(n_407), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_629), .Y(n_708) );
OAI22xp5_ASAP7_75t_L g709 ( .A1(n_629), .A2(n_83), .B1(n_407), .B2(n_92), .Y(n_709) );
AOI22xp33_ASAP7_75t_SL g710 ( .A1(n_607), .A2(n_407), .B1(n_96), .B2(n_97), .Y(n_710) );
INVx2_ASAP7_75t_L g711 ( .A(n_671), .Y(n_711) );
OAI221xp5_ASAP7_75t_L g712 ( .A1(n_655), .A2(n_598), .B1(n_584), .B2(n_621), .C(n_622), .Y(n_712) );
OAI211xp5_ASAP7_75t_L g713 ( .A1(n_687), .A2(n_601), .B(n_638), .C(n_626), .Y(n_713) );
AOI22xp5_ASAP7_75t_L g714 ( .A1(n_689), .A2(n_615), .B1(n_637), .B2(n_612), .Y(n_714) );
HB1xp67_ASAP7_75t_L g715 ( .A(n_670), .Y(n_715) );
HB1xp67_ASAP7_75t_L g716 ( .A(n_670), .Y(n_716) );
OAI33xp33_ASAP7_75t_L g717 ( .A1(n_684), .A2(n_639), .A3(n_624), .B1(n_640), .B2(n_585), .B3(n_103), .Y(n_717) );
AOI22xp33_ASAP7_75t_L g718 ( .A1(n_688), .A2(n_585), .B1(n_640), .B2(n_632), .Y(n_718) );
INVx2_ASAP7_75t_L g719 ( .A(n_658), .Y(n_719) );
AOI211xp5_ASAP7_75t_L g720 ( .A1(n_699), .A2(n_641), .B(n_632), .C(n_588), .Y(n_720) );
AOI22xp33_ASAP7_75t_L g721 ( .A1(n_688), .A2(n_641), .B1(n_632), .B2(n_588), .Y(n_721) );
AOI211xp5_ASAP7_75t_SL g722 ( .A1(n_684), .A2(n_567), .B(n_564), .C(n_100), .Y(n_722) );
OAI33xp33_ASAP7_75t_L g723 ( .A1(n_701), .A2(n_91), .A3(n_99), .B1(n_101), .B2(n_104), .B3(n_105), .Y(n_723) );
AOI33xp33_ASAP7_75t_L g724 ( .A1(n_706), .A2(n_106), .A3(n_108), .B1(n_111), .B2(n_113), .B3(n_115), .Y(n_724) );
OAI221xp5_ASAP7_75t_L g725 ( .A1(n_667), .A2(n_567), .B1(n_564), .B2(n_118), .C(n_119), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_650), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_657), .Y(n_727) );
AOI22xp33_ASAP7_75t_L g728 ( .A1(n_661), .A2(n_567), .B1(n_116), .B2(n_122), .Y(n_728) );
AND2x4_ASAP7_75t_L g729 ( .A(n_696), .B(n_127), .Y(n_729) );
HB1xp67_ASAP7_75t_L g730 ( .A(n_708), .Y(n_730) );
NAND2xp5_ASAP7_75t_SL g731 ( .A(n_647), .B(n_132), .Y(n_731) );
AOI221xp5_ASAP7_75t_L g732 ( .A1(n_674), .A2(n_133), .B1(n_134), .B2(n_136), .C(n_137), .Y(n_732) );
AOI22xp33_ASAP7_75t_L g733 ( .A1(n_644), .A2(n_138), .B1(n_140), .B2(n_141), .Y(n_733) );
AND2x4_ASAP7_75t_L g734 ( .A(n_696), .B(n_144), .Y(n_734) );
NOR2x1_ASAP7_75t_L g735 ( .A(n_702), .B(n_146), .Y(n_735) );
INVx2_ASAP7_75t_L g736 ( .A(n_683), .Y(n_736) );
NOR2xp33_ASAP7_75t_L g737 ( .A(n_659), .B(n_149), .Y(n_737) );
INVx2_ASAP7_75t_L g738 ( .A(n_664), .Y(n_738) );
AOI22xp33_ASAP7_75t_SL g739 ( .A1(n_690), .A2(n_151), .B1(n_152), .B2(n_154), .Y(n_739) );
NOR2xp33_ASAP7_75t_L g740 ( .A(n_677), .B(n_156), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_679), .B(n_223), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_691), .Y(n_742) );
OR2x6_ASAP7_75t_L g743 ( .A(n_675), .B(n_157), .Y(n_743) );
AOI221xp5_ASAP7_75t_L g744 ( .A1(n_676), .A2(n_159), .B1(n_161), .B2(n_162), .C(n_164), .Y(n_744) );
AO21x2_ASAP7_75t_L g745 ( .A1(n_681), .A2(n_168), .B(n_172), .Y(n_745) );
AOI22xp33_ASAP7_75t_L g746 ( .A1(n_648), .A2(n_173), .B1(n_174), .B2(n_178), .Y(n_746) );
AND2x2_ASAP7_75t_L g747 ( .A(n_662), .B(n_180), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_692), .Y(n_748) );
OA21x2_ASAP7_75t_L g749 ( .A1(n_682), .A2(n_187), .B(n_189), .Y(n_749) );
AO21x2_ASAP7_75t_L g750 ( .A1(n_694), .A2(n_192), .B(n_195), .Y(n_750) );
INVx2_ASAP7_75t_L g751 ( .A(n_673), .Y(n_751) );
INVx2_ASAP7_75t_L g752 ( .A(n_673), .Y(n_752) );
BUFx6f_ASAP7_75t_L g753 ( .A(n_696), .Y(n_753) );
INVx2_ASAP7_75t_L g754 ( .A(n_673), .Y(n_754) );
OA21x2_ASAP7_75t_L g755 ( .A1(n_646), .A2(n_196), .B(n_197), .Y(n_755) );
AOI22xp33_ASAP7_75t_L g756 ( .A1(n_707), .A2(n_199), .B1(n_201), .B2(n_202), .Y(n_756) );
AND2x2_ASAP7_75t_L g757 ( .A(n_680), .B(n_203), .Y(n_757) );
INVx2_ASAP7_75t_L g758 ( .A(n_675), .Y(n_758) );
AOI22xp33_ASAP7_75t_L g759 ( .A1(n_707), .A2(n_205), .B1(n_207), .B2(n_209), .Y(n_759) );
HB1xp67_ASAP7_75t_L g760 ( .A(n_703), .Y(n_760) );
AOI22xp33_ASAP7_75t_SL g761 ( .A1(n_695), .A2(n_216), .B1(n_217), .B2(n_709), .Y(n_761) );
NAND2xp33_ASAP7_75t_R g762 ( .A(n_703), .B(n_693), .Y(n_762) );
HB1xp67_ASAP7_75t_L g763 ( .A(n_649), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_700), .B(n_697), .Y(n_764) );
BUFx2_ASAP7_75t_L g765 ( .A(n_665), .Y(n_765) );
OR2x6_ASAP7_75t_L g766 ( .A(n_656), .B(n_653), .Y(n_766) );
INVx2_ASAP7_75t_L g767 ( .A(n_698), .Y(n_767) );
INVx2_ASAP7_75t_L g768 ( .A(n_660), .Y(n_768) );
AOI22xp33_ASAP7_75t_L g769 ( .A1(n_669), .A2(n_686), .B1(n_672), .B2(n_705), .Y(n_769) );
INVx1_ASAP7_75t_L g770 ( .A(n_704), .Y(n_770) );
OAI211xp5_ASAP7_75t_L g771 ( .A1(n_642), .A2(n_668), .B(n_672), .C(n_652), .Y(n_771) );
AND2x2_ASAP7_75t_L g772 ( .A(n_668), .B(n_652), .Y(n_772) );
OAI211xp5_ASAP7_75t_L g773 ( .A1(n_666), .A2(n_710), .B(n_643), .C(n_685), .Y(n_773) );
INVx2_ASAP7_75t_L g774 ( .A(n_738), .Y(n_774) );
INVx4_ASAP7_75t_L g775 ( .A(n_753), .Y(n_775) );
INVxp67_ASAP7_75t_L g776 ( .A(n_765), .Y(n_776) );
AND2x2_ASAP7_75t_L g777 ( .A(n_726), .B(n_645), .Y(n_777) );
BUFx2_ASAP7_75t_L g778 ( .A(n_760), .Y(n_778) );
INVx1_ASAP7_75t_L g779 ( .A(n_727), .Y(n_779) );
AND2x2_ASAP7_75t_L g780 ( .A(n_719), .B(n_663), .Y(n_780) );
INVx2_ASAP7_75t_L g781 ( .A(n_738), .Y(n_781) );
OAI21xp33_ASAP7_75t_SL g782 ( .A1(n_743), .A2(n_654), .B(n_651), .Y(n_782) );
INVx1_ASAP7_75t_L g783 ( .A(n_715), .Y(n_783) );
INVx1_ASAP7_75t_L g784 ( .A(n_716), .Y(n_784) );
INVx1_ASAP7_75t_L g785 ( .A(n_716), .Y(n_785) );
INVx1_ASAP7_75t_L g786 ( .A(n_730), .Y(n_786) );
AND2x2_ASAP7_75t_L g787 ( .A(n_736), .B(n_678), .Y(n_787) );
AND4x1_ASAP7_75t_L g788 ( .A(n_722), .B(n_724), .C(n_720), .D(n_721), .Y(n_788) );
INVx2_ASAP7_75t_L g789 ( .A(n_711), .Y(n_789) );
INVx1_ASAP7_75t_L g790 ( .A(n_742), .Y(n_790) );
INVx1_ASAP7_75t_L g791 ( .A(n_748), .Y(n_791) );
INVxp67_ASAP7_75t_SL g792 ( .A(n_762), .Y(n_792) );
INVx2_ASAP7_75t_L g793 ( .A(n_711), .Y(n_793) );
AOI211x1_ASAP7_75t_SL g794 ( .A1(n_758), .A2(n_764), .B(n_741), .C(n_767), .Y(n_794) );
INVx2_ASAP7_75t_L g795 ( .A(n_751), .Y(n_795) );
INVx1_ASAP7_75t_L g796 ( .A(n_751), .Y(n_796) );
AND2x2_ASAP7_75t_SL g797 ( .A(n_729), .B(n_734), .Y(n_797) );
NOR2x1_ASAP7_75t_L g798 ( .A(n_743), .B(n_734), .Y(n_798) );
AND2x2_ASAP7_75t_L g799 ( .A(n_772), .B(n_763), .Y(n_799) );
AOI221xp5_ASAP7_75t_L g800 ( .A1(n_770), .A2(n_769), .B1(n_712), .B2(n_717), .C(n_773), .Y(n_800) );
INVx1_ASAP7_75t_L g801 ( .A(n_752), .Y(n_801) );
OAI22xp5_ASAP7_75t_L g802 ( .A1(n_743), .A2(n_714), .B1(n_769), .B2(n_728), .Y(n_802) );
AND2x2_ASAP7_75t_L g803 ( .A(n_763), .B(n_754), .Y(n_803) );
INVx1_ASAP7_75t_L g804 ( .A(n_729), .Y(n_804) );
AND2x2_ASAP7_75t_L g805 ( .A(n_752), .B(n_754), .Y(n_805) );
AOI221xp5_ASAP7_75t_L g806 ( .A1(n_737), .A2(n_740), .B1(n_713), .B2(n_723), .C(n_725), .Y(n_806) );
INVx2_ASAP7_75t_L g807 ( .A(n_755), .Y(n_807) );
OR2x2_ASAP7_75t_L g808 ( .A(n_766), .B(n_718), .Y(n_808) );
INVx1_ASAP7_75t_L g809 ( .A(n_735), .Y(n_809) );
AND2x2_ASAP7_75t_L g810 ( .A(n_766), .B(n_747), .Y(n_810) );
AND2x2_ASAP7_75t_L g811 ( .A(n_766), .B(n_757), .Y(n_811) );
OAI31xp33_ASAP7_75t_SL g812 ( .A1(n_731), .A2(n_771), .A3(n_737), .B(n_761), .Y(n_812) );
AND2x2_ASAP7_75t_L g813 ( .A(n_724), .B(n_745), .Y(n_813) );
OAI211xp5_ASAP7_75t_L g814 ( .A1(n_728), .A2(n_739), .B(n_733), .C(n_746), .Y(n_814) );
AOI33xp33_ASAP7_75t_L g815 ( .A1(n_756), .A2(n_759), .A3(n_733), .B1(n_746), .B2(n_732), .B3(n_744), .Y(n_815) );
INVx2_ASAP7_75t_L g816 ( .A(n_755), .Y(n_816) );
INVx2_ASAP7_75t_SL g817 ( .A(n_768), .Y(n_817) );
AND2x2_ASAP7_75t_L g818 ( .A(n_750), .B(n_749), .Y(n_818) );
AND2x2_ASAP7_75t_L g819 ( .A(n_726), .B(n_727), .Y(n_819) );
INVx2_ASAP7_75t_SL g820 ( .A(n_753), .Y(n_820) );
INVx1_ASAP7_75t_L g821 ( .A(n_715), .Y(n_821) );
AND2x2_ASAP7_75t_L g822 ( .A(n_799), .B(n_803), .Y(n_822) );
NOR2x1_ASAP7_75t_L g823 ( .A(n_798), .B(n_775), .Y(n_823) );
INVx1_ASAP7_75t_L g824 ( .A(n_796), .Y(n_824) );
HB1xp67_ASAP7_75t_L g825 ( .A(n_778), .Y(n_825) );
INVx2_ASAP7_75t_L g826 ( .A(n_795), .Y(n_826) );
INVx1_ASAP7_75t_L g827 ( .A(n_801), .Y(n_827) );
INVx2_ASAP7_75t_L g828 ( .A(n_795), .Y(n_828) );
INVx1_ASAP7_75t_L g829 ( .A(n_786), .Y(n_829) );
INVx3_ASAP7_75t_L g830 ( .A(n_807), .Y(n_830) );
AND2x2_ASAP7_75t_L g831 ( .A(n_819), .B(n_777), .Y(n_831) );
INVx2_ASAP7_75t_L g832 ( .A(n_805), .Y(n_832) );
AND2x2_ASAP7_75t_L g833 ( .A(n_783), .B(n_784), .Y(n_833) );
NAND2xp5_ASAP7_75t_L g834 ( .A(n_790), .B(n_791), .Y(n_834) );
AND4x1_ASAP7_75t_L g835 ( .A(n_812), .B(n_800), .C(n_806), .D(n_815), .Y(n_835) );
INVx1_ASAP7_75t_L g836 ( .A(n_785), .Y(n_836) );
AND2x2_ASAP7_75t_L g837 ( .A(n_785), .B(n_821), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_779), .Y(n_838) );
AND2x4_ASAP7_75t_L g839 ( .A(n_817), .B(n_808), .Y(n_839) );
INVx1_ASAP7_75t_L g840 ( .A(n_789), .Y(n_840) );
AOI21xp5_ASAP7_75t_L g841 ( .A1(n_797), .A2(n_782), .B(n_814), .Y(n_841) );
INVx1_ASAP7_75t_L g842 ( .A(n_789), .Y(n_842) );
INVx1_ASAP7_75t_L g843 ( .A(n_793), .Y(n_843) );
AND2x4_ASAP7_75t_L g844 ( .A(n_792), .B(n_774), .Y(n_844) );
AND2x4_ASAP7_75t_L g845 ( .A(n_774), .B(n_781), .Y(n_845) );
AND2x2_ASAP7_75t_L g846 ( .A(n_810), .B(n_811), .Y(n_846) );
AND2x2_ASAP7_75t_L g847 ( .A(n_810), .B(n_811), .Y(n_847) );
INVx1_ASAP7_75t_L g848 ( .A(n_781), .Y(n_848) );
INVx3_ASAP7_75t_L g849 ( .A(n_807), .Y(n_849) );
AND2x2_ASAP7_75t_L g850 ( .A(n_813), .B(n_780), .Y(n_850) );
NAND2xp5_ASAP7_75t_L g851 ( .A(n_802), .B(n_804), .Y(n_851) );
AND2x2_ASAP7_75t_SL g852 ( .A(n_788), .B(n_818), .Y(n_852) );
AND2x2_ASAP7_75t_L g853 ( .A(n_850), .B(n_816), .Y(n_853) );
INVx2_ASAP7_75t_L g854 ( .A(n_828), .Y(n_854) );
INVx1_ASAP7_75t_L g855 ( .A(n_824), .Y(n_855) );
HB1xp67_ASAP7_75t_L g856 ( .A(n_825), .Y(n_856) );
A2O1A1Ixp33_ASAP7_75t_L g857 ( .A1(n_841), .A2(n_776), .B(n_815), .C(n_787), .Y(n_857) );
NAND2xp5_ASAP7_75t_L g858 ( .A(n_831), .B(n_794), .Y(n_858) );
NAND3xp33_ASAP7_75t_L g859 ( .A(n_835), .B(n_809), .C(n_787), .Y(n_859) );
AND2x2_ASAP7_75t_L g860 ( .A(n_850), .B(n_816), .Y(n_860) );
AND2x4_ASAP7_75t_L g861 ( .A(n_839), .B(n_775), .Y(n_861) );
INVx2_ASAP7_75t_SL g862 ( .A(n_823), .Y(n_862) );
AND2x2_ASAP7_75t_SL g863 ( .A(n_852), .B(n_820), .Y(n_863) );
AND2x2_ASAP7_75t_L g864 ( .A(n_822), .B(n_832), .Y(n_864) );
AO21x1_ASAP7_75t_L g865 ( .A1(n_851), .A2(n_838), .B(n_834), .Y(n_865) );
AND2x2_ASAP7_75t_L g866 ( .A(n_846), .B(n_847), .Y(n_866) );
NAND3xp33_ASAP7_75t_L g867 ( .A(n_835), .B(n_852), .C(n_836), .Y(n_867) );
INVxp67_ASAP7_75t_L g868 ( .A(n_856), .Y(n_868) );
AND2x2_ASAP7_75t_L g869 ( .A(n_866), .B(n_839), .Y(n_869) );
NAND2xp33_ASAP7_75t_L g870 ( .A(n_857), .B(n_827), .Y(n_870) );
NOR2xp33_ASAP7_75t_L g871 ( .A(n_859), .B(n_829), .Y(n_871) );
XNOR2xp5_ASAP7_75t_L g872 ( .A(n_867), .B(n_833), .Y(n_872) );
NAND2xp5_ASAP7_75t_L g873 ( .A(n_858), .B(n_837), .Y(n_873) );
AND2x2_ASAP7_75t_L g874 ( .A(n_864), .B(n_844), .Y(n_874) );
INVx1_ASAP7_75t_L g875 ( .A(n_855), .Y(n_875) );
OAI22xp5_ASAP7_75t_L g876 ( .A1(n_863), .A2(n_826), .B1(n_848), .B2(n_840), .Y(n_876) );
NAND2xp5_ASAP7_75t_SL g877 ( .A(n_865), .B(n_845), .Y(n_877) );
OAI221xp5_ASAP7_75t_L g878 ( .A1(n_862), .A2(n_830), .B1(n_849), .B2(n_843), .C(n_842), .Y(n_878) );
AOI222xp33_ASAP7_75t_L g879 ( .A1(n_870), .A2(n_873), .B1(n_877), .B2(n_871), .C1(n_872), .C2(n_868), .Y(n_879) );
AND2x2_ASAP7_75t_L g880 ( .A(n_869), .B(n_874), .Y(n_880) );
NAND4xp25_ASAP7_75t_L g881 ( .A(n_879), .B(n_876), .C(n_878), .D(n_861), .Y(n_881) );
AND4x1_ASAP7_75t_L g882 ( .A(n_881), .B(n_880), .C(n_860), .D(n_853), .Y(n_882) );
AND2x2_ASAP7_75t_L g883 ( .A(n_882), .B(n_875), .Y(n_883) );
INVx2_ASAP7_75t_L g884 ( .A(n_883), .Y(n_884) );
INVx2_ASAP7_75t_L g885 ( .A(n_884), .Y(n_885) );
INVx1_ASAP7_75t_L g886 ( .A(n_885), .Y(n_886) );
INVx1_ASAP7_75t_L g887 ( .A(n_886), .Y(n_887) );
AOI21xp5_ASAP7_75t_L g888 ( .A1(n_887), .A2(n_854), .B(n_848), .Y(n_888) );
endmodule