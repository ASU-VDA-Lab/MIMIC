module fake_jpeg_21464_n_100 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_100);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_100;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_7),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_8),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx4f_ASAP7_75t_SL g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx11_ASAP7_75t_SL g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_21),
.B(n_0),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_24),
.B(n_4),
.Y(n_53)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_21),
.B(n_1),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_27),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_12),
.B(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_29),
.Y(n_37)
);

INVx6_ASAP7_75t_SL g29 ( 
.A(n_22),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_31),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_17),
.B(n_2),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_12),
.B(n_14),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_34),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_17),
.B(n_2),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_24),
.A2(n_20),
.B1(n_18),
.B2(n_14),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_47),
.Y(n_59)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_41),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_13),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_13),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_45),
.Y(n_57)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_18),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_26),
.A2(n_28),
.B1(n_25),
.B2(n_20),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_29),
.A2(n_16),
.B1(n_15),
.B2(n_23),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_48),
.B(n_50),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_24),
.A2(n_16),
.B1(n_23),
.B2(n_7),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_33),
.B(n_16),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_52),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_33),
.B(n_4),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_10),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

AO21x1_ASAP7_75t_L g70 ( 
.A1(n_56),
.A2(n_63),
.B(n_66),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_61),
.B(n_67),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_6),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_6),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_65),
.B(n_53),
.C(n_47),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_71),
.C(n_72),
.Y(n_81)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_54),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_59),
.A2(n_49),
.B(n_35),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_59),
.B(n_36),
.C(n_38),
.Y(n_72)
);

NOR3xp33_ASAP7_75t_SL g73 ( 
.A(n_57),
.B(n_64),
.C(n_55),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_73),
.B(n_75),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_49),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_50),
.Y(n_76)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_76),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_9),
.Y(n_77)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_77),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_SL g79 ( 
.A(n_71),
.B(n_66),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_72),
.C(n_68),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_60),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_82),
.B(n_60),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_83),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_86),
.B(n_88),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_83),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_73),
.C(n_78),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_89),
.B(n_90),
.C(n_80),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_91),
.A2(n_93),
.B(n_94),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_87),
.B(n_82),
.C(n_84),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_88),
.B(n_85),
.C(n_56),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_92),
.A2(n_70),
.B(n_74),
.Y(n_96)
);

BUFx24_ASAP7_75t_SL g97 ( 
.A(n_96),
.Y(n_97)
);

A2O1A1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_95),
.A2(n_63),
.B(n_9),
.C(n_43),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_98),
.B(n_97),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_39),
.Y(n_100)
);


endmodule