module fake_netlist_6_699_n_1792 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1792);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1792;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1371;
wire n_1285;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_297;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_1764;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1373;
wire n_1292;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_146),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_1),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_36),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_41),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_131),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_66),
.Y(n_168)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_160),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_154),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_35),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_5),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_113),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_50),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_57),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_114),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_31),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_157),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_11),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_148),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_125),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_4),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_147),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_15),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_90),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_19),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_31),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_110),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_77),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_3),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_139),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_56),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_133),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_104),
.Y(n_194)
);

INVxp67_ASAP7_75t_SL g195 ( 
.A(n_156),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_12),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_94),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_111),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_65),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_63),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_52),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_88),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_129),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_42),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_116),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_95),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_79),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_13),
.Y(n_208)
);

BUFx10_ASAP7_75t_L g209 ( 
.A(n_1),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_123),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_57),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_102),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_25),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_83),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_65),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_71),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_75),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_74),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_161),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_55),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_100),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_55),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_106),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_69),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_47),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_30),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_122),
.Y(n_227)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_121),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_120),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_23),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_98),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_28),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_109),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_127),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_58),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_118),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_27),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_137),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_145),
.Y(n_239)
);

INVxp67_ASAP7_75t_SL g240 ( 
.A(n_81),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_91),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_32),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_153),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_101),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_130),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_134),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_84),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_23),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_34),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_35),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_33),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_48),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_16),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_2),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_44),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_33),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_17),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_80),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_24),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_67),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_119),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_26),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_159),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_128),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_158),
.Y(n_265)
);

BUFx2_ASAP7_75t_SL g266 ( 
.A(n_30),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_140),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_93),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_76),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_18),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_34),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_45),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_0),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_150),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g275 ( 
.A(n_46),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_68),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_92),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_6),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_26),
.Y(n_279)
);

CKINVDCx14_ASAP7_75t_R g280 ( 
.A(n_126),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_39),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_52),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_11),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_62),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_47),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_89),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_59),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_70),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_144),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_67),
.Y(n_290)
);

BUFx10_ASAP7_75t_L g291 ( 
.A(n_10),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_97),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_32),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_107),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_115),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_51),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_4),
.Y(n_297)
);

BUFx10_ASAP7_75t_L g298 ( 
.A(n_105),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_20),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_40),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_53),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_99),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_63),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_132),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_18),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_39),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_82),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_96),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_48),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_42),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_61),
.Y(n_311)
);

CKINVDCx14_ASAP7_75t_R g312 ( 
.A(n_117),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_151),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_256),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_256),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_256),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_163),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_256),
.Y(n_318)
);

INVxp67_ASAP7_75t_SL g319 ( 
.A(n_250),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_167),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_203),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_207),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_308),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_187),
.B(n_2),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_174),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_256),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_170),
.Y(n_327)
);

CKINVDCx14_ASAP7_75t_R g328 ( 
.A(n_280),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_173),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_180),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_210),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_181),
.Y(n_332)
);

CKINVDCx16_ASAP7_75t_R g333 ( 
.A(n_281),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_256),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_250),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_188),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_238),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_174),
.Y(n_338)
);

INVxp33_ASAP7_75t_SL g339 ( 
.A(n_165),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_191),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_202),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_206),
.Y(n_342)
);

CKINVDCx16_ASAP7_75t_R g343 ( 
.A(n_281),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_250),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_164),
.Y(n_345)
);

INVxp33_ASAP7_75t_SL g346 ( 
.A(n_166),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_214),
.Y(n_347)
);

INVxp67_ASAP7_75t_SL g348 ( 
.A(n_228),
.Y(n_348)
);

CKINVDCx16_ASAP7_75t_R g349 ( 
.A(n_310),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_164),
.Y(n_350)
);

BUFx2_ASAP7_75t_L g351 ( 
.A(n_187),
.Y(n_351)
);

OAI21x1_ASAP7_75t_L g352 ( 
.A1(n_169),
.A2(n_3),
.B(n_5),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_247),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_247),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_204),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_204),
.Y(n_356)
);

BUFx3_ASAP7_75t_L g357 ( 
.A(n_298),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_187),
.Y(n_358)
);

INVxp67_ASAP7_75t_SL g359 ( 
.A(n_179),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_176),
.B(n_6),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_179),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_216),
.Y(n_362)
);

OR2x2_ASAP7_75t_L g363 ( 
.A(n_184),
.B(n_7),
.Y(n_363)
);

INVxp67_ASAP7_75t_SL g364 ( 
.A(n_267),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_282),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_312),
.Y(n_366)
);

INVxp67_ASAP7_75t_SL g367 ( 
.A(n_184),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_218),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_219),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_221),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_282),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_223),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_282),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_231),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_236),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_239),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_243),
.Y(n_377)
);

HB1xp67_ASAP7_75t_L g378 ( 
.A(n_310),
.Y(n_378)
);

INVxp33_ASAP7_75t_SL g379 ( 
.A(n_168),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_208),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_244),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_308),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_245),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_246),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_176),
.B(n_7),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_208),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_258),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_215),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_215),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_261),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_321),
.A2(n_171),
.B1(n_259),
.B2(n_220),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_323),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_314),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_319),
.B(n_263),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_323),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_314),
.Y(n_396)
);

BUFx3_ASAP7_75t_L g397 ( 
.A(n_315),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_315),
.Y(n_398)
);

HB1xp67_ASAP7_75t_L g399 ( 
.A(n_378),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_316),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_316),
.Y(n_401)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_323),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_318),
.Y(n_403)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_382),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_318),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_326),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_382),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_326),
.Y(n_408)
);

AND2x4_ASAP7_75t_SL g409 ( 
.A(n_368),
.B(n_298),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_322),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_382),
.Y(n_411)
);

BUFx3_ASAP7_75t_L g412 ( 
.A(n_334),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_334),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_319),
.B(n_264),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_335),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_335),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_344),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_344),
.Y(n_418)
);

NOR2x1_ASAP7_75t_L g419 ( 
.A(n_345),
.B(n_169),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_352),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_352),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_345),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_358),
.B(n_265),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_350),
.Y(n_424)
);

AND2x4_ASAP7_75t_L g425 ( 
.A(n_324),
.B(n_169),
.Y(n_425)
);

BUFx3_ASAP7_75t_L g426 ( 
.A(n_358),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_352),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_365),
.B(n_269),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_350),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_355),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g431 ( 
.A(n_351),
.Y(n_431)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_351),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_355),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_324),
.B(n_169),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_356),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_356),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_380),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_380),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_369),
.Y(n_439)
);

INVx2_ASAP7_75t_SL g440 ( 
.A(n_365),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_386),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_386),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_388),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_388),
.Y(n_444)
);

AND2x6_ASAP7_75t_L g445 ( 
.A(n_360),
.B(n_308),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_371),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_371),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_373),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_373),
.B(n_313),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_363),
.Y(n_450)
);

NAND2x1_ASAP7_75t_L g451 ( 
.A(n_385),
.B(n_194),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_359),
.Y(n_452)
);

OA21x2_ASAP7_75t_L g453 ( 
.A1(n_325),
.A2(n_222),
.B(n_220),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_359),
.B(n_276),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_SL g455 ( 
.A(n_333),
.B(n_209),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_367),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_363),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_367),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_325),
.Y(n_459)
);

CKINVDCx16_ASAP7_75t_R g460 ( 
.A(n_333),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_338),
.Y(n_461)
);

OA21x2_ASAP7_75t_L g462 ( 
.A1(n_338),
.A2(n_230),
.B(n_222),
.Y(n_462)
);

INVx3_ASAP7_75t_L g463 ( 
.A(n_357),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_361),
.Y(n_464)
);

NAND2xp33_ASAP7_75t_SL g465 ( 
.A(n_451),
.B(n_366),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_452),
.B(n_339),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_442),
.Y(n_467)
);

AOI22xp33_ASAP7_75t_L g468 ( 
.A1(n_445),
.A2(n_348),
.B1(n_364),
.B2(n_230),
.Y(n_468)
);

INVx3_ASAP7_75t_L g469 ( 
.A(n_407),
.Y(n_469)
);

BUFx3_ASAP7_75t_L g470 ( 
.A(n_426),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_463),
.B(n_394),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_463),
.B(n_317),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_410),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_448),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_450),
.B(n_357),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_463),
.B(n_320),
.Y(n_476)
);

INVx2_ASAP7_75t_SL g477 ( 
.A(n_431),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_391),
.B(n_331),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_452),
.B(n_346),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_455),
.B(n_327),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_448),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_448),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_463),
.B(n_329),
.Y(n_483)
);

NAND2xp33_ASAP7_75t_SL g484 ( 
.A(n_451),
.B(n_353),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_392),
.Y(n_485)
);

NAND3xp33_ASAP7_75t_L g486 ( 
.A(n_451),
.B(n_183),
.C(n_178),
.Y(n_486)
);

BUFx3_ASAP7_75t_L g487 ( 
.A(n_426),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_426),
.Y(n_488)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_407),
.Y(n_489)
);

INVx4_ASAP7_75t_L g490 ( 
.A(n_407),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_463),
.B(n_330),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_463),
.B(n_332),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_450),
.B(n_357),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_413),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_452),
.B(n_379),
.Y(n_495)
);

AOI22xp33_ASAP7_75t_SL g496 ( 
.A1(n_455),
.A2(n_354),
.B1(n_343),
.B2(n_349),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_426),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_397),
.Y(n_498)
);

BUFx4f_ASAP7_75t_L g499 ( 
.A(n_453),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_456),
.B(n_336),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_442),
.Y(n_501)
);

BUFx3_ASAP7_75t_L g502 ( 
.A(n_397),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_397),
.Y(n_503)
);

BUFx4f_ASAP7_75t_L g504 ( 
.A(n_453),
.Y(n_504)
);

AND2x2_ASAP7_75t_L g505 ( 
.A(n_450),
.B(n_361),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_392),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_413),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_413),
.Y(n_508)
);

INVx3_ASAP7_75t_L g509 ( 
.A(n_407),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_456),
.B(n_340),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_456),
.B(n_341),
.Y(n_511)
);

OR2x6_ASAP7_75t_L g512 ( 
.A(n_450),
.B(n_266),
.Y(n_512)
);

INVx4_ASAP7_75t_L g513 ( 
.A(n_407),
.Y(n_513)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_407),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_413),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_394),
.B(n_342),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_414),
.B(n_347),
.Y(n_517)
);

AND3x2_ASAP7_75t_L g518 ( 
.A(n_399),
.B(n_262),
.C(n_234),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_392),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_392),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_397),
.Y(n_521)
);

AOI22xp33_ASAP7_75t_L g522 ( 
.A1(n_445),
.A2(n_272),
.B1(n_290),
.B2(n_284),
.Y(n_522)
);

INVxp67_ASAP7_75t_SL g523 ( 
.A(n_458),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_432),
.B(n_362),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_442),
.Y(n_525)
);

OR2x6_ASAP7_75t_L g526 ( 
.A(n_457),
.B(n_266),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_414),
.B(n_377),
.Y(n_527)
);

INVx5_ASAP7_75t_L g528 ( 
.A(n_407),
.Y(n_528)
);

INVx3_ASAP7_75t_L g529 ( 
.A(n_407),
.Y(n_529)
);

AO22x2_ASAP7_75t_L g530 ( 
.A1(n_425),
.A2(n_271),
.B1(n_235),
.B2(n_242),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g531 ( 
.A1(n_445),
.A2(n_275),
.B1(n_343),
.B2(n_349),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_412),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_458),
.B(n_381),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_412),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_407),
.Y(n_535)
);

OR2x2_ASAP7_75t_L g536 ( 
.A(n_431),
.B(n_383),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_458),
.B(n_384),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_425),
.B(n_387),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_432),
.B(n_390),
.Y(n_539)
);

BUFx3_ASAP7_75t_L g540 ( 
.A(n_412),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_442),
.Y(n_541)
);

OAI21xp33_ASAP7_75t_SL g542 ( 
.A1(n_457),
.A2(n_242),
.B(n_235),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_395),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_395),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_412),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_457),
.B(n_370),
.Y(n_546)
);

OAI22xp33_ASAP7_75t_L g547 ( 
.A1(n_454),
.A2(n_211),
.B1(n_186),
.B2(n_190),
.Y(n_547)
);

BUFx3_ASAP7_75t_L g548 ( 
.A(n_425),
.Y(n_548)
);

INVx2_ASAP7_75t_SL g549 ( 
.A(n_425),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_425),
.B(n_328),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_440),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_440),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_395),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_440),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_395),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_457),
.B(n_372),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_440),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_438),
.Y(n_558)
);

AND2x6_ASAP7_75t_L g559 ( 
.A(n_420),
.B(n_194),
.Y(n_559)
);

BUFx3_ASAP7_75t_L g560 ( 
.A(n_425),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_393),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_438),
.Y(n_562)
);

BUFx2_ASAP7_75t_L g563 ( 
.A(n_399),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_411),
.Y(n_564)
);

INVx1_ASAP7_75t_SL g565 ( 
.A(n_410),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_438),
.Y(n_566)
);

OR2x2_ASAP7_75t_L g567 ( 
.A(n_454),
.B(n_389),
.Y(n_567)
);

AOI22xp33_ASAP7_75t_L g568 ( 
.A1(n_445),
.A2(n_271),
.B1(n_272),
.B2(n_311),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_449),
.B(n_389),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_441),
.Y(n_570)
);

BUFx3_ASAP7_75t_L g571 ( 
.A(n_453),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_441),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_423),
.B(n_374),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_402),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_434),
.B(n_286),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_402),
.Y(n_576)
);

INVx4_ASAP7_75t_SL g577 ( 
.A(n_420),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_441),
.Y(n_578)
);

INVx3_ASAP7_75t_L g579 ( 
.A(n_411),
.Y(n_579)
);

NAND2xp33_ASAP7_75t_R g580 ( 
.A(n_439),
.B(n_172),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_464),
.B(n_375),
.Y(n_581)
);

AOI22xp33_ASAP7_75t_L g582 ( 
.A1(n_445),
.A2(n_284),
.B1(n_249),
.B2(n_311),
.Y(n_582)
);

INVx2_ASAP7_75t_SL g583 ( 
.A(n_434),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_443),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_393),
.Y(n_585)
);

INVx5_ASAP7_75t_L g586 ( 
.A(n_411),
.Y(n_586)
);

NAND3xp33_ASAP7_75t_L g587 ( 
.A(n_453),
.B(n_183),
.C(n_178),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_464),
.B(n_376),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_402),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_434),
.B(n_288),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_402),
.Y(n_591)
);

OAI21xp33_ASAP7_75t_SL g592 ( 
.A1(n_434),
.A2(n_254),
.B(n_249),
.Y(n_592)
);

INVx4_ASAP7_75t_L g593 ( 
.A(n_411),
.Y(n_593)
);

XOR2x2_ASAP7_75t_L g594 ( 
.A(n_391),
.B(n_8),
.Y(n_594)
);

BUFx3_ASAP7_75t_L g595 ( 
.A(n_453),
.Y(n_595)
);

INVx1_ASAP7_75t_SL g596 ( 
.A(n_439),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_443),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_393),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_396),
.Y(n_599)
);

CKINVDCx20_ASAP7_75t_R g600 ( 
.A(n_460),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_449),
.B(n_185),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_396),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_396),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_423),
.B(n_337),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_398),
.Y(n_605)
);

INVx3_ASAP7_75t_L g606 ( 
.A(n_411),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_398),
.Y(n_607)
);

BUFx4f_ASAP7_75t_L g608 ( 
.A(n_453),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_443),
.Y(n_609)
);

BUFx4f_ASAP7_75t_L g610 ( 
.A(n_453),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_446),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_442),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_446),
.Y(n_613)
);

NOR2x1p5_ASAP7_75t_L g614 ( 
.A(n_464),
.B(n_459),
.Y(n_614)
);

NOR2xp67_ASAP7_75t_L g615 ( 
.A(n_486),
.B(n_428),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_583),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_583),
.B(n_445),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_500),
.B(n_460),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_558),
.Y(n_619)
);

AOI22xp5_ASAP7_75t_L g620 ( 
.A1(n_573),
.A2(n_445),
.B1(n_428),
.B2(n_409),
.Y(n_620)
);

OAI221xp5_ASAP7_75t_L g621 ( 
.A1(n_468),
.A2(n_461),
.B1(n_459),
.B2(n_462),
.C(n_299),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_510),
.B(n_445),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_548),
.Y(n_623)
);

HB1xp67_ASAP7_75t_L g624 ( 
.A(n_563),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_511),
.B(n_445),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_558),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_562),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_562),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_533),
.B(n_445),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_549),
.B(n_420),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_523),
.B(n_445),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_566),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_475),
.B(n_445),
.Y(n_633)
);

INVx2_ASAP7_75t_SL g634 ( 
.A(n_614),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_549),
.B(n_420),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_548),
.Y(n_636)
);

AOI22xp5_ASAP7_75t_SL g637 ( 
.A1(n_478),
.A2(n_232),
.B1(n_226),
.B2(n_225),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_566),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_499),
.B(n_420),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_499),
.B(n_420),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_475),
.B(n_462),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_570),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_548),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_570),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_572),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_560),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_560),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_493),
.B(n_462),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_572),
.Y(n_649)
);

AOI22xp5_ASAP7_75t_L g650 ( 
.A1(n_604),
.A2(n_409),
.B1(n_195),
.B2(n_240),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_578),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_493),
.B(n_462),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_516),
.B(n_409),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_499),
.B(n_420),
.Y(n_654)
);

AOI22xp33_ASAP7_75t_L g655 ( 
.A1(n_571),
.A2(n_595),
.B1(n_587),
.B2(n_560),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_498),
.Y(n_656)
);

BUFx6f_ASAP7_75t_L g657 ( 
.A(n_571),
.Y(n_657)
);

HB1xp67_ASAP7_75t_L g658 ( 
.A(n_563),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_517),
.B(n_462),
.Y(n_659)
);

OR2x2_ASAP7_75t_L g660 ( 
.A(n_477),
.B(n_567),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_527),
.B(n_462),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_504),
.B(n_608),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_578),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_537),
.B(n_462),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_584),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_498),
.Y(n_666)
);

INVx4_ASAP7_75t_L g667 ( 
.A(n_577),
.Y(n_667)
);

AOI22xp33_ASAP7_75t_L g668 ( 
.A1(n_571),
.A2(n_420),
.B1(n_421),
.B2(n_427),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_575),
.B(n_420),
.Y(n_669)
);

BUFx6f_ASAP7_75t_L g670 ( 
.A(n_470),
.Y(n_670)
);

NAND3xp33_ASAP7_75t_SL g671 ( 
.A(n_531),
.B(n_177),
.C(n_175),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_590),
.B(n_421),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_471),
.B(n_421),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_503),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_466),
.B(n_479),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_503),
.Y(n_676)
);

NOR2xp67_ASAP7_75t_L g677 ( 
.A(n_486),
.B(n_459),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_495),
.B(n_421),
.Y(n_678)
);

NOR2xp67_ASAP7_75t_L g679 ( 
.A(n_536),
.B(n_567),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_569),
.B(n_461),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_521),
.Y(n_681)
);

INVx1_ASAP7_75t_SL g682 ( 
.A(n_473),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_505),
.B(n_421),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_584),
.Y(n_684)
);

NOR3xp33_ASAP7_75t_L g685 ( 
.A(n_546),
.B(n_461),
.C(n_449),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_505),
.B(n_421),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_504),
.B(n_421),
.Y(n_687)
);

OR2x6_ASAP7_75t_L g688 ( 
.A(n_530),
.B(n_449),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_536),
.B(n_524),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_551),
.B(n_421),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_597),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_521),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_551),
.B(n_421),
.Y(n_693)
);

AOI22xp33_ASAP7_75t_L g694 ( 
.A1(n_595),
.A2(n_427),
.B1(n_234),
.B2(n_419),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_552),
.B(n_427),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_539),
.B(n_182),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_581),
.B(n_192),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_504),
.B(n_608),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_R g699 ( 
.A(n_580),
.B(n_289),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_608),
.B(n_610),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_597),
.Y(n_701)
);

INVxp67_ASAP7_75t_L g702 ( 
.A(n_477),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_552),
.B(n_427),
.Y(n_703)
);

OR2x6_ASAP7_75t_L g704 ( 
.A(n_530),
.B(n_185),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_532),
.Y(n_705)
);

AOI22xp5_ASAP7_75t_L g706 ( 
.A1(n_484),
.A2(n_307),
.B1(n_304),
.B2(n_295),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_554),
.B(n_427),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_532),
.Y(n_708)
);

AOI22xp33_ASAP7_75t_L g709 ( 
.A1(n_595),
.A2(n_427),
.B1(n_419),
.B2(n_233),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_534),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_554),
.B(n_557),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_557),
.B(n_427),
.Y(n_712)
);

INVxp33_ASAP7_75t_L g713 ( 
.A(n_569),
.Y(n_713)
);

INVx5_ASAP7_75t_L g714 ( 
.A(n_559),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_609),
.B(n_427),
.Y(n_715)
);

INVxp67_ASAP7_75t_L g716 ( 
.A(n_556),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_534),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_609),
.B(n_427),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_545),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_610),
.B(n_577),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_561),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_488),
.B(n_446),
.Y(n_722)
);

AOI22xp5_ASAP7_75t_L g723 ( 
.A1(n_465),
.A2(n_292),
.B1(n_294),
.B2(n_302),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_488),
.B(n_497),
.Y(n_724)
);

NAND2xp33_ASAP7_75t_L g725 ( 
.A(n_559),
.B(n_189),
.Y(n_725)
);

AOI22xp5_ASAP7_75t_L g726 ( 
.A1(n_531),
.A2(n_538),
.B1(n_512),
.B2(n_526),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_545),
.Y(n_727)
);

NAND2xp33_ASAP7_75t_L g728 ( 
.A(n_559),
.B(n_189),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_561),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_610),
.B(n_442),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_577),
.B(n_442),
.Y(n_731)
);

INVx3_ASAP7_75t_L g732 ( 
.A(n_502),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_585),
.Y(n_733)
);

NAND2xp33_ASAP7_75t_L g734 ( 
.A(n_559),
.B(n_193),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_497),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_474),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_SL g737 ( 
.A(n_596),
.B(n_298),
.Y(n_737)
);

OAI22xp5_ASAP7_75t_L g738 ( 
.A1(n_512),
.A2(n_229),
.B1(n_313),
.B2(n_302),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_474),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_598),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_588),
.B(n_196),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_481),
.B(n_447),
.Y(n_742)
);

INVxp67_ASAP7_75t_L g743 ( 
.A(n_565),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_577),
.B(n_442),
.Y(n_744)
);

AOI221xp5_ASAP7_75t_L g745 ( 
.A1(n_547),
.A2(n_306),
.B1(n_305),
.B2(n_301),
.C(n_300),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_481),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_480),
.B(n_199),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_577),
.B(n_442),
.Y(n_748)
);

NOR2x1p5_ASAP7_75t_L g749 ( 
.A(n_550),
.B(n_200),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_472),
.B(n_201),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_476),
.B(n_213),
.Y(n_751)
);

AOI21xp5_ASAP7_75t_L g752 ( 
.A1(n_483),
.A2(n_419),
.B(n_446),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_598),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_482),
.B(n_447),
.Y(n_754)
);

OAI22xp33_ASAP7_75t_L g755 ( 
.A1(n_512),
.A2(n_229),
.B1(n_197),
.B2(n_198),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_482),
.B(n_447),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_601),
.B(n_447),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_601),
.B(n_398),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_614),
.B(n_400),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_470),
.B(n_400),
.Y(n_760)
);

INVxp67_ASAP7_75t_L g761 ( 
.A(n_496),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_470),
.B(n_400),
.Y(n_762)
);

BUFx8_ASAP7_75t_L g763 ( 
.A(n_600),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_491),
.B(n_429),
.Y(n_764)
);

AND2x4_ASAP7_75t_L g765 ( 
.A(n_487),
.B(n_193),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_492),
.B(n_429),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_512),
.B(n_237),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_487),
.B(n_401),
.Y(n_768)
);

AOI22xp33_ASAP7_75t_L g769 ( 
.A1(n_587),
.A2(n_582),
.B1(n_522),
.B2(n_568),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_599),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_487),
.B(n_429),
.Y(n_771)
);

OR2x2_ASAP7_75t_L g772 ( 
.A(n_526),
.B(n_254),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_526),
.B(n_248),
.Y(n_773)
);

AOI22xp5_ASAP7_75t_L g774 ( 
.A1(n_526),
.A2(n_217),
.B1(n_197),
.B2(n_277),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_592),
.B(n_429),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_592),
.B(n_429),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_526),
.B(n_251),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_502),
.B(n_429),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_502),
.Y(n_779)
);

OAI221xp5_ASAP7_75t_L g780 ( 
.A1(n_542),
.A2(n_290),
.B1(n_278),
.B2(n_283),
.C(n_293),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_599),
.Y(n_781)
);

AOI22xp33_ASAP7_75t_L g782 ( 
.A1(n_530),
.A2(n_212),
.B1(n_198),
.B2(n_205),
.Y(n_782)
);

OAI22xp5_ASAP7_75t_L g783 ( 
.A1(n_675),
.A2(n_540),
.B1(n_530),
.B2(n_602),
.Y(n_783)
);

AOI21xp5_ASAP7_75t_L g784 ( 
.A1(n_668),
.A2(n_673),
.B(n_672),
.Y(n_784)
);

CKINVDCx10_ASAP7_75t_R g785 ( 
.A(n_763),
.Y(n_785)
);

AOI21xp5_ASAP7_75t_L g786 ( 
.A1(n_669),
.A2(n_513),
.B(n_490),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_679),
.B(n_518),
.Y(n_787)
);

OAI21xp5_ASAP7_75t_L g788 ( 
.A1(n_678),
.A2(n_559),
.B(n_613),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_616),
.B(n_540),
.Y(n_789)
);

NOR2xp67_ASAP7_75t_L g790 ( 
.A(n_743),
.B(n_542),
.Y(n_790)
);

OAI21xp5_ASAP7_75t_L g791 ( 
.A1(n_659),
.A2(n_559),
.B(n_611),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_616),
.Y(n_792)
);

AOI21xp5_ASAP7_75t_L g793 ( 
.A1(n_683),
.A2(n_513),
.B(n_490),
.Y(n_793)
);

AOI21xp5_ASAP7_75t_L g794 ( 
.A1(n_686),
.A2(n_513),
.B(n_490),
.Y(n_794)
);

AND2x4_ASAP7_75t_L g795 ( 
.A(n_634),
.B(n_540),
.Y(n_795)
);

O2A1O1Ixp33_ASAP7_75t_L g796 ( 
.A1(n_621),
.A2(n_607),
.B(n_602),
.C(n_605),
.Y(n_796)
);

O2A1O1Ixp33_ASAP7_75t_L g797 ( 
.A1(n_661),
.A2(n_607),
.B(n_603),
.C(n_605),
.Y(n_797)
);

AOI21xp5_ASAP7_75t_L g798 ( 
.A1(n_639),
.A2(n_513),
.B(n_490),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_619),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_619),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_750),
.B(n_559),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_639),
.A2(n_593),
.B(n_501),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_713),
.B(n_603),
.Y(n_803)
);

OAI321xp33_ASAP7_75t_L g804 ( 
.A1(n_745),
.A2(n_283),
.A3(n_278),
.B1(n_293),
.B2(n_296),
.C(n_297),
.Y(n_804)
);

AND2x4_ASAP7_75t_L g805 ( 
.A(n_634),
.B(n_623),
.Y(n_805)
);

AOI21xp5_ASAP7_75t_L g806 ( 
.A1(n_640),
.A2(n_687),
.B(n_654),
.Y(n_806)
);

INVx3_ASAP7_75t_L g807 ( 
.A(n_670),
.Y(n_807)
);

A2O1A1Ixp33_ASAP7_75t_L g808 ( 
.A1(n_697),
.A2(n_224),
.B(n_217),
.C(n_212),
.Y(n_808)
);

INVxp67_ASAP7_75t_L g809 ( 
.A(n_660),
.Y(n_809)
);

O2A1O1Ixp33_ASAP7_75t_L g810 ( 
.A1(n_664),
.A2(n_613),
.B(n_611),
.C(n_268),
.Y(n_810)
);

NOR3xp33_ASAP7_75t_L g811 ( 
.A(n_761),
.B(n_224),
.C(n_205),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_751),
.B(n_469),
.Y(n_812)
);

AOI33xp33_ASAP7_75t_L g813 ( 
.A1(n_680),
.A2(n_305),
.A3(n_306),
.B1(n_301),
.B2(n_300),
.B3(n_299),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_R g814 ( 
.A(n_671),
.B(n_252),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_680),
.B(n_469),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_626),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_677),
.B(n_469),
.Y(n_817)
);

BUFx2_ASAP7_75t_L g818 ( 
.A(n_624),
.Y(n_818)
);

AOI21xp5_ASAP7_75t_L g819 ( 
.A1(n_640),
.A2(n_593),
.B(n_501),
.Y(n_819)
);

AOI22xp5_ASAP7_75t_L g820 ( 
.A1(n_620),
.A2(n_689),
.B1(n_653),
.B2(n_618),
.Y(n_820)
);

OAI21xp5_ASAP7_75t_L g821 ( 
.A1(n_641),
.A2(n_507),
.B(n_494),
.Y(n_821)
);

AOI21x1_ASAP7_75t_L g822 ( 
.A1(n_731),
.A2(n_507),
.B(n_494),
.Y(n_822)
);

AOI22xp5_ASAP7_75t_L g823 ( 
.A1(n_615),
.A2(n_535),
.B1(n_606),
.B2(n_514),
.Y(n_823)
);

O2A1O1Ixp5_ASAP7_75t_L g824 ( 
.A1(n_775),
.A2(n_515),
.B(n_508),
.C(n_489),
.Y(n_824)
);

BUFx6f_ASAP7_75t_L g825 ( 
.A(n_657),
.Y(n_825)
);

O2A1O1Ixp33_ASAP7_75t_L g826 ( 
.A1(n_713),
.A2(n_274),
.B(n_241),
.C(n_268),
.Y(n_826)
);

OAI21xp5_ASAP7_75t_L g827 ( 
.A1(n_648),
.A2(n_515),
.B(n_508),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_736),
.B(n_739),
.Y(n_828)
);

INVx3_ASAP7_75t_L g829 ( 
.A(n_670),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_746),
.B(n_469),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_627),
.Y(n_831)
);

INVx11_ASAP7_75t_L g832 ( 
.A(n_763),
.Y(n_832)
);

OAI21xp5_ASAP7_75t_L g833 ( 
.A1(n_652),
.A2(n_520),
.B(n_519),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_628),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_657),
.B(n_667),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_694),
.B(n_489),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_655),
.B(n_732),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_732),
.B(n_685),
.Y(n_838)
);

AND2x2_ASAP7_75t_SL g839 ( 
.A(n_782),
.B(n_227),
.Y(n_839)
);

A2O1A1Ixp33_ASAP7_75t_L g840 ( 
.A1(n_741),
.A2(n_233),
.B(n_227),
.C(n_241),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_654),
.A2(n_593),
.B(n_541),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_732),
.B(n_489),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_628),
.Y(n_843)
);

HB1xp67_ASAP7_75t_L g844 ( 
.A(n_658),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_657),
.B(n_467),
.Y(n_845)
);

INVx3_ASAP7_75t_L g846 ( 
.A(n_670),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_687),
.A2(n_593),
.B(n_541),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_630),
.A2(n_612),
.B(n_467),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_630),
.A2(n_612),
.B(n_467),
.Y(n_849)
);

OAI21xp5_ASAP7_75t_L g850 ( 
.A1(n_633),
.A2(n_543),
.B(n_553),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_632),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_709),
.B(n_489),
.Y(n_852)
);

OAI21xp33_ASAP7_75t_L g853 ( 
.A1(n_696),
.A2(n_594),
.B(n_260),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_759),
.B(n_509),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_716),
.B(n_253),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_657),
.B(n_467),
.Y(n_856)
);

INVxp67_ASAP7_75t_L g857 ( 
.A(n_772),
.Y(n_857)
);

BUFx6f_ASAP7_75t_L g858 ( 
.A(n_657),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_632),
.B(n_509),
.Y(n_859)
);

OAI21xp5_ASAP7_75t_L g860 ( 
.A1(n_617),
.A2(n_543),
.B(n_555),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_702),
.B(n_255),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_635),
.A2(n_612),
.B(n_467),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_699),
.Y(n_863)
);

OAI21xp5_ASAP7_75t_L g864 ( 
.A1(n_631),
.A2(n_544),
.B(n_519),
.Y(n_864)
);

INVx1_ASAP7_75t_SL g865 ( 
.A(n_682),
.Y(n_865)
);

BUFx6f_ASAP7_75t_L g866 ( 
.A(n_670),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_638),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_638),
.B(n_509),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_L g869 ( 
.A(n_767),
.B(n_257),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_SL g870 ( 
.A(n_667),
.B(n_467),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_642),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_642),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_644),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_763),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_644),
.Y(n_875)
);

AOI22xp5_ASAP7_75t_L g876 ( 
.A1(n_726),
.A2(n_564),
.B1(n_606),
.B2(n_509),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_645),
.Y(n_877)
);

BUFx12f_ASAP7_75t_L g878 ( 
.A(n_749),
.Y(n_878)
);

OAI321xp33_ASAP7_75t_L g879 ( 
.A1(n_650),
.A2(n_747),
.A3(n_780),
.B1(n_723),
.B2(n_777),
.C(n_773),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_635),
.A2(n_612),
.B(n_541),
.Y(n_880)
);

O2A1O1Ixp33_ASAP7_75t_L g881 ( 
.A1(n_772),
.A2(n_738),
.B(n_755),
.C(n_775),
.Y(n_881)
);

NAND2x1p5_ASAP7_75t_L g882 ( 
.A(n_667),
.B(n_514),
.Y(n_882)
);

NOR3xp33_ASAP7_75t_L g883 ( 
.A(n_662),
.B(n_270),
.C(n_273),
.Y(n_883)
);

A2O1A1Ixp33_ASAP7_75t_L g884 ( 
.A1(n_622),
.A2(n_514),
.B(n_606),
.C(n_535),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_645),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_SL g886 ( 
.A(n_714),
.B(n_501),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_737),
.B(n_298),
.Y(n_887)
);

O2A1O1Ixp5_ASAP7_75t_L g888 ( 
.A1(n_776),
.A2(n_514),
.B(n_606),
.C(n_529),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_690),
.A2(n_612),
.B(n_501),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_649),
.B(n_529),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_L g891 ( 
.A(n_636),
.B(n_279),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_651),
.B(n_529),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_651),
.B(n_529),
.Y(n_893)
);

A2O1A1Ixp33_ASAP7_75t_L g894 ( 
.A1(n_625),
.A2(n_535),
.B(n_579),
.C(n_564),
.Y(n_894)
);

OAI21xp5_ASAP7_75t_L g895 ( 
.A1(n_629),
.A2(n_520),
.B(n_544),
.Y(n_895)
);

OAI21xp5_ASAP7_75t_L g896 ( 
.A1(n_730),
.A2(n_553),
.B(n_555),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_SL g897 ( 
.A(n_688),
.B(n_209),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_714),
.B(n_501),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_693),
.A2(n_612),
.B(n_501),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_695),
.A2(n_525),
.B(n_541),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_663),
.B(n_535),
.Y(n_901)
);

NOR3xp33_ASAP7_75t_L g902 ( 
.A(n_662),
.B(n_303),
.C(n_309),
.Y(n_902)
);

A2O1A1Ixp33_ASAP7_75t_L g903 ( 
.A1(n_769),
.A2(n_564),
.B(n_579),
.C(n_591),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_665),
.B(n_684),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_637),
.B(n_209),
.Y(n_905)
);

BUFx6f_ASAP7_75t_L g906 ( 
.A(n_688),
.Y(n_906)
);

INVx2_ASAP7_75t_SL g907 ( 
.A(n_765),
.Y(n_907)
);

INVxp67_ASAP7_75t_L g908 ( 
.A(n_765),
.Y(n_908)
);

BUFx4f_ASAP7_75t_L g909 ( 
.A(n_688),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_703),
.A2(n_525),
.B(n_541),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_707),
.A2(n_541),
.B(n_525),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_665),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_643),
.B(n_285),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_684),
.Y(n_914)
);

CKINVDCx10_ASAP7_75t_R g915 ( 
.A(n_704),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_691),
.B(n_579),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_691),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_701),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_701),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_712),
.A2(n_525),
.B(n_579),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_715),
.A2(n_525),
.B(n_528),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_718),
.A2(n_730),
.B(n_757),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_758),
.B(n_485),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_711),
.B(n_485),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_646),
.B(n_485),
.Y(n_925)
);

INVx3_ASAP7_75t_L g926 ( 
.A(n_647),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_698),
.B(n_700),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_698),
.A2(n_525),
.B(n_528),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_656),
.B(n_506),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_700),
.A2(n_586),
.B(n_528),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_764),
.A2(n_586),
.B(n_528),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_666),
.B(n_506),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_674),
.B(n_506),
.Y(n_933)
);

OAI22xp5_ASAP7_75t_L g934 ( 
.A1(n_688),
.A2(n_591),
.B1(n_589),
.B2(n_574),
.Y(n_934)
);

AND2x4_ASAP7_75t_L g935 ( 
.A(n_779),
.B(n_765),
.Y(n_935)
);

INVxp67_ASAP7_75t_L g936 ( 
.A(n_704),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_764),
.A2(n_586),
.B(n_528),
.Y(n_937)
);

O2A1O1Ixp33_ASAP7_75t_L g938 ( 
.A1(n_776),
.A2(n_676),
.B(n_681),
.C(n_692),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_705),
.B(n_574),
.Y(n_939)
);

OAI21xp5_ASAP7_75t_L g940 ( 
.A1(n_752),
.A2(n_591),
.B(n_589),
.Y(n_940)
);

OR2x6_ASAP7_75t_L g941 ( 
.A(n_704),
.B(n_720),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_766),
.A2(n_586),
.B(n_528),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_708),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_710),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_766),
.A2(n_586),
.B(n_589),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_724),
.A2(n_586),
.B(n_576),
.Y(n_946)
);

O2A1O1Ixp33_ASAP7_75t_L g947 ( 
.A1(n_717),
.A2(n_405),
.B(n_406),
.C(n_401),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_SL g948 ( 
.A(n_704),
.B(n_209),
.Y(n_948)
);

BUFx6f_ASAP7_75t_L g949 ( 
.A(n_714),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_714),
.A2(n_576),
.B(n_574),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_719),
.B(n_576),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_714),
.A2(n_404),
.B(n_402),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_727),
.B(n_735),
.Y(n_953)
);

NOR2xp33_ASAP7_75t_L g954 ( 
.A(n_720),
.B(n_287),
.Y(n_954)
);

OAI21xp5_ASAP7_75t_L g955 ( 
.A1(n_731),
.A2(n_401),
.B(n_403),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_721),
.B(n_429),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_729),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_760),
.A2(n_402),
.B(n_404),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_762),
.A2(n_404),
.B(n_411),
.Y(n_959)
);

NAND2x1_ASAP7_75t_L g960 ( 
.A(n_729),
.B(n_404),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_L g961 ( 
.A(n_706),
.B(n_8),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_768),
.A2(n_404),
.B(n_411),
.Y(n_962)
);

AND2x2_ASAP7_75t_L g963 ( 
.A(n_774),
.B(n_733),
.Y(n_963)
);

NAND2x1p5_ASAP7_75t_L g964 ( 
.A(n_771),
.B(n_778),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_799),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_784),
.A2(n_748),
.B(n_744),
.Y(n_966)
);

O2A1O1Ixp33_ASAP7_75t_SL g967 ( 
.A1(n_808),
.A2(n_744),
.B(n_748),
.C(n_771),
.Y(n_967)
);

AND2x4_ASAP7_75t_L g968 ( 
.A(n_906),
.B(n_733),
.Y(n_968)
);

O2A1O1Ixp33_ASAP7_75t_L g969 ( 
.A1(n_961),
.A2(n_725),
.B(n_728),
.C(n_734),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_SL g970 ( 
.A(n_820),
.B(n_740),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_SL g971 ( 
.A(n_879),
.B(n_740),
.Y(n_971)
);

O2A1O1Ixp33_ASAP7_75t_L g972 ( 
.A1(n_961),
.A2(n_725),
.B(n_728),
.C(n_734),
.Y(n_972)
);

XOR2x2_ASAP7_75t_SL g973 ( 
.A(n_853),
.B(n_291),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_801),
.A2(n_778),
.B(n_722),
.Y(n_974)
);

INVx3_ASAP7_75t_L g975 ( 
.A(n_866),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_803),
.B(n_753),
.Y(n_976)
);

A2O1A1Ixp33_ASAP7_75t_SL g977 ( 
.A1(n_869),
.A2(n_954),
.B(n_811),
.C(n_902),
.Y(n_977)
);

OAI22xp5_ASAP7_75t_L g978 ( 
.A1(n_839),
.A2(n_770),
.B1(n_753),
.B2(n_781),
.Y(n_978)
);

OAI22xp5_ASAP7_75t_L g979 ( 
.A1(n_839),
.A2(n_837),
.B1(n_909),
.B2(n_941),
.Y(n_979)
);

A2O1A1Ixp33_ASAP7_75t_L g980 ( 
.A1(n_869),
.A2(n_781),
.B(n_770),
.C(n_756),
.Y(n_980)
);

BUFx6f_ASAP7_75t_L g981 ( 
.A(n_906),
.Y(n_981)
);

A2O1A1Ixp33_ASAP7_75t_SL g982 ( 
.A1(n_954),
.A2(n_754),
.B(n_742),
.C(n_444),
.Y(n_982)
);

AOI21x1_ASAP7_75t_L g983 ( 
.A1(n_922),
.A2(n_403),
.B(n_405),
.Y(n_983)
);

BUFx6f_ASAP7_75t_L g984 ( 
.A(n_906),
.Y(n_984)
);

HB1xp67_ASAP7_75t_L g985 ( 
.A(n_844),
.Y(n_985)
);

INVx4_ASAP7_75t_L g986 ( 
.A(n_825),
.Y(n_986)
);

OAI22xp33_ASAP7_75t_L g987 ( 
.A1(n_948),
.A2(n_433),
.B1(n_430),
.B2(n_422),
.Y(n_987)
);

BUFx6f_ASAP7_75t_L g988 ( 
.A(n_906),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_803),
.B(n_403),
.Y(n_989)
);

AND2x4_ASAP7_75t_L g990 ( 
.A(n_805),
.B(n_430),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_815),
.B(n_405),
.Y(n_991)
);

AND2x6_ASAP7_75t_L g992 ( 
.A(n_927),
.B(n_406),
.Y(n_992)
);

O2A1O1Ixp33_ASAP7_75t_L g993 ( 
.A1(n_811),
.A2(n_444),
.B(n_437),
.C(n_408),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_816),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_843),
.Y(n_995)
);

OAI22xp5_ASAP7_75t_L g996 ( 
.A1(n_909),
.A2(n_941),
.B1(n_908),
.B2(n_828),
.Y(n_996)
);

BUFx2_ASAP7_75t_L g997 ( 
.A(n_818),
.Y(n_997)
);

BUFx6f_ASAP7_75t_L g998 ( 
.A(n_866),
.Y(n_998)
);

OAI21xp33_ASAP7_75t_SL g999 ( 
.A1(n_927),
.A2(n_444),
.B(n_437),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_792),
.B(n_406),
.Y(n_1000)
);

INVxp67_ASAP7_75t_L g1001 ( 
.A(n_844),
.Y(n_1001)
);

CKINVDCx8_ASAP7_75t_R g1002 ( 
.A(n_785),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_800),
.Y(n_1003)
);

OR2x2_ASAP7_75t_L g1004 ( 
.A(n_865),
.B(n_415),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_867),
.B(n_408),
.Y(n_1005)
);

A2O1A1Ixp33_ASAP7_75t_SL g1006 ( 
.A1(n_883),
.A2(n_408),
.B(n_418),
.C(n_415),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_812),
.A2(n_404),
.B(n_411),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_871),
.Y(n_1008)
);

INVx4_ASAP7_75t_L g1009 ( 
.A(n_825),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_872),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_877),
.B(n_418),
.Y(n_1011)
);

OR2x2_ASAP7_75t_L g1012 ( 
.A(n_809),
.B(n_418),
.Y(n_1012)
);

O2A1O1Ixp33_ASAP7_75t_L g1013 ( 
.A1(n_840),
.A2(n_415),
.B(n_435),
.C(n_424),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_836),
.A2(n_411),
.B(n_417),
.Y(n_1014)
);

NAND3xp33_ASAP7_75t_L g1015 ( 
.A(n_855),
.B(n_436),
.C(n_435),
.Y(n_1015)
);

OAI22xp5_ASAP7_75t_L g1016 ( 
.A1(n_941),
.A2(n_436),
.B1(n_435),
.B2(n_424),
.Y(n_1016)
);

OAI21x1_ASAP7_75t_L g1017 ( 
.A1(n_920),
.A2(n_436),
.B(n_435),
.Y(n_1017)
);

HB1xp67_ASAP7_75t_L g1018 ( 
.A(n_857),
.Y(n_1018)
);

INVx2_ASAP7_75t_SL g1019 ( 
.A(n_787),
.Y(n_1019)
);

OAI22xp5_ASAP7_75t_L g1020 ( 
.A1(n_908),
.A2(n_436),
.B1(n_424),
.B2(n_417),
.Y(n_1020)
);

AOI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_883),
.A2(n_424),
.B1(n_429),
.B2(n_417),
.Y(n_1021)
);

BUFx3_ASAP7_75t_L g1022 ( 
.A(n_878),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_786),
.A2(n_417),
.B(n_416),
.Y(n_1023)
);

HB1xp67_ASAP7_75t_L g1024 ( 
.A(n_857),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_R g1025 ( 
.A(n_863),
.B(n_874),
.Y(n_1025)
);

OAI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_806),
.A2(n_416),
.B(n_429),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_832),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_793),
.A2(n_416),
.B(n_162),
.Y(n_1028)
);

AOI22xp33_ASAP7_75t_L g1029 ( 
.A1(n_902),
.A2(n_291),
.B1(n_416),
.B2(n_12),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_831),
.Y(n_1030)
);

OAI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_852),
.A2(n_124),
.B(n_155),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_885),
.B(n_152),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_834),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_851),
.Y(n_1034)
);

A2O1A1Ixp33_ASAP7_75t_L g1035 ( 
.A1(n_881),
.A2(n_291),
.B(n_10),
.C(n_13),
.Y(n_1035)
);

AOI22xp5_ASAP7_75t_L g1036 ( 
.A1(n_897),
.A2(n_291),
.B1(n_149),
.B2(n_143),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_SL g1037 ( 
.A(n_790),
.B(n_825),
.Y(n_1037)
);

A2O1A1Ixp33_ASAP7_75t_L g1038 ( 
.A1(n_938),
.A2(n_9),
.B(n_14),
.C(n_15),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_794),
.A2(n_142),
.B(n_141),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_873),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_SL g1041 ( 
.A(n_825),
.B(n_858),
.Y(n_1041)
);

NOR2xp67_ASAP7_75t_SL g1042 ( 
.A(n_949),
.B(n_14),
.Y(n_1042)
);

NOR3xp33_ASAP7_75t_L g1043 ( 
.A(n_887),
.B(n_16),
.C(n_17),
.Y(n_1043)
);

BUFx3_ASAP7_75t_L g1044 ( 
.A(n_805),
.Y(n_1044)
);

INVx4_ASAP7_75t_L g1045 ( 
.A(n_858),
.Y(n_1045)
);

BUFx6f_ASAP7_75t_L g1046 ( 
.A(n_866),
.Y(n_1046)
);

AOI22xp33_ASAP7_75t_L g1047 ( 
.A1(n_936),
.A2(n_935),
.B1(n_907),
.B2(n_814),
.Y(n_1047)
);

BUFx12f_ASAP7_75t_L g1048 ( 
.A(n_866),
.Y(n_1048)
);

INVx3_ASAP7_75t_L g1049 ( 
.A(n_858),
.Y(n_1049)
);

BUFx6f_ASAP7_75t_SL g1050 ( 
.A(n_795),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_912),
.B(n_138),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_915),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_914),
.Y(n_1053)
);

AOI22xp5_ASAP7_75t_L g1054 ( 
.A1(n_936),
.A2(n_136),
.B1(n_135),
.B2(n_112),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_875),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_835),
.A2(n_798),
.B(n_845),
.Y(n_1056)
);

AND2x6_ASAP7_75t_L g1057 ( 
.A(n_858),
.B(n_108),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_835),
.A2(n_103),
.B(n_87),
.Y(n_1058)
);

A2O1A1Ixp33_ASAP7_75t_L g1059 ( 
.A1(n_855),
.A2(n_19),
.B(n_20),
.C(n_21),
.Y(n_1059)
);

OAI22x1_ASAP7_75t_L g1060 ( 
.A1(n_905),
.A2(n_21),
.B1(n_22),
.B2(n_24),
.Y(n_1060)
);

AND2x2_ASAP7_75t_L g1061 ( 
.A(n_809),
.B(n_861),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_845),
.A2(n_86),
.B(n_85),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_917),
.Y(n_1063)
);

OAI21xp33_ASAP7_75t_L g1064 ( 
.A1(n_861),
.A2(n_22),
.B(n_25),
.Y(n_1064)
);

NOR2xp33_ASAP7_75t_SL g1065 ( 
.A(n_935),
.B(n_78),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_919),
.B(n_73),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_856),
.A2(n_72),
.B(n_29),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_904),
.B(n_27),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_918),
.B(n_29),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_923),
.B(n_953),
.Y(n_1070)
);

BUFx3_ASAP7_75t_L g1071 ( 
.A(n_795),
.Y(n_1071)
);

O2A1O1Ixp5_ASAP7_75t_SL g1072 ( 
.A1(n_783),
.A2(n_36),
.B(n_37),
.C(n_38),
.Y(n_1072)
);

BUFx3_ASAP7_75t_L g1073 ( 
.A(n_943),
.Y(n_1073)
);

OAI22xp5_ASAP7_75t_SL g1074 ( 
.A1(n_944),
.A2(n_38),
.B1(n_40),
.B2(n_43),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_838),
.B(n_43),
.Y(n_1075)
);

AOI21x1_ASAP7_75t_L g1076 ( 
.A1(n_889),
.A2(n_910),
.B(n_900),
.Y(n_1076)
);

OR2x2_ASAP7_75t_L g1077 ( 
.A(n_891),
.B(n_45),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_957),
.Y(n_1078)
);

AOI21x1_ASAP7_75t_L g1079 ( 
.A1(n_899),
.A2(n_46),
.B(n_49),
.Y(n_1079)
);

OR2x6_ASAP7_75t_L g1080 ( 
.A(n_807),
.B(n_49),
.Y(n_1080)
);

NOR3xp33_ASAP7_75t_L g1081 ( 
.A(n_804),
.B(n_50),
.C(n_51),
.Y(n_1081)
);

OAI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_888),
.A2(n_53),
.B(n_54),
.Y(n_1082)
);

NOR2xp33_ASAP7_75t_L g1083 ( 
.A(n_891),
.B(n_913),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_SL g1084 ( 
.A(n_814),
.B(n_913),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_SL g1085 ( 
.A(n_926),
.B(n_59),
.Y(n_1085)
);

NAND2x1p5_ASAP7_75t_L g1086 ( 
.A(n_949),
.B(n_60),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_807),
.Y(n_1087)
);

INVx3_ASAP7_75t_L g1088 ( 
.A(n_829),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_856),
.A2(n_60),
.B(n_61),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_924),
.B(n_62),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_926),
.B(n_64),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_SL g1092 ( 
.A(n_963),
.B(n_64),
.Y(n_1092)
);

NAND2xp33_ASAP7_75t_SL g1093 ( 
.A(n_813),
.B(n_949),
.Y(n_1093)
);

OAI22xp5_ASAP7_75t_L g1094 ( 
.A1(n_876),
.A2(n_964),
.B1(n_823),
.B2(n_789),
.Y(n_1094)
);

A2O1A1Ixp33_ASAP7_75t_L g1095 ( 
.A1(n_826),
.A2(n_810),
.B(n_888),
.C(n_796),
.Y(n_1095)
);

AND2x4_ASAP7_75t_L g1096 ( 
.A(n_829),
.B(n_846),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_925),
.Y(n_1097)
);

AND2x2_ASAP7_75t_L g1098 ( 
.A(n_846),
.B(n_964),
.Y(n_1098)
);

INVx1_ASAP7_75t_SL g1099 ( 
.A(n_939),
.Y(n_1099)
);

NOR2x1_ASAP7_75t_L g1100 ( 
.A(n_886),
.B(n_898),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_949),
.A2(n_791),
.B(n_842),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_951),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_788),
.A2(n_911),
.B(n_827),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_821),
.A2(n_895),
.B(n_940),
.Y(n_1104)
);

INVx3_ASAP7_75t_L g1105 ( 
.A(n_882),
.Y(n_1105)
);

OAI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_884),
.A2(n_894),
.B(n_903),
.Y(n_1106)
);

O2A1O1Ixp33_ASAP7_75t_L g1107 ( 
.A1(n_934),
.A2(n_947),
.B(n_854),
.C(n_830),
.Y(n_1107)
);

AOI22xp5_ASAP7_75t_L g1108 ( 
.A1(n_817),
.A2(n_898),
.B1(n_886),
.B2(n_870),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_SL g1109 ( 
.A(n_929),
.B(n_932),
.Y(n_1109)
);

AOI22x1_ASAP7_75t_L g1110 ( 
.A1(n_848),
.A2(n_849),
.B1(n_862),
.B2(n_880),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_SL g1111 ( 
.A(n_933),
.B(n_901),
.Y(n_1111)
);

A2O1A1Ixp33_ASAP7_75t_L g1112 ( 
.A1(n_797),
.A2(n_824),
.B(n_819),
.C(n_802),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_859),
.B(n_868),
.Y(n_1113)
);

INVx3_ASAP7_75t_L g1114 ( 
.A(n_882),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_833),
.A2(n_841),
.B(n_847),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_864),
.A2(n_850),
.B(n_860),
.Y(n_1116)
);

BUFx12f_ASAP7_75t_L g1117 ( 
.A(n_1027),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_1104),
.A2(n_870),
.B(n_921),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_965),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_1099),
.B(n_916),
.Y(n_1120)
);

INVx3_ASAP7_75t_SL g1121 ( 
.A(n_1052),
.Y(n_1121)
);

NAND2x1p5_ASAP7_75t_L g1122 ( 
.A(n_997),
.B(n_960),
.Y(n_1122)
);

A2O1A1Ixp33_ASAP7_75t_L g1123 ( 
.A1(n_977),
.A2(n_824),
.B(n_946),
.C(n_958),
.Y(n_1123)
);

INVx1_ASAP7_75t_SL g1124 ( 
.A(n_985),
.Y(n_1124)
);

OA22x2_ASAP7_75t_L g1125 ( 
.A1(n_1074),
.A2(n_955),
.B1(n_896),
.B2(n_956),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_1061),
.B(n_890),
.Y(n_1126)
);

OAI21xp5_ASAP7_75t_SL g1127 ( 
.A1(n_1029),
.A2(n_892),
.B(n_893),
.Y(n_1127)
);

AND2x4_ASAP7_75t_L g1128 ( 
.A(n_1071),
.B(n_822),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_1070),
.B(n_962),
.Y(n_1129)
);

O2A1O1Ixp33_ASAP7_75t_L g1130 ( 
.A1(n_1084),
.A2(n_956),
.B(n_959),
.C(n_945),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_1104),
.A2(n_928),
.B(n_930),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_994),
.Y(n_1132)
);

NAND2x1p5_ASAP7_75t_L g1133 ( 
.A(n_981),
.B(n_950),
.Y(n_1133)
);

OAI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_970),
.A2(n_931),
.B(n_937),
.Y(n_1134)
);

OAI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_1106),
.A2(n_942),
.B(n_952),
.Y(n_1135)
);

INVx3_ASAP7_75t_L g1136 ( 
.A(n_1096),
.Y(n_1136)
);

OAI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_971),
.A2(n_999),
.B(n_1103),
.Y(n_1137)
);

OAI22xp5_ASAP7_75t_L g1138 ( 
.A1(n_1070),
.A2(n_979),
.B1(n_1073),
.B2(n_1102),
.Y(n_1138)
);

BUFx3_ASAP7_75t_L g1139 ( 
.A(n_1022),
.Y(n_1139)
);

NOR2xp33_ASAP7_75t_L g1140 ( 
.A(n_1001),
.B(n_1018),
.Y(n_1140)
);

A2O1A1Ixp33_ASAP7_75t_L g1141 ( 
.A1(n_969),
.A2(n_972),
.B(n_1077),
.C(n_1031),
.Y(n_1141)
);

OAI21x1_ASAP7_75t_L g1142 ( 
.A1(n_1017),
.A2(n_1076),
.B(n_1056),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_995),
.Y(n_1143)
);

OAI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_1103),
.A2(n_1095),
.B(n_974),
.Y(n_1144)
);

OAI22xp5_ASAP7_75t_L g1145 ( 
.A1(n_979),
.A2(n_1047),
.B1(n_996),
.B2(n_1108),
.Y(n_1145)
);

AND2x6_ASAP7_75t_L g1146 ( 
.A(n_1098),
.B(n_981),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1008),
.Y(n_1147)
);

AOI221x1_ASAP7_75t_L g1148 ( 
.A1(n_1035),
.A2(n_1064),
.B1(n_1038),
.B2(n_1081),
.C(n_1082),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_SL g1149 ( 
.A(n_973),
.B(n_1019),
.Y(n_1149)
);

A2O1A1Ixp33_ASAP7_75t_L g1150 ( 
.A1(n_1075),
.A2(n_1107),
.B(n_1116),
.C(n_1093),
.Y(n_1150)
);

O2A1O1Ixp5_ASAP7_75t_L g1151 ( 
.A1(n_1028),
.A2(n_1075),
.B(n_1037),
.C(n_982),
.Y(n_1151)
);

OAI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_1116),
.A2(n_966),
.B(n_980),
.Y(n_1152)
);

BUFx6f_ASAP7_75t_L g1153 ( 
.A(n_1048),
.Y(n_1153)
);

OAI21x1_ASAP7_75t_L g1154 ( 
.A1(n_1110),
.A2(n_1101),
.B(n_1023),
.Y(n_1154)
);

BUFx10_ASAP7_75t_L g1155 ( 
.A(n_1050),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_1115),
.A2(n_1112),
.B(n_1109),
.Y(n_1156)
);

INVx8_ASAP7_75t_L g1157 ( 
.A(n_998),
.Y(n_1157)
);

AO31x2_ASAP7_75t_L g1158 ( 
.A1(n_1115),
.A2(n_1094),
.A3(n_1016),
.B(n_978),
.Y(n_1158)
);

BUFx10_ASAP7_75t_L g1159 ( 
.A(n_1050),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1097),
.B(n_976),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_1113),
.A2(n_1111),
.B(n_1094),
.Y(n_1161)
);

OAI21x1_ASAP7_75t_L g1162 ( 
.A1(n_983),
.A2(n_1014),
.B(n_1026),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1113),
.A2(n_976),
.B(n_991),
.Y(n_1163)
);

AND2x4_ASAP7_75t_L g1164 ( 
.A(n_1044),
.B(n_981),
.Y(n_1164)
);

OA21x2_ASAP7_75t_L g1165 ( 
.A1(n_989),
.A2(n_1090),
.B(n_1007),
.Y(n_1165)
);

OA21x2_ASAP7_75t_L g1166 ( 
.A1(n_989),
.A2(n_1090),
.B(n_1068),
.Y(n_1166)
);

AND2x4_ASAP7_75t_L g1167 ( 
.A(n_984),
.B(n_988),
.Y(n_1167)
);

AO31x2_ASAP7_75t_L g1168 ( 
.A1(n_1016),
.A2(n_978),
.A3(n_996),
.B(n_1020),
.Y(n_1168)
);

OAI21x1_ASAP7_75t_SL g1169 ( 
.A1(n_1089),
.A2(n_1067),
.B(n_1058),
.Y(n_1169)
);

AND2x4_ASAP7_75t_L g1170 ( 
.A(n_984),
.B(n_988),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_991),
.A2(n_967),
.B(n_1039),
.Y(n_1171)
);

INVxp67_ASAP7_75t_SL g1172 ( 
.A(n_1024),
.Y(n_1172)
);

OR2x2_ASAP7_75t_L g1173 ( 
.A(n_1004),
.B(n_1012),
.Y(n_1173)
);

NAND3xp33_ASAP7_75t_SL g1174 ( 
.A(n_1043),
.B(n_1059),
.C(n_1036),
.Y(n_1174)
);

OA21x2_ASAP7_75t_L g1175 ( 
.A1(n_1068),
.A2(n_1015),
.B(n_1005),
.Y(n_1175)
);

HB1xp67_ASAP7_75t_L g1176 ( 
.A(n_1087),
.Y(n_1176)
);

OAI21x1_ASAP7_75t_L g1177 ( 
.A1(n_1032),
.A2(n_1066),
.B(n_1051),
.Y(n_1177)
);

NOR2xp33_ASAP7_75t_L g1178 ( 
.A(n_1092),
.B(n_990),
.Y(n_1178)
);

OAI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1072),
.A2(n_1021),
.B(n_1020),
.Y(n_1179)
);

BUFx2_ASAP7_75t_L g1180 ( 
.A(n_984),
.Y(n_1180)
);

NAND2x1p5_ASAP7_75t_L g1181 ( 
.A(n_988),
.B(n_1009),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1032),
.A2(n_1051),
.B(n_1066),
.Y(n_1182)
);

O2A1O1Ixp33_ASAP7_75t_SL g1183 ( 
.A1(n_1006),
.A2(n_1085),
.B(n_1069),
.C(n_1041),
.Y(n_1183)
);

INVx2_ASAP7_75t_SL g1184 ( 
.A(n_1025),
.Y(n_1184)
);

NAND3xp33_ASAP7_75t_L g1185 ( 
.A(n_1091),
.B(n_1069),
.C(n_1065),
.Y(n_1185)
);

OAI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_992),
.A2(n_993),
.B(n_1011),
.Y(n_1186)
);

OAI21x1_ASAP7_75t_SL g1187 ( 
.A1(n_1079),
.A2(n_1062),
.B(n_1054),
.Y(n_1187)
);

OR2x2_ASAP7_75t_L g1188 ( 
.A(n_1003),
.B(n_1030),
.Y(n_1188)
);

BUFx6f_ASAP7_75t_L g1189 ( 
.A(n_998),
.Y(n_1189)
);

BUFx12f_ASAP7_75t_L g1190 ( 
.A(n_1080),
.Y(n_1190)
);

A2O1A1Ixp33_ASAP7_75t_L g1191 ( 
.A1(n_1010),
.A2(n_1053),
.B(n_1063),
.C(n_968),
.Y(n_1191)
);

AOI221x1_ASAP7_75t_L g1192 ( 
.A1(n_1060),
.A2(n_1005),
.B1(n_1011),
.B2(n_1000),
.C(n_1078),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_987),
.A2(n_1100),
.B(n_1105),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1105),
.A2(n_1114),
.B(n_1000),
.Y(n_1194)
);

AOI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_1114),
.A2(n_968),
.B(n_1096),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1088),
.A2(n_1045),
.B(n_986),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1033),
.B(n_1055),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1088),
.A2(n_986),
.B(n_1045),
.Y(n_1198)
);

AO31x2_ASAP7_75t_L g1199 ( 
.A1(n_1034),
.A2(n_1040),
.A3(n_1009),
.B(n_992),
.Y(n_1199)
);

O2A1O1Ixp33_ASAP7_75t_SL g1200 ( 
.A1(n_1049),
.A2(n_975),
.B(n_1013),
.C(n_1042),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_975),
.Y(n_1201)
);

NAND3xp33_ASAP7_75t_L g1202 ( 
.A(n_1080),
.B(n_998),
.C(n_1046),
.Y(n_1202)
);

OAI21x1_ASAP7_75t_L g1203 ( 
.A1(n_1049),
.A2(n_1086),
.B(n_992),
.Y(n_1203)
);

AND2x2_ASAP7_75t_L g1204 ( 
.A(n_1086),
.B(n_1046),
.Y(n_1204)
);

AOI22xp5_ASAP7_75t_L g1205 ( 
.A1(n_992),
.A2(n_1057),
.B1(n_1046),
.B2(n_1002),
.Y(n_1205)
);

HB1xp67_ASAP7_75t_L g1206 ( 
.A(n_992),
.Y(n_1206)
);

OAI21x1_ASAP7_75t_L g1207 ( 
.A1(n_1057),
.A2(n_1017),
.B(n_1076),
.Y(n_1207)
);

BUFx6f_ASAP7_75t_L g1208 ( 
.A(n_1057),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1057),
.B(n_1083),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1057),
.B(n_1083),
.Y(n_1210)
);

AND2x2_ASAP7_75t_L g1211 ( 
.A(n_1061),
.B(n_679),
.Y(n_1211)
);

OAI21x1_ASAP7_75t_L g1212 ( 
.A1(n_1017),
.A2(n_1076),
.B(n_1056),
.Y(n_1212)
);

AOI221xp5_ASAP7_75t_SL g1213 ( 
.A1(n_1064),
.A2(n_1035),
.B1(n_675),
.B2(n_745),
.C(n_1083),
.Y(n_1213)
);

OAI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1083),
.A2(n_1106),
.B(n_678),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1083),
.B(n_675),
.Y(n_1215)
);

A2O1A1Ixp33_ASAP7_75t_L g1216 ( 
.A1(n_1083),
.A2(n_675),
.B(n_820),
.C(n_869),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1104),
.A2(n_668),
.B(n_667),
.Y(n_1217)
);

OAI22x1_ASAP7_75t_L g1218 ( 
.A1(n_1083),
.A2(n_675),
.B1(n_478),
.B2(n_1092),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1083),
.B(n_675),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_1025),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1083),
.B(n_675),
.Y(n_1221)
);

BUFx3_ASAP7_75t_L g1222 ( 
.A(n_997),
.Y(n_1222)
);

AO21x2_ASAP7_75t_L g1223 ( 
.A1(n_1104),
.A2(n_1115),
.B(n_1116),
.Y(n_1223)
);

AO31x2_ASAP7_75t_L g1224 ( 
.A1(n_1104),
.A2(n_1112),
.A3(n_1115),
.B(n_1103),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_SL g1225 ( 
.A(n_1083),
.B(n_679),
.Y(n_1225)
);

OR2x2_ASAP7_75t_L g1226 ( 
.A(n_997),
.B(n_565),
.Y(n_1226)
);

AOI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1104),
.A2(n_668),
.B(n_667),
.Y(n_1227)
);

A2O1A1Ixp33_ASAP7_75t_L g1228 ( 
.A1(n_1083),
.A2(n_675),
.B(n_820),
.C(n_869),
.Y(n_1228)
);

NOR2x1_ASAP7_75t_R g1229 ( 
.A(n_1027),
.B(n_439),
.Y(n_1229)
);

AO21x1_ASAP7_75t_L g1230 ( 
.A1(n_1083),
.A2(n_820),
.B(n_675),
.Y(n_1230)
);

OAI21x1_ASAP7_75t_L g1231 ( 
.A1(n_1017),
.A2(n_1076),
.B(n_1056),
.Y(n_1231)
);

A2O1A1Ixp33_ASAP7_75t_L g1232 ( 
.A1(n_1083),
.A2(n_675),
.B(n_820),
.C(n_869),
.Y(n_1232)
);

OR2x6_ASAP7_75t_L g1233 ( 
.A(n_1048),
.B(n_906),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1104),
.A2(n_668),
.B(n_667),
.Y(n_1234)
);

OAI21x1_ASAP7_75t_L g1235 ( 
.A1(n_1017),
.A2(n_1076),
.B(n_1056),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1083),
.B(n_675),
.Y(n_1236)
);

INVx1_ASAP7_75t_SL g1237 ( 
.A(n_997),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_SL g1238 ( 
.A(n_1083),
.B(n_679),
.Y(n_1238)
);

OAI21x1_ASAP7_75t_L g1239 ( 
.A1(n_1017),
.A2(n_1076),
.B(n_1056),
.Y(n_1239)
);

AO32x2_ASAP7_75t_L g1240 ( 
.A1(n_979),
.A2(n_996),
.A3(n_1094),
.B1(n_1016),
.B2(n_783),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1104),
.A2(n_668),
.B(n_667),
.Y(n_1241)
);

AOI22xp5_ASAP7_75t_L g1242 ( 
.A1(n_1083),
.A2(n_675),
.B1(n_961),
.B2(n_853),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_965),
.Y(n_1243)
);

NAND2x1p5_ASAP7_75t_L g1244 ( 
.A(n_997),
.B(n_825),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1104),
.A2(n_668),
.B(n_667),
.Y(n_1245)
);

NOR2x1_ASAP7_75t_SL g1246 ( 
.A(n_1037),
.B(n_941),
.Y(n_1246)
);

INVx2_ASAP7_75t_SL g1247 ( 
.A(n_997),
.Y(n_1247)
);

O2A1O1Ixp33_ASAP7_75t_SL g1248 ( 
.A1(n_977),
.A2(n_1035),
.B(n_1083),
.C(n_1038),
.Y(n_1248)
);

BUFx3_ASAP7_75t_L g1249 ( 
.A(n_997),
.Y(n_1249)
);

AO21x2_ASAP7_75t_L g1250 ( 
.A1(n_1104),
.A2(n_1115),
.B(n_1116),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1104),
.A2(n_668),
.B(n_667),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1083),
.B(n_675),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_L g1253 ( 
.A1(n_1017),
.A2(n_1076),
.B(n_1056),
.Y(n_1253)
);

O2A1O1Ixp33_ASAP7_75t_SL g1254 ( 
.A1(n_977),
.A2(n_1035),
.B(n_1083),
.C(n_1038),
.Y(n_1254)
);

A2O1A1Ixp33_ASAP7_75t_L g1255 ( 
.A1(n_1083),
.A2(n_675),
.B(n_820),
.C(n_869),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1104),
.A2(n_668),
.B(n_667),
.Y(n_1256)
);

AOI22xp5_ASAP7_75t_L g1257 ( 
.A1(n_1083),
.A2(n_675),
.B1(n_961),
.B2(n_853),
.Y(n_1257)
);

AO32x2_ASAP7_75t_L g1258 ( 
.A1(n_979),
.A2(n_996),
.A3(n_1094),
.B1(n_1016),
.B2(n_783),
.Y(n_1258)
);

AOI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1104),
.A2(n_668),
.B(n_667),
.Y(n_1259)
);

AO32x2_ASAP7_75t_L g1260 ( 
.A1(n_979),
.A2(n_996),
.A3(n_1094),
.B1(n_1016),
.B2(n_783),
.Y(n_1260)
);

AO31x2_ASAP7_75t_L g1261 ( 
.A1(n_1104),
.A2(n_1112),
.A3(n_1115),
.B(n_1103),
.Y(n_1261)
);

AOI31xp67_ASAP7_75t_L g1262 ( 
.A1(n_971),
.A2(n_820),
.A3(n_970),
.B(n_1021),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1104),
.A2(n_668),
.B(n_667),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_965),
.Y(n_1264)
);

NOR2xp33_ASAP7_75t_L g1265 ( 
.A(n_1083),
.B(n_675),
.Y(n_1265)
);

AOI22xp5_ASAP7_75t_L g1266 ( 
.A1(n_1083),
.A2(n_675),
.B1(n_961),
.B2(n_853),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1188),
.Y(n_1267)
);

AOI22xp33_ASAP7_75t_L g1268 ( 
.A1(n_1265),
.A2(n_1230),
.B1(n_1242),
.B2(n_1257),
.Y(n_1268)
);

CKINVDCx6p67_ASAP7_75t_R g1269 ( 
.A(n_1121),
.Y(n_1269)
);

OAI22xp33_ASAP7_75t_L g1270 ( 
.A1(n_1242),
.A2(n_1266),
.B1(n_1257),
.B2(n_1236),
.Y(n_1270)
);

BUFx3_ASAP7_75t_L g1271 ( 
.A(n_1222),
.Y(n_1271)
);

AOI22xp33_ASAP7_75t_SL g1272 ( 
.A1(n_1215),
.A2(n_1221),
.B1(n_1252),
.B2(n_1219),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1266),
.B(n_1216),
.Y(n_1273)
);

CKINVDCx20_ASAP7_75t_R g1274 ( 
.A(n_1220),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_1117),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1228),
.B(n_1232),
.Y(n_1276)
);

AOI22xp33_ASAP7_75t_SL g1277 ( 
.A1(n_1214),
.A2(n_1145),
.B1(n_1125),
.B2(n_1190),
.Y(n_1277)
);

BUFx2_ASAP7_75t_L g1278 ( 
.A(n_1249),
.Y(n_1278)
);

AOI22xp33_ASAP7_75t_SL g1279 ( 
.A1(n_1214),
.A2(n_1208),
.B1(n_1185),
.B2(n_1255),
.Y(n_1279)
);

AOI22xp33_ASAP7_75t_SL g1280 ( 
.A1(n_1208),
.A2(n_1185),
.B1(n_1209),
.B2(n_1210),
.Y(n_1280)
);

BUFx8_ASAP7_75t_L g1281 ( 
.A(n_1153),
.Y(n_1281)
);

INVx6_ASAP7_75t_L g1282 ( 
.A(n_1155),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_1174),
.A2(n_1218),
.B1(n_1211),
.B2(n_1225),
.Y(n_1283)
);

CKINVDCx6p67_ASAP7_75t_R g1284 ( 
.A(n_1139),
.Y(n_1284)
);

INVx6_ASAP7_75t_L g1285 ( 
.A(n_1155),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1132),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1173),
.B(n_1120),
.Y(n_1287)
);

AOI22xp33_ASAP7_75t_L g1288 ( 
.A1(n_1178),
.A2(n_1238),
.B1(n_1149),
.B2(n_1138),
.Y(n_1288)
);

CKINVDCx11_ASAP7_75t_R g1289 ( 
.A(n_1159),
.Y(n_1289)
);

INVx6_ASAP7_75t_L g1290 ( 
.A(n_1159),
.Y(n_1290)
);

AOI22xp33_ASAP7_75t_L g1291 ( 
.A1(n_1206),
.A2(n_1226),
.B1(n_1202),
.B2(n_1237),
.Y(n_1291)
);

BUFx3_ASAP7_75t_L g1292 ( 
.A(n_1247),
.Y(n_1292)
);

AOI22xp33_ASAP7_75t_L g1293 ( 
.A1(n_1202),
.A2(n_1144),
.B1(n_1208),
.B2(n_1126),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1143),
.Y(n_1294)
);

OAI22xp5_ASAP7_75t_L g1295 ( 
.A1(n_1141),
.A2(n_1172),
.B1(n_1124),
.B2(n_1191),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1144),
.A2(n_1176),
.B1(n_1187),
.B2(n_1179),
.Y(n_1296)
);

OAI22xp33_ASAP7_75t_L g1297 ( 
.A1(n_1148),
.A2(n_1205),
.B1(n_1192),
.B2(n_1160),
.Y(n_1297)
);

INVx5_ASAP7_75t_L g1298 ( 
.A(n_1157),
.Y(n_1298)
);

OAI21xp5_ASAP7_75t_SL g1299 ( 
.A1(n_1205),
.A2(n_1150),
.B(n_1179),
.Y(n_1299)
);

BUFx4f_ASAP7_75t_SL g1300 ( 
.A(n_1153),
.Y(n_1300)
);

INVxp67_ASAP7_75t_SL g1301 ( 
.A(n_1163),
.Y(n_1301)
);

INVx1_ASAP7_75t_SL g1302 ( 
.A(n_1140),
.Y(n_1302)
);

AOI22xp33_ASAP7_75t_SL g1303 ( 
.A1(n_1246),
.A2(n_1213),
.B1(n_1186),
.B2(n_1263),
.Y(n_1303)
);

BUFx6f_ASAP7_75t_L g1304 ( 
.A(n_1189),
.Y(n_1304)
);

OAI21xp5_ASAP7_75t_SL g1305 ( 
.A1(n_1186),
.A2(n_1182),
.B(n_1127),
.Y(n_1305)
);

AOI22xp33_ASAP7_75t_L g1306 ( 
.A1(n_1169),
.A2(n_1250),
.B1(n_1223),
.B2(n_1128),
.Y(n_1306)
);

BUFx2_ASAP7_75t_SL g1307 ( 
.A(n_1153),
.Y(n_1307)
);

AOI22xp33_ASAP7_75t_SL g1308 ( 
.A1(n_1213),
.A2(n_1217),
.B1(n_1227),
.B2(n_1251),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1147),
.Y(n_1309)
);

OAI22xp33_ASAP7_75t_L g1310 ( 
.A1(n_1243),
.A2(n_1264),
.B1(n_1129),
.B2(n_1127),
.Y(n_1310)
);

AOI22xp33_ASAP7_75t_L g1311 ( 
.A1(n_1223),
.A2(n_1250),
.B1(n_1128),
.B2(n_1161),
.Y(n_1311)
);

CKINVDCx11_ASAP7_75t_R g1312 ( 
.A(n_1233),
.Y(n_1312)
);

AOI22xp33_ASAP7_75t_SL g1313 ( 
.A1(n_1234),
.A2(n_1241),
.B1(n_1245),
.B2(n_1259),
.Y(n_1313)
);

CKINVDCx20_ASAP7_75t_R g1314 ( 
.A(n_1184),
.Y(n_1314)
);

OAI22xp5_ASAP7_75t_L g1315 ( 
.A1(n_1233),
.A2(n_1193),
.B1(n_1244),
.B2(n_1136),
.Y(n_1315)
);

OAI21xp5_ASAP7_75t_SL g1316 ( 
.A1(n_1156),
.A2(n_1171),
.B(n_1152),
.Y(n_1316)
);

CKINVDCx20_ASAP7_75t_R g1317 ( 
.A(n_1180),
.Y(n_1317)
);

AOI22xp33_ASAP7_75t_SL g1318 ( 
.A1(n_1256),
.A2(n_1152),
.B1(n_1137),
.B2(n_1146),
.Y(n_1318)
);

AOI22xp33_ASAP7_75t_L g1319 ( 
.A1(n_1136),
.A2(n_1166),
.B1(n_1204),
.B2(n_1146),
.Y(n_1319)
);

AOI22xp33_ASAP7_75t_L g1320 ( 
.A1(n_1166),
.A2(n_1146),
.B1(n_1164),
.B2(n_1201),
.Y(n_1320)
);

OAI22xp33_ASAP7_75t_L g1321 ( 
.A1(n_1197),
.A2(n_1233),
.B1(n_1137),
.B2(n_1122),
.Y(n_1321)
);

OAI22xp5_ASAP7_75t_L g1322 ( 
.A1(n_1164),
.A2(n_1195),
.B1(n_1194),
.B2(n_1181),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1248),
.B(n_1254),
.Y(n_1323)
);

BUFx10_ASAP7_75t_L g1324 ( 
.A(n_1167),
.Y(n_1324)
);

CKINVDCx6p67_ASAP7_75t_R g1325 ( 
.A(n_1157),
.Y(n_1325)
);

BUFx6f_ASAP7_75t_L g1326 ( 
.A(n_1157),
.Y(n_1326)
);

OAI22xp5_ASAP7_75t_SL g1327 ( 
.A1(n_1167),
.A2(n_1170),
.B1(n_1229),
.B2(n_1133),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1135),
.A2(n_1175),
.B1(n_1177),
.B2(n_1134),
.Y(n_1328)
);

AOI22xp33_ASAP7_75t_L g1329 ( 
.A1(n_1135),
.A2(n_1175),
.B1(n_1165),
.B2(n_1170),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_SL g1330 ( 
.A1(n_1240),
.A2(n_1260),
.B1(n_1258),
.B2(n_1203),
.Y(n_1330)
);

INVx2_ASAP7_75t_SL g1331 ( 
.A(n_1199),
.Y(n_1331)
);

BUFx6f_ASAP7_75t_L g1332 ( 
.A(n_1207),
.Y(n_1332)
);

AOI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1165),
.A2(n_1118),
.B1(n_1131),
.B2(n_1154),
.Y(n_1333)
);

AOI22xp33_ASAP7_75t_SL g1334 ( 
.A1(n_1240),
.A2(n_1258),
.B1(n_1260),
.B2(n_1262),
.Y(n_1334)
);

CKINVDCx20_ASAP7_75t_R g1335 ( 
.A(n_1229),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1224),
.B(n_1261),
.Y(n_1336)
);

AOI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1151),
.A2(n_1123),
.B(n_1130),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_L g1338 ( 
.A1(n_1196),
.A2(n_1198),
.B1(n_1162),
.B2(n_1253),
.Y(n_1338)
);

INVx6_ASAP7_75t_L g1339 ( 
.A(n_1200),
.Y(n_1339)
);

AOI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1142),
.A2(n_1231),
.B1(n_1235),
.B2(n_1239),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1224),
.Y(n_1341)
);

BUFx6f_ASAP7_75t_L g1342 ( 
.A(n_1240),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1261),
.Y(n_1343)
);

OAI22xp33_ASAP7_75t_L g1344 ( 
.A1(n_1258),
.A2(n_1260),
.B1(n_1158),
.B2(n_1168),
.Y(n_1344)
);

OAI22xp5_ASAP7_75t_L g1345 ( 
.A1(n_1183),
.A2(n_1158),
.B1(n_1168),
.B2(n_1212),
.Y(n_1345)
);

INVx1_ASAP7_75t_SL g1346 ( 
.A(n_1168),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1158),
.Y(n_1347)
);

BUFx6f_ASAP7_75t_L g1348 ( 
.A(n_1208),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1265),
.A2(n_1083),
.B1(n_675),
.B2(n_1230),
.Y(n_1349)
);

AOI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1216),
.A2(n_1232),
.B(n_1228),
.Y(n_1350)
);

AOI22xp33_ASAP7_75t_L g1351 ( 
.A1(n_1265),
.A2(n_1083),
.B1(n_675),
.B2(n_1230),
.Y(n_1351)
);

AOI22xp33_ASAP7_75t_L g1352 ( 
.A1(n_1265),
.A2(n_1083),
.B1(n_675),
.B2(n_1230),
.Y(n_1352)
);

INVx2_ASAP7_75t_SL g1353 ( 
.A(n_1155),
.Y(n_1353)
);

AOI22xp33_ASAP7_75t_L g1354 ( 
.A1(n_1265),
.A2(n_1083),
.B1(n_675),
.B2(n_1230),
.Y(n_1354)
);

AOI22xp5_ASAP7_75t_SL g1355 ( 
.A1(n_1265),
.A2(n_1083),
.B1(n_675),
.B2(n_478),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_1188),
.Y(n_1356)
);

OAI22xp5_ASAP7_75t_L g1357 ( 
.A1(n_1265),
.A2(n_1257),
.B1(n_1266),
.B2(n_1242),
.Y(n_1357)
);

AOI22xp33_ASAP7_75t_L g1358 ( 
.A1(n_1265),
.A2(n_1083),
.B1(n_675),
.B2(n_1230),
.Y(n_1358)
);

BUFx12f_ASAP7_75t_L g1359 ( 
.A(n_1155),
.Y(n_1359)
);

AOI22xp33_ASAP7_75t_L g1360 ( 
.A1(n_1265),
.A2(n_1083),
.B1(n_675),
.B2(n_1230),
.Y(n_1360)
);

CKINVDCx20_ASAP7_75t_R g1361 ( 
.A(n_1121),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1188),
.Y(n_1362)
);

AOI22xp5_ASAP7_75t_L g1363 ( 
.A1(n_1265),
.A2(n_1083),
.B1(n_1257),
.B2(n_1242),
.Y(n_1363)
);

CKINVDCx6p67_ASAP7_75t_R g1364 ( 
.A(n_1121),
.Y(n_1364)
);

AOI22xp33_ASAP7_75t_SL g1365 ( 
.A1(n_1265),
.A2(n_675),
.B1(n_1083),
.B2(n_455),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_1220),
.Y(n_1366)
);

CKINVDCx20_ASAP7_75t_R g1367 ( 
.A(n_1121),
.Y(n_1367)
);

INVx6_ASAP7_75t_L g1368 ( 
.A(n_1155),
.Y(n_1368)
);

CKINVDCx11_ASAP7_75t_R g1369 ( 
.A(n_1121),
.Y(n_1369)
);

INVx1_ASAP7_75t_SL g1370 ( 
.A(n_1237),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1119),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1119),
.Y(n_1372)
);

CKINVDCx20_ASAP7_75t_R g1373 ( 
.A(n_1121),
.Y(n_1373)
);

BUFx2_ASAP7_75t_L g1374 ( 
.A(n_1222),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_1220),
.Y(n_1375)
);

CKINVDCx20_ASAP7_75t_R g1376 ( 
.A(n_1121),
.Y(n_1376)
);

OAI22xp33_ASAP7_75t_L g1377 ( 
.A1(n_1242),
.A2(n_1257),
.B1(n_1266),
.B2(n_1265),
.Y(n_1377)
);

INVx1_ASAP7_75t_SL g1378 ( 
.A(n_1237),
.Y(n_1378)
);

INVxp67_ASAP7_75t_L g1379 ( 
.A(n_1140),
.Y(n_1379)
);

AOI22xp33_ASAP7_75t_L g1380 ( 
.A1(n_1265),
.A2(n_1083),
.B1(n_675),
.B2(n_1230),
.Y(n_1380)
);

BUFx2_ASAP7_75t_L g1381 ( 
.A(n_1222),
.Y(n_1381)
);

AOI22xp33_ASAP7_75t_L g1382 ( 
.A1(n_1265),
.A2(n_1083),
.B1(n_675),
.B2(n_1230),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1188),
.Y(n_1383)
);

BUFx3_ASAP7_75t_L g1384 ( 
.A(n_1222),
.Y(n_1384)
);

INVx6_ASAP7_75t_L g1385 ( 
.A(n_1155),
.Y(n_1385)
);

NAND2x1p5_ASAP7_75t_L g1386 ( 
.A(n_1208),
.B(n_825),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1119),
.Y(n_1387)
);

AOI22xp5_ASAP7_75t_L g1388 ( 
.A1(n_1265),
.A2(n_1083),
.B1(n_1257),
.B2(n_1242),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1119),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1119),
.Y(n_1390)
);

BUFx8_ASAP7_75t_L g1391 ( 
.A(n_1153),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1119),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_L g1393 ( 
.A1(n_1265),
.A2(n_1083),
.B1(n_675),
.B2(n_1230),
.Y(n_1393)
);

CKINVDCx6p67_ASAP7_75t_R g1394 ( 
.A(n_1121),
.Y(n_1394)
);

AO21x2_ASAP7_75t_L g1395 ( 
.A1(n_1337),
.A2(n_1316),
.B(n_1310),
.Y(n_1395)
);

AO31x2_ASAP7_75t_L g1396 ( 
.A1(n_1345),
.A2(n_1347),
.A3(n_1343),
.B(n_1341),
.Y(n_1396)
);

CKINVDCx8_ASAP7_75t_R g1397 ( 
.A(n_1307),
.Y(n_1397)
);

INVx1_ASAP7_75t_SL g1398 ( 
.A(n_1302),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1342),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1272),
.B(n_1287),
.Y(n_1400)
);

HB1xp67_ASAP7_75t_L g1401 ( 
.A(n_1370),
.Y(n_1401)
);

INVx2_ASAP7_75t_L g1402 ( 
.A(n_1286),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1342),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1342),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1294),
.Y(n_1405)
);

INVxp67_ASAP7_75t_L g1406 ( 
.A(n_1378),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1336),
.Y(n_1407)
);

AOI21x1_ASAP7_75t_L g1408 ( 
.A1(n_1350),
.A2(n_1276),
.B(n_1273),
.Y(n_1408)
);

OAI21xp5_ASAP7_75t_L g1409 ( 
.A1(n_1363),
.A2(n_1388),
.B(n_1357),
.Y(n_1409)
);

OR2x2_ASAP7_75t_L g1410 ( 
.A(n_1346),
.B(n_1296),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1331),
.Y(n_1411)
);

CKINVDCx20_ASAP7_75t_R g1412 ( 
.A(n_1361),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1301),
.Y(n_1413)
);

OA21x2_ASAP7_75t_L g1414 ( 
.A1(n_1305),
.A2(n_1333),
.B(n_1299),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1309),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_1332),
.Y(n_1416)
);

INVx2_ASAP7_75t_SL g1417 ( 
.A(n_1282),
.Y(n_1417)
);

INVx3_ASAP7_75t_L g1418 ( 
.A(n_1332),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1330),
.B(n_1334),
.Y(n_1419)
);

INVx3_ASAP7_75t_L g1420 ( 
.A(n_1332),
.Y(n_1420)
);

INVx3_ASAP7_75t_L g1421 ( 
.A(n_1332),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1371),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1372),
.Y(n_1423)
);

AND2x4_ASAP7_75t_L g1424 ( 
.A(n_1319),
.B(n_1306),
.Y(n_1424)
);

BUFx2_ASAP7_75t_L g1425 ( 
.A(n_1295),
.Y(n_1425)
);

OAI21x1_ASAP7_75t_L g1426 ( 
.A1(n_1340),
.A2(n_1338),
.B(n_1328),
.Y(n_1426)
);

INVx3_ASAP7_75t_L g1427 ( 
.A(n_1339),
.Y(n_1427)
);

OAI22x1_ASAP7_75t_SL g1428 ( 
.A1(n_1275),
.A2(n_1335),
.B1(n_1376),
.B2(n_1373),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1387),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1389),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1390),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1272),
.B(n_1354),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1392),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1330),
.Y(n_1434)
);

OA21x2_ASAP7_75t_L g1435 ( 
.A1(n_1329),
.A2(n_1311),
.B(n_1323),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1344),
.Y(n_1436)
);

AO21x2_ASAP7_75t_L g1437 ( 
.A1(n_1310),
.A2(n_1297),
.B(n_1377),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1344),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1334),
.Y(n_1439)
);

HB1xp67_ASAP7_75t_L g1440 ( 
.A(n_1267),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1318),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1318),
.Y(n_1442)
);

INVx3_ASAP7_75t_L g1443 ( 
.A(n_1339),
.Y(n_1443)
);

INVxp67_ASAP7_75t_L g1444 ( 
.A(n_1278),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1268),
.B(n_1277),
.Y(n_1445)
);

INVx2_ASAP7_75t_SL g1446 ( 
.A(n_1282),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1277),
.B(n_1280),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1280),
.B(n_1279),
.Y(n_1448)
);

AND2x4_ASAP7_75t_L g1449 ( 
.A(n_1320),
.B(n_1348),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1279),
.B(n_1303),
.Y(n_1450)
);

OR2x2_ASAP7_75t_L g1451 ( 
.A(n_1283),
.B(n_1377),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1358),
.B(n_1360),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1303),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1283),
.B(n_1356),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1362),
.B(n_1383),
.Y(n_1455)
);

INVx3_ASAP7_75t_L g1456 ( 
.A(n_1339),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1297),
.Y(n_1457)
);

INVx2_ASAP7_75t_SL g1458 ( 
.A(n_1282),
.Y(n_1458)
);

OAI21xp5_ASAP7_75t_L g1459 ( 
.A1(n_1380),
.A2(n_1382),
.B(n_1393),
.Y(n_1459)
);

INVx2_ASAP7_75t_SL g1460 ( 
.A(n_1285),
.Y(n_1460)
);

AOI22xp33_ASAP7_75t_L g1461 ( 
.A1(n_1365),
.A2(n_1270),
.B1(n_1349),
.B2(n_1351),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1308),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1308),
.Y(n_1463)
);

BUFx8_ASAP7_75t_L g1464 ( 
.A(n_1374),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1313),
.B(n_1293),
.Y(n_1465)
);

OAI21x1_ASAP7_75t_L g1466 ( 
.A1(n_1322),
.A2(n_1315),
.B(n_1386),
.Y(n_1466)
);

NOR2xp33_ASAP7_75t_L g1467 ( 
.A(n_1355),
.B(n_1379),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1313),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1321),
.Y(n_1469)
);

OR2x2_ASAP7_75t_L g1470 ( 
.A(n_1270),
.B(n_1288),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1321),
.Y(n_1471)
);

AOI21xp5_ASAP7_75t_L g1472 ( 
.A1(n_1349),
.A2(n_1351),
.B(n_1352),
.Y(n_1472)
);

OR2x2_ASAP7_75t_L g1473 ( 
.A(n_1291),
.B(n_1379),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1327),
.Y(n_1474)
);

AND2x4_ASAP7_75t_L g1475 ( 
.A(n_1298),
.B(n_1353),
.Y(n_1475)
);

OR2x2_ASAP7_75t_L g1476 ( 
.A(n_1381),
.B(n_1292),
.Y(n_1476)
);

HB1xp67_ASAP7_75t_L g1477 ( 
.A(n_1304),
.Y(n_1477)
);

INVx2_ASAP7_75t_SL g1478 ( 
.A(n_1285),
.Y(n_1478)
);

OR2x2_ASAP7_75t_L g1479 ( 
.A(n_1271),
.B(n_1384),
.Y(n_1479)
);

OAI21xp5_ASAP7_75t_L g1480 ( 
.A1(n_1317),
.A2(n_1314),
.B(n_1298),
.Y(n_1480)
);

AOI22xp5_ASAP7_75t_L g1481 ( 
.A1(n_1312),
.A2(n_1289),
.B1(n_1368),
.B2(n_1290),
.Y(n_1481)
);

AND2x4_ASAP7_75t_SL g1482 ( 
.A(n_1412),
.B(n_1269),
.Y(n_1482)
);

OR2x2_ASAP7_75t_L g1483 ( 
.A(n_1473),
.B(n_1394),
.Y(n_1483)
);

OA21x2_ASAP7_75t_L g1484 ( 
.A1(n_1426),
.A2(n_1324),
.B(n_1366),
.Y(n_1484)
);

A2O1A1Ixp33_ASAP7_75t_L g1485 ( 
.A1(n_1409),
.A2(n_1298),
.B(n_1326),
.C(n_1375),
.Y(n_1485)
);

BUFx6f_ASAP7_75t_L g1486 ( 
.A(n_1397),
.Y(n_1486)
);

O2A1O1Ixp33_ASAP7_75t_SL g1487 ( 
.A1(n_1432),
.A2(n_1367),
.B(n_1274),
.C(n_1300),
.Y(n_1487)
);

AO21x2_ASAP7_75t_L g1488 ( 
.A1(n_1472),
.A2(n_1324),
.B(n_1368),
.Y(n_1488)
);

AOI21xp5_ASAP7_75t_L g1489 ( 
.A1(n_1395),
.A2(n_1326),
.B(n_1325),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1415),
.Y(n_1490)
);

A2O1A1Ixp33_ASAP7_75t_L g1491 ( 
.A1(n_1459),
.A2(n_1326),
.B(n_1368),
.C(n_1290),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1440),
.B(n_1385),
.Y(n_1492)
);

OR2x2_ASAP7_75t_L g1493 ( 
.A(n_1473),
.B(n_1364),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1454),
.B(n_1385),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1455),
.B(n_1284),
.Y(n_1495)
);

NOR3xp33_ASAP7_75t_SL g1496 ( 
.A(n_1467),
.B(n_1480),
.C(n_1400),
.Y(n_1496)
);

AND2x2_ASAP7_75t_SL g1497 ( 
.A(n_1425),
.B(n_1369),
.Y(n_1497)
);

A2O1A1Ixp33_ASAP7_75t_L g1498 ( 
.A1(n_1425),
.A2(n_1281),
.B(n_1391),
.C(n_1359),
.Y(n_1498)
);

NOR2xp33_ASAP7_75t_L g1499 ( 
.A(n_1398),
.B(n_1281),
.Y(n_1499)
);

NOR2xp33_ASAP7_75t_L g1500 ( 
.A(n_1406),
.B(n_1391),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1441),
.B(n_1442),
.Y(n_1501)
);

NOR2x1_ASAP7_75t_SL g1502 ( 
.A(n_1395),
.B(n_1413),
.Y(n_1502)
);

A2O1A1Ixp33_ASAP7_75t_L g1503 ( 
.A1(n_1461),
.A2(n_1451),
.B(n_1450),
.C(n_1470),
.Y(n_1503)
);

AOI221xp5_ASAP7_75t_SL g1504 ( 
.A1(n_1445),
.A2(n_1450),
.B1(n_1447),
.B2(n_1448),
.C(n_1457),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1415),
.Y(n_1505)
);

AOI221xp5_ASAP7_75t_L g1506 ( 
.A1(n_1452),
.A2(n_1445),
.B1(n_1457),
.B2(n_1448),
.C(n_1451),
.Y(n_1506)
);

OR2x2_ASAP7_75t_L g1507 ( 
.A(n_1468),
.B(n_1399),
.Y(n_1507)
);

OA21x2_ASAP7_75t_L g1508 ( 
.A1(n_1426),
.A2(n_1469),
.B(n_1471),
.Y(n_1508)
);

AOI221xp5_ASAP7_75t_L g1509 ( 
.A1(n_1468),
.A2(n_1447),
.B1(n_1453),
.B2(n_1463),
.C(n_1462),
.Y(n_1509)
);

AND2x4_ASAP7_75t_L g1510 ( 
.A(n_1403),
.B(n_1404),
.Y(n_1510)
);

AOI22xp33_ASAP7_75t_L g1511 ( 
.A1(n_1470),
.A2(n_1465),
.B1(n_1437),
.B2(n_1453),
.Y(n_1511)
);

OAI22xp5_ASAP7_75t_L g1512 ( 
.A1(n_1474),
.A2(n_1462),
.B1(n_1463),
.B2(n_1439),
.Y(n_1512)
);

AOI22xp5_ASAP7_75t_L g1513 ( 
.A1(n_1437),
.A2(n_1465),
.B1(n_1474),
.B2(n_1395),
.Y(n_1513)
);

OR2x2_ASAP7_75t_L g1514 ( 
.A(n_1403),
.B(n_1404),
.Y(n_1514)
);

O2A1O1Ixp33_ASAP7_75t_L g1515 ( 
.A1(n_1437),
.A2(n_1471),
.B(n_1444),
.C(n_1401),
.Y(n_1515)
);

INVx1_ASAP7_75t_SL g1516 ( 
.A(n_1477),
.Y(n_1516)
);

AOI22xp5_ASAP7_75t_L g1517 ( 
.A1(n_1414),
.A2(n_1481),
.B1(n_1424),
.B2(n_1410),
.Y(n_1517)
);

OAI221xp5_ASAP7_75t_L g1518 ( 
.A1(n_1481),
.A2(n_1408),
.B1(n_1414),
.B2(n_1476),
.C(n_1427),
.Y(n_1518)
);

OAI21xp5_ASAP7_75t_L g1519 ( 
.A1(n_1408),
.A2(n_1414),
.B(n_1466),
.Y(n_1519)
);

OR2x6_ASAP7_75t_L g1520 ( 
.A(n_1449),
.B(n_1424),
.Y(n_1520)
);

CKINVDCx5p33_ASAP7_75t_R g1521 ( 
.A(n_1428),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1402),
.B(n_1405),
.Y(n_1522)
);

AO32x2_ASAP7_75t_L g1523 ( 
.A1(n_1434),
.A2(n_1460),
.A3(n_1458),
.B1(n_1478),
.B2(n_1417),
.Y(n_1523)
);

AOI221xp5_ASAP7_75t_L g1524 ( 
.A1(n_1436),
.A2(n_1438),
.B1(n_1434),
.B2(n_1419),
.C(n_1439),
.Y(n_1524)
);

NOR2xp33_ASAP7_75t_L g1525 ( 
.A(n_1479),
.B(n_1476),
.Y(n_1525)
);

AOI22xp5_ASAP7_75t_L g1526 ( 
.A1(n_1424),
.A2(n_1410),
.B1(n_1449),
.B2(n_1443),
.Y(n_1526)
);

OAI21x1_ASAP7_75t_L g1527 ( 
.A1(n_1418),
.A2(n_1420),
.B(n_1421),
.Y(n_1527)
);

NAND3xp33_ASAP7_75t_L g1528 ( 
.A(n_1464),
.B(n_1456),
.C(n_1443),
.Y(n_1528)
);

A2O1A1Ixp33_ASAP7_75t_L g1529 ( 
.A1(n_1427),
.A2(n_1443),
.B(n_1456),
.C(n_1449),
.Y(n_1529)
);

AOI21xp5_ASAP7_75t_SL g1530 ( 
.A1(n_1475),
.A2(n_1458),
.B(n_1446),
.Y(n_1530)
);

AO32x2_ASAP7_75t_L g1531 ( 
.A1(n_1417),
.A2(n_1446),
.A3(n_1478),
.B1(n_1460),
.B2(n_1419),
.Y(n_1531)
);

OAI21xp33_ASAP7_75t_L g1532 ( 
.A1(n_1511),
.A2(n_1436),
.B(n_1438),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1490),
.Y(n_1533)
);

OR2x2_ASAP7_75t_L g1534 ( 
.A(n_1508),
.B(n_1396),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1531),
.B(n_1396),
.Y(n_1535)
);

OR2x2_ASAP7_75t_L g1536 ( 
.A(n_1508),
.B(n_1396),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1505),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1531),
.B(n_1396),
.Y(n_1538)
);

OAI211xp5_ASAP7_75t_L g1539 ( 
.A1(n_1513),
.A2(n_1422),
.B(n_1430),
.C(n_1429),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1531),
.B(n_1396),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1519),
.B(n_1396),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1519),
.B(n_1407),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1523),
.B(n_1411),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1523),
.B(n_1411),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1523),
.B(n_1411),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1522),
.Y(n_1546)
);

AND2x4_ASAP7_75t_L g1547 ( 
.A(n_1527),
.B(n_1418),
.Y(n_1547)
);

NAND4xp25_ASAP7_75t_L g1548 ( 
.A(n_1506),
.B(n_1429),
.C(n_1433),
.D(n_1431),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1520),
.B(n_1435),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1520),
.B(n_1435),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1513),
.B(n_1423),
.Y(n_1551)
);

BUFx2_ASAP7_75t_L g1552 ( 
.A(n_1484),
.Y(n_1552)
);

OR2x2_ASAP7_75t_L g1553 ( 
.A(n_1507),
.B(n_1435),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1502),
.B(n_1416),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1514),
.Y(n_1555)
);

AND2x4_ASAP7_75t_L g1556 ( 
.A(n_1547),
.B(n_1510),
.Y(n_1556)
);

NAND2x1_ASAP7_75t_L g1557 ( 
.A(n_1543),
.B(n_1530),
.Y(n_1557)
);

AO21x2_ASAP7_75t_L g1558 ( 
.A1(n_1541),
.A2(n_1515),
.B(n_1517),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1535),
.B(n_1484),
.Y(n_1559)
);

NOR2xp33_ASAP7_75t_L g1560 ( 
.A(n_1548),
.B(n_1483),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1543),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1537),
.Y(n_1562)
);

HB1xp67_ASAP7_75t_L g1563 ( 
.A(n_1543),
.Y(n_1563)
);

BUFx2_ASAP7_75t_L g1564 ( 
.A(n_1547),
.Y(n_1564)
);

AOI221xp5_ASAP7_75t_L g1565 ( 
.A1(n_1532),
.A2(n_1504),
.B1(n_1509),
.B2(n_1503),
.C(n_1512),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1535),
.B(n_1526),
.Y(n_1566)
);

OR2x2_ASAP7_75t_L g1567 ( 
.A(n_1553),
.B(n_1534),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1537),
.Y(n_1568)
);

OR2x2_ASAP7_75t_L g1569 ( 
.A(n_1553),
.B(n_1516),
.Y(n_1569)
);

INVx4_ASAP7_75t_L g1570 ( 
.A(n_1547),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1538),
.B(n_1517),
.Y(n_1571)
);

AOI221xp5_ASAP7_75t_SL g1572 ( 
.A1(n_1548),
.A2(n_1524),
.B1(n_1512),
.B2(n_1518),
.C(n_1491),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1538),
.B(n_1540),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1540),
.B(n_1501),
.Y(n_1574)
);

OAI211xp5_ASAP7_75t_L g1575 ( 
.A1(n_1539),
.A2(n_1504),
.B(n_1496),
.C(n_1485),
.Y(n_1575)
);

HB1xp67_ASAP7_75t_L g1576 ( 
.A(n_1544),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1546),
.B(n_1525),
.Y(n_1577)
);

OR2x2_ASAP7_75t_L g1578 ( 
.A(n_1534),
.B(n_1488),
.Y(n_1578)
);

BUFx3_ASAP7_75t_L g1579 ( 
.A(n_1554),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1533),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1533),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1549),
.B(n_1529),
.Y(n_1582)
);

INVx1_ASAP7_75t_SL g1583 ( 
.A(n_1545),
.Y(n_1583)
);

OAI21xp5_ASAP7_75t_SL g1584 ( 
.A1(n_1539),
.A2(n_1498),
.B(n_1482),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1571),
.B(n_1555),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1562),
.Y(n_1586)
);

INVx2_ASAP7_75t_SL g1587 ( 
.A(n_1557),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1573),
.B(n_1549),
.Y(n_1588)
);

AND2x6_ASAP7_75t_SL g1589 ( 
.A(n_1560),
.B(n_1499),
.Y(n_1589)
);

AND2x4_ASAP7_75t_L g1590 ( 
.A(n_1570),
.B(n_1549),
.Y(n_1590)
);

INVx2_ASAP7_75t_SL g1591 ( 
.A(n_1557),
.Y(n_1591)
);

OA21x2_ASAP7_75t_L g1592 ( 
.A1(n_1564),
.A2(n_1552),
.B(n_1536),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1580),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1562),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1562),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1573),
.B(n_1550),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1573),
.B(n_1550),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1561),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1568),
.Y(n_1599)
);

NAND3xp33_ASAP7_75t_SL g1600 ( 
.A(n_1565),
.B(n_1521),
.C(n_1493),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1571),
.B(n_1555),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1571),
.B(n_1546),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1580),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1580),
.B(n_1551),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1581),
.B(n_1551),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1568),
.Y(n_1606)
);

HB1xp67_ASAP7_75t_L g1607 ( 
.A(n_1581),
.Y(n_1607)
);

INVxp67_ASAP7_75t_L g1608 ( 
.A(n_1560),
.Y(n_1608)
);

HB1xp67_ASAP7_75t_L g1609 ( 
.A(n_1581),
.Y(n_1609)
);

INVx1_ASAP7_75t_SL g1610 ( 
.A(n_1569),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1574),
.B(n_1542),
.Y(n_1611)
);

NOR2xp33_ASAP7_75t_L g1612 ( 
.A(n_1575),
.B(n_1497),
.Y(n_1612)
);

AOI22xp5_ASAP7_75t_L g1613 ( 
.A1(n_1600),
.A2(n_1565),
.B1(n_1575),
.B2(n_1572),
.Y(n_1613)
);

INVx2_ASAP7_75t_SL g1614 ( 
.A(n_1607),
.Y(n_1614)
);

AOI32xp33_ASAP7_75t_L g1615 ( 
.A1(n_1612),
.A2(n_1566),
.A3(n_1559),
.B1(n_1582),
.B2(n_1572),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1588),
.B(n_1582),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1607),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1592),
.Y(n_1618)
);

INVx2_ASAP7_75t_SL g1619 ( 
.A(n_1609),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1609),
.Y(n_1620)
);

AND2x4_ASAP7_75t_L g1621 ( 
.A(n_1587),
.B(n_1579),
.Y(n_1621)
);

OR2x2_ASAP7_75t_L g1622 ( 
.A(n_1610),
.B(n_1567),
.Y(n_1622)
);

BUFx2_ASAP7_75t_L g1623 ( 
.A(n_1587),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1608),
.B(n_1577),
.Y(n_1624)
);

NOR2xp33_ASAP7_75t_L g1625 ( 
.A(n_1612),
.B(n_1428),
.Y(n_1625)
);

AND2x2_ASAP7_75t_SL g1626 ( 
.A(n_1592),
.B(n_1552),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1588),
.B(n_1582),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1593),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1588),
.B(n_1582),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1593),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1603),
.Y(n_1631)
);

HB1xp67_ASAP7_75t_L g1632 ( 
.A(n_1585),
.Y(n_1632)
);

AOI22xp5_ASAP7_75t_L g1633 ( 
.A1(n_1600),
.A2(n_1608),
.B1(n_1584),
.B2(n_1558),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1596),
.B(n_1556),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1603),
.Y(n_1635)
);

INVx1_ASAP7_75t_SL g1636 ( 
.A(n_1589),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1586),
.Y(n_1637)
);

INVxp67_ASAP7_75t_L g1638 ( 
.A(n_1604),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_SL g1639 ( 
.A(n_1602),
.B(n_1577),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1602),
.B(n_1566),
.Y(n_1640)
);

INVxp67_ASAP7_75t_L g1641 ( 
.A(n_1604),
.Y(n_1641)
);

AOI22xp5_ASAP7_75t_L g1642 ( 
.A1(n_1589),
.A2(n_1584),
.B1(n_1558),
.B2(n_1532),
.Y(n_1642)
);

NOR2xp33_ASAP7_75t_SL g1643 ( 
.A(n_1610),
.B(n_1528),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1592),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1586),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1586),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1594),
.Y(n_1647)
);

INVx1_ASAP7_75t_SL g1648 ( 
.A(n_1585),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1596),
.B(n_1597),
.Y(n_1649)
);

HB1xp67_ASAP7_75t_L g1650 ( 
.A(n_1601),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1601),
.B(n_1566),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1592),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1596),
.B(n_1556),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1592),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1594),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1616),
.B(n_1597),
.Y(n_1656)
);

OR2x2_ASAP7_75t_L g1657 ( 
.A(n_1651),
.B(n_1605),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1628),
.Y(n_1658)
);

OR2x2_ASAP7_75t_L g1659 ( 
.A(n_1640),
.B(n_1605),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1615),
.B(n_1613),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1628),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1616),
.B(n_1627),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1615),
.B(n_1574),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1613),
.B(n_1574),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1627),
.B(n_1597),
.Y(n_1665)
);

INVxp67_ASAP7_75t_L g1666 ( 
.A(n_1636),
.Y(n_1666)
);

NOR2xp33_ASAP7_75t_SL g1667 ( 
.A(n_1625),
.B(n_1486),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1624),
.B(n_1574),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1630),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1626),
.Y(n_1670)
);

CKINVDCx20_ASAP7_75t_L g1671 ( 
.A(n_1642),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1629),
.B(n_1649),
.Y(n_1672)
);

OAI21xp33_ASAP7_75t_L g1673 ( 
.A1(n_1633),
.A2(n_1541),
.B(n_1559),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1629),
.B(n_1587),
.Y(n_1674)
);

OR2x2_ASAP7_75t_L g1675 ( 
.A(n_1648),
.B(n_1611),
.Y(n_1675)
);

NOR2x1_ASAP7_75t_L g1676 ( 
.A(n_1623),
.B(n_1557),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1639),
.B(n_1611),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1638),
.B(n_1563),
.Y(n_1678)
);

CKINVDCx16_ASAP7_75t_R g1679 ( 
.A(n_1633),
.Y(n_1679)
);

INVx2_ASAP7_75t_L g1680 ( 
.A(n_1626),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1649),
.B(n_1591),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1634),
.B(n_1591),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1634),
.B(n_1591),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1653),
.B(n_1590),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1630),
.Y(n_1685)
);

OAI33xp33_ASAP7_75t_L g1686 ( 
.A1(n_1617),
.A2(n_1578),
.A3(n_1606),
.B1(n_1594),
.B2(n_1595),
.B3(n_1599),
.Y(n_1686)
);

OR2x2_ASAP7_75t_L g1687 ( 
.A(n_1632),
.B(n_1598),
.Y(n_1687)
);

AND2x4_ASAP7_75t_L g1688 ( 
.A(n_1614),
.B(n_1590),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1653),
.B(n_1590),
.Y(n_1689)
);

OR2x2_ASAP7_75t_L g1690 ( 
.A(n_1650),
.B(n_1598),
.Y(n_1690)
);

INVx2_ASAP7_75t_L g1691 ( 
.A(n_1626),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_1688),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1658),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1658),
.Y(n_1694)
);

AOI21xp33_ASAP7_75t_SL g1695 ( 
.A1(n_1679),
.A2(n_1642),
.B(n_1558),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1661),
.Y(n_1696)
);

INVx2_ASAP7_75t_SL g1697 ( 
.A(n_1688),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1666),
.B(n_1641),
.Y(n_1698)
);

HB1xp67_ASAP7_75t_L g1699 ( 
.A(n_1661),
.Y(n_1699)
);

NOR2xp33_ASAP7_75t_L g1700 ( 
.A(n_1660),
.B(n_1643),
.Y(n_1700)
);

OAI21xp33_ASAP7_75t_L g1701 ( 
.A1(n_1660),
.A2(n_1622),
.B(n_1541),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1669),
.Y(n_1702)
);

NAND2x1_ASAP7_75t_L g1703 ( 
.A(n_1676),
.B(n_1623),
.Y(n_1703)
);

AOI22xp5_ASAP7_75t_L g1704 ( 
.A1(n_1679),
.A2(n_1671),
.B1(n_1673),
.B2(n_1667),
.Y(n_1704)
);

AOI22xp33_ASAP7_75t_L g1705 ( 
.A1(n_1671),
.A2(n_1558),
.B1(n_1552),
.B2(n_1559),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1662),
.B(n_1556),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1669),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1662),
.B(n_1672),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1685),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1685),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_SL g1711 ( 
.A(n_1667),
.B(n_1621),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1664),
.B(n_1622),
.Y(n_1712)
);

OR2x2_ASAP7_75t_L g1713 ( 
.A(n_1664),
.B(n_1558),
.Y(n_1713)
);

OR2x6_ASAP7_75t_L g1714 ( 
.A(n_1670),
.B(n_1486),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1672),
.Y(n_1715)
);

NOR2x1p5_ASAP7_75t_L g1716 ( 
.A(n_1663),
.B(n_1486),
.Y(n_1716)
);

OAI22xp5_ASAP7_75t_L g1717 ( 
.A1(n_1663),
.A2(n_1583),
.B1(n_1563),
.B2(n_1576),
.Y(n_1717)
);

AOI32xp33_ASAP7_75t_L g1718 ( 
.A1(n_1700),
.A2(n_1673),
.A3(n_1670),
.B1(n_1680),
.B2(n_1691),
.Y(n_1718)
);

AOI22xp33_ASAP7_75t_SL g1719 ( 
.A1(n_1700),
.A2(n_1691),
.B1(n_1680),
.B2(n_1670),
.Y(n_1719)
);

A2O1A1Ixp33_ASAP7_75t_L g1720 ( 
.A1(n_1704),
.A2(n_1691),
.B(n_1680),
.C(n_1676),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1715),
.B(n_1656),
.Y(n_1721)
);

O2A1O1Ixp33_ASAP7_75t_SL g1722 ( 
.A1(n_1703),
.A2(n_1619),
.B(n_1614),
.C(n_1617),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1699),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1699),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1693),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1698),
.B(n_1656),
.Y(n_1726)
);

AOI22xp5_ASAP7_75t_L g1727 ( 
.A1(n_1705),
.A2(n_1674),
.B1(n_1686),
.B2(n_1677),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1708),
.B(n_1665),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1694),
.Y(n_1729)
);

OAI22xp33_ASAP7_75t_L g1730 ( 
.A1(n_1695),
.A2(n_1677),
.B1(n_1675),
.B2(n_1668),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1696),
.Y(n_1731)
);

AOI21xp33_ASAP7_75t_L g1732 ( 
.A1(n_1705),
.A2(n_1675),
.B(n_1659),
.Y(n_1732)
);

OAI22xp5_ASAP7_75t_L g1733 ( 
.A1(n_1711),
.A2(n_1678),
.B1(n_1618),
.B2(n_1644),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1702),
.Y(n_1734)
);

OR2x2_ASAP7_75t_L g1735 ( 
.A(n_1712),
.B(n_1668),
.Y(n_1735)
);

AOI221xp5_ASAP7_75t_L g1736 ( 
.A1(n_1701),
.A2(n_1678),
.B1(n_1674),
.B2(n_1665),
.C(n_1688),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1708),
.B(n_1681),
.Y(n_1737)
);

OAI21xp5_ASAP7_75t_L g1738 ( 
.A1(n_1720),
.A2(n_1711),
.B(n_1713),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1719),
.B(n_1716),
.Y(n_1739)
);

AOI221xp5_ASAP7_75t_L g1740 ( 
.A1(n_1718),
.A2(n_1717),
.B1(n_1710),
.B2(n_1709),
.C(n_1707),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1723),
.Y(n_1741)
);

AOI21xp33_ASAP7_75t_SL g1742 ( 
.A1(n_1730),
.A2(n_1714),
.B(n_1697),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1724),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1721),
.Y(n_1744)
);

INVxp67_ASAP7_75t_SL g1745 ( 
.A(n_1733),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1728),
.Y(n_1746)
);

AOI211xp5_ASAP7_75t_L g1747 ( 
.A1(n_1722),
.A2(n_1697),
.B(n_1692),
.C(n_1487),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1737),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1745),
.B(n_1726),
.Y(n_1749)
);

NOR3xp33_ASAP7_75t_L g1750 ( 
.A(n_1739),
.B(n_1729),
.C(n_1725),
.Y(n_1750)
);

NAND4xp25_ASAP7_75t_L g1751 ( 
.A(n_1747),
.B(n_1732),
.C(n_1736),
.D(n_1727),
.Y(n_1751)
);

INVxp67_ASAP7_75t_L g1752 ( 
.A(n_1745),
.Y(n_1752)
);

OAI211xp5_ASAP7_75t_SL g1753 ( 
.A1(n_1738),
.A2(n_1734),
.B(n_1731),
.C(n_1735),
.Y(n_1753)
);

NOR2x1_ASAP7_75t_L g1754 ( 
.A(n_1741),
.B(n_1714),
.Y(n_1754)
);

NAND3xp33_ASAP7_75t_L g1755 ( 
.A(n_1742),
.B(n_1733),
.C(n_1714),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1748),
.B(n_1692),
.Y(n_1756)
);

NOR3xp33_ASAP7_75t_L g1757 ( 
.A(n_1746),
.B(n_1744),
.C(n_1748),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1743),
.B(n_1681),
.Y(n_1758)
);

INVxp67_ASAP7_75t_SL g1759 ( 
.A(n_1754),
.Y(n_1759)
);

OAI211xp5_ASAP7_75t_SL g1760 ( 
.A1(n_1749),
.A2(n_1740),
.B(n_1500),
.C(n_1657),
.Y(n_1760)
);

AOI321xp33_ASAP7_75t_L g1761 ( 
.A1(n_1750),
.A2(n_1688),
.A3(n_1682),
.B1(n_1683),
.B2(n_1706),
.C(n_1689),
.Y(n_1761)
);

NOR3xp33_ASAP7_75t_L g1762 ( 
.A(n_1751),
.B(n_1659),
.C(n_1657),
.Y(n_1762)
);

OAI21xp5_ASAP7_75t_SL g1763 ( 
.A1(n_1755),
.A2(n_1683),
.B(n_1682),
.Y(n_1763)
);

INVxp33_ASAP7_75t_SL g1764 ( 
.A(n_1757),
.Y(n_1764)
);

OAI21xp5_ASAP7_75t_SL g1765 ( 
.A1(n_1760),
.A2(n_1752),
.B(n_1753),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1759),
.B(n_1763),
.Y(n_1766)
);

INVx2_ASAP7_75t_L g1767 ( 
.A(n_1761),
.Y(n_1767)
);

NOR2xp67_ASAP7_75t_L g1768 ( 
.A(n_1764),
.B(n_1758),
.Y(n_1768)
);

OAI22xp5_ASAP7_75t_L g1769 ( 
.A1(n_1762),
.A2(n_1756),
.B1(n_1619),
.B2(n_1621),
.Y(n_1769)
);

OAI311xp33_ASAP7_75t_L g1770 ( 
.A1(n_1763),
.A2(n_1690),
.A3(n_1687),
.B1(n_1689),
.C1(n_1684),
.Y(n_1770)
);

AOI211xp5_ASAP7_75t_L g1771 ( 
.A1(n_1760),
.A2(n_1684),
.B(n_1687),
.C(n_1690),
.Y(n_1771)
);

AOI22xp5_ASAP7_75t_L g1772 ( 
.A1(n_1767),
.A2(n_1620),
.B1(n_1621),
.B2(n_1590),
.Y(n_1772)
);

AOI22xp5_ASAP7_75t_L g1773 ( 
.A1(n_1765),
.A2(n_1620),
.B1(n_1621),
.B2(n_1590),
.Y(n_1773)
);

XNOR2xp5_ASAP7_75t_L g1774 ( 
.A(n_1768),
.B(n_1528),
.Y(n_1774)
);

NAND5xp2_ASAP7_75t_L g1775 ( 
.A(n_1766),
.B(n_1489),
.C(n_1495),
.D(n_1492),
.E(n_1494),
.Y(n_1775)
);

NOR2x1_ASAP7_75t_L g1776 ( 
.A(n_1769),
.B(n_1631),
.Y(n_1776)
);

OR2x2_ASAP7_75t_L g1777 ( 
.A(n_1772),
.B(n_1770),
.Y(n_1777)
);

OAI221xp5_ASAP7_75t_L g1778 ( 
.A1(n_1773),
.A2(n_1771),
.B1(n_1618),
.B2(n_1644),
.C(n_1654),
.Y(n_1778)
);

NAND3xp33_ASAP7_75t_L g1779 ( 
.A(n_1774),
.B(n_1654),
.C(n_1652),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1777),
.Y(n_1780)
);

HB1xp67_ASAP7_75t_L g1781 ( 
.A(n_1780),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1781),
.Y(n_1782)
);

CKINVDCx20_ASAP7_75t_R g1783 ( 
.A(n_1781),
.Y(n_1783)
);

AND3x2_ASAP7_75t_L g1784 ( 
.A(n_1782),
.B(n_1776),
.C(n_1775),
.Y(n_1784)
);

AOI22xp5_ASAP7_75t_L g1785 ( 
.A1(n_1783),
.A2(n_1778),
.B1(n_1779),
.B2(n_1652),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1784),
.B(n_1631),
.Y(n_1786)
);

INVxp67_ASAP7_75t_L g1787 ( 
.A(n_1785),
.Y(n_1787)
);

OR5x1_ASAP7_75t_L g1788 ( 
.A(n_1787),
.B(n_1655),
.C(n_1647),
.D(n_1646),
.E(n_1645),
.Y(n_1788)
);

AO21x2_ASAP7_75t_L g1789 ( 
.A1(n_1788),
.A2(n_1786),
.B(n_1655),
.Y(n_1789)
);

HB1xp67_ASAP7_75t_L g1790 ( 
.A(n_1789),
.Y(n_1790)
);

OAI221xp5_ASAP7_75t_R g1791 ( 
.A1(n_1790),
.A2(n_1635),
.B1(n_1646),
.B2(n_1645),
.C(n_1637),
.Y(n_1791)
);

AOI211xp5_ASAP7_75t_L g1792 ( 
.A1(n_1791),
.A2(n_1635),
.B(n_1637),
.C(n_1647),
.Y(n_1792)
);


endmodule