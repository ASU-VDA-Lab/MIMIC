module fake_jpeg_21680_n_152 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_152);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_152;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_40),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g44 ( 
.A(n_27),
.Y(n_44)
);

INVx6_ASAP7_75t_SL g45 ( 
.A(n_36),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_20),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_9),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_17),
.Y(n_52)
);

BUFx8_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_10),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_4),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_32),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_7),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_7),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_41),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_33),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_6),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_12),
.Y(n_72)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

INVx3_ASAP7_75t_SL g88 ( 
.A(n_74),
.Y(n_88)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_75),
.B(n_78),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_77),
.B(n_56),
.Y(n_81)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_79),
.B(n_55),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_55),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_80),
.A2(n_77),
.B1(n_73),
.B2(n_44),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_84),
.Y(n_93)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_76),
.Y(n_82)
);

INVx3_ASAP7_75t_SL g94 ( 
.A(n_82),
.Y(n_94)
);

O2A1O1Ixp33_ASAP7_75t_SL g97 ( 
.A1(n_86),
.A2(n_90),
.B(n_70),
.C(n_65),
.Y(n_97)
);

BUFx16f_ASAP7_75t_L g87 ( 
.A(n_80),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_87),
.B(n_89),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_74),
.B(n_63),
.Y(n_89)
);

NAND3xp33_ASAP7_75t_SL g90 ( 
.A(n_80),
.B(n_71),
.C(n_64),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_87),
.B(n_44),
.C(n_47),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_92),
.B(n_99),
.C(n_61),
.Y(n_113)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_95),
.B(n_101),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_97),
.A2(n_98),
.B1(n_91),
.B2(n_96),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_85),
.A2(n_54),
.B1(n_66),
.B2(n_48),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_90),
.B(n_56),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_88),
.A2(n_72),
.B1(n_69),
.B2(n_46),
.Y(n_100)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_100),
.Y(n_107)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_91),
.Y(n_101)
);

INVx2_ASAP7_75t_SL g102 ( 
.A(n_88),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_102),
.B(n_103),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_82),
.Y(n_103)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_94),
.Y(n_104)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_99),
.A2(n_50),
.B1(n_58),
.B2(n_60),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_105),
.A2(n_111),
.B1(n_5),
.B2(n_8),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_93),
.B(n_68),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_108),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_96),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_109),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_102),
.A2(n_67),
.B1(n_62),
.B2(n_43),
.Y(n_111)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_103),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_112),
.B(n_115),
.Y(n_127)
);

OR2x2_ASAP7_75t_SL g121 ( 
.A(n_113),
.B(n_114),
.Y(n_121)
);

AND2x2_ASAP7_75t_SL g114 ( 
.A(n_95),
.B(n_48),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_100),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_93),
.B(n_52),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_116),
.B(n_119),
.Y(n_126)
);

MAJx2_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_49),
.C(n_23),
.Y(n_117)
);

A2O1A1Ixp33_ASAP7_75t_L g128 ( 
.A1(n_117),
.A2(n_3),
.B(n_4),
.C(n_5),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_99),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_120),
.A2(n_107),
.B1(n_126),
.B2(n_123),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_110),
.B(n_45),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_124),
.B(n_128),
.Y(n_137)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_110),
.Y(n_125)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_125),
.Y(n_134)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_118),
.Y(n_129)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_129),
.Y(n_136)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_118),
.Y(n_130)
);

INVx1_ASAP7_75t_SL g138 ( 
.A(n_130),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_131),
.B(n_13),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_132),
.A2(n_133),
.B1(n_135),
.B2(n_121),
.Y(n_140)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_122),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_132),
.B(n_126),
.Y(n_139)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_139),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_141),
.A2(n_140),
.B1(n_136),
.B2(n_138),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_142),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_134),
.C(n_114),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_127),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_145),
.A2(n_138),
.B1(n_119),
.B2(n_127),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_137),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_147),
.A2(n_14),
.B(n_15),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_148),
.B(n_16),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_19),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_150),
.A2(n_21),
.B1(n_25),
.B2(n_29),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_31),
.Y(n_152)
);


endmodule