module fake_jpeg_181_n_224 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_224);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_224;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

INVx2_ASAP7_75t_L g14 ( 
.A(n_13),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_11),
.B(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_36),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_37),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_38),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_39),
.Y(n_98)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_40),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_41),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_21),
.B(n_1),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_42),
.B(n_46),
.Y(n_78)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_43),
.Y(n_107)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_25),
.B(n_3),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_48),
.Y(n_109)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_49),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_33),
.B(n_12),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_65),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_51),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_54),
.Y(n_99)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_55),
.Y(n_86)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_56),
.Y(n_112)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_57),
.Y(n_93)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_59),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_28),
.B(n_4),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_60),
.B(n_63),
.Y(n_97)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_14),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_62),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_16),
.B(n_26),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_67),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_33),
.B(n_4),
.Y(n_65)
);

AOI21xp33_ASAP7_75t_L g66 ( 
.A1(n_15),
.A2(n_4),
.B(n_5),
.Y(n_66)
);

OR2x4_ASAP7_75t_L g106 ( 
.A(n_66),
.B(n_7),
.Y(n_106)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_15),
.Y(n_67)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_18),
.Y(n_68)
);

BUFx12_ASAP7_75t_L g94 ( 
.A(n_68),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_18),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_70),
.Y(n_90)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_22),
.Y(n_70)
);

INVx6_ASAP7_75t_SL g71 ( 
.A(n_23),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_71),
.B(n_73),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_72),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_27),
.Y(n_73)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_27),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_74),
.B(n_75),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_31),
.B(n_5),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_76),
.A2(n_58),
.B1(n_62),
.B2(n_56),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g121 ( 
.A(n_87),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_45),
.A2(n_47),
.B1(n_51),
.B2(n_37),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_101),
.A2(n_102),
.B1(n_105),
.B2(n_113),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_42),
.A2(n_31),
.B1(n_29),
.B2(n_30),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_38),
.A2(n_30),
.B1(n_6),
.B2(n_7),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_106),
.B(n_6),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_54),
.A2(n_5),
.B1(n_6),
.B2(n_69),
.Y(n_113)
);

INVx2_ASAP7_75t_SL g114 ( 
.A(n_112),
.Y(n_114)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_114),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_81),
.A2(n_75),
.B1(n_60),
.B2(n_73),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_115),
.B(n_122),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_81),
.B(n_76),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_116),
.B(n_125),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_108),
.A2(n_65),
.B(n_46),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_117),
.A2(n_93),
.B(n_84),
.Y(n_155)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_83),
.Y(n_118)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_118),
.Y(n_143)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_89),
.Y(n_119)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_119),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_79),
.Y(n_123)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_123),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_97),
.B(n_63),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_124),
.B(n_126),
.Y(n_150)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_103),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_80),
.B(n_72),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_90),
.B(n_39),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_127),
.B(n_128),
.Y(n_156)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_92),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_107),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_129),
.B(n_131),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_95),
.B(n_41),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_130),
.B(n_132),
.C(n_139),
.Y(n_145)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_88),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_78),
.B(n_52),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_96),
.B(n_64),
.Y(n_133)
);

BUFx24_ASAP7_75t_SL g154 ( 
.A(n_133),
.Y(n_154)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_134),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_105),
.A2(n_113),
.B1(n_101),
.B2(n_87),
.Y(n_135)
);

AO22x1_ASAP7_75t_L g151 ( 
.A1(n_135),
.A2(n_137),
.B1(n_85),
.B2(n_86),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_82),
.B(n_77),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_136),
.Y(n_157)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_110),
.Y(n_137)
);

OAI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_110),
.A2(n_79),
.B1(n_98),
.B2(n_111),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_138),
.A2(n_130),
.B1(n_116),
.B2(n_121),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_99),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_91),
.B(n_111),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_140),
.B(n_104),
.C(n_91),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_141),
.A2(n_160),
.B1(n_119),
.B2(n_117),
.Y(n_167)
);

O2A1O1Ixp33_ASAP7_75t_SL g144 ( 
.A1(n_121),
.A2(n_93),
.B(n_89),
.C(n_85),
.Y(n_144)
);

A2O1A1Ixp33_ASAP7_75t_L g165 ( 
.A1(n_144),
.A2(n_131),
.B(n_129),
.C(n_134),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_151),
.A2(n_123),
.B1(n_141),
.B2(n_158),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_155),
.A2(n_114),
.B(n_120),
.Y(n_166)
);

AO22x1_ASAP7_75t_L g158 ( 
.A1(n_135),
.A2(n_85),
.B1(n_98),
.B2(n_100),
.Y(n_158)
);

NAND2x1_ASAP7_75t_L g162 ( 
.A(n_158),
.B(n_116),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_159),
.B(n_114),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_127),
.A2(n_94),
.B1(n_99),
.B2(n_140),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_145),
.B(n_125),
.C(n_118),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_161),
.B(n_163),
.Y(n_182)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_162),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_145),
.B(n_132),
.C(n_128),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_164),
.B(n_146),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_165),
.A2(n_167),
.B1(n_146),
.B2(n_160),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_166),
.A2(n_172),
.B(n_146),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_156),
.B(n_137),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_168),
.B(n_174),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_150),
.B(n_94),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_169),
.B(n_171),
.Y(n_184)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_143),
.Y(n_170)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_170),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_152),
.Y(n_171)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_143),
.Y(n_173)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_173),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_156),
.B(n_159),
.Y(n_174)
);

AO21x2_ASAP7_75t_SL g175 ( 
.A1(n_144),
.A2(n_158),
.B(n_151),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_175),
.B(n_162),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_167),
.A2(n_151),
.B1(n_155),
.B2(n_148),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_176),
.A2(n_183),
.B1(n_177),
.B2(n_186),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_178),
.B(n_164),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_180),
.B(n_181),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_168),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_161),
.B(n_157),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_185),
.Y(n_189)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_186),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_182),
.B(n_174),
.C(n_163),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_191),
.B(n_182),
.C(n_177),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_192),
.A2(n_194),
.B1(n_195),
.B2(n_175),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_184),
.Y(n_193)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_193),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_183),
.A2(n_175),
.B1(n_165),
.B2(n_166),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_179),
.A2(n_172),
.B1(n_175),
.B2(n_162),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_179),
.Y(n_197)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_197),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_198),
.B(n_187),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_200),
.B(n_202),
.C(n_190),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_201),
.B(n_203),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_198),
.B(n_180),
.C(n_176),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_194),
.A2(n_187),
.B1(n_188),
.B2(n_154),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_204),
.B(n_191),
.Y(n_207)
);

MAJx2_ASAP7_75t_L g214 ( 
.A(n_207),
.B(n_209),
.C(n_202),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_199),
.Y(n_208)
);

NOR3xp33_ASAP7_75t_L g211 ( 
.A(n_208),
.B(n_188),
.C(n_153),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_205),
.A2(n_189),
.B(n_192),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_210),
.B(n_203),
.C(n_196),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_211),
.B(n_212),
.C(n_196),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_206),
.B(n_200),
.Y(n_213)
);

MAJx2_ASAP7_75t_L g216 ( 
.A(n_213),
.B(n_214),
.C(n_204),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_215),
.B(n_216),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_211),
.B(n_206),
.C(n_195),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_217),
.B(n_142),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_218),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_216),
.A2(n_142),
.B(n_147),
.Y(n_219)
);

BUFx24_ASAP7_75t_SL g221 ( 
.A(n_219),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_222),
.A2(n_220),
.B(n_149),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_223),
.B(n_221),
.Y(n_224)
);


endmodule