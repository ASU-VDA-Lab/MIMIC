module fake_jpeg_21694_n_326 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_326);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_326;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_0),
.B(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx4f_ASAP7_75t_SL g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx6f_ASAP7_75t_SL g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_20),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_36),
.B(n_39),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_20),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_20),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_45),
.Y(n_60)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_19),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_41),
.A2(n_22),
.B1(n_25),
.B2(n_18),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_47),
.A2(n_48),
.B1(n_55),
.B2(n_61),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_41),
.A2(n_22),
.B1(n_35),
.B2(n_18),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_22),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_32),
.Y(n_69)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx6_ASAP7_75t_SL g68 ( 
.A(n_53),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_35),
.A2(n_18),
.B1(n_25),
.B2(n_23),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_35),
.A2(n_25),
.B1(n_23),
.B2(n_28),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_56),
.A2(n_17),
.B1(n_30),
.B2(n_33),
.Y(n_76)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_45),
.A2(n_23),
.B1(n_31),
.B2(n_29),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_36),
.A2(n_40),
.B1(n_39),
.B2(n_23),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_62),
.A2(n_31),
.B1(n_42),
.B2(n_44),
.Y(n_94)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_36),
.B(n_29),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_28),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_60),
.B(n_45),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_67),
.B(n_74),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_69),
.B(n_72),
.Y(n_99)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

INVx3_ASAP7_75t_SL g111 ( 
.A(n_70),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_52),
.B(n_38),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_71),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_46),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_40),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_73),
.B(n_77),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_51),
.B(n_39),
.Y(n_74)
);

AOI22x1_ASAP7_75t_L g75 ( 
.A1(n_62),
.A2(n_43),
.B1(n_37),
.B2(n_44),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_75),
.A2(n_42),
.B1(n_33),
.B2(n_32),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_76),
.A2(n_82),
.B1(n_57),
.B2(n_66),
.Y(n_109)
);

BUFx24_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_51),
.B(n_38),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_80),
.B(n_89),
.Y(n_108)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_61),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_85),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_50),
.A2(n_17),
.B1(n_30),
.B2(n_19),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_83),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_59),
.Y(n_85)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_88),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_65),
.B(n_38),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_90),
.B(n_63),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_91),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_55),
.Y(n_92)
);

BUFx24_ASAP7_75t_SL g113 ( 
.A(n_92),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_52),
.B(n_44),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_37),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_L g120 ( 
.A1(n_94),
.A2(n_42),
.B1(n_32),
.B2(n_26),
.Y(n_120)
);

OAI21xp33_ASAP7_75t_L g98 ( 
.A1(n_67),
.A2(n_46),
.B(n_50),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_98),
.A2(n_106),
.B(n_79),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_78),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_100),
.B(n_115),
.Y(n_142)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_101),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_73),
.B(n_64),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_103),
.B(n_105),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_77),
.B(n_32),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_48),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_109),
.A2(n_118),
.B1(n_70),
.B2(n_79),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_74),
.B(n_32),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_112),
.B(n_114),
.Y(n_141)
);

A2O1A1Ixp33_ASAP7_75t_L g114 ( 
.A1(n_93),
.A2(n_66),
.B(n_49),
.C(n_33),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_78),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_116),
.B(n_117),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_89),
.B(n_63),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_88),
.A2(n_58),
.B1(n_53),
.B2(n_49),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_119),
.A2(n_120),
.B1(n_71),
.B2(n_72),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_80),
.B(n_34),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_122),
.B(n_123),
.C(n_124),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_71),
.B(n_69),
.C(n_81),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_71),
.B(n_34),
.C(n_27),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_106),
.A2(n_75),
.B1(n_87),
.B2(n_94),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_125),
.A2(n_126),
.B1(n_127),
.B2(n_132),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_106),
.A2(n_87),
.B1(n_75),
.B2(n_90),
.Y(n_126)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_101),
.Y(n_129)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_129),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_119),
.A2(n_84),
.B1(n_70),
.B2(n_88),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_133),
.A2(n_118),
.B1(n_100),
.B2(n_117),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_102),
.A2(n_84),
.B1(n_86),
.B2(n_68),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_134),
.A2(n_145),
.B1(n_149),
.B2(n_133),
.Y(n_168)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_110),
.Y(n_135)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_135),
.Y(n_165)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_110),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_136),
.Y(n_176)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_114),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_137),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_102),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_139),
.B(n_140),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_103),
.Y(n_140)
);

MAJx2_ASAP7_75t_L g143 ( 
.A(n_123),
.B(n_21),
.C(n_79),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_143),
.B(n_124),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_144),
.B(n_147),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_109),
.A2(n_86),
.B1(n_68),
.B2(n_91),
.Y(n_145)
);

NAND2xp33_ASAP7_75t_SL g146 ( 
.A(n_114),
.B(n_91),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_146),
.A2(n_96),
.B(n_115),
.Y(n_158)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_95),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_95),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_148),
.B(n_97),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_96),
.A2(n_26),
.B1(n_34),
.B2(n_27),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g150 ( 
.A(n_98),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_150),
.B(n_97),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_130),
.B(n_123),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_151),
.B(n_152),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_130),
.B(n_108),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_135),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_153),
.B(n_148),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_131),
.B(n_108),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_154),
.B(n_156),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_139),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_157),
.B(n_163),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_158),
.A2(n_169),
.B(n_159),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_143),
.B(n_107),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_160),
.B(n_162),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_150),
.A2(n_113),
.B1(n_124),
.B2(n_116),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_131),
.B(n_99),
.Y(n_163)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_164),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_166),
.A2(n_168),
.B1(n_170),
.B2(n_175),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_141),
.B(n_99),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_167),
.B(n_171),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_141),
.A2(n_112),
.B(n_107),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_137),
.A2(n_122),
.B1(n_105),
.B2(n_104),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_140),
.B(n_104),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_145),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_173),
.B(n_174),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_132),
.A2(n_111),
.B1(n_26),
.B2(n_83),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_144),
.B(n_21),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_177),
.B(n_149),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_164),
.Y(n_179)
);

OR2x2_ASAP7_75t_L g218 ( 
.A(n_179),
.B(n_181),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_157),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_165),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_183),
.B(n_187),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_159),
.Y(n_186)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_186),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_165),
.Y(n_187)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_189),
.Y(n_216)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_172),
.Y(n_190)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_190),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_161),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_192),
.B(n_194),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_170),
.B(n_138),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_193),
.B(n_200),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_161),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_195),
.B(n_177),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_197),
.B(n_111),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_171),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_198),
.B(n_199),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_178),
.B(n_142),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_176),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_173),
.A2(n_125),
.B1(n_126),
.B2(n_146),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_201),
.A2(n_204),
.B1(n_10),
.B2(n_16),
.Y(n_227)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_166),
.Y(n_202)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_202),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_155),
.A2(n_129),
.B1(n_128),
.B2(n_134),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_175),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_205),
.Y(n_217)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_153),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_206),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_158),
.A2(n_136),
.B(n_143),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_207),
.A2(n_156),
.B(n_160),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_202),
.A2(n_128),
.B1(n_169),
.B2(n_167),
.Y(n_208)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_208),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_210),
.B(n_188),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_211),
.A2(n_219),
.B(n_195),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_185),
.A2(n_162),
.B1(n_152),
.B2(n_154),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_212),
.A2(n_228),
.B1(n_231),
.B2(n_204),
.Y(n_238)
);

BUFx5_ASAP7_75t_L g214 ( 
.A(n_190),
.Y(n_214)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_214),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_198),
.A2(n_151),
.B1(n_163),
.B2(n_147),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_181),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_220),
.B(n_183),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_224),
.B(n_207),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_185),
.A2(n_111),
.B1(n_26),
.B2(n_21),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_225),
.A2(n_227),
.B1(n_188),
.B2(n_199),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_180),
.B(n_111),
.C(n_121),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_226),
.B(n_232),
.C(n_203),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_184),
.A2(n_83),
.B1(n_121),
.B2(n_95),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_184),
.A2(n_121),
.B1(n_1),
.B2(n_2),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_180),
.B(n_15),
.C(n_14),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_233),
.B(n_235),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_218),
.A2(n_196),
.B(n_179),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_234),
.B(n_250),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_226),
.B(n_203),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_220),
.B(n_200),
.Y(n_236)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_236),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_237),
.B(n_239),
.C(n_244),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_238),
.A2(n_249),
.B1(n_253),
.B2(n_227),
.Y(n_269)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_240),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_214),
.B(n_230),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_241),
.B(n_243),
.Y(n_264)
);

BUFx2_ASAP7_75t_L g258 ( 
.A(n_242),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_211),
.B(n_182),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_212),
.B(n_182),
.C(n_191),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_245),
.B(n_247),
.C(n_210),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_222),
.B(n_196),
.Y(n_246)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_246),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_219),
.B(n_191),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_223),
.A2(n_201),
.B1(n_197),
.B2(n_194),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_218),
.A2(n_192),
.B(n_187),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_222),
.B(n_206),
.Y(n_251)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_251),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_217),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_248),
.A2(n_223),
.B1(n_217),
.B2(n_224),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_257),
.B(n_260),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_252),
.B(n_216),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_238),
.B(n_216),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_262),
.B(n_268),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_263),
.B(n_235),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_244),
.A2(n_249),
.B(n_215),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_265),
.A2(n_250),
.B(n_234),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_233),
.A2(n_213),
.B1(n_209),
.B2(n_215),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_269),
.A2(n_229),
.B1(n_228),
.B2(n_221),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_237),
.B(n_209),
.C(n_213),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_270),
.B(n_13),
.C(n_11),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_271),
.A2(n_276),
.B1(n_0),
.B2(n_1),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_SL g272 ( 
.A(n_255),
.B(n_243),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_272),
.B(n_275),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_256),
.B(n_221),
.Y(n_273)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_273),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_274),
.A2(n_278),
.B1(n_0),
.B2(n_1),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_259),
.A2(n_265),
.B(n_261),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_257),
.A2(n_229),
.B(n_247),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_277),
.B(n_279),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_269),
.A2(n_239),
.B1(n_231),
.B2(n_245),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_266),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_232),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_282),
.B(n_284),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_264),
.A2(n_15),
.B(n_14),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_283),
.A2(n_11),
.B(n_9),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_270),
.B(n_11),
.C(n_10),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_285),
.B(n_284),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_281),
.A2(n_258),
.B1(n_268),
.B2(n_254),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_286),
.B(n_272),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_287),
.B(n_285),
.Y(n_300)
);

FAx1_ASAP7_75t_SL g289 ( 
.A(n_271),
.B(n_255),
.CI(n_263),
.CON(n_289),
.SN(n_289)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_289),
.B(n_291),
.Y(n_307)
);

AND2x4_ASAP7_75t_L g290 ( 
.A(n_276),
.B(n_258),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_290),
.B(n_297),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_280),
.B(n_254),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_292),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_295),
.B(n_274),
.Y(n_302)
);

A2O1A1Ixp33_ASAP7_75t_L g298 ( 
.A1(n_277),
.A2(n_8),
.B(n_2),
.C(n_3),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_298),
.A2(n_1),
.B(n_2),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_300),
.B(n_303),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_301),
.B(n_302),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_288),
.B(n_278),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_296),
.B(n_275),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_304),
.B(n_303),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_305),
.A2(n_295),
.B1(n_290),
.B2(n_286),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_306),
.A2(n_290),
.B1(n_293),
.B2(n_289),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_296),
.B(n_5),
.Y(n_308)
);

AOI21xp33_ASAP7_75t_L g312 ( 
.A1(n_308),
.A2(n_298),
.B(n_290),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_307),
.B(n_294),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_309),
.A2(n_311),
.B(n_312),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_310),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_314),
.B(n_299),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_299),
.A2(n_5),
.B(n_6),
.Y(n_315)
);

AOI21x1_ASAP7_75t_L g320 ( 
.A1(n_315),
.A2(n_6),
.B(n_7),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_317),
.A2(n_320),
.B1(n_316),
.B2(n_7),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_318),
.B(n_313),
.C(n_316),
.Y(n_321)
);

AO21x1_ASAP7_75t_L g323 ( 
.A1(n_321),
.A2(n_322),
.B(n_319),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_6),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_8),
.C(n_6),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_L g326 ( 
.A1(n_325),
.A2(n_7),
.B1(n_8),
.B2(n_220),
.Y(n_326)
);


endmodule