module fake_jpeg_29119_n_59 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_59);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_59;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_51;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_6),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

BUFx5_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

INVx6_ASAP7_75t_SL g11 ( 
.A(n_4),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g16 ( 
.A(n_7),
.B(n_5),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_16),
.B(n_7),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_18),
.B(n_19),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_16),
.B(n_1),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_8),
.B(n_3),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_20),
.B(n_21),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_8),
.B(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_22),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_9),
.A2(n_1),
.B(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_23),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_L g28 ( 
.A1(n_21),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_28)
);

OAI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_28),
.A2(n_15),
.B1(n_13),
.B2(n_17),
.Y(n_35)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_10),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_12),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_25),
.C(n_24),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_31),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_14),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_35),
.Y(n_40)
);

OR2x2_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_9),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_34),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_26),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_37),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_27),
.B(n_12),
.Y(n_37)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g44 ( 
.A(n_43),
.B(n_30),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_43),
.C(n_41),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_39),
.B(n_24),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_45),
.B(n_48),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_40),
.A2(n_31),
.B1(n_33),
.B2(n_13),
.Y(n_46)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_38),
.A2(n_15),
.B1(n_17),
.B2(n_29),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_49),
.A2(n_51),
.B1(n_10),
.B2(n_11),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_29),
.C(n_38),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_52),
.A2(n_46),
.B1(n_47),
.B2(n_17),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_53),
.B(n_11),
.Y(n_56)
);

XOR2xp5_ASAP7_75t_L g55 ( 
.A(n_54),
.B(n_50),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_55),
.B(n_56),
.C(n_53),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_2),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_2),
.Y(n_59)
);


endmodule