module fake_jpeg_6626_n_137 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_137);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_137;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_11),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_SL g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_13),
.B(n_0),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_26),
.B(n_30),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_31),
.Y(n_39)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

CKINVDCx6p67_ASAP7_75t_R g36 ( 
.A(n_29),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_17),
.B(n_0),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_33),
.Y(n_44)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_40),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_25),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_38),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_33),
.B(n_25),
.Y(n_38)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_43),
.Y(n_50)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_27),
.B(n_18),
.Y(n_45)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_36),
.A2(n_24),
.B1(n_19),
.B2(n_16),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_46),
.A2(n_40),
.B1(n_15),
.B2(n_21),
.Y(n_67)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_53),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_41),
.A2(n_24),
.B1(n_19),
.B2(n_22),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_52),
.A2(n_44),
.B1(n_42),
.B2(n_15),
.Y(n_72)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_37),
.B(n_13),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_54),
.B(n_56),
.Y(n_64)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_55),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_35),
.B(n_22),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_58),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_42),
.Y(n_69)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_60),
.B(n_63),
.Y(n_88)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_68),
.Y(n_85)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_67),
.A2(n_72),
.B1(n_1),
.B2(n_5),
.Y(n_89)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_51),
.A2(n_21),
.B(n_35),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_71),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_39),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_34),
.Y(n_73)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_73),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_56),
.A2(n_20),
.B(n_31),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_74),
.B(n_47),
.C(n_20),
.Y(n_76)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_76),
.B(n_73),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_68),
.A2(n_53),
.B1(n_48),
.B2(n_47),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_84),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_34),
.C(n_31),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_83),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_28),
.C(n_58),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_72),
.A2(n_28),
.B1(n_58),
.B2(n_20),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_66),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_86),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_64),
.A2(n_20),
.B1(n_2),
.B2(n_3),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_87),
.B(n_8),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_89),
.A2(n_63),
.B1(n_61),
.B2(n_75),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_78),
.A2(n_80),
.B(n_82),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_92),
.A2(n_98),
.B(n_1),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_93),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_94),
.A2(n_95),
.B1(n_101),
.B2(n_62),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_83),
.Y(n_95)
);

AOI322xp5_ASAP7_75t_L g96 ( 
.A1(n_80),
.A2(n_85),
.A3(n_74),
.B1(n_77),
.B2(n_79),
.C1(n_60),
.C2(n_84),
.Y(n_96)
);

INVx13_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

AOI21x1_ASAP7_75t_L g98 ( 
.A1(n_88),
.A2(n_73),
.B(n_86),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_81),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_99),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_85),
.Y(n_100)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_100),
.Y(n_102)
);

A2O1A1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_98),
.A2(n_66),
.B(n_65),
.C(n_6),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_103),
.B(n_109),
.Y(n_117)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_104),
.B(n_105),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_107),
.B(n_94),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_97),
.B(n_92),
.Y(n_108)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_108),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_97),
.A2(n_1),
.B1(n_5),
.B2(n_6),
.Y(n_109)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_109),
.Y(n_113)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_102),
.Y(n_114)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_114),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_115),
.B(n_118),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_117),
.A2(n_103),
.B(n_104),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_108),
.B(n_95),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_119),
.B(n_120),
.Y(n_126)
);

OAI21x1_ASAP7_75t_L g120 ( 
.A1(n_116),
.A2(n_105),
.B(n_107),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_112),
.A2(n_113),
.B(n_111),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_123),
.B(n_124),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_115),
.B(n_111),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_121),
.A2(n_114),
.B1(n_102),
.B2(n_118),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_125),
.B(n_128),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_122),
.B(n_106),
.Y(n_128)
);

OAI31xp67_ASAP7_75t_L g129 ( 
.A1(n_122),
.A2(n_110),
.A3(n_91),
.B(n_7),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_129),
.A2(n_91),
.B1(n_8),
.B2(n_11),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_127),
.B(n_110),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_130),
.B(n_132),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_131),
.B(n_126),
.Y(n_134)
);

NAND3xp33_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_129),
.C(n_130),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_133),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_136),
.A2(n_6),
.B(n_7),
.Y(n_137)
);


endmodule