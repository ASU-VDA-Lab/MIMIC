module fake_jpeg_16477_n_61 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_61);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_61;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVx2_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_0),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

INVx11_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

BUFx16f_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_0),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_18),
.B(n_20),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_8),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_19),
.A2(n_10),
.B1(n_15),
.B2(n_14),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_22),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_8),
.B(n_16),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_23),
.B(n_24),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_16),
.B(n_2),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_24),
.B(n_15),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_29),
.B(n_14),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g30 ( 
.A1(n_18),
.A2(n_17),
.B1(n_11),
.B2(n_19),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_30),
.A2(n_31),
.B1(n_23),
.B2(n_11),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_32),
.A2(n_35),
.B1(n_13),
.B2(n_9),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_27),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_33),
.B(n_34),
.Y(n_42)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g35 ( 
.A1(n_31),
.A2(n_17),
.B(n_21),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_SL g36 ( 
.A1(n_28),
.A2(n_30),
.B(n_29),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_21),
.C(n_20),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_37),
.A2(n_40),
.B1(n_13),
.B2(n_9),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_22),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_38),
.B(n_39),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_22),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_26),
.B(n_10),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_25),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_39),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_44),
.Y(n_49)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g50 ( 
.A1(n_46),
.A2(n_35),
.B(n_32),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_L g53 ( 
.A1(n_50),
.A2(n_43),
.B(n_41),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_49),
.A2(n_46),
.B1(n_42),
.B2(n_36),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g54 ( 
.A(n_52),
.B(n_53),
.Y(n_54)
);

NAND3xp33_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_41),
.C(n_48),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_55),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_54),
.A2(n_47),
.B1(n_25),
.B2(n_7),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_57),
.Y(n_58)
);

INVxp33_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

OAI221xp5_ASAP7_75t_L g60 ( 
.A1(n_59),
.A2(n_56),
.B1(n_25),
.B2(n_4),
.C(n_3),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g61 ( 
.A(n_60),
.B(n_4),
.Y(n_61)
);


endmodule