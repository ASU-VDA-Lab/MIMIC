module fake_aes_6372_n_36 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_36);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_36;
wire n_20;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
CKINVDCx5p33_ASAP7_75t_R g11 ( .A(n_9), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_7), .Y(n_12) );
INVx2_ASAP7_75t_L g13 ( .A(n_1), .Y(n_13) );
CKINVDCx20_ASAP7_75t_R g14 ( .A(n_3), .Y(n_14) );
NAND2xp5_ASAP7_75t_SL g15 ( .A(n_2), .B(n_3), .Y(n_15) );
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_8), .Y(n_16) );
AND3x1_ASAP7_75t_L g17 ( .A(n_10), .B(n_7), .C(n_5), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_13), .Y(n_18) );
OAI22xp5_ASAP7_75t_L g19 ( .A1(n_17), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_19) );
NOR2xp33_ASAP7_75t_L g20 ( .A(n_12), .B(n_0), .Y(n_20) );
AOI22xp5_ASAP7_75t_L g21 ( .A1(n_17), .A2(n_4), .B1(n_5), .B2(n_6), .Y(n_21) );
INVx3_ASAP7_75t_SL g22 ( .A(n_18), .Y(n_22) );
OA21x2_ASAP7_75t_L g23 ( .A1(n_20), .A2(n_13), .B(n_12), .Y(n_23) );
OAI211xp5_ASAP7_75t_L g24 ( .A1(n_21), .A2(n_13), .B(n_15), .C(n_14), .Y(n_24) );
AND2x6_ASAP7_75t_L g25 ( .A(n_22), .B(n_19), .Y(n_25) );
AND2x4_ASAP7_75t_SL g26 ( .A(n_22), .B(n_15), .Y(n_26) );
AND2x2_ASAP7_75t_L g27 ( .A(n_26), .B(n_23), .Y(n_27) );
AND2x2_ASAP7_75t_L g28 ( .A(n_25), .B(n_24), .Y(n_28) );
INVx2_ASAP7_75t_L g29 ( .A(n_27), .Y(n_29) );
OAI22xp5_ASAP7_75t_SL g30 ( .A1(n_28), .A2(n_25), .B1(n_11), .B2(n_16), .Y(n_30) );
AND2x2_ASAP7_75t_SL g31 ( .A(n_30), .B(n_23), .Y(n_31) );
NAND2xp5_ASAP7_75t_L g32 ( .A(n_29), .B(n_25), .Y(n_32) );
OR2x6_ASAP7_75t_L g33 ( .A(n_32), .B(n_23), .Y(n_33) );
INVxp67_ASAP7_75t_SL g34 ( .A(n_31), .Y(n_34) );
AOI22xp33_ASAP7_75t_SL g35 ( .A1(n_34), .A2(n_31), .B1(n_4), .B2(n_6), .Y(n_35) );
AOI22xp33_ASAP7_75t_L g36 ( .A1(n_35), .A2(n_33), .B1(n_34), .B2(n_31), .Y(n_36) );
endmodule