module real_jpeg_5435_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_104;
wire n_153;
wire n_64;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_113;
wire n_155;
wire n_120;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_134;
wire n_72;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

INVx8_ASAP7_75t_L g63 ( 
.A(n_0),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_1),
.B(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_2),
.B(n_32),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_2),
.B(n_48),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_2),
.B(n_42),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_3),
.B(n_54),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_3),
.B(n_79),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_3),
.B(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_3),
.B(n_48),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_3),
.B(n_45),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_5),
.B(n_45),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_5),
.B(n_60),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_5),
.B(n_129),
.Y(n_128)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_6),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_7),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_7),
.Y(n_129)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_9),
.B(n_23),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_9),
.B(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_9),
.B(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_9),
.B(n_109),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_9),
.B(n_134),
.Y(n_133)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_11),
.B(n_36),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_11),
.B(n_68),
.Y(n_67)
);

AND2x6_ASAP7_75t_SL g27 ( 
.A(n_12),
.B(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_12),
.B(n_76),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_12),
.B(n_54),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_12),
.B(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_12),
.B(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_12),
.B(n_138),
.Y(n_137)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_13),
.Y(n_92)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_13),
.Y(n_115)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_102),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_100),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_82),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_18),
.B(n_82),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_50),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_37),
.Y(n_19)
);

XNOR2x1_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_29),
.Y(n_20)
);

XNOR2x1_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_27),
.Y(n_21)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_26),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_34),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_30),
.A2(n_31),
.B1(n_34),
.B2(n_35),
.Y(n_38)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_33),
.Y(n_110)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_39),
.C(n_43),
.Y(n_37)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_38),
.B(n_39),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_41),
.Y(n_39)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_43),
.B(n_84),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_47),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_44),
.B(n_47),
.Y(n_145)
);

BUFx8_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

XOR2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_64),
.Y(n_50)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_59),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_58),
.Y(n_52)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_61),
.Y(n_96)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_63),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_66),
.B1(n_72),
.B2(n_73),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_69),
.Y(n_66)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_71),
.Y(n_120)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_73),
.Y(n_72)
);

MAJx2_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_78),
.C(n_80),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_74),
.A2(n_75),
.B1(n_80),
.B2(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_78),
.B(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_80),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_85),
.C(n_97),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_83),
.B(n_155),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_85),
.B(n_97),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_88),
.C(n_93),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_87),
.B(n_89),
.Y(n_148)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_92),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_93),
.B(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

OAI21x1_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_151),
.B(n_156),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_142),
.B(n_150),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_122),
.B(n_141),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_116),
.B(n_121),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_107),
.B(n_112),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_107),
.B(n_112),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_111),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_117),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_108),
.B(n_111),
.Y(n_123)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_124),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_123),
.B(n_124),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_126),
.B1(n_130),
.B2(n_131),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_125),
.B(n_133),
.C(n_136),
.Y(n_149)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_SL g126 ( 
.A(n_127),
.B(n_128),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_127),
.B(n_128),
.Y(n_146)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_133),
.B1(n_136),
.B2(n_137),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_143),
.B(n_149),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_143),
.B(n_149),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_147),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_145),
.B(n_146),
.C(n_153),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_147),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_154),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_152),
.B(n_154),
.Y(n_156)
);


endmodule