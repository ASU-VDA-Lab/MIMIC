module fake_aes_8167_n_717 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_717);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_717;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_307;
wire n_191;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_420;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_195;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g81 ( .A(n_59), .Y(n_81) );
INVxp67_ASAP7_75t_SL g82 ( .A(n_52), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_31), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_74), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_12), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_64), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_60), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_15), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_15), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_33), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_43), .Y(n_91) );
INVx2_ASAP7_75t_L g92 ( .A(n_65), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_8), .Y(n_93) );
CKINVDCx20_ASAP7_75t_R g94 ( .A(n_24), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_30), .Y(n_95) );
INVx2_ASAP7_75t_L g96 ( .A(n_47), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_49), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_18), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_69), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_32), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_57), .Y(n_101) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_10), .Y(n_102) );
INVxp33_ASAP7_75t_SL g103 ( .A(n_29), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_2), .Y(n_104) );
INVxp33_ASAP7_75t_SL g105 ( .A(n_44), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_20), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_73), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_5), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_46), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_2), .Y(n_110) );
BUFx3_ASAP7_75t_L g111 ( .A(n_54), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_72), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_7), .Y(n_113) );
INVxp67_ASAP7_75t_SL g114 ( .A(n_25), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_20), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_26), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_75), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_8), .Y(n_118) );
INVxp33_ASAP7_75t_L g119 ( .A(n_58), .Y(n_119) );
INVxp67_ASAP7_75t_L g120 ( .A(n_3), .Y(n_120) );
INVxp67_ASAP7_75t_SL g121 ( .A(n_36), .Y(n_121) );
BUFx3_ASAP7_75t_L g122 ( .A(n_7), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_28), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_48), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_39), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_38), .Y(n_126) );
BUFx2_ASAP7_75t_L g127 ( .A(n_23), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_55), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_67), .Y(n_129) );
AND2x2_ASAP7_75t_L g130 ( .A(n_127), .B(n_0), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_92), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_81), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_81), .Y(n_133) );
CKINVDCx20_ASAP7_75t_R g134 ( .A(n_94), .Y(n_134) );
BUFx8_ASAP7_75t_L g135 ( .A(n_127), .Y(n_135) );
HB1xp67_ASAP7_75t_L g136 ( .A(n_122), .Y(n_136) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_111), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_92), .Y(n_138) );
CKINVDCx16_ASAP7_75t_R g139 ( .A(n_122), .Y(n_139) );
INVx3_ASAP7_75t_L g140 ( .A(n_83), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_103), .Y(n_141) );
CKINVDCx20_ASAP7_75t_R g142 ( .A(n_102), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_96), .Y(n_143) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_111), .Y(n_144) );
BUFx2_ASAP7_75t_L g145 ( .A(n_120), .Y(n_145) );
BUFx3_ASAP7_75t_L g146 ( .A(n_96), .Y(n_146) );
INVxp67_ASAP7_75t_L g147 ( .A(n_85), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_83), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_105), .Y(n_149) );
CKINVDCx16_ASAP7_75t_R g150 ( .A(n_106), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_84), .Y(n_151) );
NAND2xp5_ASAP7_75t_SL g152 ( .A(n_119), .B(n_0), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_84), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_86), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_86), .Y(n_155) );
NAND2xp33_ASAP7_75t_L g156 ( .A(n_129), .B(n_35), .Y(n_156) );
CKINVDCx5p33_ASAP7_75t_R g157 ( .A(n_109), .Y(n_157) );
BUFx2_ASAP7_75t_L g158 ( .A(n_85), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_87), .Y(n_159) );
CKINVDCx20_ASAP7_75t_R g160 ( .A(n_88), .Y(n_160) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_87), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_90), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_90), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_88), .B(n_1), .Y(n_164) );
CKINVDCx16_ASAP7_75t_R g165 ( .A(n_91), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_91), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_95), .Y(n_167) );
CKINVDCx5p33_ASAP7_75t_R g168 ( .A(n_112), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_95), .Y(n_169) );
AND2x4_ASAP7_75t_L g170 ( .A(n_89), .B(n_1), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_97), .Y(n_171) );
CKINVDCx20_ASAP7_75t_R g172 ( .A(n_89), .Y(n_172) );
INVx3_ASAP7_75t_L g173 ( .A(n_97), .Y(n_173) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_135), .B(n_116), .Y(n_174) );
INVx1_ASAP7_75t_SL g175 ( .A(n_139), .Y(n_175) );
INVx3_ASAP7_75t_L g176 ( .A(n_170), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_137), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_136), .B(n_117), .Y(n_178) );
BUFx2_ASAP7_75t_L g179 ( .A(n_135), .Y(n_179) );
AND2x2_ASAP7_75t_L g180 ( .A(n_136), .B(n_118), .Y(n_180) );
AND2x2_ASAP7_75t_L g181 ( .A(n_130), .B(n_118), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_161), .Y(n_182) );
AND2x4_ASAP7_75t_L g183 ( .A(n_158), .B(n_93), .Y(n_183) );
INVxp67_ASAP7_75t_L g184 ( .A(n_135), .Y(n_184) );
AND3x4_ASAP7_75t_L g185 ( .A(n_170), .B(n_114), .C(n_110), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_161), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_161), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_161), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_161), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_161), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_137), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_141), .B(n_129), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_137), .Y(n_193) );
OAI22xp5_ASAP7_75t_SL g194 ( .A1(n_134), .A2(n_104), .B1(n_98), .B2(n_93), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_137), .Y(n_195) );
INVx3_ASAP7_75t_L g196 ( .A(n_170), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_135), .B(n_128), .Y(n_197) );
INVx3_ASAP7_75t_L g198 ( .A(n_170), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_161), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_140), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_140), .Y(n_201) );
OR2x6_ASAP7_75t_L g202 ( .A(n_130), .B(n_98), .Y(n_202) );
AND2x2_ASAP7_75t_L g203 ( .A(n_130), .B(n_104), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_140), .Y(n_204) );
NAND2x1_ASAP7_75t_L g205 ( .A(n_170), .B(n_128), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_137), .Y(n_206) );
INVx4_ASAP7_75t_L g207 ( .A(n_140), .Y(n_207) );
AO22x2_ASAP7_75t_L g208 ( .A1(n_132), .A2(n_126), .B1(n_125), .B2(n_124), .Y(n_208) );
BUFx6f_ASAP7_75t_L g209 ( .A(n_137), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_137), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_140), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_144), .Y(n_212) );
AND2x6_ASAP7_75t_L g213 ( .A(n_173), .B(n_126), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_144), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_173), .Y(n_215) );
OAI22xp5_ASAP7_75t_L g216 ( .A1(n_165), .A2(n_108), .B1(n_113), .B2(n_115), .Y(n_216) );
NAND3xp33_ASAP7_75t_L g217 ( .A(n_135), .B(n_125), .C(n_124), .Y(n_217) );
CKINVDCx20_ASAP7_75t_R g218 ( .A(n_142), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_144), .Y(n_219) );
INVx8_ASAP7_75t_L g220 ( .A(n_173), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_173), .Y(n_221) );
AND2x4_ASAP7_75t_L g222 ( .A(n_158), .B(n_107), .Y(n_222) );
AO22x2_ASAP7_75t_L g223 ( .A1(n_132), .A2(n_123), .B1(n_107), .B2(n_101), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_139), .B(n_123), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_173), .Y(n_225) );
INVx2_ASAP7_75t_SL g226 ( .A(n_145), .Y(n_226) );
INVx4_ASAP7_75t_SL g227 ( .A(n_144), .Y(n_227) );
AND2x2_ASAP7_75t_L g228 ( .A(n_147), .B(n_101), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_155), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g230 ( .A(n_149), .B(n_100), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_155), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_165), .B(n_100), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_155), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_163), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_229), .Y(n_235) );
AND2x2_ASAP7_75t_L g236 ( .A(n_183), .B(n_145), .Y(n_236) );
NOR3xp33_ASAP7_75t_SL g237 ( .A(n_194), .B(n_150), .C(n_168), .Y(n_237) );
NOR3xp33_ASAP7_75t_SL g238 ( .A(n_194), .B(n_150), .C(n_157), .Y(n_238) );
CKINVDCx6p67_ASAP7_75t_R g239 ( .A(n_179), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_226), .B(n_147), .Y(n_240) );
OAI22xp33_ASAP7_75t_L g241 ( .A1(n_202), .A2(n_172), .B1(n_160), .B2(n_164), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_229), .Y(n_242) );
INVx1_ASAP7_75t_SL g243 ( .A(n_179), .Y(n_243) );
INVx3_ASAP7_75t_L g244 ( .A(n_207), .Y(n_244) );
NOR2xp33_ASAP7_75t_SL g245 ( .A(n_220), .B(n_171), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_226), .B(n_133), .Y(n_246) );
BUFx6f_ASAP7_75t_L g247 ( .A(n_220), .Y(n_247) );
INVx4_ASAP7_75t_L g248 ( .A(n_220), .Y(n_248) );
BUFx3_ASAP7_75t_L g249 ( .A(n_231), .Y(n_249) );
NAND3xp33_ASAP7_75t_L g250 ( .A(n_192), .B(n_152), .C(n_156), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_231), .Y(n_251) );
AND2x4_ASAP7_75t_L g252 ( .A(n_202), .B(n_152), .Y(n_252) );
AND2x4_ASAP7_75t_L g253 ( .A(n_202), .B(n_171), .Y(n_253) );
BUFx2_ASAP7_75t_L g254 ( .A(n_175), .Y(n_254) );
NAND2xp33_ASAP7_75t_SL g255 ( .A(n_185), .B(n_164), .Y(n_255) );
AND2x2_ASAP7_75t_L g256 ( .A(n_183), .B(n_148), .Y(n_256) );
AOI21xp33_ASAP7_75t_L g257 ( .A1(n_205), .A2(n_148), .B(n_133), .Y(n_257) );
NOR3xp33_ASAP7_75t_SL g258 ( .A(n_216), .B(n_153), .C(n_159), .Y(n_258) );
NOR2x1p5_ASAP7_75t_L g259 ( .A(n_183), .B(n_151), .Y(n_259) );
INVx2_ASAP7_75t_L g260 ( .A(n_207), .Y(n_260) );
NOR2xp33_ASAP7_75t_R g261 ( .A(n_218), .B(n_162), .Y(n_261) );
CKINVDCx5p33_ASAP7_75t_R g262 ( .A(n_202), .Y(n_262) );
OR2x2_ASAP7_75t_L g263 ( .A(n_232), .B(n_154), .Y(n_263) );
BUFx10_ASAP7_75t_L g264 ( .A(n_222), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_207), .B(n_151), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_222), .B(n_162), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_233), .Y(n_267) );
BUFx2_ASAP7_75t_L g268 ( .A(n_202), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_233), .Y(n_269) );
AND2x6_ASAP7_75t_L g270 ( .A(n_176), .B(n_99), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_234), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_234), .Y(n_272) );
AND2x4_ASAP7_75t_L g273 ( .A(n_184), .B(n_159), .Y(n_273) );
BUFx12f_ASAP7_75t_L g274 ( .A(n_183), .Y(n_274) );
NOR2xp33_ASAP7_75t_L g275 ( .A(n_230), .B(n_154), .Y(n_275) );
OR2x6_ASAP7_75t_L g276 ( .A(n_222), .B(n_153), .Y(n_276) );
A2O1A1Ixp33_ASAP7_75t_L g277 ( .A1(n_176), .A2(n_198), .B(n_196), .C(n_205), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_200), .Y(n_278) );
NOR3xp33_ASAP7_75t_SL g279 ( .A(n_224), .B(n_82), .C(n_121), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_200), .Y(n_280) );
NOR2xp33_ASAP7_75t_L g281 ( .A(n_222), .B(n_169), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_228), .B(n_169), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_228), .B(n_169), .Y(n_283) );
OR2x6_ASAP7_75t_L g284 ( .A(n_174), .B(n_167), .Y(n_284) );
AND2x2_ASAP7_75t_L g285 ( .A(n_181), .B(n_146), .Y(n_285) );
AOI22xp5_ASAP7_75t_L g286 ( .A1(n_185), .A2(n_167), .B1(n_166), .B2(n_163), .Y(n_286) );
INVx4_ASAP7_75t_L g287 ( .A(n_220), .Y(n_287) );
A2O1A1Ixp33_ASAP7_75t_L g288 ( .A1(n_176), .A2(n_167), .B(n_166), .C(n_163), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_220), .B(n_166), .Y(n_289) );
AND2x4_ASAP7_75t_L g290 ( .A(n_181), .B(n_146), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_208), .Y(n_291) );
NAND3xp33_ASAP7_75t_SL g292 ( .A(n_185), .B(n_99), .C(n_131), .Y(n_292) );
INVx1_ASAP7_75t_SL g293 ( .A(n_213), .Y(n_293) );
AOI22xp5_ASAP7_75t_L g294 ( .A1(n_197), .A2(n_146), .B1(n_143), .B2(n_138), .Y(n_294) );
BUFx6f_ASAP7_75t_L g295 ( .A(n_213), .Y(n_295) );
NOR2xp33_ASAP7_75t_R g296 ( .A(n_196), .B(n_41), .Y(n_296) );
CKINVDCx11_ASAP7_75t_R g297 ( .A(n_209), .Y(n_297) );
NAND3xp33_ASAP7_75t_SL g298 ( .A(n_217), .B(n_131), .C(n_138), .Y(n_298) );
INVx6_ASAP7_75t_L g299 ( .A(n_213), .Y(n_299) );
INVx3_ASAP7_75t_L g300 ( .A(n_196), .Y(n_300) );
AND2x4_ASAP7_75t_L g301 ( .A(n_203), .B(n_143), .Y(n_301) );
BUFx3_ASAP7_75t_L g302 ( .A(n_247), .Y(n_302) );
AND2x4_ASAP7_75t_L g303 ( .A(n_248), .B(n_203), .Y(n_303) );
AOI21xp5_ASAP7_75t_L g304 ( .A1(n_277), .A2(n_198), .B(n_225), .Y(n_304) );
AND2x2_ASAP7_75t_L g305 ( .A(n_276), .B(n_180), .Y(n_305) );
HB1xp67_ASAP7_75t_L g306 ( .A(n_276), .Y(n_306) );
AOI21xp5_ASAP7_75t_L g307 ( .A1(n_265), .A2(n_198), .B(n_225), .Y(n_307) );
NOR2x1_ASAP7_75t_SL g308 ( .A(n_276), .B(n_201), .Y(n_308) );
AOI21xp5_ASAP7_75t_L g309 ( .A1(n_265), .A2(n_204), .B(n_211), .Y(n_309) );
OAI22xp5_ASAP7_75t_L g310 ( .A1(n_253), .A2(n_208), .B1(n_223), .B2(n_178), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_278), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_253), .B(n_180), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_300), .Y(n_313) );
BUFx2_ASAP7_75t_L g314 ( .A(n_274), .Y(n_314) );
BUFx2_ASAP7_75t_L g315 ( .A(n_248), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_300), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_285), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_280), .Y(n_318) );
OR2x6_ASAP7_75t_L g319 ( .A(n_268), .B(n_208), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_249), .Y(n_320) );
BUFx2_ASAP7_75t_L g321 ( .A(n_287), .Y(n_321) );
AOI21xp5_ASAP7_75t_L g322 ( .A1(n_266), .A2(n_201), .B(n_221), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_290), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_290), .Y(n_324) );
BUFx3_ASAP7_75t_L g325 ( .A(n_247), .Y(n_325) );
NAND2x1p5_ASAP7_75t_L g326 ( .A(n_287), .B(n_204), .Y(n_326) );
NOR2x1_ASAP7_75t_SL g327 ( .A(n_295), .B(n_247), .Y(n_327) );
AOI22xp5_ASAP7_75t_L g328 ( .A1(n_255), .A2(n_223), .B1(n_208), .B2(n_213), .Y(n_328) );
OAI22xp33_ASAP7_75t_L g329 ( .A1(n_262), .A2(n_215), .B1(n_211), .B2(n_221), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_235), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_242), .Y(n_331) );
BUFx3_ASAP7_75t_L g332 ( .A(n_239), .Y(n_332) );
AND3x1_ASAP7_75t_SL g333 ( .A(n_238), .B(n_3), .C(n_4), .Y(n_333) );
OR2x6_ASAP7_75t_L g334 ( .A(n_299), .B(n_223), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_256), .B(n_223), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_251), .Y(n_336) );
BUFx2_ASAP7_75t_L g337 ( .A(n_254), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_266), .B(n_213), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_275), .B(n_213), .Y(n_339) );
BUFx6f_ASAP7_75t_L g340 ( .A(n_295), .Y(n_340) );
OAI22xp5_ASAP7_75t_L g341 ( .A1(n_291), .A2(n_215), .B1(n_138), .B2(n_143), .Y(n_341) );
INVx3_ASAP7_75t_L g342 ( .A(n_244), .Y(n_342) );
INVxp67_ASAP7_75t_L g343 ( .A(n_236), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_267), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_271), .Y(n_345) );
NOR2xp33_ASAP7_75t_R g346 ( .A(n_292), .B(n_213), .Y(n_346) );
INVx1_ASAP7_75t_SL g347 ( .A(n_261), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_263), .B(n_131), .Y(n_348) );
INVxp67_ASAP7_75t_SL g349 ( .A(n_295), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_240), .B(n_144), .Y(n_350) );
INVx3_ASAP7_75t_L g351 ( .A(n_244), .Y(n_351) );
AOI21xp5_ASAP7_75t_L g352 ( .A1(n_257), .A2(n_182), .B(n_186), .Y(n_352) );
AND2x4_ASAP7_75t_L g353 ( .A(n_259), .B(n_227), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_269), .Y(n_354) );
AOI22xp5_ASAP7_75t_L g355 ( .A1(n_292), .A2(n_144), .B1(n_182), .B2(n_186), .Y(n_355) );
NOR2xp33_ASAP7_75t_L g356 ( .A(n_343), .B(n_241), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_317), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_330), .Y(n_358) );
INVx2_ASAP7_75t_SL g359 ( .A(n_315), .Y(n_359) );
INVx3_ASAP7_75t_L g360 ( .A(n_326), .Y(n_360) );
NOR2xp67_ASAP7_75t_SL g361 ( .A(n_340), .B(n_299), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_330), .Y(n_362) );
AOI22xp5_ASAP7_75t_L g363 ( .A1(n_334), .A2(n_243), .B1(n_252), .B2(n_273), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_331), .Y(n_364) );
AOI21xp5_ASAP7_75t_L g365 ( .A1(n_339), .A2(n_245), .B(n_257), .Y(n_365) );
AND2x2_ASAP7_75t_SL g366 ( .A(n_315), .B(n_245), .Y(n_366) );
INVx2_ASAP7_75t_L g367 ( .A(n_311), .Y(n_367) );
INVx4_ASAP7_75t_L g368 ( .A(n_334), .Y(n_368) );
OAI22xp33_ASAP7_75t_L g369 ( .A1(n_334), .A2(n_243), .B1(n_286), .B2(n_282), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_303), .B(n_252), .Y(n_370) );
OR2x2_ASAP7_75t_L g371 ( .A(n_337), .B(n_282), .Y(n_371) );
OAI22xp5_ASAP7_75t_L g372 ( .A1(n_334), .A2(n_273), .B1(n_283), .B2(n_281), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_331), .Y(n_373) );
OAI22xp5_ASAP7_75t_L g374 ( .A1(n_319), .A2(n_283), .B1(n_289), .B2(n_246), .Y(n_374) );
BUFx2_ASAP7_75t_SL g375 ( .A(n_321), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_303), .B(n_264), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_311), .Y(n_377) );
NAND2xp33_ASAP7_75t_SL g378 ( .A(n_346), .B(n_296), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_336), .Y(n_379) );
CKINVDCx20_ASAP7_75t_R g380 ( .A(n_337), .Y(n_380) );
OAI21xp5_ASAP7_75t_L g381 ( .A1(n_307), .A2(n_288), .B(n_250), .Y(n_381) );
AO31x2_ASAP7_75t_L g382 ( .A1(n_310), .A2(n_214), .A3(n_210), .B(n_177), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_336), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_303), .B(n_264), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g385 ( .A1(n_305), .A2(n_270), .B1(n_301), .B2(n_284), .Y(n_385) );
NAND2x1_ASAP7_75t_L g386 ( .A(n_340), .B(n_270), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_312), .B(n_258), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_305), .B(n_301), .Y(n_388) );
OAI22xp5_ASAP7_75t_L g389 ( .A1(n_319), .A2(n_289), .B1(n_272), .B2(n_284), .Y(n_389) );
OAI21x1_ASAP7_75t_SL g390 ( .A1(n_368), .A2(n_308), .B(n_328), .Y(n_390) );
OAI22xp5_ASAP7_75t_L g391 ( .A1(n_372), .A2(n_319), .B1(n_335), .B2(n_348), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_373), .B(n_344), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_373), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_367), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_383), .B(n_319), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_371), .B(n_323), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_367), .Y(n_397) );
OAI22xp5_ASAP7_75t_L g398 ( .A1(n_369), .A2(n_354), .B1(n_344), .B2(n_306), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_377), .Y(n_399) );
OAI22xp5_ASAP7_75t_L g400 ( .A1(n_368), .A2(n_354), .B1(n_321), .B2(n_345), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g401 ( .A1(n_356), .A2(n_374), .B1(n_387), .B2(n_380), .Y(n_401) );
NAND3xp33_ASAP7_75t_L g402 ( .A(n_381), .B(n_350), .C(n_238), .Y(n_402) );
OA21x2_ASAP7_75t_L g403 ( .A1(n_365), .A2(n_304), .B(n_352), .Y(n_403) );
CKINVDCx11_ASAP7_75t_R g404 ( .A(n_380), .Y(n_404) );
OAI22xp33_ASAP7_75t_L g405 ( .A1(n_363), .A2(n_347), .B1(n_332), .B2(n_314), .Y(n_405) );
AND2x4_ASAP7_75t_L g406 ( .A(n_360), .B(n_308), .Y(n_406) );
AO21x1_ASAP7_75t_L g407 ( .A1(n_389), .A2(n_341), .B(n_338), .Y(n_407) );
NAND3xp33_ASAP7_75t_L g408 ( .A(n_385), .B(n_355), .C(n_237), .Y(n_408) );
OAI211xp5_ASAP7_75t_SL g409 ( .A1(n_357), .A2(n_279), .B(n_324), .C(n_294), .Y(n_409) );
AOI221xp5_ASAP7_75t_L g410 ( .A1(n_388), .A2(n_314), .B1(n_329), .B2(n_332), .C(n_322), .Y(n_410) );
INVx3_ASAP7_75t_L g411 ( .A(n_360), .Y(n_411) );
AOI22xp33_ASAP7_75t_SL g412 ( .A1(n_375), .A2(n_270), .B1(n_333), .B2(n_320), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_368), .A2(n_270), .B1(n_284), .B2(n_353), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_383), .B(n_345), .Y(n_414) );
AOI22xp33_ASAP7_75t_L g415 ( .A1(n_375), .A2(n_270), .B1(n_353), .B2(n_313), .Y(n_415) );
OAI22xp5_ASAP7_75t_L g416 ( .A1(n_366), .A2(n_318), .B1(n_326), .B2(n_325), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_358), .Y(n_417) );
AOI22xp33_ASAP7_75t_SL g418 ( .A1(n_366), .A2(n_326), .B1(n_353), .B2(n_327), .Y(n_418) );
OR2x2_ASAP7_75t_L g419 ( .A(n_393), .B(n_371), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_394), .Y(n_420) );
INVxp67_ASAP7_75t_L g421 ( .A(n_414), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_414), .B(n_393), .Y(n_422) );
OAI33xp33_ASAP7_75t_L g423 ( .A1(n_405), .A2(n_362), .A3(n_379), .B1(n_364), .B2(n_370), .B3(n_187), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_401), .B(n_376), .Y(n_424) );
OAI322xp33_ASAP7_75t_L g425 ( .A1(n_417), .A2(n_144), .A3(n_359), .B1(n_377), .B2(n_313), .C1(n_316), .C2(n_187), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_396), .B(n_417), .Y(n_426) );
OAI33xp33_ASAP7_75t_L g427 ( .A1(n_398), .A2(n_199), .A3(n_188), .B1(n_189), .B2(n_190), .B3(n_316), .Y(n_427) );
AOI22xp5_ASAP7_75t_L g428 ( .A1(n_391), .A2(n_376), .B1(n_384), .B2(n_359), .Y(n_428) );
OAI22xp5_ASAP7_75t_L g429 ( .A1(n_391), .A2(n_360), .B1(n_384), .B2(n_386), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_394), .B(n_318), .Y(n_430) );
AOI22xp5_ASAP7_75t_L g431 ( .A1(n_410), .A2(n_378), .B1(n_298), .B2(n_342), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_394), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_397), .Y(n_433) );
OAI22xp33_ASAP7_75t_L g434 ( .A1(n_400), .A2(n_386), .B1(n_325), .B2(n_302), .Y(n_434) );
OAI22xp5_ASAP7_75t_L g435 ( .A1(n_398), .A2(n_302), .B1(n_378), .B2(n_299), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_397), .B(n_382), .Y(n_436) );
NAND2xp33_ASAP7_75t_R g437 ( .A(n_406), .B(n_411), .Y(n_437) );
AOI31xp33_ASAP7_75t_L g438 ( .A1(n_412), .A2(n_418), .A3(n_416), .B(n_400), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_392), .B(n_382), .Y(n_439) );
NOR5xp2_ASAP7_75t_SL g440 ( .A(n_416), .B(n_4), .C(n_5), .D(n_6), .E(n_9), .Y(n_440) );
AOI22xp5_ASAP7_75t_L g441 ( .A1(n_408), .A2(n_298), .B1(n_342), .B2(n_351), .Y(n_441) );
BUFx3_ASAP7_75t_L g442 ( .A(n_404), .Y(n_442) );
AND2x4_ASAP7_75t_L g443 ( .A(n_406), .B(n_382), .Y(n_443) );
OAI31xp33_ASAP7_75t_L g444 ( .A1(n_408), .A2(n_351), .A3(n_342), .B(n_293), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_397), .B(n_382), .Y(n_445) );
NAND3xp33_ASAP7_75t_L g446 ( .A(n_402), .B(n_297), .C(n_209), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_399), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_399), .B(n_382), .Y(n_448) );
BUFx2_ASAP7_75t_L g449 ( .A(n_406), .Y(n_449) );
OAI22xp33_ASAP7_75t_L g450 ( .A1(n_392), .A2(n_351), .B1(n_340), .B2(n_293), .Y(n_450) );
AO21x2_ASAP7_75t_L g451 ( .A1(n_407), .A2(n_210), .B(n_191), .Y(n_451) );
NAND4xp25_ASAP7_75t_L g452 ( .A(n_402), .B(n_199), .C(n_188), .D(n_189), .Y(n_452) );
OAI21xp5_ASAP7_75t_L g453 ( .A1(n_409), .A2(n_309), .B(n_349), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_433), .Y(n_454) );
NAND3xp33_ASAP7_75t_L g455 ( .A(n_452), .B(n_399), .C(n_395), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_433), .Y(n_456) );
AOI221xp5_ASAP7_75t_L g457 ( .A1(n_438), .A2(n_395), .B1(n_407), .B2(n_390), .C(n_413), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_447), .Y(n_458) );
INVx5_ASAP7_75t_L g459 ( .A(n_430), .Y(n_459) );
OAI21xp5_ASAP7_75t_SL g460 ( .A1(n_428), .A2(n_415), .B(n_406), .Y(n_460) );
OR2x2_ASAP7_75t_L g461 ( .A(n_439), .B(n_411), .Y(n_461) );
INVx4_ASAP7_75t_L g462 ( .A(n_449), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_447), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_436), .Y(n_464) );
AND2x4_ASAP7_75t_L g465 ( .A(n_443), .B(n_411), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_436), .Y(n_466) );
NOR4xp25_ASAP7_75t_L g467 ( .A(n_426), .B(n_411), .C(n_9), .D(n_10), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_445), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_445), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_422), .B(n_403), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_448), .Y(n_471) );
INVx4_ASAP7_75t_L g472 ( .A(n_449), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_422), .B(n_390), .Y(n_473) );
HB1xp67_ASAP7_75t_L g474 ( .A(n_421), .Y(n_474) );
HB1xp67_ASAP7_75t_L g475 ( .A(n_430), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_448), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_420), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_420), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_432), .B(n_403), .Y(n_479) );
OAI31xp33_ASAP7_75t_L g480 ( .A1(n_429), .A2(n_6), .A3(n_11), .B(n_12), .Y(n_480) );
NOR3xp33_ASAP7_75t_L g481 ( .A(n_423), .B(n_177), .C(n_219), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_432), .B(n_403), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_443), .B(n_403), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_443), .Y(n_484) );
BUFx2_ASAP7_75t_L g485 ( .A(n_434), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_419), .B(n_327), .Y(n_486) );
INVx2_ASAP7_75t_L g487 ( .A(n_451), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_419), .B(n_11), .Y(n_488) );
OAI22xp5_ASAP7_75t_L g489 ( .A1(n_424), .A2(n_431), .B1(n_446), .B2(n_435), .Y(n_489) );
INVx6_ASAP7_75t_L g490 ( .A(n_442), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_451), .B(n_13), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_451), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_441), .B(n_13), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_441), .B(n_14), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_453), .B(n_14), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_425), .Y(n_496) );
AND2x4_ASAP7_75t_L g497 ( .A(n_437), .B(n_209), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_444), .B(n_16), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_442), .B(n_16), .Y(n_499) );
AOI33xp33_ASAP7_75t_L g500 ( .A1(n_440), .A2(n_190), .A3(n_191), .B1(n_193), .B2(n_195), .B3(n_206), .Y(n_500) );
INVx3_ASAP7_75t_L g501 ( .A(n_427), .Y(n_501) );
OAI33xp33_ASAP7_75t_L g502 ( .A1(n_440), .A2(n_17), .A3(n_18), .B1(n_19), .B2(n_21), .B3(n_22), .Y(n_502) );
AND2x4_ASAP7_75t_L g503 ( .A(n_450), .B(n_209), .Y(n_503) );
OAI33xp33_ASAP7_75t_L g504 ( .A1(n_488), .A2(n_17), .A3(n_19), .B1(n_21), .B2(n_22), .B3(n_23), .Y(n_504) );
NAND2xp33_ASAP7_75t_SL g505 ( .A(n_500), .B(n_361), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_474), .B(n_24), .Y(n_506) );
AND2x4_ASAP7_75t_L g507 ( .A(n_484), .B(n_209), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_479), .Y(n_508) );
OR2x2_ASAP7_75t_L g509 ( .A(n_466), .B(n_25), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_475), .B(n_219), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_454), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_464), .B(n_214), .Y(n_512) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_457), .A2(n_361), .B1(n_212), .B2(n_206), .Y(n_513) );
OAI21xp33_ASAP7_75t_L g514 ( .A1(n_467), .A2(n_212), .B(n_195), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_466), .B(n_193), .Y(n_515) );
NAND2xp33_ASAP7_75t_R g516 ( .A(n_499), .B(n_27), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_454), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_456), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_464), .B(n_34), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_464), .B(n_37), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_456), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_458), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_468), .B(n_40), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_458), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_468), .B(n_42), .Y(n_525) );
OR2x2_ASAP7_75t_L g526 ( .A(n_471), .B(n_45), .Y(n_526) );
INVx2_ASAP7_75t_L g527 ( .A(n_479), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_463), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_471), .B(n_50), .Y(n_529) );
BUFx2_ASAP7_75t_L g530 ( .A(n_462), .Y(n_530) );
INVx2_ASAP7_75t_SL g531 ( .A(n_459), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_468), .B(n_51), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_469), .B(n_53), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_488), .B(n_56), .Y(n_534) );
OAI31xp33_ASAP7_75t_L g535 ( .A1(n_480), .A2(n_61), .A3(n_62), .B(n_63), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_469), .B(n_66), .Y(n_536) );
OR2x2_ASAP7_75t_L g537 ( .A(n_469), .B(n_68), .Y(n_537) );
NAND3xp33_ASAP7_75t_L g538 ( .A(n_467), .B(n_340), .C(n_260), .Y(n_538) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_490), .B(n_70), .Y(n_539) );
HB1xp67_ASAP7_75t_L g540 ( .A(n_459), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_463), .Y(n_541) );
INVxp67_ASAP7_75t_L g542 ( .A(n_499), .Y(n_542) );
HB1xp67_ASAP7_75t_L g543 ( .A(n_459), .Y(n_543) );
NOR2xp33_ASAP7_75t_L g544 ( .A(n_490), .B(n_71), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_477), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_476), .B(n_76), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_476), .B(n_77), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_476), .B(n_78), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_477), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_470), .B(n_79), .Y(n_550) );
INVxp67_ASAP7_75t_L g551 ( .A(n_455), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_478), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_478), .Y(n_553) );
INVxp67_ASAP7_75t_SL g554 ( .A(n_486), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_470), .B(n_80), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_486), .B(n_227), .Y(n_556) );
NOR2xp33_ASAP7_75t_R g557 ( .A(n_490), .B(n_340), .Y(n_557) );
INVx2_ASAP7_75t_L g558 ( .A(n_482), .Y(n_558) );
NAND4xp75_ASAP7_75t_SL g559 ( .A(n_480), .B(n_227), .C(n_493), .D(n_494), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_484), .B(n_227), .Y(n_560) );
NOR2xp33_ASAP7_75t_R g561 ( .A(n_490), .B(n_459), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_482), .Y(n_562) );
AOI21xp33_ASAP7_75t_L g563 ( .A1(n_551), .A2(n_498), .B(n_495), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_554), .B(n_493), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_517), .Y(n_565) );
INVx2_ASAP7_75t_L g566 ( .A(n_508), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_517), .Y(n_567) );
OAI22xp5_ASAP7_75t_L g568 ( .A1(n_542), .A2(n_460), .B1(n_490), .B2(n_455), .Y(n_568) );
AOI21xp5_ASAP7_75t_L g569 ( .A1(n_514), .A2(n_502), .B(n_460), .Y(n_569) );
NAND2xp5_ASAP7_75t_SL g570 ( .A(n_561), .B(n_497), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_508), .B(n_494), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_530), .B(n_465), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_508), .B(n_491), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_518), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_527), .B(n_491), .Y(n_575) );
AOI21xp33_ASAP7_75t_SL g576 ( .A1(n_516), .A2(n_498), .B(n_489), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_527), .B(n_461), .Y(n_577) );
INVx2_ASAP7_75t_L g578 ( .A(n_527), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_518), .Y(n_579) );
OAI22xp5_ASAP7_75t_L g580 ( .A1(n_530), .A2(n_457), .B1(n_472), .B2(n_462), .Y(n_580) );
INVx2_ASAP7_75t_L g581 ( .A(n_558), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_558), .B(n_465), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_521), .Y(n_583) );
AOI21xp33_ASAP7_75t_L g584 ( .A1(n_506), .A2(n_495), .B(n_489), .Y(n_584) );
AOI221xp5_ASAP7_75t_L g585 ( .A1(n_504), .A2(n_502), .B1(n_473), .B2(n_485), .C(n_496), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_521), .Y(n_586) );
NOR2xp33_ASAP7_75t_L g587 ( .A(n_509), .B(n_485), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_522), .Y(n_588) );
AOI22xp5_ASAP7_75t_L g589 ( .A1(n_505), .A2(n_473), .B1(n_496), .B2(n_501), .Y(n_589) );
AND2x4_ASAP7_75t_L g590 ( .A(n_531), .B(n_465), .Y(n_590) );
OAI32xp33_ASAP7_75t_L g591 ( .A1(n_540), .A2(n_472), .A3(n_462), .B1(n_501), .B2(n_461), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_522), .Y(n_592) );
HB1xp67_ASAP7_75t_L g593 ( .A(n_543), .Y(n_593) );
AO21x1_ASAP7_75t_SL g594 ( .A1(n_526), .A2(n_459), .B(n_462), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_524), .Y(n_595) );
OAI21xp5_ASAP7_75t_SL g596 ( .A1(n_535), .A2(n_497), .B(n_465), .Y(n_596) );
A2O1A1Ixp33_ASAP7_75t_L g597 ( .A1(n_535), .A2(n_501), .B(n_497), .C(n_503), .Y(n_597) );
INVxp67_ASAP7_75t_SL g598 ( .A(n_509), .Y(n_598) );
NOR2xp33_ASAP7_75t_L g599 ( .A(n_534), .B(n_501), .Y(n_599) );
OAI22xp5_ASAP7_75t_SL g600 ( .A1(n_531), .A2(n_472), .B1(n_459), .B2(n_497), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_558), .B(n_483), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_524), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_528), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_528), .Y(n_604) );
NOR2xp33_ASAP7_75t_L g605 ( .A(n_541), .B(n_472), .Y(n_605) );
OA21x2_ASAP7_75t_L g606 ( .A1(n_538), .A2(n_492), .B(n_487), .Y(n_606) );
AND2x2_ASAP7_75t_L g607 ( .A(n_562), .B(n_483), .Y(n_607) );
OAI22xp33_ASAP7_75t_L g608 ( .A1(n_526), .A2(n_459), .B1(n_503), .B2(n_492), .Y(n_608) );
NAND4xp25_ASAP7_75t_L g609 ( .A(n_538), .B(n_481), .C(n_503), .D(n_487), .Y(n_609) );
AOI21xp5_ASAP7_75t_L g610 ( .A1(n_514), .A2(n_503), .B(n_487), .Y(n_610) );
AOI22xp5_ASAP7_75t_L g611 ( .A1(n_513), .A2(n_555), .B1(n_550), .B2(n_539), .Y(n_611) );
OR2x2_ASAP7_75t_L g612 ( .A(n_562), .B(n_511), .Y(n_612) );
AND2x2_ASAP7_75t_L g613 ( .A(n_562), .B(n_555), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_541), .B(n_511), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_545), .Y(n_615) );
INVx2_ASAP7_75t_L g616 ( .A(n_545), .Y(n_616) );
INVx2_ASAP7_75t_L g617 ( .A(n_566), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_616), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_616), .Y(n_619) );
INVxp33_ASAP7_75t_SL g620 ( .A(n_568), .Y(n_620) );
XNOR2xp5_ASAP7_75t_L g621 ( .A(n_570), .B(n_559), .Y(n_621) );
INVxp67_ASAP7_75t_L g622 ( .A(n_593), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_598), .B(n_553), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_598), .B(n_553), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_584), .A2(n_550), .B1(n_507), .B2(n_544), .Y(n_625) );
NOR2xp33_ASAP7_75t_L g626 ( .A(n_576), .B(n_587), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_607), .B(n_552), .Y(n_627) );
AND2x2_ASAP7_75t_L g628 ( .A(n_582), .B(n_552), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_612), .Y(n_629) );
AND2x2_ASAP7_75t_L g630 ( .A(n_613), .B(n_549), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_566), .Y(n_631) );
INVx2_ASAP7_75t_L g632 ( .A(n_578), .Y(n_632) );
INVx1_ASAP7_75t_SL g633 ( .A(n_570), .Y(n_633) );
BUFx2_ASAP7_75t_L g634 ( .A(n_593), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_587), .B(n_549), .Y(n_635) );
INVx1_ASAP7_75t_SL g636 ( .A(n_590), .Y(n_636) );
INVx1_ASAP7_75t_SL g637 ( .A(n_590), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_565), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_567), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_574), .Y(n_640) );
NAND2xp5_ASAP7_75t_SL g641 ( .A(n_597), .B(n_557), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_564), .B(n_512), .Y(n_642) );
OAI21xp5_ASAP7_75t_L g643 ( .A1(n_597), .A2(n_532), .B(n_536), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_571), .B(n_512), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_579), .Y(n_645) );
NAND2xp5_ASAP7_75t_SL g646 ( .A(n_600), .B(n_537), .Y(n_646) );
AND2x2_ASAP7_75t_L g647 ( .A(n_581), .B(n_507), .Y(n_647) );
NAND2xp33_ASAP7_75t_SL g648 ( .A(n_580), .B(n_537), .Y(n_648) );
AND2x2_ASAP7_75t_L g649 ( .A(n_601), .B(n_507), .Y(n_649) );
NAND3xp33_ASAP7_75t_L g650 ( .A(n_585), .B(n_529), .C(n_525), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_583), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_586), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_573), .B(n_507), .Y(n_653) );
INVx1_ASAP7_75t_SL g654 ( .A(n_572), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_575), .B(n_533), .Y(n_655) );
OAI31xp33_ASAP7_75t_L g656 ( .A1(n_620), .A2(n_596), .A3(n_608), .B(n_563), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_623), .Y(n_657) );
NOR2x1_ASAP7_75t_L g658 ( .A(n_641), .B(n_609), .Y(n_658) );
XNOR2x1_ASAP7_75t_SL g659 ( .A(n_621), .B(n_594), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_624), .Y(n_660) );
AOI21xp5_ASAP7_75t_L g661 ( .A1(n_621), .A2(n_569), .B(n_591), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_638), .Y(n_662) );
AND2x2_ASAP7_75t_L g663 ( .A(n_636), .B(n_577), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_638), .Y(n_664) );
OAI22xp33_ASAP7_75t_L g665 ( .A1(n_633), .A2(n_611), .B1(n_589), .B2(n_608), .Y(n_665) );
AOI211xp5_ASAP7_75t_L g666 ( .A1(n_626), .A2(n_599), .B(n_605), .C(n_602), .Y(n_666) );
INVxp67_ASAP7_75t_L g667 ( .A(n_634), .Y(n_667) );
NOR2x1_ASAP7_75t_L g668 ( .A(n_634), .B(n_605), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_639), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_639), .Y(n_670) );
AND2x2_ASAP7_75t_L g671 ( .A(n_636), .B(n_604), .Y(n_671) );
AOI321xp33_ASAP7_75t_L g672 ( .A1(n_625), .A2(n_599), .A3(n_588), .B1(n_603), .B2(n_595), .C(n_592), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_640), .Y(n_673) );
XOR2x2_ASAP7_75t_L g674 ( .A(n_646), .B(n_614), .Y(n_674) );
XNOR2x2_ASAP7_75t_L g675 ( .A(n_650), .B(n_610), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_640), .Y(n_676) );
NAND3xp33_ASAP7_75t_L g677 ( .A(n_650), .B(n_615), .C(n_606), .Y(n_677) );
XNOR2x2_ASAP7_75t_L g678 ( .A(n_643), .B(n_533), .Y(n_678) );
XOR2xp5_ASAP7_75t_L g679 ( .A(n_642), .B(n_510), .Y(n_679) );
AOI322xp5_ASAP7_75t_L g680 ( .A1(n_658), .A2(n_648), .A3(n_637), .B1(n_654), .B2(n_627), .C1(n_635), .C2(n_630), .Y(n_680) );
NOR4xp75_ASAP7_75t_L g681 ( .A(n_659), .B(n_653), .C(n_644), .D(n_655), .Y(n_681) );
OAI222xp33_ASAP7_75t_L g682 ( .A1(n_661), .A2(n_665), .B1(n_668), .B2(n_637), .C1(n_667), .C2(n_678), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_662), .Y(n_683) );
AOI22xp5_ASAP7_75t_L g684 ( .A1(n_674), .A2(n_649), .B1(n_629), .B2(n_622), .Y(n_684) );
NAND3xp33_ASAP7_75t_L g685 ( .A(n_656), .B(n_652), .C(n_651), .Y(n_685) );
INVxp67_ASAP7_75t_SL g686 ( .A(n_667), .Y(n_686) );
AOI221x1_ASAP7_75t_L g687 ( .A1(n_677), .A2(n_652), .B1(n_651), .B2(n_645), .C(n_629), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_657), .B(n_627), .Y(n_688) );
AOI21xp5_ASAP7_75t_L g689 ( .A1(n_674), .A2(n_649), .B(n_632), .Y(n_689) );
AOI22xp5_ASAP7_75t_L g690 ( .A1(n_665), .A2(n_647), .B1(n_628), .B2(n_630), .Y(n_690) );
INVx1_ASAP7_75t_SL g691 ( .A(n_679), .Y(n_691) );
AOI21xp33_ASAP7_75t_SL g692 ( .A1(n_659), .A2(n_645), .B(n_631), .Y(n_692) );
A2O1A1Ixp33_ASAP7_75t_L g693 ( .A1(n_672), .A2(n_628), .B(n_647), .C(n_632), .Y(n_693) );
AOI21xp5_ASAP7_75t_L g694 ( .A1(n_666), .A2(n_631), .B(n_617), .Y(n_694) );
OAI221xp5_ASAP7_75t_L g695 ( .A1(n_660), .A2(n_619), .B1(n_618), .B2(n_617), .C(n_546), .Y(n_695) );
AOI32xp33_ASAP7_75t_L g696 ( .A1(n_678), .A2(n_547), .A3(n_519), .B1(n_520), .B2(n_523), .Y(n_696) );
OAI221xp5_ASAP7_75t_L g697 ( .A1(n_664), .A2(n_619), .B1(n_618), .B2(n_515), .C(n_556), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_669), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_670), .Y(n_699) );
NAND4xp75_ASAP7_75t_L g700 ( .A(n_675), .B(n_671), .C(n_663), .D(n_523), .Y(n_700) );
AOI22xp5_ASAP7_75t_L g701 ( .A1(n_673), .A2(n_519), .B1(n_520), .B2(n_525), .Y(n_701) );
AOI211xp5_ASAP7_75t_SL g702 ( .A1(n_675), .A2(n_532), .B(n_536), .C(n_547), .Y(n_702) );
AOI221xp5_ASAP7_75t_L g703 ( .A1(n_676), .A2(n_548), .B1(n_560), .B2(n_606), .C(n_626), .Y(n_703) );
OAI211xp5_ASAP7_75t_SL g704 ( .A1(n_680), .A2(n_690), .B(n_691), .C(n_684), .Y(n_704) );
BUFx2_ASAP7_75t_L g705 ( .A(n_686), .Y(n_705) );
CKINVDCx5p33_ASAP7_75t_R g706 ( .A(n_689), .Y(n_706) );
INVx2_ASAP7_75t_L g707 ( .A(n_683), .Y(n_707) );
CKINVDCx5p33_ASAP7_75t_R g708 ( .A(n_685), .Y(n_708) );
NOR4xp25_ASAP7_75t_L g709 ( .A(n_704), .B(n_682), .C(n_693), .D(n_699), .Y(n_709) );
OAI322xp33_ASAP7_75t_L g710 ( .A1(n_708), .A2(n_692), .A3(n_694), .B1(n_682), .B2(n_695), .C1(n_698), .C2(n_688), .Y(n_710) );
OAI322xp33_ASAP7_75t_L g711 ( .A1(n_706), .A2(n_697), .A3(n_700), .B1(n_681), .B2(n_687), .C1(n_701), .C2(n_702), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_710), .Y(n_712) );
INVx2_ASAP7_75t_L g713 ( .A(n_709), .Y(n_713) );
AOI22xp5_ASAP7_75t_L g714 ( .A1(n_712), .A2(n_705), .B1(n_700), .B2(n_707), .Y(n_714) );
INVx1_ASAP7_75t_L g715 ( .A(n_713), .Y(n_715) );
AOI322xp5_ASAP7_75t_L g716 ( .A1(n_715), .A2(n_713), .A3(n_707), .B1(n_711), .B2(n_703), .C1(n_696), .C2(n_548), .Y(n_716) );
AOI21xp5_ASAP7_75t_L g717 ( .A1(n_716), .A2(n_714), .B(n_606), .Y(n_717) );
endmodule