module fake_jpeg_12879_n_71 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_71);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_71;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_55;
wire n_27;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_65;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_11;
wire n_62;
wire n_25;
wire n_31;
wire n_17;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

BUFx10_ASAP7_75t_L g10 ( 
.A(n_7),
.Y(n_10)
);

INVx13_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

INVx3_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

OR2x2_ASAP7_75t_L g13 ( 
.A(n_8),
.B(n_9),
.Y(n_13)
);

BUFx10_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

OR2x2_ASAP7_75t_L g21 ( 
.A(n_18),
.B(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

INVx2_ASAP7_75t_SL g23 ( 
.A(n_19),
.Y(n_23)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

AOI21xp33_ASAP7_75t_SL g24 ( 
.A1(n_10),
.A2(n_0),
.B(n_2),
.Y(n_24)
);

OR2x2_ASAP7_75t_L g38 ( 
.A(n_24),
.B(n_14),
.Y(n_38)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_12),
.B(n_13),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_13),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_23),
.A2(n_12),
.B1(n_14),
.B2(n_10),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_30),
.A2(n_37),
.B(n_38),
.Y(n_48)
);

NOR2xp67_ASAP7_75t_R g47 ( 
.A(n_33),
.B(n_38),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_20),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_21),
.B(n_20),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_23),
.A2(n_14),
.B1(n_16),
.B2(n_15),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_34),
.A2(n_22),
.B1(n_28),
.B2(n_26),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_40),
.A2(n_46),
.B(n_32),
.Y(n_51)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_45),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_39),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_36),
.A2(n_25),
.B1(n_14),
.B2(n_17),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_47),
.B(n_33),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_11),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_51),
.A2(n_48),
.B1(n_40),
.B2(n_42),
.Y(n_54)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_53),
.B(n_43),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_57),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_35),
.C(n_27),
.Y(n_56)
);

XOR2xp5_ASAP7_75t_L g60 ( 
.A(n_56),
.B(n_58),
.Y(n_60)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_27),
.C(n_11),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_59),
.Y(n_61)
);

OA21x2_ASAP7_75t_L g64 ( 
.A1(n_62),
.A2(n_50),
.B(n_52),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_64),
.A2(n_65),
.B(n_61),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_63),
.B(n_2),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_66),
.B(n_67),
.Y(n_68)
);

MAJx2_ASAP7_75t_L g67 ( 
.A(n_64),
.B(n_60),
.C(n_4),
.Y(n_67)
);

NAND4xp25_ASAP7_75t_L g69 ( 
.A(n_68),
.B(n_0),
.C(n_9),
.D(n_66),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_69),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g71 ( 
.A(n_70),
.Y(n_71)
);


endmodule