module fake_ibex_1094_n_1324 (n_151, n_147, n_85, n_167, n_128, n_208, n_234, n_84, n_64, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_205, n_204, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_237, n_29, n_143, n_106, n_177, n_203, n_148, n_2, n_76, n_233, n_8, n_118, n_224, n_183, n_67, n_229, n_9, n_209, n_164, n_38, n_198, n_124, n_37, n_110, n_193, n_47, n_169, n_108, n_217, n_10, n_82, n_21, n_27, n_165, n_242, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_191, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_180, n_194, n_122, n_223, n_116, n_240, n_61, n_201, n_14, n_0, n_239, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_226, n_46, n_80, n_172, n_215, n_49, n_40, n_66, n_17, n_74, n_90, n_235, n_176, n_58, n_192, n_43, n_140, n_216, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_206, n_221, n_166, n_195, n_163, n_212, n_26, n_188, n_200, n_114, n_199, n_236, n_34, n_97, n_102, n_197, n_181, n_15, n_131, n_123, n_24, n_52, n_189, n_99, n_135, n_105, n_156, n_126, n_187, n_1, n_154, n_182, n_111, n_196, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_222, n_107, n_115, n_149, n_186, n_227, n_50, n_11, n_92, n_144, n_170, n_213, n_101, n_190, n_113, n_138, n_230, n_96, n_185, n_241, n_68, n_117, n_214, n_238, n_79, n_81, n_35, n_159, n_202, n_231, n_158, n_211, n_218, n_132, n_174, n_210, n_157, n_219, n_160, n_220, n_225, n_184, n_31, n_56, n_23, n_146, n_232, n_91, n_207, n_54, n_19, n_228, n_1324);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_208;
input n_234;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_205;
input n_204;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_237;
input n_29;
input n_143;
input n_106;
input n_177;
input n_203;
input n_148;
input n_2;
input n_76;
input n_233;
input n_8;
input n_118;
input n_224;
input n_183;
input n_67;
input n_229;
input n_9;
input n_209;
input n_164;
input n_38;
input n_198;
input n_124;
input n_37;
input n_110;
input n_193;
input n_47;
input n_169;
input n_108;
input n_217;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_242;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_191;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_180;
input n_194;
input n_122;
input n_223;
input n_116;
input n_240;
input n_61;
input n_201;
input n_14;
input n_0;
input n_239;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_226;
input n_46;
input n_80;
input n_172;
input n_215;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_235;
input n_176;
input n_58;
input n_192;
input n_43;
input n_140;
input n_216;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_206;
input n_221;
input n_166;
input n_195;
input n_163;
input n_212;
input n_26;
input n_188;
input n_200;
input n_114;
input n_199;
input n_236;
input n_34;
input n_97;
input n_102;
input n_197;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_189;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_187;
input n_1;
input n_154;
input n_182;
input n_111;
input n_196;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_222;
input n_107;
input n_115;
input n_149;
input n_186;
input n_227;
input n_50;
input n_11;
input n_92;
input n_144;
input n_170;
input n_213;
input n_101;
input n_190;
input n_113;
input n_138;
input n_230;
input n_96;
input n_185;
input n_241;
input n_68;
input n_117;
input n_214;
input n_238;
input n_79;
input n_81;
input n_35;
input n_159;
input n_202;
input n_231;
input n_158;
input n_211;
input n_218;
input n_132;
input n_174;
input n_210;
input n_157;
input n_219;
input n_160;
input n_220;
input n_225;
input n_184;
input n_31;
input n_56;
input n_23;
input n_146;
input n_232;
input n_91;
input n_207;
input n_54;
input n_19;
input n_228;

output n_1324;

wire n_1084;
wire n_1295;
wire n_507;
wire n_992;
wire n_766;
wire n_1110;
wire n_273;
wire n_309;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_446;
wire n_452;
wire n_1234;
wire n_773;
wire n_821;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_957;
wire n_678;
wire n_969;
wire n_1125;
wire n_733;
wire n_312;
wire n_622;
wire n_1226;
wire n_1034;
wire n_872;
wire n_457;
wire n_494;
wire n_930;
wire n_1044;
wire n_1134;
wire n_911;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_1233;
wire n_1045;
wire n_500;
wire n_963;
wire n_376;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_280;
wire n_375;
wire n_667;
wire n_884;
wire n_850;
wire n_879;
wire n_723;
wire n_1144;
wire n_346;
wire n_1268;
wire n_739;
wire n_853;
wire n_504;
wire n_948;
wire n_875;
wire n_1307;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_671;
wire n_989;
wire n_829;
wire n_825;
wire n_939;
wire n_655;
wire n_306;
wire n_550;
wire n_641;
wire n_557;
wire n_527;
wire n_893;
wire n_496;
wire n_434;
wire n_1258;
wire n_835;
wire n_1195;
wire n_824;
wire n_441;
wire n_694;
wire n_523;
wire n_787;
wire n_614;
wire n_431;
wire n_1130;
wire n_1228;
wire n_321;
wire n_1081;
wire n_279;
wire n_374;
wire n_538;
wire n_1155;
wire n_1292;
wire n_459;
wire n_518;
wire n_852;
wire n_1133;
wire n_904;
wire n_355;
wire n_448;
wire n_646;
wire n_466;
wire n_1030;
wire n_1094;
wire n_715;
wire n_530;
wire n_1214;
wire n_1274;
wire n_420;
wire n_769;
wire n_857;
wire n_765;
wire n_1070;
wire n_777;
wire n_331;
wire n_917;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1313;
wire n_352;
wire n_558;
wire n_666;
wire n_1071;
wire n_793;
wire n_937;
wire n_973;
wire n_1038;
wire n_618;
wire n_1269;
wire n_662;
wire n_979;
wire n_1309;
wire n_1316;
wire n_1215;
wire n_629;
wire n_573;
wire n_359;
wire n_262;
wire n_433;
wire n_439;
wire n_1007;
wire n_643;
wire n_1276;
wire n_841;
wire n_772;
wire n_810;
wire n_338;
wire n_369;
wire n_1301;
wire n_257;
wire n_869;
wire n_718;
wire n_554;
wire n_553;
wire n_1078;
wire n_1219;
wire n_713;
wire n_307;
wire n_1252;
wire n_1170;
wire n_605;
wire n_539;
wire n_630;
wire n_567;
wire n_745;
wire n_447;
wire n_562;
wire n_564;
wire n_1322;
wire n_1305;
wire n_795;
wire n_592;
wire n_1248;
wire n_762;
wire n_308;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_397;
wire n_894;
wire n_1118;
wire n_692;
wire n_709;
wire n_1296;
wire n_499;
wire n_702;
wire n_971;
wire n_451;
wire n_906;
wire n_1093;
wire n_978;
wire n_579;
wire n_899;
wire n_1019;
wire n_902;
wire n_1250;
wire n_1190;
wire n_1304;
wire n_744;
wire n_314;
wire n_563;
wire n_881;
wire n_734;
wire n_1073;
wire n_1108;
wire n_382;
wire n_1239;
wire n_1209;
wire n_288;
wire n_379;
wire n_551;
wire n_729;
wire n_603;
wire n_422;
wire n_324;
wire n_391;
wire n_820;
wire n_805;
wire n_670;
wire n_1132;
wire n_892;
wire n_390;
wire n_544;
wire n_1281;
wire n_695;
wire n_639;
wire n_482;
wire n_282;
wire n_870;
wire n_1298;
wire n_609;
wire n_1040;
wire n_476;
wire n_1159;
wire n_1154;
wire n_345;
wire n_455;
wire n_1243;
wire n_1121;
wire n_693;
wire n_406;
wire n_606;
wire n_737;
wire n_462;
wire n_1235;
wire n_1003;
wire n_889;
wire n_435;
wire n_396;
wire n_252;
wire n_816;
wire n_1058;
wire n_399;
wire n_823;
wire n_657;
wire n_1156;
wire n_1293;
wire n_749;
wire n_819;
wire n_822;
wire n_1042;
wire n_743;
wire n_754;
wire n_395;
wire n_1319;
wire n_389;
wire n_1041;
wire n_1090;
wire n_1196;
wire n_330;
wire n_1182;
wire n_1271;
wire n_1031;
wire n_372;
wire n_256;
wire n_981;
wire n_350;
wire n_398;
wire n_583;
wire n_1015;
wire n_663;
wire n_1152;
wire n_371;
wire n_974;
wire n_1036;
wire n_608;
wire n_864;
wire n_412;
wire n_959;
wire n_1106;
wire n_258;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_449;
wire n_1318;
wire n_421;
wire n_738;
wire n_1217;
wire n_1189;
wire n_761;
wire n_748;
wire n_901;
wire n_340;
wire n_1255;
wire n_1218;
wire n_1181;
wire n_1140;
wire n_1056;
wire n_1283;
wire n_840;
wire n_1203;
wire n_561;
wire n_471;
wire n_846;
wire n_1237;
wire n_859;
wire n_965;
wire n_1109;
wire n_384;
wire n_1051;
wire n_1008;
wire n_458;
wire n_1053;
wire n_1207;
wire n_310;
wire n_1076;
wire n_1032;
wire n_936;
wire n_469;
wire n_1210;
wire n_591;
wire n_1201;
wire n_1246;
wire n_732;
wire n_1236;
wire n_832;
wire n_316;
wire n_590;
wire n_325;
wire n_1184;
wire n_1013;
wire n_929;
wire n_315;
wire n_637;
wire n_1136;
wire n_1075;
wire n_1249;
wire n_574;
wire n_515;
wire n_1229;
wire n_907;
wire n_1179;
wire n_1153;
wire n_669;
wire n_521;
wire n_1117;
wire n_1273;
wire n_1083;
wire n_1014;
wire n_724;
wire n_437;
wire n_938;
wire n_1178;
wire n_474;
wire n_878;
wire n_594;
wire n_944;
wire n_623;
wire n_585;
wire n_483;
wire n_1137;
wire n_660;
wire n_524;
wire n_1200;
wire n_295;
wire n_1120;
wire n_576;
wire n_388;
wire n_1279;
wire n_290;
wire n_931;
wire n_607;
wire n_827;
wire n_1064;
wire n_1028;
wire n_1264;
wire n_1146;
wire n_358;
wire n_488;
wire n_705;
wire n_429;
wire n_267;
wire n_1009;
wire n_1260;
wire n_589;
wire n_472;
wire n_347;
wire n_847;
wire n_413;
wire n_1069;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_679;
wire n_696;
wire n_837;
wire n_640;
wire n_954;
wire n_363;
wire n_725;
wire n_596;
wire n_351;
wire n_456;
wire n_998;
wire n_1115;
wire n_801;
wire n_1046;
wire n_882;
wire n_942;
wire n_651;
wire n_721;
wire n_365;
wire n_814;
wire n_943;
wire n_1086;
wire n_444;
wire n_986;
wire n_495;
wire n_411;
wire n_927;
wire n_615;
wire n_803;
wire n_1087;
wire n_757;
wire n_712;
wire n_650;
wire n_409;
wire n_332;
wire n_517;
wire n_817;
wire n_555;
wire n_337;
wire n_951;
wire n_272;
wire n_468;
wire n_780;
wire n_502;
wire n_633;
wire n_532;
wire n_726;
wire n_863;
wire n_597;
wire n_285;
wire n_1128;
wire n_1266;
wire n_1300;
wire n_291;
wire n_318;
wire n_268;
wire n_807;
wire n_741;
wire n_430;
wire n_486;
wire n_997;
wire n_891;
wire n_303;
wire n_717;
wire n_668;
wire n_871;
wire n_266;
wire n_485;
wire n_1315;
wire n_811;
wire n_808;
wire n_250;
wire n_945;
wire n_460;
wire n_461;
wire n_903;
wire n_1095;
wire n_1265;
wire n_1048;
wire n_774;
wire n_588;
wire n_1251;
wire n_1247;
wire n_528;
wire n_260;
wire n_836;
wire n_1263;
wire n_443;
wire n_1185;
wire n_344;
wire n_436;
wire n_1122;
wire n_628;
wire n_890;
wire n_874;
wire n_1163;
wire n_677;
wire n_964;
wire n_916;
wire n_503;
wire n_292;
wire n_895;
wire n_687;
wire n_1035;
wire n_751;
wire n_1127;
wire n_932;
wire n_380;
wire n_281;
wire n_1004;
wire n_947;
wire n_831;
wire n_778;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1104;
wire n_1011;
wire n_529;
wire n_626;
wire n_1143;
wire n_328;
wire n_418;
wire n_510;
wire n_972;
wire n_601;
wire n_610;
wire n_920;
wire n_664;
wire n_1067;
wire n_255;
wire n_994;
wire n_545;
wire n_887;
wire n_1162;
wire n_334;
wire n_634;
wire n_991;
wire n_961;
wire n_1223;
wire n_1323;
wire n_578;
wire n_432;
wire n_403;
wire n_423;
wire n_357;
wire n_1320;
wire n_996;
wire n_915;
wire n_1174;
wire n_1286;
wire n_542;
wire n_1294;
wire n_900;
wire n_377;
wire n_647;
wire n_1291;
wire n_317;
wire n_326;
wire n_270;
wire n_259;
wire n_339;
wire n_276;
wire n_348;
wire n_674;
wire n_287;
wire n_552;
wire n_251;
wire n_1112;
wire n_1267;
wire n_703;
wire n_426;
wire n_1172;
wire n_1099;
wire n_598;
wire n_508;
wire n_453;
wire n_400;
wire n_1055;
wire n_673;
wire n_798;
wire n_278;
wire n_404;
wire n_1177;
wire n_1025;
wire n_296;
wire n_690;
wire n_1225;
wire n_982;
wire n_785;
wire n_604;
wire n_977;
wire n_719;
wire n_370;
wire n_289;
wire n_716;
wire n_923;
wire n_642;
wire n_286;
wire n_933;
wire n_1037;
wire n_464;
wire n_1289;
wire n_838;
wire n_1021;
wire n_746;
wire n_1188;
wire n_261;
wire n_742;
wire n_1191;
wire n_1052;
wire n_789;
wire n_656;
wire n_602;
wire n_842;
wire n_767;
wire n_636;
wire n_1259;
wire n_490;
wire n_407;
wire n_595;
wire n_1001;
wire n_269;
wire n_570;
wire n_1224;
wire n_356;
wire n_487;
wire n_349;
wire n_454;
wire n_1017;
wire n_730;
wire n_625;
wire n_619;
wire n_1124;
wire n_611;
wire n_246;
wire n_922;
wire n_851;
wire n_993;
wire n_253;
wire n_300;
wire n_1135;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_1066;
wire n_1169;
wire n_245;
wire n_648;
wire n_571;
wire n_830;
wire n_473;
wire n_1241;
wire n_445;
wire n_1072;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_353;
wire n_826;
wire n_768;
wire n_839;
wire n_1278;
wire n_796;
wire n_797;
wire n_1006;
wire n_402;
wire n_1238;
wire n_976;
wire n_1063;
wire n_1270;
wire n_834;
wire n_935;
wire n_925;
wire n_1054;
wire n_722;
wire n_804;
wire n_484;
wire n_480;
wire n_354;
wire n_1057;
wire n_516;
wire n_329;
wire n_1149;
wire n_1176;
wire n_506;
wire n_868;
wire n_1202;
wire n_1065;
wire n_905;
wire n_975;
wire n_675;
wire n_463;
wire n_624;
wire n_520;
wire n_934;
wire n_775;
wire n_512;
wire n_950;
wire n_685;
wire n_1222;
wire n_1198;
wire n_1311;
wire n_1261;
wire n_248;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_1282;
wire n_277;
wire n_1321;
wire n_700;
wire n_360;
wire n_1107;
wire n_525;
wire n_815;
wire n_919;
wire n_535;
wire n_681;
wire n_415;
wire n_320;
wire n_247;
wire n_1139;
wire n_1018;
wire n_858;
wire n_385;
wire n_782;
wire n_616;
wire n_833;
wire n_728;
wire n_786;
wire n_362;
wire n_505;
wire n_501;
wire n_752;
wire n_958;
wire n_1175;
wire n_1221;
wire n_284;
wire n_1047;
wire n_792;
wire n_1314;
wire n_575;
wire n_313;
wire n_1242;
wire n_1119;
wire n_1085;
wire n_419;
wire n_885;
wire n_513;
wire n_877;
wire n_311;
wire n_1088;
wire n_896;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_1288;
wire n_302;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_393;
wire n_428;
wire n_697;
wire n_1105;
wire n_912;
wire n_424;
wire n_701;
wire n_995;
wire n_1000;
wire n_298;
wire n_1256;
wire n_587;
wire n_1303;
wire n_764;
wire n_1206;
wire n_855;
wire n_812;
wire n_1050;
wire n_599;
wire n_1060;
wire n_756;
wire n_1257;
wire n_274;
wire n_387;
wire n_688;
wire n_946;
wire n_707;
wire n_1097;
wire n_293;
wire n_341;
wire n_621;
wire n_956;
wire n_790;
wire n_586;
wire n_638;
wire n_304;
wire n_593;
wire n_1212;
wire n_1199;
wire n_249;
wire n_478;
wire n_336;
wire n_861;
wire n_1131;
wire n_547;
wire n_727;
wire n_1077;
wire n_828;
wire n_753;
wire n_645;
wire n_747;
wire n_1147;
wire n_1098;
wire n_584;
wire n_1187;
wire n_698;
wire n_1061;
wire n_682;
wire n_327;
wire n_1302;
wire n_383;
wire n_886;
wire n_1010;
wire n_883;
wire n_417;
wire n_755;
wire n_265;
wire n_1029;
wire n_470;
wire n_770;
wire n_941;
wire n_1245;
wire n_1317;
wire n_243;
wire n_632;
wire n_373;
wire n_854;
wire n_244;
wire n_343;
wire n_714;
wire n_1297;
wire n_323;
wire n_740;
wire n_386;
wire n_549;
wire n_533;
wire n_898;
wire n_928;
wire n_333;
wire n_1285;
wire n_967;
wire n_736;
wire n_1103;
wire n_1161;
wire n_465;
wire n_1068;
wire n_617;
wire n_301;
wire n_914;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1197;
wire n_1168;
wire n_865;
wire n_569;
wire n_600;
wire n_1192;
wire n_1290;
wire n_987;
wire n_750;
wire n_1299;
wire n_665;
wire n_1101;
wire n_367;
wire n_880;
wire n_654;
wire n_731;
wire n_1166;
wire n_758;
wire n_720;
wire n_710;
wire n_1023;
wire n_568;
wire n_813;
wire n_1211;
wire n_1284;
wire n_1116;
wire n_791;
wire n_543;
wire n_580;
wire n_1082;
wire n_1213;
wire n_980;
wire n_1193;
wire n_849;
wire n_1074;
wire n_759;
wire n_953;
wire n_1180;
wire n_536;
wire n_1220;
wire n_467;
wire n_427;
wire n_1262;
wire n_442;
wire n_438;
wire n_1012;
wire n_689;
wire n_960;
wire n_1022;
wire n_676;
wire n_1240;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_560;
wire n_910;
wire n_635;
wire n_844;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_335;
wire n_263;
wire n_966;
wire n_299;
wire n_949;
wire n_704;
wire n_924;
wire n_477;
wire n_699;
wire n_368;
wire n_918;
wire n_672;
wire n_1039;
wire n_401;
wire n_1043;
wire n_735;
wire n_305;
wire n_566;
wire n_416;
wire n_581;
wire n_1089;
wire n_392;
wire n_1049;
wire n_548;
wire n_1158;
wire n_763;
wire n_940;
wire n_546;
wire n_788;
wire n_410;
wire n_1160;
wire n_658;
wire n_1216;
wire n_1026;
wire n_283;
wire n_366;
wire n_1033;
wire n_627;
wire n_990;
wire n_322;
wire n_888;
wire n_582;
wire n_653;
wire n_1205;
wire n_843;
wire n_1059;
wire n_799;
wire n_691;
wire n_522;
wire n_479;
wire n_534;
wire n_511;
wire n_381;
wire n_1002;
wire n_1111;
wire n_405;
wire n_1310;
wire n_612;
wire n_955;
wire n_440;
wire n_342;
wire n_414;
wire n_378;
wire n_952;
wire n_264;
wire n_1145;
wire n_537;
wire n_1113;
wire n_913;
wire n_509;
wire n_1164;
wire n_1277;
wire n_1016;
wire n_680;
wire n_809;
wire n_856;
wire n_779;
wire n_294;
wire n_1280;
wire n_493;
wire n_519;
wire n_408;
wire n_361;
wire n_319;
wire n_1091;
wire n_1287;
wire n_860;
wire n_661;
wire n_848;
wire n_683;
wire n_1194;
wire n_1150;
wire n_620;
wire n_450;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_644;
wire n_577;
wire n_970;
wire n_491;
wire n_297;
wire n_921;
wire n_489;
wire n_254;
wire n_908;
wire n_565;
wire n_1123;
wire n_1272;
wire n_271;
wire n_984;
wire n_394;
wire n_364;
wire n_988;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_492;
wire n_649;
wire n_866;
wire n_559;
wire n_425;

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_195),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_20),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_175),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_227),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_129),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_228),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_169),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_104),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_186),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_209),
.Y(n_252)
);

INVxp33_ASAP7_75t_L g253 ( 
.A(n_98),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_217),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_118),
.Y(n_255)
);

INVx2_ASAP7_75t_SL g256 ( 
.A(n_192),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_164),
.Y(n_257)
);

BUFx2_ASAP7_75t_SL g258 ( 
.A(n_137),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_190),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_160),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_238),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_22),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_20),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_106),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_1),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_149),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_145),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_135),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_35),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_64),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_24),
.Y(n_271)
);

CKINVDCx14_ASAP7_75t_R g272 ( 
.A(n_232),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_142),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_47),
.Y(n_274)
);

BUFx10_ASAP7_75t_L g275 ( 
.A(n_117),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_50),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_147),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_220),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_97),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_28),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_139),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_184),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_221),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_34),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g285 ( 
.A(n_125),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_185),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_140),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_230),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_154),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_65),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_7),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_90),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_21),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_87),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_61),
.Y(n_295)
);

BUFx5_ASAP7_75t_L g296 ( 
.A(n_201),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_119),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_91),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_116),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_151),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_59),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_210),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_8),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_191),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_22),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_65),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_92),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_178),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_193),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_166),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_133),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_208),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_136),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_156),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_152),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_4),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_225),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_219),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_93),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_237),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_159),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_206),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_37),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_115),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_42),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_30),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_163),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_229),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_126),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_233),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_122),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_242),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_43),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_181),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_82),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_197),
.Y(n_336)
);

INVx2_ASAP7_75t_SL g337 ( 
.A(n_25),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_189),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_27),
.Y(n_339)
);

INVxp67_ASAP7_75t_SL g340 ( 
.A(n_53),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_194),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_188),
.Y(n_342)
);

NOR2xp67_ASAP7_75t_L g343 ( 
.A(n_153),
.B(n_72),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_110),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_67),
.Y(n_345)
);

HB1xp67_ASAP7_75t_L g346 ( 
.A(n_114),
.Y(n_346)
);

INVxp67_ASAP7_75t_SL g347 ( 
.A(n_59),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_95),
.Y(n_348)
);

INVx1_ASAP7_75t_SL g349 ( 
.A(n_2),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_111),
.B(n_146),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_171),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_86),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_33),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_53),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_207),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_143),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_212),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_72),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_226),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_162),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_196),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_168),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_13),
.Y(n_363)
);

CKINVDCx16_ASAP7_75t_R g364 ( 
.A(n_11),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_157),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_112),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_216),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_205),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_74),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_148),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_102),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_10),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_10),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_39),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_83),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_234),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_113),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_96),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_19),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_222),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_57),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_211),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_66),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_33),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_69),
.Y(n_385)
);

CKINVDCx14_ASAP7_75t_R g386 ( 
.A(n_123),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_18),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_158),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_57),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_30),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_203),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_231),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_48),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_58),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_177),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_37),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_128),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_80),
.Y(n_398)
);

CKINVDCx14_ASAP7_75t_R g399 ( 
.A(n_69),
.Y(n_399)
);

BUFx3_ASAP7_75t_L g400 ( 
.A(n_88),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_172),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_81),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_75),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_199),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_70),
.Y(n_405)
);

INVx1_ASAP7_75t_SL g406 ( 
.A(n_180),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_170),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_99),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_121),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_52),
.Y(n_410)
);

BUFx2_ASAP7_75t_L g411 ( 
.A(n_17),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_331),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_346),
.Y(n_413)
);

BUFx8_ASAP7_75t_L g414 ( 
.A(n_411),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_354),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_251),
.Y(n_416)
);

INVx5_ASAP7_75t_L g417 ( 
.A(n_251),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_399),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_251),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_403),
.B(n_0),
.Y(n_420)
);

BUFx12f_ASAP7_75t_L g421 ( 
.A(n_275),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_337),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_244),
.Y(n_423)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_275),
.Y(n_424)
);

INVx5_ASAP7_75t_L g425 ( 
.A(n_251),
.Y(n_425)
);

BUFx12f_ASAP7_75t_L g426 ( 
.A(n_275),
.Y(n_426)
);

BUFx2_ASAP7_75t_L g427 ( 
.A(n_399),
.Y(n_427)
);

INVx6_ASAP7_75t_L g428 ( 
.A(n_296),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_327),
.Y(n_429)
);

AND2x4_ASAP7_75t_L g430 ( 
.A(n_256),
.B(n_0),
.Y(n_430)
);

OAI22x1_ASAP7_75t_R g431 ( 
.A1(n_325),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_296),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_296),
.Y(n_433)
);

AND2x6_ASAP7_75t_L g434 ( 
.A(n_400),
.B(n_84),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_296),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_253),
.B(n_3),
.Y(n_436)
);

OA21x2_ASAP7_75t_L g437 ( 
.A1(n_259),
.A2(n_89),
.B(n_85),
.Y(n_437)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_265),
.Y(n_438)
);

INVx2_ASAP7_75t_SL g439 ( 
.A(n_400),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_327),
.Y(n_440)
);

CKINVDCx6p67_ASAP7_75t_R g441 ( 
.A(n_258),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_270),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_272),
.Y(n_443)
);

BUFx8_ASAP7_75t_SL g444 ( 
.A(n_325),
.Y(n_444)
);

OAI22x1_ASAP7_75t_L g445 ( 
.A1(n_340),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_253),
.B(n_5),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g447 ( 
.A(n_364),
.B(n_6),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_271),
.Y(n_448)
);

BUFx8_ASAP7_75t_L g449 ( 
.A(n_296),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_327),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_373),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_280),
.Y(n_452)
);

INVx5_ASAP7_75t_L g453 ( 
.A(n_330),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_296),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_284),
.Y(n_455)
);

AND2x6_ASAP7_75t_L g456 ( 
.A(n_259),
.B(n_94),
.Y(n_456)
);

AND2x4_ASAP7_75t_L g457 ( 
.A(n_300),
.B(n_7),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_300),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_313),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_290),
.Y(n_460)
);

HB1xp67_ASAP7_75t_L g461 ( 
.A(n_262),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_313),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_330),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_272),
.B(n_386),
.Y(n_464)
);

INVx3_ASAP7_75t_L g465 ( 
.A(n_265),
.Y(n_465)
);

OA21x2_ASAP7_75t_L g466 ( 
.A1(n_315),
.A2(n_101),
.B(n_100),
.Y(n_466)
);

BUFx8_ASAP7_75t_L g467 ( 
.A(n_315),
.Y(n_467)
);

OA21x2_ASAP7_75t_L g468 ( 
.A1(n_332),
.A2(n_105),
.B(n_103),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_291),
.B(n_8),
.Y(n_469)
);

OAI22x1_ASAP7_75t_L g470 ( 
.A1(n_347),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_470)
);

BUFx2_ASAP7_75t_L g471 ( 
.A(n_263),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_293),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_332),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_265),
.Y(n_474)
);

AND2x4_ASAP7_75t_L g475 ( 
.A(n_344),
.B(n_9),
.Y(n_475)
);

HB1xp67_ASAP7_75t_L g476 ( 
.A(n_269),
.Y(n_476)
);

AND2x4_ASAP7_75t_L g477 ( 
.A(n_348),
.B(n_13),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_348),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_360),
.Y(n_479)
);

INVx5_ASAP7_75t_L g480 ( 
.A(n_330),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_360),
.Y(n_481)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_265),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_L g483 ( 
.A1(n_326),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_243),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_330),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_334),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_334),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_339),
.Y(n_488)
);

BUFx8_ASAP7_75t_SL g489 ( 
.A(n_384),
.Y(n_489)
);

CKINVDCx8_ASAP7_75t_R g490 ( 
.A(n_274),
.Y(n_490)
);

INVx5_ASAP7_75t_L g491 ( 
.A(n_334),
.Y(n_491)
);

OA21x2_ASAP7_75t_L g492 ( 
.A1(n_376),
.A2(n_108),
.B(n_107),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_334),
.Y(n_493)
);

INVx3_ASAP7_75t_L g494 ( 
.A(n_303),
.Y(n_494)
);

INVx5_ASAP7_75t_L g495 ( 
.A(n_336),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_376),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_243),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_497)
);

NOR2x1_ASAP7_75t_L g498 ( 
.A(n_410),
.B(n_109),
.Y(n_498)
);

BUFx6f_ASAP7_75t_L g499 ( 
.A(n_336),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_L g500 ( 
.A1(n_385),
.A2(n_21),
.B1(n_23),
.B2(n_24),
.Y(n_500)
);

INVx3_ASAP7_75t_L g501 ( 
.A(n_303),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_336),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_336),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_387),
.Y(n_504)
);

AND2x4_ASAP7_75t_L g505 ( 
.A(n_408),
.B(n_390),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_393),
.Y(n_506)
);

OAI22x1_ASAP7_75t_L g507 ( 
.A1(n_394),
.A2(n_23),
.B1(n_26),
.B2(n_27),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_384),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_246),
.A2(n_26),
.B1(n_28),
.B2(n_29),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_457),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_457),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_432),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_475),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_475),
.Y(n_514)
);

NOR2x1p5_ASAP7_75t_L g515 ( 
.A(n_421),
.B(n_402),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_424),
.B(n_283),
.Y(n_516)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_475),
.Y(n_517)
);

BUFx3_ASAP7_75t_L g518 ( 
.A(n_434),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_449),
.B(n_408),
.Y(n_519)
);

OR2x2_ASAP7_75t_L g520 ( 
.A(n_415),
.B(n_349),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_433),
.Y(n_521)
);

BUFx10_ASAP7_75t_L g522 ( 
.A(n_443),
.Y(n_522)
);

INVx2_ASAP7_75t_SL g523 ( 
.A(n_427),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_424),
.B(n_397),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_435),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_427),
.B(n_386),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_464),
.B(n_295),
.Y(n_527)
);

INVxp33_ASAP7_75t_SL g528 ( 
.A(n_418),
.Y(n_528)
);

INVx3_ASAP7_75t_L g529 ( 
.A(n_477),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_435),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_477),
.Y(n_531)
);

OAI22xp33_ASAP7_75t_L g532 ( 
.A1(n_484),
.A2(n_389),
.B1(n_345),
.B2(n_276),
.Y(n_532)
);

INVx4_ASAP7_75t_L g533 ( 
.A(n_434),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_454),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_449),
.B(n_430),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_508),
.Y(n_536)
);

BUFx10_ASAP7_75t_L g537 ( 
.A(n_443),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_422),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_430),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g540 ( 
.A(n_416),
.Y(n_540)
);

INVx3_ASAP7_75t_L g541 ( 
.A(n_430),
.Y(n_541)
);

AND3x2_ASAP7_75t_L g542 ( 
.A(n_447),
.B(n_247),
.C(n_245),
.Y(n_542)
);

INVx2_ASAP7_75t_SL g543 ( 
.A(n_449),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_464),
.B(n_301),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_505),
.B(n_249),
.Y(n_545)
);

BUFx3_ASAP7_75t_L g546 ( 
.A(n_434),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_412),
.B(n_413),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_436),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_471),
.B(n_305),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_419),
.Y(n_550)
);

INVx4_ASAP7_75t_L g551 ( 
.A(n_434),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_436),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_505),
.B(n_250),
.Y(n_553)
);

INVx2_ASAP7_75t_SL g554 ( 
.A(n_467),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_446),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_471),
.B(n_254),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_419),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_451),
.B(n_306),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_419),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g560 ( 
.A(n_419),
.Y(n_560)
);

INVx2_ASAP7_75t_SL g561 ( 
.A(n_428),
.Y(n_561)
);

INVxp67_ASAP7_75t_SL g562 ( 
.A(n_467),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_423),
.B(n_255),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_429),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_429),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_442),
.B(n_257),
.Y(n_566)
);

NAND2xp33_ASAP7_75t_L g567 ( 
.A(n_456),
.B(n_357),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_429),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_458),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_429),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_458),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_440),
.Y(n_572)
);

AND2x2_ASAP7_75t_SL g573 ( 
.A(n_437),
.B(n_303),
.Y(n_573)
);

NAND2xp33_ASAP7_75t_L g574 ( 
.A(n_456),
.B(n_357),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_459),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_461),
.B(n_316),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_439),
.B(n_323),
.Y(n_577)
);

NAND2xp33_ASAP7_75t_L g578 ( 
.A(n_456),
.B(n_357),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_440),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_440),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_448),
.B(n_260),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_476),
.B(n_333),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_459),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_462),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_462),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_473),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_450),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_450),
.Y(n_588)
);

BUFx6f_ASAP7_75t_L g589 ( 
.A(n_450),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_463),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_463),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_473),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_478),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_463),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_479),
.Y(n_595)
);

INVx2_ASAP7_75t_SL g596 ( 
.A(n_428),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_479),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_481),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_485),
.Y(n_599)
);

INVx2_ASAP7_75t_SL g600 ( 
.A(n_467),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_481),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_496),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_485),
.Y(n_603)
);

CKINVDCx6p67_ASAP7_75t_R g604 ( 
.A(n_421),
.Y(n_604)
);

OR2x2_ASAP7_75t_L g605 ( 
.A(n_452),
.B(n_353),
.Y(n_605)
);

INVxp33_ASAP7_75t_SL g606 ( 
.A(n_447),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_455),
.B(n_277),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_460),
.B(n_358),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_485),
.Y(n_609)
);

INVx8_ASAP7_75t_L g610 ( 
.A(n_426),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_472),
.B(n_363),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_498),
.B(n_279),
.Y(n_612)
);

CKINVDCx6p67_ASAP7_75t_R g613 ( 
.A(n_426),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_486),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_414),
.Y(n_615)
);

OR2x6_ASAP7_75t_L g616 ( 
.A(n_445),
.B(n_470),
.Y(n_616)
);

BUFx6f_ASAP7_75t_SL g617 ( 
.A(n_456),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_487),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_490),
.B(n_369),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_487),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_488),
.B(n_372),
.Y(n_621)
);

INVx3_ASAP7_75t_L g622 ( 
.A(n_428),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_504),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_487),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_506),
.Y(n_625)
);

AO21x2_ASAP7_75t_L g626 ( 
.A1(n_469),
.A2(n_350),
.B(n_294),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_417),
.B(n_288),
.Y(n_627)
);

AOI22xp33_ASAP7_75t_L g628 ( 
.A1(n_420),
.A2(n_396),
.B1(n_405),
.B2(n_303),
.Y(n_628)
);

NAND3xp33_ASAP7_75t_L g629 ( 
.A(n_490),
.B(n_379),
.C(n_374),
.Y(n_629)
);

NAND3xp33_ASAP7_75t_L g630 ( 
.A(n_437),
.B(n_468),
.C(n_466),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_441),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_441),
.B(n_381),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_438),
.Y(n_633)
);

NAND3xp33_ASAP7_75t_L g634 ( 
.A(n_437),
.B(n_398),
.C(n_383),
.Y(n_634)
);

INVx2_ASAP7_75t_SL g635 ( 
.A(n_414),
.Y(n_635)
);

INVx2_ASAP7_75t_SL g636 ( 
.A(n_414),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_438),
.Y(n_637)
);

INVx4_ASAP7_75t_L g638 ( 
.A(n_456),
.Y(n_638)
);

OR2x2_ASAP7_75t_L g639 ( 
.A(n_438),
.B(n_396),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_493),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_417),
.B(n_297),
.Y(n_641)
);

INVx2_ASAP7_75t_SL g642 ( 
.A(n_417),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_508),
.B(n_465),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_465),
.B(n_252),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_474),
.B(n_482),
.Y(n_645)
);

INVx5_ASAP7_75t_L g646 ( 
.A(n_456),
.Y(n_646)
);

INVx3_ASAP7_75t_L g647 ( 
.A(n_474),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_493),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_493),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_474),
.B(n_299),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_499),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_499),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_425),
.B(n_302),
.Y(n_653)
);

BUFx10_ASAP7_75t_L g654 ( 
.A(n_499),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_482),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_499),
.Y(n_656)
);

NOR2x1p5_ASAP7_75t_L g657 ( 
.A(n_444),
.B(n_396),
.Y(n_657)
);

BUFx6f_ASAP7_75t_L g658 ( 
.A(n_502),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_494),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_502),
.Y(n_660)
);

BUFx6f_ASAP7_75t_SL g661 ( 
.A(n_635),
.Y(n_661)
);

OAI21xp5_ASAP7_75t_L g662 ( 
.A1(n_630),
.A2(n_468),
.B(n_466),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_538),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_543),
.B(n_554),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_543),
.B(n_600),
.Y(n_665)
);

AOI22xp5_ASAP7_75t_L g666 ( 
.A1(n_606),
.A2(n_248),
.B1(n_309),
.B2(n_246),
.Y(n_666)
);

OR2x2_ASAP7_75t_L g667 ( 
.A(n_520),
.B(n_483),
.Y(n_667)
);

INVx1_ASAP7_75t_SL g668 ( 
.A(n_610),
.Y(n_668)
);

A2O1A1Ixp33_ASAP7_75t_L g669 ( 
.A1(n_548),
.A2(n_312),
.B(n_319),
.C(n_314),
.Y(n_669)
);

AOI22xp5_ASAP7_75t_L g670 ( 
.A1(n_606),
.A2(n_309),
.B1(n_248),
.B2(n_509),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_552),
.B(n_468),
.Y(n_671)
);

INVx1_ASAP7_75t_SL g672 ( 
.A(n_610),
.Y(n_672)
);

NOR3xp33_ASAP7_75t_L g673 ( 
.A(n_532),
.B(n_500),
.C(n_497),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_555),
.B(n_492),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_539),
.B(n_492),
.Y(n_675)
);

NOR3xp33_ASAP7_75t_L g676 ( 
.A(n_629),
.B(n_335),
.C(n_329),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_626),
.B(n_492),
.Y(n_677)
);

OAI22xp5_ASAP7_75t_L g678 ( 
.A1(n_616),
.A2(n_407),
.B1(n_273),
.B2(n_389),
.Y(n_678)
);

INVx3_ASAP7_75t_L g679 ( 
.A(n_541),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_526),
.B(n_261),
.Y(n_680)
);

BUFx6f_ASAP7_75t_SL g681 ( 
.A(n_636),
.Y(n_681)
);

INVxp67_ASAP7_75t_L g682 ( 
.A(n_558),
.Y(n_682)
);

OR2x6_ASAP7_75t_L g683 ( 
.A(n_610),
.B(n_445),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_516),
.B(n_264),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_524),
.B(n_266),
.Y(n_685)
);

AOI22xp5_ASAP7_75t_L g686 ( 
.A1(n_535),
.A2(n_470),
.B1(n_507),
.B2(n_352),
.Y(n_686)
);

INVx2_ASAP7_75t_SL g687 ( 
.A(n_610),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_524),
.B(n_267),
.Y(n_688)
);

AOI22xp5_ASAP7_75t_L g689 ( 
.A1(n_535),
.A2(n_556),
.B1(n_547),
.B2(n_562),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_556),
.B(n_268),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_517),
.Y(n_691)
);

BUFx3_ASAP7_75t_L g692 ( 
.A(n_604),
.Y(n_692)
);

AND2x6_ASAP7_75t_L g693 ( 
.A(n_518),
.B(n_338),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_544),
.B(n_285),
.Y(n_694)
);

INVxp67_ASAP7_75t_L g695 ( 
.A(n_576),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_517),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_533),
.B(n_278),
.Y(n_697)
);

INVx2_ASAP7_75t_SL g698 ( 
.A(n_523),
.Y(n_698)
);

BUFx3_ASAP7_75t_L g699 ( 
.A(n_604),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_551),
.B(n_281),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_623),
.B(n_625),
.Y(n_701)
);

AOI22xp5_ASAP7_75t_L g702 ( 
.A1(n_527),
.A2(n_355),
.B1(n_361),
.B2(n_356),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_608),
.B(n_282),
.Y(n_703)
);

OR2x2_ASAP7_75t_L g704 ( 
.A(n_613),
.B(n_605),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_517),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_551),
.B(n_286),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_529),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_611),
.B(n_287),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_621),
.B(n_289),
.Y(n_709)
);

AOI22xp33_ASAP7_75t_SL g710 ( 
.A1(n_616),
.A2(n_431),
.B1(n_489),
.B2(n_444),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_545),
.B(n_553),
.Y(n_711)
);

INVx8_ASAP7_75t_L g712 ( 
.A(n_617),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_551),
.B(n_292),
.Y(n_713)
);

INVxp67_ASAP7_75t_SL g714 ( 
.A(n_546),
.Y(n_714)
);

AOI22xp5_ASAP7_75t_L g715 ( 
.A1(n_582),
.A2(n_377),
.B1(n_365),
.B2(n_368),
.Y(n_715)
);

AOI22xp5_ASAP7_75t_L g716 ( 
.A1(n_631),
.A2(n_370),
.B1(n_375),
.B2(n_382),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_613),
.B(n_405),
.Y(n_717)
);

AOI22xp5_ASAP7_75t_L g718 ( 
.A1(n_632),
.A2(n_388),
.B1(n_392),
.B2(n_343),
.Y(n_718)
);

BUFx5_ASAP7_75t_L g719 ( 
.A(n_573),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_626),
.B(n_298),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_545),
.B(n_304),
.Y(n_721)
);

INVx2_ASAP7_75t_SL g722 ( 
.A(n_515),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_510),
.B(n_307),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_549),
.B(n_406),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_511),
.B(n_308),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_638),
.B(n_310),
.Y(n_726)
);

OR2x2_ASAP7_75t_L g727 ( 
.A(n_643),
.B(n_489),
.Y(n_727)
);

A2O1A1Ixp33_ASAP7_75t_L g728 ( 
.A1(n_529),
.A2(n_494),
.B(n_501),
.C(n_311),
.Y(n_728)
);

NOR2x1p5_ASAP7_75t_L g729 ( 
.A(n_615),
.B(n_317),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_619),
.B(n_318),
.Y(n_730)
);

INVx1_ASAP7_75t_SL g731 ( 
.A(n_528),
.Y(n_731)
);

INVxp67_ASAP7_75t_L g732 ( 
.A(n_615),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_513),
.B(n_320),
.Y(n_733)
);

BUFx8_ASAP7_75t_L g734 ( 
.A(n_657),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_514),
.B(n_321),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_569),
.Y(n_736)
);

NAND3xp33_ASAP7_75t_L g737 ( 
.A(n_634),
.B(n_324),
.C(n_322),
.Y(n_737)
);

AOI22xp5_ASAP7_75t_L g738 ( 
.A1(n_519),
.A2(n_378),
.B1(n_341),
.B2(n_342),
.Y(n_738)
);

INVxp33_ASAP7_75t_L g739 ( 
.A(n_563),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_571),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_575),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_522),
.B(n_328),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_647),
.Y(n_743)
);

AND2x2_ASAP7_75t_L g744 ( 
.A(n_522),
.B(n_351),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_583),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_584),
.Y(n_746)
);

INVx1_ASAP7_75t_SL g747 ( 
.A(n_528),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_585),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_577),
.B(n_359),
.Y(n_749)
);

CKINVDCx20_ASAP7_75t_R g750 ( 
.A(n_536),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_531),
.B(n_366),
.Y(n_751)
);

AND2x4_ASAP7_75t_L g752 ( 
.A(n_542),
.B(n_367),
.Y(n_752)
);

HB1xp67_ASAP7_75t_L g753 ( 
.A(n_536),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_586),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_563),
.B(n_371),
.Y(n_755)
);

BUFx6f_ASAP7_75t_L g756 ( 
.A(n_573),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_537),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_566),
.B(n_380),
.Y(n_758)
);

AOI22xp33_ASAP7_75t_L g759 ( 
.A1(n_581),
.A2(n_494),
.B1(n_501),
.B2(n_409),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_537),
.B(n_391),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_581),
.B(n_401),
.Y(n_761)
);

O2A1O1Ixp33_ASAP7_75t_L g762 ( 
.A1(n_616),
.A2(n_501),
.B(n_404),
.C(n_32),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_639),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_607),
.B(n_425),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_592),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_607),
.B(n_425),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_616),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_612),
.B(n_357),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_593),
.Y(n_769)
);

BUFx6f_ASAP7_75t_L g770 ( 
.A(n_646),
.Y(n_770)
);

BUFx6f_ASAP7_75t_L g771 ( 
.A(n_646),
.Y(n_771)
);

NOR3xp33_ASAP7_75t_L g772 ( 
.A(n_644),
.B(n_29),
.C(n_31),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_595),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_597),
.Y(n_774)
);

INVx2_ASAP7_75t_SL g775 ( 
.A(n_598),
.Y(n_775)
);

AOI22xp5_ASAP7_75t_L g776 ( 
.A1(n_650),
.A2(n_362),
.B1(n_395),
.B2(n_495),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_601),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_602),
.Y(n_778)
);

BUFx10_ASAP7_75t_L g779 ( 
.A(n_650),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_561),
.B(n_453),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_596),
.B(n_453),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_596),
.B(n_480),
.Y(n_782)
);

AND2x2_ASAP7_75t_SL g783 ( 
.A(n_567),
.B(n_31),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_645),
.Y(n_784)
);

A2O1A1Ixp33_ASAP7_75t_L g785 ( 
.A1(n_512),
.A2(n_503),
.B(n_495),
.C(n_491),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_622),
.B(n_480),
.Y(n_786)
);

AOI22xp5_ASAP7_75t_L g787 ( 
.A1(n_617),
.A2(n_495),
.B1(n_491),
.B2(n_36),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_622),
.B(n_491),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_521),
.Y(n_789)
);

INVx8_ASAP7_75t_L g790 ( 
.A(n_622),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_525),
.B(n_34),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_525),
.Y(n_792)
);

CKINVDCx11_ASAP7_75t_R g793 ( 
.A(n_654),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_530),
.B(n_36),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_627),
.B(n_120),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_627),
.B(n_124),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_534),
.B(n_127),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_633),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_628),
.B(n_38),
.Y(n_799)
);

NOR2x1_ASAP7_75t_R g800 ( 
.A(n_692),
.B(n_641),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_731),
.B(n_38),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_671),
.A2(n_578),
.B(n_574),
.Y(n_802)
);

A2O1A1Ixp33_ASAP7_75t_L g803 ( 
.A1(n_663),
.A2(n_578),
.B(n_653),
.C(n_637),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_691),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_682),
.B(n_642),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_689),
.B(n_655),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_739),
.B(n_659),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_695),
.B(n_39),
.Y(n_808)
);

INVxp67_ASAP7_75t_SL g809 ( 
.A(n_666),
.Y(n_809)
);

BUFx3_ASAP7_75t_L g810 ( 
.A(n_793),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_701),
.B(n_40),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_668),
.B(n_654),
.Y(n_812)
);

OAI21xp5_ASAP7_75t_L g813 ( 
.A1(n_677),
.A2(n_557),
.B(n_550),
.Y(n_813)
);

BUFx2_ASAP7_75t_L g814 ( 
.A(n_672),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_775),
.B(n_41),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_711),
.B(n_724),
.Y(n_816)
);

AND2x2_ASAP7_75t_SL g817 ( 
.A(n_783),
.B(n_41),
.Y(n_817)
);

AND2x4_ASAP7_75t_L g818 ( 
.A(n_687),
.B(n_42),
.Y(n_818)
);

OAI22xp5_ASAP7_75t_L g819 ( 
.A1(n_667),
.A2(n_660),
.B1(n_656),
.B2(n_652),
.Y(n_819)
);

NOR3xp33_ASAP7_75t_L g820 ( 
.A(n_678),
.B(n_564),
.C(n_559),
.Y(n_820)
);

O2A1O1Ixp33_ASAP7_75t_L g821 ( 
.A1(n_669),
.A2(n_565),
.B(n_568),
.C(n_570),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_715),
.B(n_44),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_702),
.B(n_44),
.Y(n_823)
);

OAI21xp5_ASAP7_75t_L g824 ( 
.A1(n_662),
.A2(n_568),
.B(n_565),
.Y(n_824)
);

OAI21xp33_ASAP7_75t_L g825 ( 
.A1(n_731),
.A2(n_580),
.B(n_579),
.Y(n_825)
);

AOI22xp33_ASAP7_75t_L g826 ( 
.A1(n_673),
.A2(n_603),
.B1(n_651),
.B2(n_649),
.Y(n_826)
);

CKINVDCx6p67_ASAP7_75t_R g827 ( 
.A(n_699),
.Y(n_827)
);

INVx8_ASAP7_75t_L g828 ( 
.A(n_661),
.Y(n_828)
);

OAI321xp33_ASAP7_75t_L g829 ( 
.A1(n_686),
.A2(n_609),
.A3(n_651),
.B1(n_649),
.B2(n_648),
.C(n_640),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_720),
.A2(n_588),
.B(n_587),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_696),
.Y(n_831)
);

NOR3xp33_ASAP7_75t_L g832 ( 
.A(n_678),
.B(n_591),
.C(n_588),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_694),
.B(n_45),
.Y(n_833)
);

AOI21x1_ASAP7_75t_L g834 ( 
.A1(n_720),
.A2(n_594),
.B(n_591),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_704),
.B(n_730),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_698),
.B(n_46),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_705),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_742),
.B(n_46),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_723),
.A2(n_733),
.B(n_725),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_744),
.B(n_47),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_779),
.B(n_48),
.Y(n_841)
);

INVx4_ASAP7_75t_L g842 ( 
.A(n_712),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_779),
.B(n_49),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_735),
.A2(n_599),
.B(n_624),
.Y(n_844)
);

BUFx2_ASAP7_75t_L g845 ( 
.A(n_750),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_735),
.A2(n_599),
.B(n_620),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_690),
.B(n_49),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_755),
.B(n_51),
.Y(n_848)
);

BUFx4f_ASAP7_75t_L g849 ( 
.A(n_683),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_707),
.Y(n_850)
);

NOR2xp33_ASAP7_75t_L g851 ( 
.A(n_732),
.B(n_51),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_679),
.Y(n_852)
);

OAI21xp5_ASAP7_75t_L g853 ( 
.A1(n_784),
.A2(n_618),
.B(n_658),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_758),
.B(n_52),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_761),
.B(n_54),
.Y(n_855)
);

OAI22xp5_ASAP7_75t_L g856 ( 
.A1(n_756),
.A2(n_54),
.B1(n_55),
.B2(n_56),
.Y(n_856)
);

AOI21x1_ASAP7_75t_L g857 ( 
.A1(n_797),
.A2(n_658),
.B(n_614),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_680),
.B(n_55),
.Y(n_858)
);

NAND3xp33_ASAP7_75t_L g859 ( 
.A(n_772),
.B(n_590),
.C(n_589),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_736),
.B(n_740),
.Y(n_860)
);

HB1xp67_ASAP7_75t_L g861 ( 
.A(n_757),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_741),
.B(n_56),
.Y(n_862)
);

O2A1O1Ixp33_ASAP7_75t_L g863 ( 
.A1(n_762),
.A2(n_58),
.B(n_60),
.C(n_61),
.Y(n_863)
);

AOI21x1_ASAP7_75t_L g864 ( 
.A1(n_797),
.A2(n_590),
.B(n_589),
.Y(n_864)
);

AOI22xp5_ASAP7_75t_L g865 ( 
.A1(n_670),
.A2(n_589),
.B1(n_572),
.B2(n_560),
.Y(n_865)
);

BUFx6f_ASAP7_75t_L g866 ( 
.A(n_770),
.Y(n_866)
);

NOR2x1p5_ASAP7_75t_L g867 ( 
.A(n_727),
.B(n_62),
.Y(n_867)
);

HB1xp67_ASAP7_75t_L g868 ( 
.A(n_753),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_697),
.A2(n_706),
.B(n_700),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_745),
.B(n_62),
.Y(n_870)
);

BUFx12f_ASAP7_75t_L g871 ( 
.A(n_734),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_746),
.B(n_63),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_748),
.Y(n_873)
);

BUFx6f_ASAP7_75t_L g874 ( 
.A(n_770),
.Y(n_874)
);

BUFx6f_ASAP7_75t_L g875 ( 
.A(n_771),
.Y(n_875)
);

AOI21xp33_ASAP7_75t_L g876 ( 
.A1(n_737),
.A2(n_63),
.B(n_66),
.Y(n_876)
);

NOR2x1_ASAP7_75t_L g877 ( 
.A(n_729),
.B(n_540),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_754),
.B(n_67),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_765),
.B(n_68),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_769),
.Y(n_880)
);

NOR3xp33_ASAP7_75t_L g881 ( 
.A(n_710),
.B(n_70),
.C(n_71),
.Y(n_881)
);

NOR3xp33_ASAP7_75t_L g882 ( 
.A(n_664),
.B(n_71),
.C(n_73),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_713),
.A2(n_714),
.B(n_726),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_777),
.B(n_73),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_R g885 ( 
.A(n_661),
.B(n_74),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_773),
.B(n_76),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_774),
.B(n_76),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_778),
.B(n_77),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_722),
.B(n_77),
.Y(n_889)
);

AOI22xp33_ASAP7_75t_L g890 ( 
.A1(n_756),
.A2(n_78),
.B1(n_79),
.B2(n_80),
.Y(n_890)
);

OAI22xp5_ASAP7_75t_L g891 ( 
.A1(n_763),
.A2(n_78),
.B1(n_79),
.B2(n_81),
.Y(n_891)
);

OAI22xp5_ASAP7_75t_L g892 ( 
.A1(n_789),
.A2(n_130),
.B1(n_131),
.B2(n_132),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_L g893 ( 
.A(n_681),
.B(n_134),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_703),
.B(n_241),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_708),
.A2(n_138),
.B(n_141),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_709),
.A2(n_144),
.B(n_150),
.Y(n_896)
);

OR2x6_ASAP7_75t_L g897 ( 
.A(n_683),
.B(n_155),
.Y(n_897)
);

INVx3_ASAP7_75t_L g898 ( 
.A(n_790),
.Y(n_898)
);

HB1xp67_ASAP7_75t_L g899 ( 
.A(n_681),
.Y(n_899)
);

BUFx6f_ASAP7_75t_L g900 ( 
.A(n_771),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_665),
.B(n_161),
.Y(n_901)
);

BUFx8_ASAP7_75t_L g902 ( 
.A(n_752),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_751),
.A2(n_766),
.B(n_764),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_749),
.A2(n_165),
.B(n_167),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_794),
.Y(n_905)
);

BUFx2_ASAP7_75t_L g906 ( 
.A(n_734),
.Y(n_906)
);

AOI22xp5_ASAP7_75t_L g907 ( 
.A1(n_716),
.A2(n_173),
.B1(n_174),
.B2(n_176),
.Y(n_907)
);

O2A1O1Ixp33_ASAP7_75t_L g908 ( 
.A1(n_728),
.A2(n_240),
.B(n_182),
.C(n_183),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_684),
.A2(n_179),
.B(n_187),
.Y(n_909)
);

INVx3_ASAP7_75t_L g910 ( 
.A(n_790),
.Y(n_910)
);

BUFx6f_ASAP7_75t_L g911 ( 
.A(n_712),
.Y(n_911)
);

INVx4_ASAP7_75t_L g912 ( 
.A(n_712),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_752),
.B(n_239),
.Y(n_913)
);

O2A1O1Ixp33_ASAP7_75t_L g914 ( 
.A1(n_676),
.A2(n_685),
.B(n_688),
.C(n_791),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_718),
.B(n_236),
.Y(n_915)
);

A2O1A1Ixp33_ASAP7_75t_L g916 ( 
.A1(n_768),
.A2(n_198),
.B(n_200),
.C(n_202),
.Y(n_916)
);

INVx2_ASAP7_75t_SL g917 ( 
.A(n_717),
.Y(n_917)
);

AND2x2_ASAP7_75t_SL g918 ( 
.A(n_799),
.B(n_204),
.Y(n_918)
);

NOR2xp67_ASAP7_75t_L g919 ( 
.A(n_767),
.B(n_738),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_721),
.B(n_235),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_L g921 ( 
.A(n_760),
.B(n_213),
.Y(n_921)
);

OAI21xp5_ASAP7_75t_L g922 ( 
.A1(n_792),
.A2(n_214),
.B(n_215),
.Y(n_922)
);

OAI22xp5_ASAP7_75t_L g923 ( 
.A1(n_787),
.A2(n_218),
.B1(n_223),
.B2(n_224),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_816),
.B(n_719),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_835),
.B(n_759),
.Y(n_925)
);

OAI21xp5_ASAP7_75t_L g926 ( 
.A1(n_813),
.A2(n_796),
.B(n_795),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_880),
.B(n_719),
.Y(n_927)
);

NAND2x1p5_ASAP7_75t_L g928 ( 
.A(n_842),
.B(n_743),
.Y(n_928)
);

AO31x2_ASAP7_75t_L g929 ( 
.A1(n_916),
.A2(n_785),
.A3(n_781),
.B(n_782),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_871),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_SL g931 ( 
.A(n_814),
.B(n_776),
.Y(n_931)
);

AND2x4_ASAP7_75t_L g932 ( 
.A(n_842),
.B(n_693),
.Y(n_932)
);

OAI21x1_ASAP7_75t_L g933 ( 
.A1(n_824),
.A2(n_798),
.B(n_780),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_860),
.B(n_788),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_804),
.B(n_786),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_831),
.B(n_837),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_850),
.B(n_918),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_SL g938 ( 
.A1(n_897),
.A2(n_818),
.B(n_922),
.Y(n_938)
);

OAI21xp5_ASAP7_75t_L g939 ( 
.A1(n_806),
.A2(n_830),
.B(n_853),
.Y(n_939)
);

OAI21x1_ASAP7_75t_SL g940 ( 
.A1(n_922),
.A2(n_811),
.B(n_847),
.Y(n_940)
);

OAI21x1_ASAP7_75t_SL g941 ( 
.A1(n_841),
.A2(n_843),
.B(n_848),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_808),
.B(n_818),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_817),
.B(n_867),
.Y(n_943)
);

BUFx2_ASAP7_75t_L g944 ( 
.A(n_897),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_L g945 ( 
.A(n_868),
.B(n_845),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_862),
.Y(n_946)
);

INVx2_ASAP7_75t_SL g947 ( 
.A(n_828),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_801),
.B(n_807),
.Y(n_948)
);

OAI22xp5_ASAP7_75t_L g949 ( 
.A1(n_897),
.A2(n_870),
.B1(n_872),
.B2(n_878),
.Y(n_949)
);

AO21x2_ASAP7_75t_L g950 ( 
.A1(n_859),
.A2(n_829),
.B(n_803),
.Y(n_950)
);

OAI21x1_ASAP7_75t_SL g951 ( 
.A1(n_854),
.A2(n_855),
.B(n_912),
.Y(n_951)
);

OAI21xp5_ASAP7_75t_L g952 ( 
.A1(n_909),
.A2(n_903),
.B(n_896),
.Y(n_952)
);

CKINVDCx16_ASAP7_75t_R g953 ( 
.A(n_810),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_879),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_858),
.B(n_838),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_840),
.B(n_865),
.Y(n_956)
);

NAND3xp33_ASAP7_75t_SL g957 ( 
.A(n_881),
.B(n_885),
.C(n_863),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_894),
.A2(n_846),
.B(n_844),
.Y(n_958)
);

AO21x2_ASAP7_75t_L g959 ( 
.A1(n_829),
.A2(n_895),
.B(n_904),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_919),
.B(n_917),
.Y(n_960)
);

INVx1_ASAP7_75t_SL g961 ( 
.A(n_827),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_828),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_884),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_920),
.A2(n_883),
.B(n_869),
.Y(n_964)
);

OAI22xp5_ASAP7_75t_L g965 ( 
.A1(n_833),
.A2(n_849),
.B1(n_886),
.B2(n_888),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_836),
.B(n_913),
.Y(n_966)
);

NAND3xp33_ASAP7_75t_L g967 ( 
.A(n_876),
.B(n_882),
.C(n_832),
.Y(n_967)
);

NOR2x1_ASAP7_75t_L g968 ( 
.A(n_912),
.B(n_906),
.Y(n_968)
);

INVx4_ASAP7_75t_L g969 ( 
.A(n_828),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_851),
.B(n_805),
.Y(n_970)
);

AND2x2_ASAP7_75t_L g971 ( 
.A(n_861),
.B(n_911),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_L g972 ( 
.A(n_899),
.B(n_800),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_911),
.B(n_910),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_887),
.Y(n_974)
);

NAND3xp33_ASAP7_75t_L g975 ( 
.A(n_820),
.B(n_908),
.C(n_890),
.Y(n_975)
);

OAI21xp5_ASAP7_75t_L g976 ( 
.A1(n_821),
.A2(n_826),
.B(n_819),
.Y(n_976)
);

OAI21xp33_ASAP7_75t_L g977 ( 
.A1(n_815),
.A2(n_889),
.B(n_825),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_898),
.B(n_910),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_891),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_898),
.B(n_877),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_915),
.B(n_901),
.Y(n_981)
);

NOR2xp67_ASAP7_75t_L g982 ( 
.A(n_893),
.B(n_921),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_812),
.B(n_856),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_923),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_907),
.B(n_923),
.Y(n_985)
);

NOR2x1_ASAP7_75t_SL g986 ( 
.A(n_866),
.B(n_875),
.Y(n_986)
);

OR2x6_ASAP7_75t_L g987 ( 
.A(n_902),
.B(n_874),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_900),
.B(n_902),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_SL g989 ( 
.A(n_814),
.B(n_668),
.Y(n_989)
);

AO31x2_ASAP7_75t_L g990 ( 
.A1(n_802),
.A2(n_677),
.A3(n_674),
.B(n_671),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_839),
.A2(n_675),
.B(n_677),
.Y(n_991)
);

OAI21xp5_ASAP7_75t_L g992 ( 
.A1(n_802),
.A2(n_677),
.B(n_839),
.Y(n_992)
);

AND2x2_ASAP7_75t_L g993 ( 
.A(n_835),
.B(n_809),
.Y(n_993)
);

BUFx8_ASAP7_75t_L g994 ( 
.A(n_871),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_839),
.A2(n_675),
.B(n_677),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_839),
.A2(n_675),
.B(n_677),
.Y(n_996)
);

BUFx2_ASAP7_75t_L g997 ( 
.A(n_814),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_816),
.B(n_606),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_816),
.B(n_606),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_839),
.A2(n_675),
.B(n_677),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_839),
.A2(n_675),
.B(n_677),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_871),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_816),
.B(n_606),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_839),
.A2(n_675),
.B(n_677),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_816),
.B(n_606),
.Y(n_1005)
);

BUFx5_ASAP7_75t_L g1006 ( 
.A(n_852),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_839),
.A2(n_675),
.B(n_677),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_816),
.B(n_606),
.Y(n_1008)
);

OAI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_802),
.A2(n_677),
.B(n_839),
.Y(n_1009)
);

AOI22xp5_ASAP7_75t_L g1010 ( 
.A1(n_817),
.A2(n_918),
.B1(n_673),
.B2(n_809),
.Y(n_1010)
);

NAND2x1p5_ASAP7_75t_L g1011 ( 
.A(n_842),
.B(n_912),
.Y(n_1011)
);

NOR2xp67_ASAP7_75t_L g1012 ( 
.A(n_871),
.B(n_635),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_839),
.B(n_873),
.Y(n_1013)
);

A2O1A1Ixp33_ASAP7_75t_L g1014 ( 
.A1(n_839),
.A2(n_914),
.B(n_816),
.C(n_905),
.Y(n_1014)
);

AOI21x1_ASAP7_75t_L g1015 ( 
.A1(n_857),
.A2(n_864),
.B(n_834),
.Y(n_1015)
);

O2A1O1Ixp33_ASAP7_75t_L g1016 ( 
.A1(n_822),
.A2(n_669),
.B(n_823),
.C(n_816),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_816),
.B(n_606),
.Y(n_1017)
);

AO32x2_ASAP7_75t_L g1018 ( 
.A1(n_923),
.A2(n_891),
.A3(n_856),
.B1(n_819),
.B2(n_892),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_816),
.B(n_606),
.Y(n_1019)
);

BUFx2_ASAP7_75t_L g1020 ( 
.A(n_814),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_816),
.B(n_606),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_839),
.A2(n_675),
.B(n_677),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_L g1023 ( 
.A(n_809),
.B(n_606),
.Y(n_1023)
);

BUFx5_ASAP7_75t_L g1024 ( 
.A(n_852),
.Y(n_1024)
);

OAI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_802),
.A2(n_677),
.B(n_839),
.Y(n_1025)
);

NAND3xp33_ASAP7_75t_SL g1026 ( 
.A(n_881),
.B(n_747),
.C(n_731),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_816),
.B(n_606),
.Y(n_1027)
);

INVxp67_ASAP7_75t_L g1028 ( 
.A(n_814),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_839),
.A2(n_675),
.B(n_677),
.Y(n_1029)
);

OR2x2_ASAP7_75t_L g1030 ( 
.A(n_809),
.B(n_666),
.Y(n_1030)
);

NAND2x1p5_ASAP7_75t_L g1031 ( 
.A(n_842),
.B(n_912),
.Y(n_1031)
);

OAI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_802),
.A2(n_677),
.B(n_839),
.Y(n_1032)
);

OAI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_918),
.A2(n_817),
.B1(n_897),
.B2(n_905),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_873),
.Y(n_1034)
);

INVx5_ASAP7_75t_L g1035 ( 
.A(n_897),
.Y(n_1035)
);

NAND2x1p5_ASAP7_75t_L g1036 ( 
.A(n_842),
.B(n_912),
.Y(n_1036)
);

BUFx2_ASAP7_75t_L g1037 ( 
.A(n_814),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_816),
.B(n_606),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_839),
.B(n_873),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_816),
.B(n_606),
.Y(n_1040)
);

OAI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_802),
.A2(n_677),
.B(n_839),
.Y(n_1041)
);

OAI22xp5_ASAP7_75t_L g1042 ( 
.A1(n_918),
.A2(n_817),
.B1(n_897),
.B2(n_905),
.Y(n_1042)
);

AOI21x1_ASAP7_75t_L g1043 ( 
.A1(n_857),
.A2(n_864),
.B(n_834),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_873),
.Y(n_1044)
);

BUFx3_ASAP7_75t_L g1045 ( 
.A(n_994),
.Y(n_1045)
);

INVx1_ASAP7_75t_SL g1046 ( 
.A(n_971),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_994),
.Y(n_1047)
);

INVxp67_ASAP7_75t_L g1048 ( 
.A(n_997),
.Y(n_1048)
);

OAI22xp5_ASAP7_75t_L g1049 ( 
.A1(n_1033),
.A2(n_1042),
.B1(n_1035),
.B2(n_1010),
.Y(n_1049)
);

OAI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_1014),
.A2(n_1016),
.B(n_967),
.Y(n_1050)
);

NOR2x1_ASAP7_75t_SL g1051 ( 
.A(n_987),
.B(n_1035),
.Y(n_1051)
);

OAI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_967),
.A2(n_955),
.B(n_998),
.Y(n_1052)
);

OAI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_1033),
.A2(n_1042),
.B1(n_1035),
.B2(n_1010),
.Y(n_1053)
);

INVxp67_ASAP7_75t_L g1054 ( 
.A(n_1020),
.Y(n_1054)
);

OAI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_955),
.A2(n_1003),
.B(n_999),
.Y(n_1055)
);

OR2x2_ASAP7_75t_L g1056 ( 
.A(n_1030),
.B(n_993),
.Y(n_1056)
);

AOI22xp33_ASAP7_75t_L g1057 ( 
.A1(n_1023),
.A2(n_957),
.B1(n_985),
.B2(n_943),
.Y(n_1057)
);

AND2x2_ASAP7_75t_L g1058 ( 
.A(n_1037),
.B(n_925),
.Y(n_1058)
);

AOI22xp33_ASAP7_75t_L g1059 ( 
.A1(n_979),
.A2(n_1026),
.B1(n_944),
.B2(n_949),
.Y(n_1059)
);

AOI221xp5_ASAP7_75t_L g1060 ( 
.A1(n_1005),
.A2(n_1038),
.B1(n_1008),
.B2(n_1040),
.C(n_1017),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_958),
.A2(n_940),
.B(n_991),
.Y(n_1061)
);

INVx3_ASAP7_75t_L g1062 ( 
.A(n_1011),
.Y(n_1062)
);

OAI22xp5_ASAP7_75t_L g1063 ( 
.A1(n_938),
.A2(n_949),
.B1(n_937),
.B2(n_1039),
.Y(n_1063)
);

AOI22xp33_ASAP7_75t_L g1064 ( 
.A1(n_946),
.A2(n_954),
.B1(n_963),
.B2(n_937),
.Y(n_1064)
);

AND2x4_ASAP7_75t_SL g1065 ( 
.A(n_969),
.B(n_987),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_995),
.A2(n_1000),
.B(n_996),
.Y(n_1066)
);

CKINVDCx14_ASAP7_75t_R g1067 ( 
.A(n_930),
.Y(n_1067)
);

INVx4_ASAP7_75t_L g1068 ( 
.A(n_987),
.Y(n_1068)
);

AO221x2_ASAP7_75t_L g1069 ( 
.A1(n_965),
.A2(n_936),
.B1(n_942),
.B2(n_1044),
.C(n_1034),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_1001),
.A2(n_1007),
.B(n_1004),
.Y(n_1070)
);

INVx3_ASAP7_75t_L g1071 ( 
.A(n_1011),
.Y(n_1071)
);

BUFx3_ASAP7_75t_L g1072 ( 
.A(n_969),
.Y(n_1072)
);

OAI21x1_ASAP7_75t_SL g1073 ( 
.A1(n_986),
.A2(n_951),
.B(n_941),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_L g1074 ( 
.A(n_1019),
.B(n_1021),
.Y(n_1074)
);

A2O1A1Ixp33_ASAP7_75t_L g1075 ( 
.A1(n_965),
.A2(n_977),
.B(n_974),
.C(n_970),
.Y(n_1075)
);

AO21x2_ASAP7_75t_L g1076 ( 
.A1(n_992),
.A2(n_1041),
.B(n_1025),
.Y(n_1076)
);

OR2x2_ASAP7_75t_L g1077 ( 
.A(n_1027),
.B(n_1028),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_1022),
.A2(n_1029),
.B(n_1013),
.Y(n_1078)
);

INVx1_ASAP7_75t_SL g1079 ( 
.A(n_961),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_952),
.A2(n_964),
.B(n_1025),
.Y(n_1080)
);

OAI221xp5_ASAP7_75t_L g1081 ( 
.A1(n_948),
.A2(n_966),
.B1(n_945),
.B2(n_934),
.C(n_960),
.Y(n_1081)
);

AO21x2_ASAP7_75t_L g1082 ( 
.A1(n_992),
.A2(n_1009),
.B(n_1032),
.Y(n_1082)
);

OR2x6_ASAP7_75t_L g1083 ( 
.A(n_1031),
.B(n_1036),
.Y(n_1083)
);

BUFx2_ASAP7_75t_L g1084 ( 
.A(n_1031),
.Y(n_1084)
);

INVxp67_ASAP7_75t_L g1085 ( 
.A(n_989),
.Y(n_1085)
);

AND2x4_ASAP7_75t_L g1086 ( 
.A(n_932),
.B(n_988),
.Y(n_1086)
);

BUFx4_ASAP7_75t_SL g1087 ( 
.A(n_1002),
.Y(n_1087)
);

AOI221xp5_ASAP7_75t_L g1088 ( 
.A1(n_972),
.A2(n_976),
.B1(n_935),
.B2(n_939),
.C(n_977),
.Y(n_1088)
);

BUFx2_ASAP7_75t_L g1089 ( 
.A(n_962),
.Y(n_1089)
);

INVx2_ASAP7_75t_SL g1090 ( 
.A(n_968),
.Y(n_1090)
);

CKINVDCx6p67_ASAP7_75t_R g1091 ( 
.A(n_953),
.Y(n_1091)
);

NAND3xp33_ASAP7_75t_SL g1092 ( 
.A(n_981),
.B(n_976),
.C(n_956),
.Y(n_1092)
);

AOI21xp33_ASAP7_75t_SL g1093 ( 
.A1(n_947),
.A2(n_928),
.B(n_932),
.Y(n_1093)
);

OAI22xp5_ASAP7_75t_L g1094 ( 
.A1(n_975),
.A2(n_924),
.B1(n_982),
.B2(n_983),
.Y(n_1094)
);

AO21x2_ASAP7_75t_L g1095 ( 
.A1(n_950),
.A2(n_959),
.B(n_926),
.Y(n_1095)
);

AO21x2_ASAP7_75t_L g1096 ( 
.A1(n_950),
.A2(n_959),
.B(n_933),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_990),
.Y(n_1097)
);

OR2x6_ASAP7_75t_L g1098 ( 
.A(n_1012),
.B(n_973),
.Y(n_1098)
);

AOI22xp5_ASAP7_75t_L g1099 ( 
.A1(n_961),
.A2(n_931),
.B1(n_927),
.B2(n_978),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_980),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_1006),
.B(n_1024),
.Y(n_1101)
);

NOR2xp33_ASAP7_75t_L g1102 ( 
.A(n_1006),
.B(n_1024),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_929),
.Y(n_1103)
);

NOR3xp33_ASAP7_75t_L g1104 ( 
.A(n_1018),
.B(n_1042),
.C(n_1033),
.Y(n_1104)
);

AOI22xp5_ASAP7_75t_L g1105 ( 
.A1(n_929),
.A2(n_508),
.B1(n_1023),
.B2(n_606),
.Y(n_1105)
);

OAI22xp5_ASAP7_75t_L g1106 ( 
.A1(n_1033),
.A2(n_1042),
.B1(n_1035),
.B2(n_817),
.Y(n_1106)
);

NAND2x1p5_ASAP7_75t_L g1107 ( 
.A(n_1035),
.B(n_969),
.Y(n_1107)
);

OAI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_1014),
.A2(n_839),
.B(n_1016),
.Y(n_1108)
);

AOI221xp5_ASAP7_75t_L g1109 ( 
.A1(n_1033),
.A2(n_1042),
.B1(n_673),
.B2(n_1023),
.C(n_532),
.Y(n_1109)
);

AO21x2_ASAP7_75t_L g1110 ( 
.A1(n_940),
.A2(n_1043),
.B(n_1015),
.Y(n_1110)
);

OAI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_1014),
.A2(n_839),
.B(n_1016),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_994),
.Y(n_1112)
);

AOI22xp5_ASAP7_75t_L g1113 ( 
.A1(n_1023),
.A2(n_508),
.B1(n_606),
.B2(n_1033),
.Y(n_1113)
);

INVxp67_ASAP7_75t_SL g1114 ( 
.A(n_1033),
.Y(n_1114)
);

AND2x4_ASAP7_75t_L g1115 ( 
.A(n_1035),
.B(n_969),
.Y(n_1115)
);

AOI22xp33_ASAP7_75t_L g1116 ( 
.A1(n_1033),
.A2(n_1042),
.B1(n_817),
.B2(n_984),
.Y(n_1116)
);

AO21x2_ASAP7_75t_L g1117 ( 
.A1(n_940),
.A2(n_1043),
.B(n_1015),
.Y(n_1117)
);

O2A1O1Ixp33_ASAP7_75t_SL g1118 ( 
.A1(n_1014),
.A2(n_1042),
.B(n_1033),
.C(n_1039),
.Y(n_1118)
);

AOI221xp5_ASAP7_75t_L g1119 ( 
.A1(n_1033),
.A2(n_1042),
.B1(n_673),
.B2(n_1023),
.C(n_532),
.Y(n_1119)
);

OAI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_1014),
.A2(n_839),
.B(n_1016),
.Y(n_1120)
);

OAI22xp5_ASAP7_75t_L g1121 ( 
.A1(n_1033),
.A2(n_1042),
.B1(n_1035),
.B2(n_817),
.Y(n_1121)
);

INVx3_ASAP7_75t_L g1122 ( 
.A(n_1011),
.Y(n_1122)
);

INVx3_ASAP7_75t_L g1123 ( 
.A(n_1011),
.Y(n_1123)
);

BUFx3_ASAP7_75t_L g1124 ( 
.A(n_994),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_958),
.A2(n_1014),
.B(n_940),
.Y(n_1125)
);

INVx1_ASAP7_75t_SL g1126 ( 
.A(n_971),
.Y(n_1126)
);

AO21x2_ASAP7_75t_L g1127 ( 
.A1(n_940),
.A2(n_1043),
.B(n_1015),
.Y(n_1127)
);

BUFx4f_ASAP7_75t_SL g1128 ( 
.A(n_1045),
.Y(n_1128)
);

OAI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_1075),
.A2(n_1052),
.B(n_1057),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_1097),
.Y(n_1130)
);

HB1xp67_ASAP7_75t_L g1131 ( 
.A(n_1046),
.Y(n_1131)
);

AO21x2_ASAP7_75t_L g1132 ( 
.A1(n_1125),
.A2(n_1080),
.B(n_1061),
.Y(n_1132)
);

INVx2_ASAP7_75t_SL g1133 ( 
.A(n_1083),
.Y(n_1133)
);

BUFx2_ASAP7_75t_L g1134 ( 
.A(n_1101),
.Y(n_1134)
);

OR2x2_ASAP7_75t_L g1135 ( 
.A(n_1056),
.B(n_1114),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1074),
.B(n_1060),
.Y(n_1136)
);

OAI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_1057),
.A2(n_1119),
.B(n_1109),
.Y(n_1137)
);

BUFx3_ASAP7_75t_L g1138 ( 
.A(n_1072),
.Y(n_1138)
);

OR2x2_ASAP7_75t_L g1139 ( 
.A(n_1114),
.B(n_1049),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1076),
.Y(n_1140)
);

HB1xp67_ASAP7_75t_L g1141 ( 
.A(n_1126),
.Y(n_1141)
);

CKINVDCx14_ASAP7_75t_R g1142 ( 
.A(n_1067),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1076),
.Y(n_1143)
);

HB1xp67_ASAP7_75t_L g1144 ( 
.A(n_1083),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1082),
.Y(n_1145)
);

INVxp67_ASAP7_75t_L g1146 ( 
.A(n_1084),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1050),
.Y(n_1147)
);

HB1xp67_ASAP7_75t_L g1148 ( 
.A(n_1048),
.Y(n_1148)
);

INVx2_ASAP7_75t_SL g1149 ( 
.A(n_1065),
.Y(n_1149)
);

HB1xp67_ASAP7_75t_L g1150 ( 
.A(n_1048),
.Y(n_1150)
);

BUFx12f_ASAP7_75t_L g1151 ( 
.A(n_1047),
.Y(n_1151)
);

OAI21xp33_ASAP7_75t_L g1152 ( 
.A1(n_1116),
.A2(n_1104),
.B(n_1109),
.Y(n_1152)
);

OR2x2_ASAP7_75t_L g1153 ( 
.A(n_1049),
.B(n_1053),
.Y(n_1153)
);

AOI22xp5_ASAP7_75t_L g1154 ( 
.A1(n_1119),
.A2(n_1121),
.B1(n_1106),
.B2(n_1116),
.Y(n_1154)
);

AO21x2_ASAP7_75t_L g1155 ( 
.A1(n_1066),
.A2(n_1070),
.B(n_1120),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1074),
.B(n_1060),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1069),
.Y(n_1157)
);

AO31x2_ASAP7_75t_L g1158 ( 
.A1(n_1078),
.A2(n_1103),
.A3(n_1070),
.B(n_1063),
.Y(n_1158)
);

HB1xp67_ASAP7_75t_L g1159 ( 
.A(n_1054),
.Y(n_1159)
);

NOR2xp33_ASAP7_75t_L g1160 ( 
.A(n_1113),
.B(n_1081),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1069),
.Y(n_1161)
);

AND2x2_ASAP7_75t_L g1162 ( 
.A(n_1064),
.B(n_1058),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1108),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1111),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1055),
.B(n_1077),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1078),
.Y(n_1166)
);

HB1xp67_ASAP7_75t_L g1167 ( 
.A(n_1054),
.Y(n_1167)
);

NOR2xp33_ASAP7_75t_L g1168 ( 
.A(n_1081),
.B(n_1068),
.Y(n_1168)
);

INVx4_ASAP7_75t_L g1169 ( 
.A(n_1107),
.Y(n_1169)
);

OR2x6_ASAP7_75t_L g1170 ( 
.A(n_1053),
.B(n_1121),
.Y(n_1170)
);

BUFx8_ASAP7_75t_SL g1171 ( 
.A(n_1112),
.Y(n_1171)
);

AND2x2_ASAP7_75t_L g1172 ( 
.A(n_1170),
.B(n_1095),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_SL g1173 ( 
.A(n_1168),
.B(n_1106),
.Y(n_1173)
);

BUFx2_ASAP7_75t_L g1174 ( 
.A(n_1134),
.Y(n_1174)
);

AND2x2_ASAP7_75t_SL g1175 ( 
.A(n_1153),
.B(n_1102),
.Y(n_1175)
);

CKINVDCx11_ASAP7_75t_R g1176 ( 
.A(n_1151),
.Y(n_1176)
);

AND2x2_ASAP7_75t_L g1177 ( 
.A(n_1170),
.B(n_1095),
.Y(n_1177)
);

BUFx2_ASAP7_75t_L g1178 ( 
.A(n_1134),
.Y(n_1178)
);

OR2x2_ASAP7_75t_L g1179 ( 
.A(n_1153),
.B(n_1063),
.Y(n_1179)
);

NOR2x1p5_ASAP7_75t_L g1180 ( 
.A(n_1169),
.B(n_1068),
.Y(n_1180)
);

AND2x2_ASAP7_75t_L g1181 ( 
.A(n_1170),
.B(n_1096),
.Y(n_1181)
);

HB1xp67_ASAP7_75t_L g1182 ( 
.A(n_1130),
.Y(n_1182)
);

AND2x2_ASAP7_75t_L g1183 ( 
.A(n_1139),
.B(n_1127),
.Y(n_1183)
);

AND2x2_ASAP7_75t_L g1184 ( 
.A(n_1163),
.B(n_1110),
.Y(n_1184)
);

OR2x2_ASAP7_75t_L g1185 ( 
.A(n_1135),
.B(n_1092),
.Y(n_1185)
);

AND2x2_ASAP7_75t_L g1186 ( 
.A(n_1164),
.B(n_1117),
.Y(n_1186)
);

INVx5_ASAP7_75t_L g1187 ( 
.A(n_1169),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1166),
.Y(n_1188)
);

AND2x2_ASAP7_75t_L g1189 ( 
.A(n_1140),
.B(n_1143),
.Y(n_1189)
);

BUFx3_ASAP7_75t_L g1190 ( 
.A(n_1169),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1145),
.Y(n_1191)
);

AOI22xp33_ASAP7_75t_L g1192 ( 
.A1(n_1137),
.A2(n_1105),
.B1(n_1092),
.B2(n_1088),
.Y(n_1192)
);

AOI22xp33_ASAP7_75t_L g1193 ( 
.A1(n_1152),
.A2(n_1059),
.B1(n_1094),
.B2(n_1100),
.Y(n_1193)
);

CKINVDCx16_ASAP7_75t_R g1194 ( 
.A(n_1142),
.Y(n_1194)
);

INVx4_ASAP7_75t_L g1195 ( 
.A(n_1187),
.Y(n_1195)
);

INVxp67_ASAP7_75t_L g1196 ( 
.A(n_1174),
.Y(n_1196)
);

AND2x2_ASAP7_75t_L g1197 ( 
.A(n_1183),
.B(n_1132),
.Y(n_1197)
);

AND2x2_ASAP7_75t_L g1198 ( 
.A(n_1183),
.B(n_1132),
.Y(n_1198)
);

AND2x2_ASAP7_75t_L g1199 ( 
.A(n_1183),
.B(n_1132),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1191),
.Y(n_1200)
);

NAND2x1_ASAP7_75t_L g1201 ( 
.A(n_1174),
.B(n_1073),
.Y(n_1201)
);

AND2x4_ASAP7_75t_L g1202 ( 
.A(n_1188),
.B(n_1155),
.Y(n_1202)
);

INVx2_ASAP7_75t_SL g1203 ( 
.A(n_1187),
.Y(n_1203)
);

OR2x2_ASAP7_75t_L g1204 ( 
.A(n_1185),
.B(n_1179),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1189),
.Y(n_1205)
);

HB1xp67_ASAP7_75t_L g1206 ( 
.A(n_1182),
.Y(n_1206)
);

AND2x2_ASAP7_75t_L g1207 ( 
.A(n_1184),
.B(n_1186),
.Y(n_1207)
);

AND2x4_ASAP7_75t_L g1208 ( 
.A(n_1188),
.B(n_1158),
.Y(n_1208)
);

NOR2xp33_ASAP7_75t_L g1209 ( 
.A(n_1173),
.B(n_1136),
.Y(n_1209)
);

OR2x2_ASAP7_75t_L g1210 ( 
.A(n_1185),
.B(n_1147),
.Y(n_1210)
);

BUFx3_ASAP7_75t_L g1211 ( 
.A(n_1187),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1189),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1189),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1205),
.B(n_1212),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_1207),
.B(n_1172),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1200),
.Y(n_1216)
);

INVx1_ASAP7_75t_SL g1217 ( 
.A(n_1211),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1200),
.Y(n_1218)
);

AND2x2_ASAP7_75t_L g1219 ( 
.A(n_1207),
.B(n_1172),
.Y(n_1219)
);

AND2x2_ASAP7_75t_L g1220 ( 
.A(n_1197),
.B(n_1181),
.Y(n_1220)
);

AND2x2_ASAP7_75t_L g1221 ( 
.A(n_1197),
.B(n_1177),
.Y(n_1221)
);

OR2x2_ASAP7_75t_L g1222 ( 
.A(n_1204),
.B(n_1185),
.Y(n_1222)
);

AND2x2_ASAP7_75t_L g1223 ( 
.A(n_1197),
.B(n_1177),
.Y(n_1223)
);

OR2x2_ASAP7_75t_L g1224 ( 
.A(n_1204),
.B(n_1178),
.Y(n_1224)
);

HB1xp67_ASAP7_75t_L g1225 ( 
.A(n_1206),
.Y(n_1225)
);

AND2x2_ASAP7_75t_L g1226 ( 
.A(n_1198),
.B(n_1177),
.Y(n_1226)
);

AND2x4_ASAP7_75t_L g1227 ( 
.A(n_1202),
.B(n_1208),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1213),
.B(n_1198),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1222),
.B(n_1213),
.Y(n_1229)
);

INVxp67_ASAP7_75t_SL g1230 ( 
.A(n_1225),
.Y(n_1230)
);

AND2x2_ASAP7_75t_L g1231 ( 
.A(n_1220),
.B(n_1198),
.Y(n_1231)
);

NAND2x1p5_ASAP7_75t_L g1232 ( 
.A(n_1217),
.B(n_1195),
.Y(n_1232)
);

O2A1O1Ixp33_ASAP7_75t_SL g1233 ( 
.A1(n_1217),
.A2(n_1203),
.B(n_1201),
.C(n_1149),
.Y(n_1233)
);

NAND2x1p5_ASAP7_75t_L g1234 ( 
.A(n_1224),
.B(n_1195),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1214),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1222),
.B(n_1199),
.Y(n_1236)
);

OR2x6_ASAP7_75t_L g1237 ( 
.A(n_1227),
.B(n_1195),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1214),
.Y(n_1238)
);

AND2x2_ASAP7_75t_L g1239 ( 
.A(n_1220),
.B(n_1199),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1216),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1216),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1218),
.Y(n_1242)
);

OAI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1225),
.A2(n_1160),
.B(n_1156),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1218),
.Y(n_1244)
);

AND2x4_ASAP7_75t_L g1245 ( 
.A(n_1227),
.B(n_1195),
.Y(n_1245)
);

OAI221xp5_ASAP7_75t_L g1246 ( 
.A1(n_1243),
.A2(n_1152),
.B1(n_1154),
.B2(n_1209),
.C(n_1192),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1235),
.Y(n_1247)
);

OAI22xp5_ASAP7_75t_L g1248 ( 
.A1(n_1237),
.A2(n_1195),
.B1(n_1194),
.B2(n_1154),
.Y(n_1248)
);

AOI22xp5_ASAP7_75t_L g1249 ( 
.A1(n_1237),
.A2(n_1209),
.B1(n_1227),
.B2(n_1173),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1238),
.B(n_1220),
.Y(n_1250)
);

NAND3xp33_ASAP7_75t_L g1251 ( 
.A(n_1230),
.B(n_1210),
.C(n_1228),
.Y(n_1251)
);

AOI22xp5_ASAP7_75t_L g1252 ( 
.A1(n_1237),
.A2(n_1227),
.B1(n_1175),
.B2(n_1199),
.Y(n_1252)
);

OR2x2_ASAP7_75t_L g1253 ( 
.A(n_1236),
.B(n_1228),
.Y(n_1253)
);

O2A1O1Ixp33_ASAP7_75t_L g1254 ( 
.A1(n_1233),
.A2(n_1118),
.B(n_1129),
.C(n_1148),
.Y(n_1254)
);

NOR2xp33_ASAP7_75t_L g1255 ( 
.A(n_1229),
.B(n_1194),
.Y(n_1255)
);

OAI22xp5_ASAP7_75t_L g1256 ( 
.A1(n_1237),
.A2(n_1203),
.B1(n_1187),
.B2(n_1190),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1240),
.Y(n_1257)
);

OR2x6_ASAP7_75t_L g1258 ( 
.A(n_1232),
.B(n_1203),
.Y(n_1258)
);

INVxp67_ASAP7_75t_L g1259 ( 
.A(n_1241),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1242),
.Y(n_1260)
);

AOI22xp5_ASAP7_75t_L g1261 ( 
.A1(n_1245),
.A2(n_1175),
.B1(n_1226),
.B2(n_1221),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1244),
.Y(n_1262)
);

INVx2_ASAP7_75t_L g1263 ( 
.A(n_1234),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1231),
.Y(n_1264)
);

NAND2x1_ASAP7_75t_L g1265 ( 
.A(n_1258),
.B(n_1245),
.Y(n_1265)
);

AND2x2_ASAP7_75t_L g1266 ( 
.A(n_1264),
.B(n_1231),
.Y(n_1266)
);

NOR3xp33_ASAP7_75t_L g1267 ( 
.A(n_1246),
.B(n_1176),
.C(n_1079),
.Y(n_1267)
);

OR2x2_ASAP7_75t_L g1268 ( 
.A(n_1253),
.B(n_1239),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1247),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1257),
.Y(n_1270)
);

OAI22xp33_ASAP7_75t_SL g1271 ( 
.A1(n_1258),
.A2(n_1234),
.B1(n_1232),
.B2(n_1245),
.Y(n_1271)
);

OAI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1254),
.A2(n_1233),
.B(n_1234),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1251),
.B(n_1239),
.Y(n_1273)
);

NOR2x1_ASAP7_75t_L g1274 ( 
.A(n_1272),
.B(n_1124),
.Y(n_1274)
);

AOI211x1_ASAP7_75t_L g1275 ( 
.A1(n_1272),
.A2(n_1248),
.B(n_1250),
.C(n_1256),
.Y(n_1275)
);

INVx2_ASAP7_75t_L g1276 ( 
.A(n_1265),
.Y(n_1276)
);

AOI22xp33_ASAP7_75t_L g1277 ( 
.A1(n_1267),
.A2(n_1252),
.B1(n_1249),
.B2(n_1255),
.Y(n_1277)
);

AOI211xp5_ASAP7_75t_L g1278 ( 
.A1(n_1271),
.A2(n_1118),
.B(n_1263),
.C(n_1261),
.Y(n_1278)
);

AOI221xp5_ASAP7_75t_L g1279 ( 
.A1(n_1273),
.A2(n_1259),
.B1(n_1262),
.B2(n_1260),
.C(n_1150),
.Y(n_1279)
);

INVxp33_ASAP7_75t_L g1280 ( 
.A(n_1266),
.Y(n_1280)
);

AOI22xp5_ASAP7_75t_L g1281 ( 
.A1(n_1269),
.A2(n_1258),
.B1(n_1175),
.B2(n_1223),
.Y(n_1281)
);

NAND4xp25_ASAP7_75t_L g1282 ( 
.A(n_1268),
.B(n_1192),
.C(n_1193),
.D(n_1165),
.Y(n_1282)
);

NAND4xp25_ASAP7_75t_L g1283 ( 
.A(n_1270),
.B(n_1193),
.C(n_1089),
.D(n_1161),
.Y(n_1283)
);

NOR3x1_ASAP7_75t_L g1284 ( 
.A(n_1283),
.B(n_1176),
.C(n_1149),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1274),
.Y(n_1285)
);

AOI221xp5_ASAP7_75t_SL g1286 ( 
.A1(n_1278),
.A2(n_1196),
.B1(n_1146),
.B2(n_1161),
.C(n_1157),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1279),
.B(n_1215),
.Y(n_1287)
);

NAND4xp25_ASAP7_75t_L g1288 ( 
.A(n_1275),
.B(n_1138),
.C(n_1115),
.D(n_1157),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1280),
.B(n_1215),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_SL g1290 ( 
.A(n_1276),
.B(n_1128),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1282),
.Y(n_1291)
);

NAND3xp33_ASAP7_75t_SL g1292 ( 
.A(n_1291),
.B(n_1277),
.C(n_1281),
.Y(n_1292)
);

NOR3xp33_ASAP7_75t_L g1293 ( 
.A(n_1288),
.B(n_1090),
.C(n_1138),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1289),
.Y(n_1294)
);

NOR3x1_ASAP7_75t_L g1295 ( 
.A(n_1290),
.B(n_1087),
.C(n_1091),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_SL g1296 ( 
.A(n_1286),
.B(n_1151),
.Y(n_1296)
);

NOR3xp33_ASAP7_75t_L g1297 ( 
.A(n_1290),
.B(n_1087),
.C(n_1115),
.Y(n_1297)
);

NOR3xp33_ASAP7_75t_L g1298 ( 
.A(n_1285),
.B(n_1093),
.C(n_1071),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1294),
.Y(n_1299)
);

AOI22xp5_ASAP7_75t_L g1300 ( 
.A1(n_1292),
.A2(n_1287),
.B1(n_1284),
.B2(n_1175),
.Y(n_1300)
);

NAND2x1p5_ASAP7_75t_L g1301 ( 
.A(n_1295),
.B(n_1171),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1296),
.Y(n_1302)
);

NAND4xp75_ASAP7_75t_L g1303 ( 
.A(n_1297),
.B(n_1051),
.C(n_1133),
.D(n_1107),
.Y(n_1303)
);

NAND4xp75_ASAP7_75t_L g1304 ( 
.A(n_1293),
.B(n_1133),
.C(n_1162),
.D(n_1099),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1298),
.B(n_1219),
.Y(n_1305)
);

INVx2_ASAP7_75t_SL g1306 ( 
.A(n_1296),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1299),
.Y(n_1307)
);

NOR2xp33_ASAP7_75t_L g1308 ( 
.A(n_1301),
.B(n_1131),
.Y(n_1308)
);

AND2x4_ASAP7_75t_L g1309 ( 
.A(n_1306),
.B(n_1159),
.Y(n_1309)
);

AO22x2_ASAP7_75t_L g1310 ( 
.A1(n_1307),
.A2(n_1299),
.B1(n_1302),
.B2(n_1304),
.Y(n_1310)
);

AND2x2_ASAP7_75t_L g1311 ( 
.A(n_1308),
.B(n_1309),
.Y(n_1311)
);

AOI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1308),
.A2(n_1300),
.B(n_1305),
.Y(n_1312)
);

AOI22xp33_ASAP7_75t_L g1313 ( 
.A1(n_1310),
.A2(n_1311),
.B1(n_1312),
.B2(n_1303),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1312),
.B(n_1167),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1314),
.Y(n_1315)
);

AO22x2_ASAP7_75t_L g1316 ( 
.A1(n_1313),
.A2(n_1062),
.B1(n_1071),
.B2(n_1123),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1314),
.Y(n_1317)
);

XNOR2xp5_ASAP7_75t_L g1318 ( 
.A(n_1316),
.B(n_1086),
.Y(n_1318)
);

AOI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1315),
.A2(n_1098),
.B(n_1085),
.Y(n_1319)
);

AOI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1317),
.A2(n_1180),
.B1(n_1086),
.B2(n_1144),
.Y(n_1320)
);

OAI22xp33_ASAP7_75t_L g1321 ( 
.A1(n_1320),
.A2(n_1098),
.B1(n_1187),
.B2(n_1141),
.Y(n_1321)
);

OA21x2_ASAP7_75t_L g1322 ( 
.A1(n_1321),
.A2(n_1319),
.B(n_1318),
.Y(n_1322)
);

XNOR2xp5_ASAP7_75t_L g1323 ( 
.A(n_1322),
.B(n_1098),
.Y(n_1323)
);

AOI22xp5_ASAP7_75t_L g1324 ( 
.A1(n_1323),
.A2(n_1180),
.B1(n_1122),
.B2(n_1062),
.Y(n_1324)
);


endmodule