module fake_jpeg_148_n_128 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_128);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_128;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

AND2x2_ASAP7_75t_L g12 ( 
.A(n_2),
.B(n_10),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_4),
.B(n_8),
.Y(n_13)
);

BUFx16f_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

HAxp5_ASAP7_75t_SL g28 ( 
.A(n_14),
.B(n_13),
.CON(n_28),
.SN(n_28)
);

A2O1A1Ixp33_ASAP7_75t_L g48 ( 
.A1(n_28),
.A2(n_18),
.B(n_24),
.C(n_19),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g29 ( 
.A1(n_13),
.A2(n_2),
.B(n_3),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_29),
.B(n_36),
.C(n_40),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_22),
.B(n_3),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_31),
.B(n_38),
.Y(n_65)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx4_ASAP7_75t_SL g54 ( 
.A(n_32),
.Y(n_54)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx4_ASAP7_75t_SL g36 ( 
.A(n_27),
.Y(n_36)
);

CKINVDCx14_ASAP7_75t_R g67 ( 
.A(n_36),
.Y(n_67)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_23),
.B(n_26),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_12),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_5),
.Y(n_58)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_43),
.B(n_12),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_46),
.B(n_49),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_39),
.A2(n_18),
.B1(n_24),
.B2(n_12),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_47),
.A2(n_57),
.B1(n_66),
.B2(n_67),
.Y(n_77)
);

NOR2xp67_ASAP7_75t_L g79 ( 
.A(n_48),
.B(n_65),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_33),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_28),
.B(n_20),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_56),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_34),
.A2(n_25),
.B1(n_17),
.B2(n_19),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_60),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_42),
.A2(n_20),
.B(n_17),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_39),
.A2(n_25),
.B1(n_2),
.B2(n_6),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_58),
.B(n_62),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_32),
.A2(n_7),
.B1(n_9),
.B2(n_11),
.Y(n_60)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_69),
.Y(n_91)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_70),
.Y(n_93)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_63),
.A2(n_30),
.B1(n_35),
.B2(n_44),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_84),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_48),
.B(n_47),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_SL g85 ( 
.A(n_76),
.B(n_57),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_77),
.A2(n_66),
.B(n_45),
.Y(n_96)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_79),
.B(n_81),
.Y(n_97)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_53),
.B(n_59),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_85),
.B(n_88),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_83),
.B(n_73),
.C(n_76),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_87),
.B(n_75),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_82),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_70),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_89),
.B(n_96),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_99),
.Y(n_107)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_91),
.Y(n_100)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_100),
.Y(n_112)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_93),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_101),
.B(n_102),
.Y(n_111)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_94),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_95),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_103),
.B(n_105),
.C(n_78),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_97),
.B(n_87),
.Y(n_104)
);

OAI32xp33_ASAP7_75t_L g110 ( 
.A1(n_104),
.A2(n_106),
.A3(n_90),
.B1(n_75),
.B2(n_101),
.Y(n_110)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_108),
.B(n_110),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_98),
.B(n_89),
.C(n_85),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_109),
.B(n_113),
.C(n_92),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_106),
.B(n_90),
.C(n_96),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_111),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_114),
.B(n_68),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_107),
.A2(n_102),
.B(n_100),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_116),
.A2(n_117),
.B(n_45),
.Y(n_121)
);

A2O1A1Ixp33_ASAP7_75t_SL g117 ( 
.A1(n_111),
.A2(n_72),
.B(n_105),
.C(n_69),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_112),
.C(n_71),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_119),
.B(n_82),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_120),
.B(n_121),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_123),
.B(n_44),
.Y(n_125)
);

OAI21xp33_ASAP7_75t_L g124 ( 
.A1(n_122),
.A2(n_115),
.B(n_117),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_124),
.B(n_125),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_45),
.C(n_61),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_61),
.Y(n_128)
);


endmodule