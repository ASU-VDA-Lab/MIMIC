module fake_jpeg_13745_n_214 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_214);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_214;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_2),
.B(n_5),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_10),
.B(n_9),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_0),
.B(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_28),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_32),
.B(n_39),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_33),
.Y(n_70)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_35),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_37),
.Y(n_85)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g39 ( 
.A(n_16),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_40),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_15),
.B(n_1),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_41),
.B(n_47),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_15),
.B(n_1),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_44),
.B(n_48),
.Y(n_75)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

INVx5_ASAP7_75t_SL g46 ( 
.A(n_28),
.Y(n_46)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_16),
.B(n_1),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_19),
.B(n_3),
.Y(n_48)
);

BUFx24_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

CKINVDCx12_ASAP7_75t_R g66 ( 
.A(n_51),
.Y(n_66)
);

INVx6_ASAP7_75t_SL g52 ( 
.A(n_29),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_52),
.B(n_18),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_14),
.Y(n_54)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_19),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_55),
.B(n_75),
.Y(n_103)
);

AND2x2_ASAP7_75t_SL g57 ( 
.A(n_43),
.B(n_29),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_57),
.B(n_36),
.Y(n_94)
);

NAND2xp33_ASAP7_75t_SL g61 ( 
.A(n_52),
.B(n_29),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_61),
.A2(n_65),
.B(n_64),
.Y(n_116)
);

OA22x2_ASAP7_75t_L g65 ( 
.A1(n_50),
.A2(n_22),
.B1(n_27),
.B2(n_26),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_35),
.A2(n_22),
.B1(n_30),
.B2(n_21),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_69),
.A2(n_90),
.B1(n_7),
.B2(n_8),
.Y(n_108)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_72),
.Y(n_106)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_36),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_49),
.A2(n_31),
.B1(n_27),
.B2(n_26),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_77),
.A2(n_82),
.B1(n_86),
.B2(n_3),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_48),
.B(n_44),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_79),
.B(n_80),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_32),
.B(n_30),
.Y(n_80)
);

INVx2_ASAP7_75t_SL g101 ( 
.A(n_81),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_49),
.A2(n_18),
.B1(n_25),
.B2(n_31),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_40),
.A2(n_22),
.B1(n_25),
.B2(n_24),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_83),
.A2(n_84),
.B1(n_57),
.B2(n_72),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_53),
.A2(n_22),
.B1(n_24),
.B2(n_21),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_46),
.A2(n_20),
.B1(n_5),
.B2(n_6),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_33),
.B(n_20),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_88),
.B(n_89),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_33),
.B(n_36),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_34),
.A2(n_11),
.B1(n_5),
.B2(n_6),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_33),
.Y(n_92)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_81),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_93),
.B(n_60),
.Y(n_120)
);

NAND2xp33_ASAP7_75t_SL g130 ( 
.A(n_94),
.B(n_102),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_95),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_83),
.A2(n_42),
.B1(n_45),
.B2(n_51),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_96),
.A2(n_119),
.B1(n_116),
.B2(n_92),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_62),
.B(n_9),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_99),
.B(n_107),
.Y(n_124)
);

OR2x4_ASAP7_75t_L g100 ( 
.A(n_61),
.B(n_3),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_100),
.B(n_103),
.Y(n_142)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_73),
.Y(n_104)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_104),
.Y(n_132)
);

OR2x6_ASAP7_75t_L g127 ( 
.A(n_105),
.B(n_113),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_55),
.B(n_6),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_108),
.A2(n_110),
.B1(n_117),
.B2(n_118),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_56),
.B(n_8),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_109),
.B(n_66),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_90),
.A2(n_65),
.B1(n_67),
.B2(n_56),
.Y(n_110)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_78),
.Y(n_111)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_111),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_78),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_112),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_67),
.A2(n_8),
.B1(n_70),
.B2(n_64),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_58),
.Y(n_115)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_115),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_116),
.A2(n_94),
.B(n_101),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_65),
.A2(n_76),
.B1(n_57),
.B2(n_59),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_65),
.A2(n_76),
.B1(n_87),
.B2(n_59),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_58),
.A2(n_87),
.B1(n_85),
.B2(n_70),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_120),
.B(n_123),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_121),
.B(n_125),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_93),
.B(n_85),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_122),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_102),
.A2(n_71),
.B1(n_73),
.B2(n_63),
.Y(n_125)
);

A2O1A1Ixp33_ASAP7_75t_L g128 ( 
.A1(n_103),
.A2(n_68),
.B(n_91),
.C(n_63),
.Y(n_128)
);

AO21x1_ASAP7_75t_L g156 ( 
.A1(n_128),
.A2(n_129),
.B(n_131),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_110),
.A2(n_71),
.B1(n_68),
.B2(n_91),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_129),
.A2(n_111),
.B1(n_112),
.B2(n_127),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_131),
.A2(n_133),
.B(n_140),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_94),
.A2(n_101),
.B(n_100),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_106),
.Y(n_135)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_135),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_109),
.B(n_107),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_137),
.B(n_112),
.C(n_143),
.Y(n_152)
);

OAI32xp33_ASAP7_75t_L g138 ( 
.A1(n_98),
.A2(n_117),
.A3(n_106),
.B1(n_118),
.B2(n_97),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_138),
.B(n_139),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_98),
.B(n_101),
.Y(n_139)
);

AOI21xp33_ASAP7_75t_SL g140 ( 
.A1(n_108),
.A2(n_114),
.B(n_104),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_115),
.B(n_114),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_141),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_147),
.A2(n_125),
.B1(n_123),
.B2(n_121),
.Y(n_165)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_135),
.Y(n_148)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_148),
.Y(n_167)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_144),
.Y(n_149)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_149),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_144),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_151),
.B(n_153),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_152),
.B(n_138),
.Y(n_163)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_132),
.Y(n_153)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_132),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_155),
.B(n_158),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_156),
.A2(n_127),
.B(n_126),
.Y(n_169)
);

INVx13_ASAP7_75t_L g157 ( 
.A(n_128),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_157),
.Y(n_173)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_134),
.Y(n_158)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_134),
.Y(n_160)
);

OAI211xp5_ASAP7_75t_L g164 ( 
.A1(n_160),
.A2(n_159),
.B(n_161),
.C(n_143),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_163),
.B(n_166),
.C(n_156),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_164),
.B(n_170),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_165),
.A2(n_174),
.B(n_176),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_152),
.B(n_130),
.C(n_133),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_169),
.A2(n_172),
.B(n_147),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_150),
.A2(n_126),
.B1(n_127),
.B2(n_142),
.Y(n_170)
);

O2A1O1Ixp33_ASAP7_75t_L g172 ( 
.A1(n_157),
.A2(n_127),
.B(n_142),
.C(n_137),
.Y(n_172)
);

AOI322xp5_ASAP7_75t_L g174 ( 
.A1(n_157),
.A2(n_124),
.A3(n_127),
.B1(n_136),
.B2(n_159),
.C1(n_145),
.C2(n_154),
.Y(n_174)
);

OAI21xp33_ASAP7_75t_L g176 ( 
.A1(n_145),
.A2(n_162),
.B(n_154),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_163),
.B(n_162),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_178),
.B(n_180),
.C(n_187),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_170),
.B(n_151),
.Y(n_179)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_179),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_168),
.B(n_146),
.Y(n_181)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_181),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_166),
.B(n_156),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_183),
.B(n_172),
.Y(n_194)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_168),
.Y(n_184)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_184),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_173),
.A2(n_127),
.B(n_148),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_185),
.A2(n_175),
.B(n_167),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_186),
.A2(n_165),
.B(n_172),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_169),
.B(n_146),
.C(n_149),
.Y(n_187)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_190),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_192),
.B(n_187),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_194),
.B(n_178),
.C(n_175),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_189),
.A2(n_177),
.B1(n_186),
.B2(n_182),
.Y(n_195)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_195),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_196),
.B(n_200),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_191),
.A2(n_180),
.B1(n_183),
.B2(n_174),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_197),
.A2(n_194),
.B(n_188),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_198),
.B(n_188),
.C(n_190),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_193),
.A2(n_167),
.B1(n_171),
.B2(n_158),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_202),
.B(n_197),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_204),
.B(n_136),
.C(n_201),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_198),
.B(n_153),
.Y(n_205)
);

OAI221xp5_ASAP7_75t_L g207 ( 
.A1(n_205),
.A2(n_171),
.B1(n_160),
.B2(n_155),
.C(n_199),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_206),
.Y(n_210)
);

INVx11_ASAP7_75t_L g209 ( 
.A(n_207),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_210),
.B(n_203),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_211),
.A2(n_209),
.B(n_208),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_212),
.B(n_204),
.C(n_210),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_213),
.B(n_209),
.Y(n_214)
);


endmodule