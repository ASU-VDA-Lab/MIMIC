module fake_jpeg_1166_n_133 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_133);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_133;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_0),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_2),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

INVx6_ASAP7_75t_SL g49 ( 
.A(n_46),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_54),
.B(n_39),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_55),
.B(n_59),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_50),
.B(n_36),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_63),
.Y(n_65)
);

AO22x1_ASAP7_75t_SL g59 ( 
.A1(n_53),
.A2(n_44),
.B1(n_34),
.B2(n_36),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_40),
.Y(n_63)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_63),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_71),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_34),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_70),
.Y(n_84)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_38),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_74),
.Y(n_85)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

BUFx8_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_35),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_73),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_45),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_82),
.C(n_6),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_76),
.A2(n_54),
.B1(n_61),
.B2(n_47),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_79),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_SL g82 ( 
.A(n_67),
.B(n_37),
.C(n_42),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_76),
.B(n_44),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_86),
.B(n_87),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_62),
.Y(n_87)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_88),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_71),
.B(n_1),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_89),
.B(n_15),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_83),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_90),
.A2(n_95),
.B1(n_93),
.B2(n_103),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_91),
.B(n_96),
.Y(n_113)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_80),
.A2(n_4),
.B(n_5),
.Y(n_95)
);

NAND3xp33_ASAP7_75t_L g107 ( 
.A(n_95),
.B(n_97),
.C(n_98),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_78),
.B(n_6),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_77),
.Y(n_99)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_99),
.Y(n_112)
);

OA22x2_ASAP7_75t_L g100 ( 
.A1(n_87),
.A2(n_81),
.B1(n_84),
.B2(n_18),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_100),
.B(n_102),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_81),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_101),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_7),
.Y(n_102)
);

OAI21xp33_ASAP7_75t_SL g103 ( 
.A1(n_83),
.A2(n_16),
.B(n_27),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_13),
.Y(n_114)
);

XOR2x2_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_14),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_106),
.B(n_110),
.C(n_114),
.Y(n_120)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_109),
.Y(n_116)
);

MAJx2_ASAP7_75t_L g110 ( 
.A(n_100),
.B(n_98),
.C(n_19),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_100),
.Y(n_111)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_111),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_99),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_115),
.Y(n_118)
);

OA22x2_ASAP7_75t_L g119 ( 
.A1(n_108),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_119),
.B(n_104),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_20),
.C(n_26),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_121),
.B(n_104),
.C(n_113),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_122),
.A2(n_123),
.B(n_124),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_119),
.B(n_113),
.Y(n_124)
);

BUFx24_ASAP7_75t_SL g125 ( 
.A(n_118),
.Y(n_125)
);

OA21x2_ASAP7_75t_SL g126 ( 
.A1(n_125),
.A2(n_117),
.B(n_112),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_126),
.B(n_107),
.Y(n_128)
);

NOR2xp67_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_120),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_129),
.A2(n_127),
.B(n_116),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_10),
.C(n_12),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_24),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_33),
.Y(n_133)
);


endmodule