module fake_jpeg_8402_n_174 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_174);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_174;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_152;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

OR2x2_ASAP7_75t_L g29 ( 
.A(n_3),
.B(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_0),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_33),
.B(n_44),
.Y(n_61)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_34),
.B(n_35),
.Y(n_52)
);

INVx6_ASAP7_75t_SL g35 ( 
.A(n_17),
.Y(n_35)
);

HB1xp67_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_40),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_0),
.Y(n_38)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_41),
.Y(n_47)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_39),
.B(n_30),
.Y(n_66)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_0),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_15),
.A2(n_23),
.B1(n_16),
.B2(n_22),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_32),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_21),
.B(n_1),
.Y(n_43)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_20),
.B(n_2),
.Y(n_44)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_46),
.B(n_37),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_48),
.B(n_67),
.Y(n_75)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_49),
.Y(n_70)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_50),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_45),
.A2(n_15),
.B1(n_23),
.B2(n_28),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_51),
.A2(n_56),
.B1(n_60),
.B2(n_20),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_33),
.A2(n_38),
.B1(n_41),
.B2(n_31),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_18),
.Y(n_59)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_34),
.A2(n_28),
.B1(n_19),
.B2(n_22),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_18),
.Y(n_63)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_27),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_64),
.B(n_4),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_66),
.B(n_27),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_42),
.B(n_19),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_68),
.Y(n_97)
);

NOR2x1_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_34),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_69),
.B(n_79),
.Y(n_101)
);

O2A1O1Ixp33_ASAP7_75t_SL g71 ( 
.A1(n_64),
.A2(n_48),
.B(n_67),
.C(n_61),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_71),
.A2(n_77),
.B1(n_81),
.B2(n_82),
.Y(n_102)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_80),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_65),
.A2(n_43),
.B(n_30),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_76),
.A2(n_79),
.B(n_88),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_65),
.A2(n_26),
.B1(n_31),
.B2(n_24),
.Y(n_77)
);

OAI21x1_ASAP7_75t_L g79 ( 
.A1(n_47),
.A2(n_32),
.B(n_21),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_49),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_61),
.A2(n_25),
.B1(n_27),
.B2(n_37),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_58),
.B(n_21),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_84),
.B(n_90),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_85),
.B(n_52),
.Y(n_108)
);

AND2x6_ASAP7_75t_L g87 ( 
.A(n_57),
.B(n_3),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_12),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_4),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_50),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_L g106 ( 
.A1(n_91),
.A2(n_55),
.B1(n_46),
.B2(n_8),
.Y(n_106)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_98),
.Y(n_117)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_69),
.Y(n_99)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_99),
.Y(n_119)
);

NOR3xp33_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_107),
.C(n_108),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_105),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_53),
.Y(n_103)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_103),
.Y(n_125)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_78),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_104),
.Y(n_114)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_69),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_106),
.A2(n_110),
.B1(n_70),
.B2(n_83),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_76),
.B(n_53),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_6),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_109),
.Y(n_121)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_97),
.A2(n_75),
.B1(n_71),
.B2(n_68),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_111),
.A2(n_122),
.B1(n_127),
.B2(n_103),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_115),
.Y(n_128)
);

MAJx2_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_75),
.C(n_71),
.Y(n_113)
);

XOR2x1_ASAP7_75t_L g138 ( 
.A(n_113),
.B(n_120),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_97),
.B(n_75),
.C(n_89),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_102),
.B(n_88),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_123),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_102),
.B(n_88),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_98),
.A2(n_87),
.B1(n_70),
.B2(n_86),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_107),
.B(n_89),
.C(n_86),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_110),
.A2(n_83),
.B1(n_54),
.B2(n_78),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_122),
.A2(n_100),
.B1(n_105),
.B2(n_99),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_129),
.A2(n_130),
.B1(n_126),
.B2(n_113),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_117),
.A2(n_96),
.B1(n_93),
.B2(n_101),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_127),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_131),
.B(n_132),
.Y(n_143)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_123),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_124),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_133),
.B(n_135),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_SL g150 ( 
.A(n_134),
.B(n_136),
.C(n_101),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_125),
.B(n_94),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_124),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_119),
.B(n_94),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_139),
.A2(n_121),
.B(n_109),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_116),
.B(n_95),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_140),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_138),
.B(n_115),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_141),
.B(n_144),
.C(n_134),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_142),
.A2(n_147),
.B1(n_150),
.B2(n_130),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_138),
.B(n_111),
.C(n_120),
.Y(n_144)
);

INVx13_ASAP7_75t_L g146 ( 
.A(n_135),
.Y(n_146)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_146),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_132),
.A2(n_131),
.B1(n_133),
.B2(n_136),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_149),
.A2(n_139),
.B(n_92),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_144),
.B(n_137),
.C(n_128),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_151),
.B(n_152),
.C(n_153),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_142),
.B(n_118),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_154),
.A2(n_156),
.B(n_148),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_141),
.B(n_129),
.C(n_108),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_155),
.B(n_157),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_150),
.B(n_92),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_158),
.B(n_148),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_159),
.B(n_160),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_157),
.A2(n_143),
.B1(n_147),
.B2(n_146),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_162),
.A2(n_149),
.B(n_155),
.Y(n_164)
);

OAI21x1_ASAP7_75t_SL g169 ( 
.A1(n_164),
.A2(n_165),
.B(n_114),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_161),
.A2(n_145),
.B1(n_153),
.B2(n_104),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_163),
.B(n_72),
.Y(n_167)
);

AOI322xp5_ASAP7_75t_L g168 ( 
.A1(n_167),
.A2(n_145),
.A3(n_163),
.B1(n_72),
.B2(n_73),
.C1(n_114),
.C2(n_54),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_168),
.B(n_170),
.C(n_10),
.Y(n_172)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_169),
.Y(n_171)
);

AOI322xp5_ASAP7_75t_L g170 ( 
.A1(n_166),
.A2(n_73),
.A3(n_10),
.B1(n_13),
.B2(n_62),
.C1(n_8),
.C2(n_7),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_13),
.C(n_6),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_173),
.B(n_171),
.Y(n_174)
);


endmodule