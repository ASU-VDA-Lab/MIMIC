module fake_ariane_1675_n_101 (n_8, n_3, n_2, n_11, n_7, n_5, n_14, n_1, n_0, n_12, n_15, n_6, n_13, n_9, n_4, n_10, n_101);

input n_8;
input n_3;
input n_2;
input n_11;
input n_7;
input n_5;
input n_14;
input n_1;
input n_0;
input n_12;
input n_15;
input n_6;
input n_13;
input n_9;
input n_4;
input n_10;

output n_101;

wire n_83;
wire n_56;
wire n_60;
wire n_64;
wire n_90;
wire n_38;
wire n_47;
wire n_18;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_34;
wire n_69;
wire n_95;
wire n_92;
wire n_98;
wire n_74;
wire n_33;
wire n_19;
wire n_40;
wire n_53;
wire n_21;
wire n_66;
wire n_71;
wire n_24;
wire n_96;
wire n_49;
wire n_20;
wire n_100;
wire n_17;
wire n_50;
wire n_62;
wire n_51;
wire n_76;
wire n_79;
wire n_26;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_72;
wire n_44;
wire n_30;
wire n_82;
wire n_31;
wire n_42;
wire n_57;
wire n_70;
wire n_85;
wire n_48;
wire n_94;
wire n_32;
wire n_37;
wire n_58;
wire n_65;
wire n_45;
wire n_52;
wire n_73;
wire n_77;
wire n_93;
wire n_23;
wire n_61;
wire n_22;
wire n_81;
wire n_87;
wire n_43;
wire n_27;
wire n_29;
wire n_41;
wire n_55;
wire n_28;
wire n_80;
wire n_97;
wire n_88;
wire n_68;
wire n_78;
wire n_39;
wire n_59;
wire n_63;
wire n_99;
wire n_16;
wire n_35;
wire n_54;
wire n_25;

CKINVDCx5p33_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVxp67_ASAP7_75t_SL g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVxp67_ASAP7_75t_SL g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx5p33_ASAP7_75t_R g25 ( 
.A(n_15),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx5p33_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_19),
.B(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

AND2x4_ASAP7_75t_L g32 ( 
.A(n_28),
.B(n_3),
.Y(n_32)
);

AND2x4_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_4),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_41),
.B(n_27),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_41),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_41),
.B(n_27),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g50 ( 
.A(n_41),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

NOR3xp33_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_26),
.C(n_30),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_L g53 ( 
.A1(n_45),
.A2(n_30),
.B1(n_16),
.B2(n_33),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_46),
.A2(n_32),
.B1(n_33),
.B2(n_48),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_42),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_36),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_56),
.B(n_44),
.Y(n_58)
);

AOI221xp5_ASAP7_75t_L g59 ( 
.A1(n_53),
.A2(n_32),
.B1(n_16),
.B2(n_52),
.C(n_54),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_57),
.A2(n_44),
.B(n_50),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_36),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_61),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_61),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_62),
.B(n_59),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_63),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_65),
.A2(n_49),
.B1(n_48),
.B2(n_46),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_70),
.B(n_65),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g73 ( 
.A(n_69),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_71),
.B(n_64),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

AND2x4_ASAP7_75t_L g77 ( 
.A(n_72),
.B(n_73),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_75),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_74),
.B(n_67),
.Y(n_79)
);

INVxp33_ASAP7_75t_L g80 ( 
.A(n_75),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_79),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_79),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_77),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_76),
.B(n_73),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_81),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_83),
.B(n_77),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_84),
.Y(n_87)
);

NOR2x1p5_ASAP7_75t_L g88 ( 
.A(n_85),
.B(n_82),
.Y(n_88)
);

NAND3xp33_ASAP7_75t_L g89 ( 
.A(n_87),
.B(n_78),
.C(n_37),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_89),
.A2(n_80),
.B1(n_78),
.B2(n_77),
.Y(n_90)
);

AOI21xp33_ASAP7_75t_L g91 ( 
.A1(n_88),
.A2(n_86),
.B(n_39),
.Y(n_91)
);

NOR2x1_ASAP7_75t_L g92 ( 
.A(n_88),
.B(n_39),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_92),
.A2(n_38),
.B1(n_66),
.B2(n_25),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_93),
.B(n_91),
.Y(n_94)
);

AOI221xp5_ASAP7_75t_L g95 ( 
.A1(n_93),
.A2(n_90),
.B1(n_23),
.B2(n_21),
.C(n_43),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_94),
.B(n_4),
.Y(n_96)
);

XNOR2x1_ASAP7_75t_L g97 ( 
.A(n_95),
.B(n_5),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_96),
.A2(n_6),
.B1(n_66),
.B2(n_67),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_L g99 ( 
.A1(n_98),
.A2(n_97),
.B1(n_71),
.B2(n_9),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_99),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_100),
.A2(n_7),
.B(n_8),
.Y(n_101)
);


endmodule