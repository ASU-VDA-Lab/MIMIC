module fake_jpeg_22813_n_268 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_268);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_268;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx3_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx4f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

CKINVDCx6p67_ASAP7_75t_R g47 ( 
.A(n_34),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_17),
.B(n_8),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_40),
.Y(n_43)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_17),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_36),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_44),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_34),
.A2(n_22),
.B1(n_28),
.B2(n_26),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_42),
.A2(n_50),
.B1(n_34),
.B2(n_37),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_22),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_39),
.A2(n_31),
.B1(n_24),
.B2(n_18),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_49),
.A2(n_18),
.B1(n_24),
.B2(n_22),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_34),
.A2(n_16),
.B1(n_26),
.B2(n_28),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_24),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_53),
.B(n_40),
.Y(n_63)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_40),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_33),
.B(n_31),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_57),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_33),
.B(n_31),
.Y(n_57)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_59),
.B(n_61),
.Y(n_91)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_56),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_60),
.B(n_71),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_62),
.B(n_44),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_63),
.B(n_66),
.Y(n_102)
);

AO22x1_ASAP7_75t_L g64 ( 
.A1(n_47),
.A2(n_36),
.B1(n_33),
.B2(n_35),
.Y(n_64)
);

AND2x4_ASAP7_75t_SL g93 ( 
.A(n_64),
.B(n_33),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx13_ASAP7_75t_L g99 ( 
.A(n_68),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_53),
.Y(n_69)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_70),
.B(n_72),
.Y(n_90)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_43),
.B(n_35),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_47),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_73),
.B(n_76),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_54),
.A2(n_39),
.B1(n_36),
.B2(n_28),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_74),
.A2(n_80),
.B1(n_83),
.B2(n_42),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_40),
.Y(n_75)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_49),
.B(n_18),
.Y(n_77)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_41),
.B(n_52),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_85),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVx13_ASAP7_75t_L g109 ( 
.A(n_79),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_44),
.A2(n_19),
.B1(n_23),
.B2(n_16),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_51),
.B(n_32),
.Y(n_81)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_55),
.A2(n_26),
.B1(n_39),
.B2(n_30),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_50),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_84),
.B(n_44),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_52),
.B(n_29),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_55),
.B(n_32),
.Y(n_86)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_92),
.A2(n_97),
.B1(n_39),
.B2(n_46),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_64),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_66),
.B(n_41),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_98),
.Y(n_120)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_103),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_65),
.B(n_41),
.Y(n_98)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_61),
.Y(n_103)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_64),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_105),
.B(n_108),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_107),
.B(n_35),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_85),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_69),
.B(n_20),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_110),
.B(n_113),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_72),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_111),
.B(n_60),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_77),
.B(n_20),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_114),
.A2(n_135),
.B(n_138),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_90),
.A2(n_78),
.B1(n_58),
.B2(n_62),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_115),
.A2(n_131),
.B1(n_92),
.B2(n_97),
.Y(n_156)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_101),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_117),
.B(n_118),
.Y(n_161)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_87),
.Y(n_118)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_121),
.Y(n_157)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_99),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_122),
.B(n_128),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_71),
.C(n_58),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_123),
.B(n_124),
.C(n_125),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_94),
.B(n_65),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_94),
.B(n_65),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_103),
.B(n_82),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g149 ( 
.A(n_126),
.Y(n_149)
);

OAI22xp33_ASAP7_75t_L g127 ( 
.A1(n_93),
.A2(n_46),
.B1(n_70),
.B2(n_73),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_127),
.A2(n_134),
.B1(n_139),
.B2(n_109),
.Y(n_168)
);

NOR3xp33_ASAP7_75t_SL g128 ( 
.A(n_108),
.B(n_58),
.C(n_63),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_89),
.B(n_76),
.Y(n_129)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_129),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_90),
.A2(n_42),
.B1(n_46),
.B2(n_80),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_91),
.Y(n_132)
);

BUFx24_ASAP7_75t_L g154 ( 
.A(n_132),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_111),
.B(n_67),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_133),
.B(n_88),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_93),
.Y(n_136)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_136),
.Y(n_142)
);

OAI21xp33_ASAP7_75t_L g137 ( 
.A1(n_100),
.A2(n_14),
.B(n_1),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_137),
.A2(n_102),
.B(n_88),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_93),
.B(n_35),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_100),
.A2(n_59),
.B1(n_33),
.B2(n_35),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_87),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_140),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_89),
.B(n_106),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_141),
.Y(n_158)
);

NOR2x1_ASAP7_75t_L g144 ( 
.A(n_128),
.B(n_113),
.Y(n_144)
);

NOR2x1_ASAP7_75t_L g175 ( 
.A(n_144),
.B(n_25),
.Y(n_175)
);

XNOR2x1_ASAP7_75t_L g145 ( 
.A(n_115),
.B(n_95),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_145),
.B(n_151),
.Y(n_181)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_147),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_136),
.A2(n_120),
.B(n_119),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_148),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_150),
.A2(n_117),
.B1(n_104),
.B2(n_30),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_120),
.A2(n_133),
.B(n_107),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_130),
.A2(n_102),
.B(n_95),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_152),
.B(n_159),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_134),
.A2(n_127),
.B1(n_105),
.B2(n_114),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_153),
.A2(n_160),
.B1(n_168),
.B2(n_139),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_156),
.A2(n_163),
.B1(n_167),
.B2(n_109),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_130),
.A2(n_113),
.B(n_97),
.Y(n_159)
);

AO22x1_ASAP7_75t_SL g160 ( 
.A1(n_114),
.A2(n_110),
.B1(n_48),
.B2(n_68),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_123),
.B(n_106),
.C(n_112),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_162),
.B(n_68),
.C(n_29),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_131),
.A2(n_138),
.B1(n_140),
.B2(n_118),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_116),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_165),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_124),
.B(n_110),
.Y(n_166)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_166),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_138),
.A2(n_96),
.B1(n_112),
.B2(n_109),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_125),
.B(n_104),
.Y(n_169)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_169),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_171),
.A2(n_172),
.B1(n_186),
.B2(n_187),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_175),
.A2(n_190),
.B(n_150),
.Y(n_198)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_161),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_176),
.B(n_182),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_177),
.B(n_191),
.C(n_162),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_142),
.B(n_160),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_178),
.A2(n_148),
.B(n_146),
.Y(n_194)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_147),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_158),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g203 ( 
.A(n_183),
.Y(n_203)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_154),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_184),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_185),
.A2(n_153),
.B1(n_160),
.B2(n_144),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_143),
.B(n_25),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_157),
.B(n_10),
.Y(n_187)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_154),
.Y(n_189)
);

NAND4xp25_ASAP7_75t_SL g204 ( 
.A(n_189),
.B(n_154),
.C(n_149),
.D(n_170),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_152),
.B(n_48),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_155),
.B(n_79),
.C(n_21),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_157),
.B(n_9),
.Y(n_193)
);

AOI322xp5_ASAP7_75t_L g210 ( 
.A1(n_193),
.A2(n_9),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.C1(n_4),
.C2(n_5),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_194),
.A2(n_179),
.B(n_190),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_172),
.A2(n_163),
.B1(n_156),
.B2(n_145),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_195),
.A2(n_206),
.B1(n_174),
.B2(n_178),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_196),
.Y(n_220)
);

NOR3xp33_ASAP7_75t_SL g226 ( 
.A(n_198),
.B(n_175),
.C(n_178),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_181),
.B(n_164),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_199),
.B(n_200),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_181),
.B(n_155),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_201),
.B(n_207),
.C(n_209),
.Y(n_214)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_204),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_185),
.A2(n_151),
.B1(n_146),
.B2(n_166),
.Y(n_205)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_205),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_179),
.A2(n_167),
.B1(n_169),
.B2(n_170),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_191),
.B(n_159),
.C(n_79),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_180),
.B(n_21),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_208),
.B(n_177),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_192),
.B(n_21),
.C(n_0),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_210),
.B(n_171),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_212),
.B(n_213),
.Y(n_239)
);

BUFx12_ASAP7_75t_L g213 ( 
.A(n_204),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_215),
.B(n_221),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_218),
.B(n_206),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_200),
.B(n_201),
.C(n_207),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_219),
.B(n_194),
.C(n_199),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_205),
.B(n_192),
.Y(n_221)
);

BUFx12f_ASAP7_75t_SL g222 ( 
.A(n_198),
.Y(n_222)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_222),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_197),
.Y(n_223)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_223),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_203),
.B(n_173),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_224),
.B(n_184),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_228),
.B(n_230),
.C(n_231),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_229),
.Y(n_248)
);

AOI322xp5_ASAP7_75t_L g231 ( 
.A1(n_222),
.A2(n_202),
.A3(n_227),
.B1(n_226),
.B2(n_220),
.C1(n_214),
.C2(n_195),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_219),
.B(n_196),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_232),
.B(n_238),
.Y(n_247)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_216),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_235),
.B(n_0),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_214),
.B(n_174),
.C(n_188),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_236),
.A2(n_238),
.B(n_213),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_217),
.B(n_188),
.C(n_209),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_237),
.B(n_221),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_233),
.A2(n_225),
.B(n_211),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_241),
.A2(n_234),
.B(n_2),
.Y(n_254)
);

AND2x6_ASAP7_75t_L g242 ( 
.A(n_237),
.B(n_213),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_243),
.B(n_247),
.C(n_230),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_236),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_244),
.B(n_249),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_245),
.B(n_248),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_239),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_250),
.B(n_252),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_251),
.B(n_255),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_246),
.B(n_232),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_254),
.A2(n_11),
.B(n_12),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_240),
.B(n_21),
.Y(n_255)
);

OAI21x1_ASAP7_75t_L g256 ( 
.A1(n_242),
.A2(n_1),
.B(n_3),
.Y(n_256)
);

NAND4xp25_ASAP7_75t_SL g257 ( 
.A(n_253),
.B(n_5),
.C(n_7),
.D(n_9),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_257),
.B(n_259),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_260),
.A2(n_253),
.B(n_13),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_261),
.A2(n_263),
.B(n_12),
.Y(n_265)
);

AOI322xp5_ASAP7_75t_L g263 ( 
.A1(n_258),
.A2(n_12),
.A3(n_13),
.B1(n_14),
.B2(n_15),
.C1(n_242),
.C2(n_256),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_262),
.Y(n_264)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_264),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_266),
.B(n_265),
.Y(n_267)
);

BUFx24_ASAP7_75t_SL g268 ( 
.A(n_267),
.Y(n_268)
);


endmodule