module fake_jpeg_22189_n_79 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_79);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_79;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

INVx1_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_3),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx14_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_15),
.B(n_0),
.Y(n_21)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_25),
.A2(n_22),
.B1(n_19),
.B2(n_13),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_30),
.B(n_33),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_24),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_31),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_21),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_34),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_28),
.Y(n_33)
);

XNOR2xp5_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_23),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_21),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_36),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_17),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_26),
.A2(n_20),
.B1(n_12),
.B2(n_11),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_37),
.B(n_29),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_39),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_37),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_28),
.Y(n_42)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_44),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_15),
.Y(n_45)
);

XOR2xp5_ASAP7_75t_L g49 ( 
.A(n_45),
.B(n_32),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_1),
.Y(n_62)
);

XOR2xp5_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_35),
.Y(n_50)
);

XOR2xp5_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_40),
.Y(n_57)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_51),
.B(n_53),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_43),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_52),
.B(n_55),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_29),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_46),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_60),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_48),
.A2(n_26),
.B1(n_45),
.B2(n_16),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_59),
.A2(n_9),
.B1(n_13),
.B2(n_10),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_16),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_51),
.A2(n_9),
.B1(n_12),
.B2(n_11),
.Y(n_61)
);

OAI21xp33_ASAP7_75t_SL g64 ( 
.A1(n_61),
.A2(n_62),
.B(n_53),
.Y(n_64)
);

NOR3xp33_ASAP7_75t_SL g63 ( 
.A(n_58),
.B(n_49),
.C(n_47),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_63),
.B(n_65),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_64),
.A2(n_67),
.B1(n_10),
.B2(n_65),
.Y(n_68)
);

INVxp67_ASAP7_75t_SL g65 ( 
.A(n_56),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_68),
.B(n_70),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_66),
.B(n_57),
.C(n_50),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g71 ( 
.A1(n_69),
.A2(n_62),
.B(n_6),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_71),
.B(n_72),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_69),
.A2(n_4),
.B(n_5),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_4),
.C(n_5),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_74),
.A2(n_75),
.B(n_7),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_76),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_77),
.A2(n_8),
.B1(n_2),
.B2(n_3),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_78),
.B(n_8),
.Y(n_79)
);


endmodule