module fake_jpeg_31757_n_108 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_29, n_12, n_8, n_15, n_7, n_108);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_108;

wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_29),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_9),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_7),
.B(n_3),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_6),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_22),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_41),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_46),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_37),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_36),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_50),
.Y(n_57)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_43),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_51),
.Y(n_54)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_46),
.B(n_42),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_0),
.Y(n_75)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_57),
.B(n_39),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_63),
.B(n_70),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_35),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_67),
.Y(n_76)
);

AND2x6_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_34),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_69),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_34),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_54),
.A2(n_0),
.B(n_1),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_68),
.A2(n_14),
.B(n_16),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_59),
.A2(n_32),
.B1(n_40),
.B2(n_2),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_40),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_75),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_L g74 ( 
.A1(n_56),
.A2(n_32),
.B1(n_1),
.B2(n_2),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_74),
.A2(n_4),
.B1(n_11),
.B2(n_13),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_77),
.A2(n_89),
.B1(n_19),
.B2(n_20),
.Y(n_90)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_4),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_81),
.B(n_84),
.Y(n_91)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_82),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_72),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_85),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_86),
.B(n_87),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_63),
.B(n_17),
.C(n_18),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_90),
.Y(n_97)
);

NAND3xp33_ASAP7_75t_L g98 ( 
.A(n_93),
.B(n_78),
.C(n_83),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_98),
.B(n_99),
.Y(n_100)
);

AOI22x1_ASAP7_75t_L g99 ( 
.A1(n_95),
.A2(n_88),
.B1(n_89),
.B2(n_83),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_97),
.B(n_96),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_100),
.C(n_93),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_102),
.B(n_76),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_103),
.B(n_92),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_104),
.A2(n_91),
.B(n_94),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_105),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_106),
.A2(n_21),
.B(n_23),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_24),
.Y(n_108)
);


endmodule