module fake_jpeg_17257_n_79 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_79);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_79;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_44;
wire n_24;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_48;
wire n_35;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

AND2x2_ASAP7_75t_L g20 ( 
.A(n_1),
.B(n_9),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_2),
.B(n_8),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx24_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_6),
.B(n_11),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_10),
.B(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

OA22x2_ASAP7_75t_L g39 ( 
.A1(n_25),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_39),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_34),
.A2(n_3),
.B1(n_5),
.B2(n_10),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_40),
.A2(n_49),
.B1(n_50),
.B2(n_51),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_20),
.B(n_11),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_43),
.Y(n_58)
);

HB1xp67_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_46),
.A2(n_47),
.B(n_48),
.Y(n_57)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_26),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_20),
.B(n_12),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_34),
.A2(n_13),
.B1(n_15),
.B2(n_38),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_21),
.A2(n_27),
.B1(n_29),
.B2(n_37),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_57),
.B(n_51),
.C(n_23),
.Y(n_62)
);

XOR2xp5_ASAP7_75t_L g69 ( 
.A(n_62),
.B(n_63),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_61),
.C(n_59),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_35),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_64),
.B(n_65),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_55),
.B(n_36),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_28),
.C(n_24),
.Y(n_66)
);

NOR3xp33_ASAP7_75t_SL g68 ( 
.A(n_66),
.B(n_28),
.C(n_39),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_68),
.Y(n_72)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_70),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_69),
.A2(n_53),
.B1(n_54),
.B2(n_40),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_71),
.B(n_69),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_67),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_74),
.B(n_75),
.Y(n_76)
);

AOI322xp5_ASAP7_75t_L g77 ( 
.A1(n_76),
.A2(n_73),
.A3(n_72),
.B1(n_71),
.B2(n_68),
.C1(n_39),
.C2(n_56),
.Y(n_77)
);

OAI221xp5_ASAP7_75t_SL g78 ( 
.A1(n_77),
.A2(n_45),
.B1(n_29),
.B2(n_27),
.C(n_60),
.Y(n_78)
);

A2O1A1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_78),
.A2(n_60),
.B(n_30),
.C(n_32),
.Y(n_79)
);


endmodule