module fake_jpeg_26888_n_59 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_59);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_59;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_47;
wire n_22;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVx8_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_5),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_4),
.B(n_3),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

BUFx3_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx10_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g17 ( 
.A(n_10),
.B(n_0),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_17),
.B(n_18),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_10),
.B(n_0),
.Y(n_18)
);

AOI21xp33_ASAP7_75t_SL g19 ( 
.A1(n_15),
.A2(n_0),
.B(n_1),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_19),
.B(n_20),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_13),
.B(n_2),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_21),
.B(n_16),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_20),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_25),
.B(n_18),
.Y(n_27)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_SL g34 ( 
.A1(n_27),
.A2(n_29),
.B(n_30),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_23),
.A2(n_19),
.B1(n_17),
.B2(n_8),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_28),
.A2(n_8),
.B1(n_11),
.B2(n_14),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_22),
.B(n_9),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

NOR2x1_ASAP7_75t_L g31 ( 
.A(n_22),
.B(n_9),
.Y(n_31)
);

AOI21xp5_ASAP7_75t_L g33 ( 
.A1(n_31),
.A2(n_25),
.B(n_14),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_36),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_SL g41 ( 
.A1(n_33),
.A2(n_37),
.B(n_12),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_31),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_28),
.A2(n_2),
.B(n_11),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_15),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_35),
.A2(n_21),
.B1(n_24),
.B2(n_8),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_39),
.B(n_40),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_38),
.A2(n_24),
.B1(n_34),
.B2(n_32),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g45 ( 
.A1(n_41),
.A2(n_12),
.B(n_13),
.Y(n_45)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_44),
.B(n_13),
.C(n_15),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_45),
.B(n_40),
.Y(n_51)
);

XOR2xp5_ASAP7_75t_L g49 ( 
.A(n_46),
.B(n_39),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_50),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_48),
.B(n_42),
.Y(n_50)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_51),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g54 ( 
.A1(n_52),
.A2(n_47),
.B(n_44),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_54),
.A2(n_55),
.B(n_6),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_52),
.B(n_4),
.Y(n_55)
);

NAND3xp33_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_6),
.C(n_2),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_57),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_53),
.Y(n_59)
);


endmodule