module real_jpeg_5627_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_507;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_17;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_1),
.A2(n_184),
.B1(n_186),
.B2(n_187),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_1),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_1),
.A2(n_186),
.B1(n_248),
.B2(n_249),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g402 ( 
.A1(n_1),
.A2(n_186),
.B1(n_403),
.B2(n_405),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g457 ( 
.A1(n_1),
.A2(n_186),
.B1(n_458),
.B2(n_463),
.Y(n_457)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_2),
.Y(n_66)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_2),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_3),
.A2(n_34),
.B1(n_36),
.B2(n_39),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_3),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_3),
.A2(n_39),
.B1(n_85),
.B2(n_101),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_3),
.A2(n_39),
.B1(n_45),
.B2(n_148),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_3),
.A2(n_39),
.B1(n_228),
.B2(n_229),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_4),
.B(n_267),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_4),
.A2(n_266),
.B(n_316),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_4),
.B(n_191),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_4),
.B(n_36),
.C(n_376),
.Y(n_375)
);

OAI22xp33_ASAP7_75t_L g379 ( 
.A1(n_4),
.A2(n_380),
.B1(n_381),
.B2(n_383),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_4),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_4),
.B(n_137),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_4),
.A2(n_25),
.B1(n_424),
.B2(n_427),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_5),
.A2(n_257),
.B1(n_283),
.B2(n_285),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_5),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_5),
.A2(n_285),
.B1(n_347),
.B2(n_348),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_5),
.A2(n_285),
.B1(n_387),
.B2(n_390),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_5),
.A2(n_285),
.B1(n_408),
.B2(n_425),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_6),
.A2(n_288),
.B1(n_290),
.B2(n_291),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_6),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_6),
.A2(n_290),
.B1(n_321),
.B2(n_325),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_6),
.A2(n_290),
.B1(n_398),
.B2(n_399),
.Y(n_397)
);

AOI22xp33_ASAP7_75t_L g413 ( 
.A1(n_6),
.A2(n_159),
.B1(n_290),
.B2(n_414),
.Y(n_413)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_7),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_8),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_8),
.Y(n_306)
);

INVx8_ASAP7_75t_L g341 ( 
.A(n_8),
.Y(n_341)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_8),
.Y(n_429)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_9),
.A2(n_73),
.B1(n_76),
.B2(n_77),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_9),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_9),
.A2(n_76),
.B1(n_104),
.B2(n_107),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_9),
.A2(n_76),
.B1(n_159),
.B2(n_164),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_9),
.A2(n_76),
.B1(n_117),
.B2(n_196),
.Y(n_195)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_10),
.Y(n_87)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_10),
.Y(n_92)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_10),
.Y(n_97)
);

BUFx5_ASAP7_75t_L g99 ( 
.A(n_10),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_10),
.Y(n_261)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_11),
.Y(n_96)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_12),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_12),
.Y(n_89)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_12),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_12),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_12),
.Y(n_185)
);

BUFx5_ASAP7_75t_L g189 ( 
.A(n_12),
.Y(n_189)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_12),
.Y(n_210)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_12),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_12),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_13),
.A2(n_43),
.B1(n_44),
.B2(n_50),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_13),
.A2(n_43),
.B1(n_139),
.B2(n_143),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_13),
.A2(n_43),
.B1(n_236),
.B2(n_238),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_13),
.A2(n_43),
.B1(n_277),
.B2(n_280),
.Y(n_276)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_14),
.Y(n_58)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_14),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_14),
.Y(n_64)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_14),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_15),
.A2(n_114),
.B1(n_116),
.B2(n_117),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_15),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_15),
.A2(n_116),
.B1(n_176),
.B2(n_178),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_15),
.A2(n_116),
.B1(n_188),
.B2(n_209),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_15),
.A2(n_116),
.B1(n_160),
.B2(n_272),
.Y(n_271)
);

MAJx2_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_507),
.C(n_511),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_505),
.B(n_509),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_495),
.B(n_504),
.Y(n_18)
);

OAI31xp33_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_215),
.A3(n_240),
.B(n_492),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_197),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_21),
.B(n_197),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_110),
.C(n_153),
.Y(n_21)
);

FAx1_ASAP7_75t_L g366 ( 
.A(n_22),
.B(n_110),
.CI(n_153),
.CON(n_366),
.SN(n_366)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_79),
.Y(n_22)
);

AOI21xp33_ASAP7_75t_L g214 ( 
.A1(n_23),
.A2(n_24),
.B(n_81),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_40),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_24),
.A2(n_80),
.B1(n_81),
.B2(n_109),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_24),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_24),
.A2(n_40),
.B1(n_80),
.B2(n_358),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_31),
.B(n_33),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_25),
.B(n_158),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_25),
.A2(n_270),
.B1(n_275),
.B2(n_276),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_25),
.A2(n_276),
.B(n_305),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g401 ( 
.A1(n_25),
.A2(n_167),
.B(n_402),
.Y(n_401)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_25),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_25),
.A2(n_413),
.B1(n_424),
.B2(n_427),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_L g452 ( 
.A1(n_25),
.A2(n_33),
.B(n_305),
.Y(n_452)
);

OR2x2_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_29),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_28),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_30),
.Y(n_418)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_33),
.Y(n_168)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_37),
.A2(n_64),
.B1(n_65),
.B2(n_67),
.Y(n_63)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_40),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_53),
.B(n_69),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_42),
.A2(n_54),
.B1(n_70),
.B2(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx3_ASAP7_75t_L g389 ( 
.A(n_47),
.Y(n_389)
);

INVx6_ASAP7_75t_L g446 ( 
.A(n_47),
.Y(n_446)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_48),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_48),
.Y(n_462)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_49),
.Y(n_180)
);

BUFx5_ASAP7_75t_L g382 ( 
.A(n_49),
.Y(n_382)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_49),
.Y(n_385)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

OA22x2_ASAP7_75t_L g119 ( 
.A1(n_52),
.A2(n_120),
.B1(n_122),
.B2(n_125),
.Y(n_119)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_52),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_53),
.B(n_151),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_53),
.A2(n_71),
.B(n_147),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_53),
.A2(n_71),
.B1(n_151),
.B2(n_175),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_53),
.A2(n_69),
.B(n_147),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g475 ( 
.A1(n_53),
.A2(n_476),
.B(n_477),
.Y(n_475)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_54),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_54),
.A2(n_70),
.B1(n_379),
.B2(n_386),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_54),
.A2(n_70),
.B1(n_386),
.B2(n_397),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_54),
.A2(n_70),
.B1(n_397),
.B2(n_457),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_63),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_57),
.B1(n_59),
.B2(n_62),
.Y(n_55)
);

INVx5_ASAP7_75t_L g374 ( 
.A(n_56),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_62),
.Y(n_391)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g280 ( 
.A(n_66),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_66),
.Y(n_404)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_66),
.Y(n_408)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_68),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_72),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_71),
.B(n_147),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_71),
.B(n_380),
.Y(n_422)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_72),
.Y(n_151)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g398 ( 
.A(n_75),
.Y(n_398)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_78),
.Y(n_177)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_81),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_100),
.B(n_102),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_82),
.B(n_212),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_82),
.A2(n_191),
.B1(n_234),
.B2(n_235),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_82),
.A2(n_191),
.B1(n_282),
.B2(n_286),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g511 ( 
.A1(n_82),
.A2(n_100),
.B(n_191),
.Y(n_511)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_83),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_83),
.A2(n_183),
.B(n_190),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_83),
.A2(n_108),
.B1(n_183),
.B2(n_287),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_83),
.A2(n_108),
.B1(n_315),
.B2(n_318),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g500 ( 
.A1(n_83),
.A2(n_501),
.B(n_502),
.Y(n_500)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_93),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_86),
.B1(n_88),
.B2(n_90),
.Y(n_84)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_92),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_93),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_97),
.B1(n_98),
.B2(n_99),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_95),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_95),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_95),
.Y(n_256)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_96),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_96),
.Y(n_142)
);

BUFx5_ASAP7_75t_L g232 ( 
.A(n_96),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_96),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_100),
.B(n_191),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g502 ( 
.A(n_102),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_108),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_103),
.Y(n_212)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_105),
.Y(n_289)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx8_ASAP7_75t_L g292 ( 
.A(n_107),
.Y(n_292)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_108),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_108),
.A2(n_208),
.B(n_211),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_145),
.B(n_152),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_111),
.B(n_145),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_118),
.B1(n_137),
.B2(n_138),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_113),
.A2(n_119),
.B(n_194),
.Y(n_193)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_114),
.Y(n_117)
);

INVx5_ASAP7_75t_L g248 ( 
.A(n_114),
.Y(n_248)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_118),
.B(n_195),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_118),
.A2(n_138),
.B(n_203),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_118),
.A2(n_226),
.B(n_247),
.Y(n_246)
);

INVx2_ASAP7_75t_SL g300 ( 
.A(n_118),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_118),
.A2(n_137),
.B1(n_346),
.B2(n_455),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_SL g498 ( 
.A1(n_118),
.A2(n_137),
.B(n_499),
.Y(n_498)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_127),
.Y(n_118)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_119),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_119),
.B(n_227),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_119),
.A2(n_300),
.B1(n_320),
.B2(n_328),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_119),
.A2(n_300),
.B1(n_320),
.B2(n_345),
.Y(n_344)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx6_ASAP7_75t_L g447 ( 
.A(n_122),
.Y(n_447)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_123),
.Y(n_136)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_124),
.Y(n_126)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_124),
.Y(n_132)
);

INVx3_ASAP7_75t_L g451 ( 
.A(n_124),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_128),
.A2(n_130),
.B1(n_133),
.B2(n_136),
.Y(n_127)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_129),
.Y(n_196)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_135),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_137),
.B(n_195),
.Y(n_204)
);

OAI21xp33_ASAP7_75t_SL g455 ( 
.A1(n_139),
.A2(n_380),
.B(n_448),
.Y(n_455)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

BUFx2_ASAP7_75t_L g347 ( 
.A(n_141),
.Y(n_347)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_142),
.Y(n_144)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_150),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g477 ( 
.A(n_146),
.Y(n_477)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

FAx1_ASAP7_75t_SL g197 ( 
.A(n_152),
.B(n_198),
.CI(n_214),
.CON(n_197),
.SN(n_197)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_181),
.C(n_192),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_154),
.B(n_360),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_172),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_155),
.A2(n_172),
.B1(n_173),
.B2(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_155),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_167),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_157),
.A2(n_271),
.B(n_337),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_158),
.Y(n_307)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

BUFx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx4_ASAP7_75t_L g426 ( 
.A(n_161),
.Y(n_426)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_162),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_163),
.Y(n_279)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g432 ( 
.A(n_165),
.B(n_433),
.Y(n_432)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_171),
.Y(n_275)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_181),
.A2(n_182),
.B1(n_192),
.B2(n_193),
.Y(n_360)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_190),
.B(n_211),
.Y(n_507)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_194),
.B(n_225),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_197),
.B(n_217),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_197),
.B(n_217),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_199),
.A2(n_200),
.B1(n_207),
.B2(n_213),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_205),
.B2(n_206),
.Y(n_200)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_201),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_201),
.A2(n_206),
.B1(n_223),
.B2(n_224),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_201),
.B(n_223),
.C(n_233),
.Y(n_503)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_202),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_202),
.B(n_206),
.C(n_207),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_204),
.A2(n_227),
.B(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_207),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_207),
.A2(n_213),
.B1(n_220),
.B2(n_221),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_207),
.B(n_218),
.C(n_221),
.Y(n_496)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_208),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_209),
.Y(n_257)
);

INVx8_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_210),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g492 ( 
.A1(n_216),
.A2(n_493),
.B(n_494),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_233),
.Y(n_221)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g499 ( 
.A(n_227),
.Y(n_499)
);

INVx8_ASAP7_75t_L g443 ( 
.A(n_228),
.Y(n_443)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx6_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_232),
.Y(n_324)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_232),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_235),
.Y(n_501)
);

INVx5_ASAP7_75t_L g284 ( 
.A(n_236),
.Y(n_284)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_237),
.Y(n_268)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

OA21x2_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_367),
.B(n_486),
.Y(n_240)
);

NAND3xp33_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_352),
.C(n_364),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_243),
.B(n_330),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g487 ( 
.A1(n_243),
.A2(n_488),
.B(n_489),
.Y(n_487)
);

NOR2xp67_ASAP7_75t_SL g243 ( 
.A(n_244),
.B(n_309),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_244),
.B(n_309),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_245),
.B(n_293),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_245),
.B(n_294),
.C(n_296),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_252),
.C(n_281),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_246),
.B(n_281),
.Y(n_311)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_247),
.Y(n_328)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_250),
.Y(n_249)
);

INVx6_ASAP7_75t_SL g250 ( 
.A(n_251),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_251),
.B(n_263),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_252),
.B(n_311),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_269),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_253),
.B(n_269),
.Y(n_333)
);

OAI32xp33_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_257),
.A3(n_258),
.B1(n_262),
.B2(n_265),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

BUFx12f_ASAP7_75t_L g349 ( 
.A(n_256),
.Y(n_349)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx8_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVxp33_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx2_ASAP7_75t_SL g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx6_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g414 ( 
.A(n_274),
.Y(n_414)
);

INVx4_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx8_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_282),
.Y(n_318)
);

INVx4_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx4_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_296),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_303),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_298),
.A2(n_299),
.B1(n_301),
.B2(n_302),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_298),
.B(n_302),
.C(n_355),
.Y(n_354)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_301),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_303),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_308),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_304),
.B(n_308),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_312),
.C(n_329),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_310),
.B(n_351),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_312),
.B(n_329),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.C(n_319),
.Y(n_312)
);

FAx1_ASAP7_75t_L g332 ( 
.A(n_313),
.B(n_314),
.CI(n_319),
.CON(n_332),
.SN(n_332)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx3_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_325),
.B(n_380),
.Y(n_448)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_350),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_331),
.B(n_350),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_333),
.C(n_334),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_332),
.B(n_484),
.Y(n_483)
);

BUFx24_ASAP7_75t_SL g512 ( 
.A(n_332),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_333),
.B(n_334),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_342),
.C(n_344),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_335),
.A2(n_336),
.B1(n_342),
.B2(n_343),
.Y(n_471)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_338),
.B(n_380),
.Y(n_433)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx8_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_SL g470 ( 
.A(n_344),
.B(n_471),
.Y(n_470)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

A2O1A1O1Ixp25_ASAP7_75t_L g486 ( 
.A1(n_352),
.A2(n_364),
.B(n_487),
.C(n_490),
.D(n_491),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_353),
.B(n_363),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_353),
.B(n_363),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_356),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_354),
.B(n_357),
.C(n_362),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_357),
.A2(n_359),
.B1(n_361),
.B2(n_362),
.Y(n_356)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_357),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_359),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_366),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_365),
.B(n_366),
.Y(n_491)
);

BUFx24_ASAP7_75t_SL g513 ( 
.A(n_366),
.Y(n_513)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_368),
.A2(n_481),
.B(n_485),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_SL g368 ( 
.A1(n_369),
.A2(n_466),
.B(n_480),
.Y(n_368)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_370),
.A2(n_437),
.B(n_465),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_SL g370 ( 
.A1(n_371),
.A2(n_409),
.B(n_436),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_392),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_372),
.B(n_392),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_378),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_373),
.B(n_378),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_375),
.Y(n_373)
);

INVx3_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx3_ASAP7_75t_SL g381 ( 
.A(n_382),
.Y(n_381)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_382),
.Y(n_464)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

BUFx3_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_385),
.Y(n_399)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

BUFx2_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_401),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_394),
.A2(n_395),
.B1(n_396),
.B2(n_400),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_394),
.B(n_400),
.C(n_401),
.Y(n_438)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx1_ASAP7_75t_SL g400 ( 
.A(n_396),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_399),
.B(n_450),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_402),
.Y(n_416)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx6_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g409 ( 
.A1(n_410),
.A2(n_420),
.B(n_435),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_419),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_411),
.B(n_419),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_412),
.A2(n_415),
.B1(n_416),
.B2(n_417),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_SL g420 ( 
.A1(n_421),
.A2(n_430),
.B(n_434),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_422),
.B(n_423),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_422),
.B(n_423),
.Y(n_434)
);

INVx4_ASAP7_75t_SL g425 ( 
.A(n_426),
.Y(n_425)
);

INVx5_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_431),
.B(n_432),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_438),
.B(n_439),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_438),
.B(n_439),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_453),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_440),
.B(n_454),
.C(n_456),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_SL g440 ( 
.A(n_441),
.B(n_452),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_441),
.B(n_452),
.Y(n_474)
);

OAI32xp33_ASAP7_75t_L g441 ( 
.A1(n_442),
.A2(n_444),
.A3(n_447),
.B1(n_448),
.B2(n_449),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx3_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVx6_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_456),
.Y(n_453)
);

INVxp67_ASAP7_75t_L g476 ( 
.A(n_457),
.Y(n_476)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_468),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_467),
.B(n_468),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_469),
.A2(n_470),
.B1(n_472),
.B2(n_473),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_469),
.B(n_475),
.C(n_478),
.Y(n_482)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_474),
.A2(n_475),
.B1(n_478),
.B2(n_479),
.Y(n_473)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_474),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_475),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_482),
.B(n_483),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_482),
.B(n_483),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_496),
.B(n_497),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_496),
.B(n_497),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_497),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_SL g510 ( 
.A(n_497),
.B(n_507),
.Y(n_510)
);

FAx1_ASAP7_75t_SL g497 ( 
.A(n_498),
.B(n_500),
.CI(n_503),
.CON(n_497),
.SN(n_497)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_506),
.B(n_508),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_507),
.Y(n_506)
);

INVxp67_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);


endmodule