module real_aes_3025_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_693;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_755;
wire n_656;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_754;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_434;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_785;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g208 ( .A(n_0), .B(n_155), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_1), .B(n_119), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_2), .B(n_139), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_3), .B(n_157), .Y(n_548) );
INVx1_ASAP7_75t_L g146 ( .A(n_4), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_5), .B(n_139), .Y(n_138) );
NAND2xp33_ASAP7_75t_SL g252 ( .A(n_6), .B(n_145), .Y(n_252) );
INVx1_ASAP7_75t_L g244 ( .A(n_7), .Y(n_244) );
CKINVDCx16_ASAP7_75t_R g119 ( .A(n_8), .Y(n_119) );
AND2x2_ASAP7_75t_L g133 ( .A(n_9), .B(n_134), .Y(n_133) );
AND2x2_ASAP7_75t_L g486 ( .A(n_10), .B(n_250), .Y(n_486) );
AND2x2_ASAP7_75t_L g550 ( .A(n_11), .B(n_184), .Y(n_550) );
INVx2_ASAP7_75t_L g135 ( .A(n_12), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_13), .B(n_157), .Y(n_532) );
CKINVDCx16_ASAP7_75t_R g111 ( .A(n_14), .Y(n_111) );
AOI221x1_ASAP7_75t_L g247 ( .A1(n_15), .A2(n_148), .B1(n_248), .B2(n_250), .C(n_251), .Y(n_247) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_16), .B(n_139), .Y(n_231) );
NAND2xp5_ASAP7_75t_SL g505 ( .A(n_17), .B(n_139), .Y(n_505) );
INVx1_ASAP7_75t_L g115 ( .A(n_18), .Y(n_115) );
AOI22xp5_ASAP7_75t_L g443 ( .A1(n_19), .A2(n_65), .B1(n_444), .B2(n_445), .Y(n_443) );
CKINVDCx20_ASAP7_75t_R g444 ( .A(n_19), .Y(n_444) );
AOI22xp33_ASAP7_75t_L g490 ( .A1(n_20), .A2(n_91), .B1(n_139), .B2(n_188), .Y(n_490) );
AOI21xp5_ASAP7_75t_L g147 ( .A1(n_21), .A2(n_148), .B(n_153), .Y(n_147) );
AOI221xp5_ASAP7_75t_SL g218 ( .A1(n_22), .A2(n_35), .B1(n_139), .B2(n_148), .C(n_219), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_23), .B(n_155), .Y(n_154) );
OR2x2_ASAP7_75t_L g136 ( .A(n_24), .B(n_90), .Y(n_136) );
OA21x2_ASAP7_75t_L g185 ( .A1(n_24), .A2(n_90), .B(n_135), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_25), .B(n_157), .Y(n_235) );
INVxp67_ASAP7_75t_L g246 ( .A(n_26), .Y(n_246) );
AND2x2_ASAP7_75t_L g179 ( .A(n_27), .B(n_169), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_28), .A2(n_148), .B(n_207), .Y(n_206) );
AO21x2_ASAP7_75t_L g527 ( .A1(n_29), .A2(n_250), .B(n_528), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_30), .B(n_157), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g545 ( .A1(n_31), .A2(n_148), .B(n_546), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_32), .B(n_157), .Y(n_521) );
AND2x2_ASAP7_75t_L g145 ( .A(n_33), .B(n_146), .Y(n_145) );
AND2x2_ASAP7_75t_L g149 ( .A(n_33), .B(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g196 ( .A(n_33), .Y(n_196) );
OR2x6_ASAP7_75t_L g113 ( .A(n_34), .B(n_114), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_36), .B(n_139), .Y(n_549) );
AOI22xp5_ASAP7_75t_L g193 ( .A1(n_37), .A2(n_82), .B1(n_148), .B2(n_194), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_38), .B(n_157), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_39), .B(n_139), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_40), .B(n_155), .Y(n_177) );
AOI21xp5_ASAP7_75t_L g481 ( .A1(n_41), .A2(n_148), .B(n_482), .Y(n_481) );
CKINVDCx20_ASAP7_75t_R g786 ( .A(n_42), .Y(n_786) );
OAI22xp5_ASAP7_75t_L g774 ( .A1(n_43), .A2(n_51), .B1(n_775), .B2(n_776), .Y(n_774) );
INVx1_ASAP7_75t_L g776 ( .A(n_43), .Y(n_776) );
AND2x2_ASAP7_75t_L g211 ( .A(n_44), .B(n_169), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_45), .B(n_155), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_46), .B(n_169), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g529 ( .A(n_47), .B(n_139), .Y(n_529) );
INVx1_ASAP7_75t_L g142 ( .A(n_48), .Y(n_142) );
INVx1_ASAP7_75t_L g152 ( .A(n_48), .Y(n_152) );
OAI22xp5_ASAP7_75t_L g125 ( .A1(n_49), .A2(n_126), .B1(n_446), .B2(n_447), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g447 ( .A(n_49), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_50), .B(n_157), .Y(n_484) );
INVx1_ASAP7_75t_L g775 ( .A(n_51), .Y(n_775) );
AND2x2_ASAP7_75t_L g496 ( .A(n_52), .B(n_169), .Y(n_496) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_53), .B(n_139), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_54), .B(n_155), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_55), .B(n_155), .Y(n_520) );
AND2x2_ASAP7_75t_L g170 ( .A(n_56), .B(n_169), .Y(n_170) );
NAND2xp5_ASAP7_75t_SL g485 ( .A(n_57), .B(n_139), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_58), .B(n_157), .Y(n_209) );
NAND2xp5_ASAP7_75t_SL g498 ( .A(n_59), .B(n_139), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_60), .A2(n_148), .B(n_519), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_61), .B(n_155), .Y(n_166) );
AND2x2_ASAP7_75t_SL g236 ( .A(n_62), .B(n_134), .Y(n_236) );
AND2x2_ASAP7_75t_L g511 ( .A(n_63), .B(n_134), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g174 ( .A1(n_64), .A2(n_148), .B(n_175), .Y(n_174) );
CKINVDCx20_ASAP7_75t_R g445 ( .A(n_65), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_66), .B(n_157), .Y(n_156) );
AND2x2_ASAP7_75t_SL g199 ( .A(n_67), .B(n_184), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_68), .B(n_155), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_69), .B(n_155), .Y(n_533) );
AOI22xp5_ASAP7_75t_L g491 ( .A1(n_70), .A2(n_93), .B1(n_148), .B2(n_194), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_71), .B(n_157), .Y(n_508) );
INVx1_ASAP7_75t_L g144 ( .A(n_72), .Y(n_144) );
INVx1_ASAP7_75t_L g150 ( .A(n_72), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_73), .B(n_155), .Y(n_547) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_74), .A2(n_148), .B(n_500), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g473 ( .A1(n_75), .A2(n_148), .B(n_474), .Y(n_473) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_76), .A2(n_148), .B(n_531), .Y(n_530) );
AND2x2_ASAP7_75t_L g523 ( .A(n_77), .B(n_134), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g488 ( .A(n_78), .B(n_169), .Y(n_488) );
AOI22xp5_ASAP7_75t_L g771 ( .A1(n_79), .A2(n_772), .B1(n_773), .B2(n_774), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_79), .Y(n_772) );
NAND2xp5_ASAP7_75t_SL g167 ( .A(n_80), .B(n_139), .Y(n_167) );
AOI22xp5_ASAP7_75t_L g187 ( .A1(n_81), .A2(n_84), .B1(n_139), .B2(n_188), .Y(n_187) );
INVx1_ASAP7_75t_L g116 ( .A(n_83), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_85), .B(n_155), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_86), .B(n_155), .Y(n_221) );
AND2x2_ASAP7_75t_L g477 ( .A(n_87), .B(n_184), .Y(n_477) );
CKINVDCx20_ASAP7_75t_R g449 ( .A(n_88), .Y(n_449) );
AOI21xp5_ASAP7_75t_L g163 ( .A1(n_89), .A2(n_148), .B(n_164), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_92), .B(n_157), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_94), .A2(n_148), .B(n_507), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_95), .B(n_157), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_96), .B(n_139), .Y(n_210) );
INVxp67_ASAP7_75t_L g249 ( .A(n_97), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_98), .B(n_157), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_99), .A2(n_148), .B(n_233), .Y(n_232) );
BUFx2_ASAP7_75t_L g510 ( .A(n_100), .Y(n_510) );
BUFx2_ASAP7_75t_L g124 ( .A(n_101), .Y(n_124) );
AOI22xp33_ASAP7_75t_SL g777 ( .A1(n_102), .A2(n_771), .B1(n_778), .B2(n_781), .Y(n_777) );
AOI21xp5_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_120), .B(n_785), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
NOR2xp33_ASAP7_75t_L g785 ( .A(n_106), .B(n_786), .Y(n_785) );
INVx2_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
NAND2xp5_ASAP7_75t_SL g107 ( .A(n_108), .B(n_117), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
BUFx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
INVxp67_ASAP7_75t_SL g123 ( .A(n_110), .Y(n_123) );
BUFx3_ASAP7_75t_L g452 ( .A(n_110), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_111), .B(n_112), .Y(n_110) );
AND2x6_ASAP7_75t_SL g461 ( .A(n_111), .B(n_113), .Y(n_461) );
OR2x6_ASAP7_75t_SL g770 ( .A(n_111), .B(n_112), .Y(n_770) );
OR2x2_ASAP7_75t_L g784 ( .A(n_111), .B(n_113), .Y(n_784) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_113), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_115), .B(n_116), .Y(n_114) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
OR2x6_ASAP7_75t_L g120 ( .A(n_121), .B(n_453), .Y(n_120) );
AO21x1_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_125), .B(n_448), .Y(n_121) );
NOR2x1_ASAP7_75t_R g122 ( .A(n_123), .B(n_124), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g455 ( .A(n_124), .Y(n_455) );
INVx2_ASAP7_75t_L g446 ( .A(n_126), .Y(n_446) );
XNOR2x1_ASAP7_75t_L g126 ( .A(n_127), .B(n_443), .Y(n_126) );
INVx3_ASAP7_75t_SL g459 ( .A(n_127), .Y(n_459) );
OAI22xp5_ASAP7_75t_SL g778 ( .A1(n_127), .A2(n_463), .B1(n_779), .B2(n_780), .Y(n_778) );
AND2x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_373), .Y(n_127) );
NOR4xp25_ASAP7_75t_SL g128 ( .A(n_129), .B(n_266), .C(n_310), .D(n_337), .Y(n_128) );
OAI221xp5_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_227), .B1(n_237), .B2(n_254), .C(n_256), .Y(n_129) );
AOI32xp33_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_180), .A3(n_200), .B1(n_212), .B2(n_223), .Y(n_130) );
NOR2xp33_ASAP7_75t_L g408 ( .A(n_131), .B(n_409), .Y(n_408) );
AOI22xp5_ASAP7_75t_L g436 ( .A1(n_131), .A2(n_379), .B1(n_437), .B2(n_440), .Y(n_436) );
AND2x4_ASAP7_75t_SL g131 ( .A(n_132), .B(n_160), .Y(n_131) );
INVx5_ASAP7_75t_L g226 ( .A(n_132), .Y(n_226) );
OR2x2_ASAP7_75t_L g255 ( .A(n_132), .B(n_225), .Y(n_255) );
AND2x4_ASAP7_75t_L g257 ( .A(n_132), .B(n_172), .Y(n_257) );
INVx2_ASAP7_75t_L g272 ( .A(n_132), .Y(n_272) );
OR2x2_ASAP7_75t_L g284 ( .A(n_132), .B(n_181), .Y(n_284) );
AND2x2_ASAP7_75t_L g291 ( .A(n_132), .B(n_171), .Y(n_291) );
AND2x2_ASAP7_75t_SL g333 ( .A(n_132), .B(n_214), .Y(n_333) );
HB1xp67_ASAP7_75t_L g390 ( .A(n_132), .Y(n_390) );
OR2x6_ASAP7_75t_L g132 ( .A(n_133), .B(n_137), .Y(n_132) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_134), .Y(n_169) );
AND2x2_ASAP7_75t_SL g134 ( .A(n_135), .B(n_136), .Y(n_134) );
AND2x4_ASAP7_75t_L g159 ( .A(n_135), .B(n_136), .Y(n_159) );
AOI21xp5_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_147), .B(n_159), .Y(n_137) );
AND2x4_ASAP7_75t_L g139 ( .A(n_140), .B(n_145), .Y(n_139) );
INVx1_ASAP7_75t_L g253 ( .A(n_140), .Y(n_253) );
AND2x4_ASAP7_75t_L g140 ( .A(n_141), .B(n_143), .Y(n_140) );
AND2x6_ASAP7_75t_L g155 ( .A(n_141), .B(n_150), .Y(n_155) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
AND2x4_ASAP7_75t_L g157 ( .A(n_143), .B(n_152), .Y(n_157) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx5_ASAP7_75t_L g158 ( .A(n_145), .Y(n_158) );
AND2x2_ASAP7_75t_L g151 ( .A(n_146), .B(n_152), .Y(n_151) );
HB1xp67_ASAP7_75t_L g191 ( .A(n_146), .Y(n_191) );
AND2x6_ASAP7_75t_L g148 ( .A(n_149), .B(n_151), .Y(n_148) );
BUFx3_ASAP7_75t_L g192 ( .A(n_149), .Y(n_192) );
INVx2_ASAP7_75t_L g198 ( .A(n_150), .Y(n_198) );
AND2x4_ASAP7_75t_L g194 ( .A(n_151), .B(n_195), .Y(n_194) );
INVx2_ASAP7_75t_L g190 ( .A(n_152), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g153 ( .A1(n_154), .A2(n_156), .B(n_158), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_155), .B(n_510), .Y(n_509) );
AOI21xp5_ASAP7_75t_L g164 ( .A1(n_158), .A2(n_165), .B(n_166), .Y(n_164) );
AOI21xp5_ASAP7_75t_L g175 ( .A1(n_158), .A2(n_176), .B(n_177), .Y(n_175) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_158), .A2(n_208), .B(n_209), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_158), .A2(n_220), .B(n_221), .Y(n_219) );
AOI21xp5_ASAP7_75t_L g233 ( .A1(n_158), .A2(n_234), .B(n_235), .Y(n_233) );
AOI21xp5_ASAP7_75t_L g474 ( .A1(n_158), .A2(n_475), .B(n_476), .Y(n_474) );
AOI21xp5_ASAP7_75t_L g482 ( .A1(n_158), .A2(n_483), .B(n_484), .Y(n_482) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_158), .A2(n_501), .B(n_502), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_158), .A2(n_508), .B(n_509), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_158), .A2(n_520), .B(n_521), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_158), .A2(n_532), .B(n_533), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g546 ( .A1(n_158), .A2(n_547), .B(n_548), .Y(n_546) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_159), .B(n_244), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_159), .B(n_246), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_159), .B(n_249), .Y(n_248) );
NOR3xp33_ASAP7_75t_L g251 ( .A(n_159), .B(n_252), .C(n_253), .Y(n_251) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_159), .A2(n_498), .B(n_499), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_159), .A2(n_529), .B(n_530), .Y(n_528) );
INVx3_ASAP7_75t_SL g285 ( .A(n_160), .Y(n_285) );
AND2x2_ASAP7_75t_L g304 ( .A(n_160), .B(n_226), .Y(n_304) );
AOI32xp33_ASAP7_75t_L g419 ( .A1(n_160), .A2(n_290), .A3(n_320), .B1(n_350), .B2(n_385), .Y(n_419) );
AND2x4_ASAP7_75t_L g160 ( .A(n_161), .B(n_171), .Y(n_160) );
AND2x2_ASAP7_75t_L g259 ( .A(n_161), .B(n_181), .Y(n_259) );
OR2x2_ASAP7_75t_L g275 ( .A(n_161), .B(n_172), .Y(n_275) );
INVx1_ASAP7_75t_L g298 ( .A(n_161), .Y(n_298) );
INVx2_ASAP7_75t_L g314 ( .A(n_161), .Y(n_314) );
AND2x2_ASAP7_75t_L g351 ( .A(n_161), .B(n_214), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_161), .B(n_172), .Y(n_370) );
HB1xp67_ASAP7_75t_L g439 ( .A(n_161), .Y(n_439) );
AO21x2_ASAP7_75t_L g161 ( .A1(n_162), .A2(n_168), .B(n_170), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_163), .B(n_167), .Y(n_162) );
AO21x2_ASAP7_75t_L g172 ( .A1(n_168), .A2(n_173), .B(n_179), .Y(n_172) );
AO21x2_ASAP7_75t_L g225 ( .A1(n_168), .A2(n_173), .B(n_179), .Y(n_225) );
AOI21x1_ASAP7_75t_L g543 ( .A1(n_168), .A2(n_544), .B(n_550), .Y(n_543) );
CKINVDCx5p33_ASAP7_75t_R g168 ( .A(n_169), .Y(n_168) );
OA21x2_ASAP7_75t_L g217 ( .A1(n_169), .A2(n_218), .B(n_222), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g471 ( .A1(n_169), .A2(n_472), .B(n_473), .Y(n_471) );
AO21x2_ASAP7_75t_L g489 ( .A1(n_169), .A2(n_490), .B(n_491), .Y(n_489) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
AND2x2_ASAP7_75t_L g406 ( .A(n_172), .B(n_181), .Y(n_406) );
HB1xp67_ASAP7_75t_L g428 ( .A(n_172), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_174), .B(n_178), .Y(n_173) );
OR2x2_ASAP7_75t_L g254 ( .A(n_180), .B(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g260 ( .A(n_180), .B(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g273 ( .A(n_180), .B(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g435 ( .A(n_180), .B(n_304), .Y(n_435) );
BUFx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
AND2x2_ASAP7_75t_L g364 ( .A(n_181), .B(n_314), .Y(n_364) );
INVx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
BUFx6f_ASAP7_75t_L g214 ( .A(n_182), .Y(n_214) );
AOI21x1_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_186), .B(n_199), .Y(n_182) );
INVx2_ASAP7_75t_SL g183 ( .A(n_184), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_184), .A2(n_231), .B(n_232), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g504 ( .A1(n_184), .A2(n_505), .B(n_506), .Y(n_504) );
BUFx4f_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
INVx3_ASAP7_75t_L g204 ( .A(n_185), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_187), .B(n_193), .Y(n_186) );
AOI22xp5_ASAP7_75t_L g242 ( .A1(n_188), .A2(n_194), .B1(n_243), .B2(n_245), .Y(n_242) );
AND2x4_ASAP7_75t_L g188 ( .A(n_189), .B(n_192), .Y(n_188) );
AND2x2_ASAP7_75t_L g189 ( .A(n_190), .B(n_191), .Y(n_189) );
NOR2x1p5_ASAP7_75t_L g195 ( .A(n_196), .B(n_197), .Y(n_195) );
INVx3_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g433 ( .A(n_200), .B(n_331), .Y(n_433) );
INVx1_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_201), .B(n_381), .Y(n_380) );
HB1xp67_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
AND2x2_ASAP7_75t_L g216 ( .A(n_202), .B(n_217), .Y(n_216) );
INVx1_ASAP7_75t_L g238 ( .A(n_202), .Y(n_238) );
AND2x2_ASAP7_75t_L g264 ( .A(n_202), .B(n_265), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_202), .B(n_240), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_202), .B(n_302), .Y(n_301) );
INVx2_ASAP7_75t_L g322 ( .A(n_202), .Y(n_322) );
OR2x2_ASAP7_75t_L g341 ( .A(n_202), .B(n_268), .Y(n_341) );
INVx1_ASAP7_75t_L g348 ( .A(n_202), .Y(n_348) );
NOR2xp33_ASAP7_75t_R g400 ( .A(n_202), .B(n_229), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_202), .B(n_241), .Y(n_404) );
INVx3_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
AOI21x1_ASAP7_75t_L g203 ( .A1(n_204), .A2(n_205), .B(n_211), .Y(n_203) );
INVx4_ASAP7_75t_L g250 ( .A(n_204), .Y(n_250) );
AO21x2_ASAP7_75t_L g479 ( .A1(n_204), .A2(n_480), .B(n_486), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_206), .B(n_210), .Y(n_205) );
AOI32xp33_ASAP7_75t_L g427 ( .A1(n_212), .A2(n_263), .A3(n_428), .B1(n_429), .B2(n_430), .Y(n_427) );
INVx3_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
OR2x2_ASAP7_75t_L g213 ( .A(n_214), .B(n_215), .Y(n_213) );
INVx2_ASAP7_75t_L g294 ( .A(n_214), .Y(n_294) );
AND2x4_ASAP7_75t_L g313 ( .A(n_214), .B(n_314), .Y(n_313) );
NOR2xp33_ASAP7_75t_L g342 ( .A(n_214), .B(n_285), .Y(n_342) );
OR2x2_ASAP7_75t_L g396 ( .A(n_214), .B(n_397), .Y(n_396) );
OR2x2_ASAP7_75t_L g354 ( .A(n_215), .B(n_355), .Y(n_354) );
OR2x2_ASAP7_75t_L g412 ( .A(n_215), .B(n_413), .Y(n_412) );
INVx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_216), .B(n_229), .Y(n_378) );
AND2x2_ASAP7_75t_L g415 ( .A(n_216), .B(n_381), .Y(n_415) );
INVx2_ASAP7_75t_L g265 ( .A(n_217), .Y(n_265) );
INVx2_ASAP7_75t_L g268 ( .A(n_217), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_217), .B(n_229), .Y(n_288) );
INVx1_ASAP7_75t_L g319 ( .A(n_217), .Y(n_319) );
OR2x2_ASAP7_75t_L g345 ( .A(n_217), .B(n_229), .Y(n_345) );
HB1xp67_ASAP7_75t_L g397 ( .A(n_217), .Y(n_397) );
BUFx3_ASAP7_75t_L g426 ( .A(n_217), .Y(n_426) );
HB1xp67_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVx2_ASAP7_75t_L g295 ( .A(n_224), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_224), .B(n_313), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_224), .B(n_384), .Y(n_383) );
AND2x4_ASAP7_75t_L g224 ( .A(n_225), .B(n_226), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_225), .B(n_298), .Y(n_297) );
OAI21xp33_ASAP7_75t_L g327 ( .A1(n_225), .A2(n_294), .B(n_312), .Y(n_327) );
OAI32xp33_ASAP7_75t_L g349 ( .A1(n_226), .A2(n_350), .A3(n_352), .B1(n_354), .B2(n_356), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_226), .B(n_313), .Y(n_422) );
HB1xp67_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
INVx1_ASAP7_75t_L g355 ( .A(n_228), .Y(n_355) );
NOR2x1p5_ASAP7_75t_L g425 ( .A(n_228), .B(n_426), .Y(n_425) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
AND2x4_ASAP7_75t_L g239 ( .A(n_229), .B(n_240), .Y(n_239) );
AND2x4_ASAP7_75t_SL g263 ( .A(n_229), .B(n_241), .Y(n_263) );
OR2x2_ASAP7_75t_L g267 ( .A(n_229), .B(n_268), .Y(n_267) );
INVx2_ASAP7_75t_L g302 ( .A(n_229), .Y(n_302) );
AND2x2_ASAP7_75t_L g320 ( .A(n_229), .B(n_321), .Y(n_320) );
OR2x2_ASAP7_75t_L g331 ( .A(n_229), .B(n_241), .Y(n_331) );
OR2x2_ASAP7_75t_L g393 ( .A(n_229), .B(n_394), .Y(n_393) );
OR2x2_ASAP7_75t_L g410 ( .A(n_229), .B(n_341), .Y(n_410) );
INVx1_ASAP7_75t_L g442 ( .A(n_229), .Y(n_442) );
OR2x6_ASAP7_75t_L g229 ( .A(n_230), .B(n_236), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_238), .B(n_239), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_238), .B(n_319), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_239), .B(n_353), .Y(n_352) );
AOI222xp33_ASAP7_75t_L g357 ( .A1(n_239), .A2(n_358), .B1(n_363), .B2(n_365), .C1(n_368), .C2(n_371), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_239), .B(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g385 ( .A(n_239), .B(n_264), .Y(n_385) );
AND2x2_ASAP7_75t_L g347 ( .A(n_240), .B(n_348), .Y(n_347) );
OR2x2_ASAP7_75t_L g362 ( .A(n_240), .B(n_267), .Y(n_362) );
INVx3_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_241), .B(n_268), .Y(n_300) );
AND2x4_ASAP7_75t_L g321 ( .A(n_241), .B(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g381 ( .A(n_241), .B(n_302), .Y(n_381) );
AND2x4_ASAP7_75t_L g241 ( .A(n_242), .B(n_247), .Y(n_241) );
INVx3_ASAP7_75t_L g516 ( .A(n_250), .Y(n_516) );
INVx1_ASAP7_75t_SL g261 ( .A(n_255), .Y(n_261) );
NAND2xp33_ASAP7_75t_SL g430 ( .A(n_255), .B(n_285), .Y(n_430) );
A2O1A1Ixp33_ASAP7_75t_L g256 ( .A1(n_257), .A2(n_258), .B(n_260), .C(n_262), .Y(n_256) );
INVx2_ASAP7_75t_SL g307 ( .A(n_257), .Y(n_307) );
AND2x2_ASAP7_75t_L g311 ( .A(n_258), .B(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_259), .B(n_307), .Y(n_306) );
O2A1O1Ixp33_ASAP7_75t_L g332 ( .A1(n_259), .A2(n_297), .B(n_333), .C(n_334), .Y(n_332) );
AND2x2_ASAP7_75t_L g409 ( .A(n_259), .B(n_390), .Y(n_409) );
AND2x2_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
AND2x4_ASAP7_75t_L g308 ( .A(n_263), .B(n_309), .Y(n_308) );
INVx1_ASAP7_75t_SL g413 ( .A(n_263), .Y(n_413) );
OAI211xp5_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_269), .B(n_276), .C(n_303), .Y(n_266) );
INVx2_ASAP7_75t_L g278 ( .A(n_267), .Y(n_278) );
OR2x2_ASAP7_75t_L g325 ( .A(n_267), .B(n_326), .Y(n_325) );
HB1xp67_ASAP7_75t_L g309 ( .A(n_268), .Y(n_309) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g270 ( .A(n_271), .B(n_273), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_271), .B(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g363 ( .A(n_271), .B(n_364), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_271), .B(n_351), .Y(n_417) );
INVx2_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AOI222xp33_ASAP7_75t_L g375 ( .A1(n_273), .A2(n_376), .B1(n_377), .B2(n_379), .C1(n_382), .C2(n_385), .Y(n_375) );
AOI221xp5_ASAP7_75t_L g338 ( .A1(n_274), .A2(n_339), .B1(n_342), .B2(n_343), .C(n_349), .Y(n_338) );
AND2x2_ASAP7_75t_L g376 ( .A(n_274), .B(n_333), .Y(n_376) );
INVx2_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
NAND2xp33_ASAP7_75t_SL g289 ( .A(n_275), .B(n_290), .Y(n_289) );
AOI221x1_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_281), .B1(n_286), .B2(n_289), .C(n_292), .Y(n_276) );
AND2x4_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
AND2x2_ASAP7_75t_L g429 ( .A(n_279), .B(n_367), .Y(n_429) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
OR2x2_ASAP7_75t_L g287 ( .A(n_280), .B(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_283), .B(n_285), .Y(n_282) );
INVx1_ASAP7_75t_SL g283 ( .A(n_284), .Y(n_283) );
OAI32xp33_ASAP7_75t_L g395 ( .A1(n_285), .A2(n_326), .A3(n_396), .B1(n_398), .B2(n_402), .Y(n_395) );
OAI21xp33_ASAP7_75t_SL g414 ( .A1(n_286), .A2(n_415), .B(n_416), .Y(n_414) );
INVx2_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AOI21xp33_ASAP7_75t_L g292 ( .A1(n_293), .A2(n_296), .B(n_299), .Y(n_292) );
OR2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_295), .Y(n_293) );
OR2x2_ASAP7_75t_L g296 ( .A(n_294), .B(n_297), .Y(n_296) );
OR2x2_ASAP7_75t_L g369 ( .A(n_294), .B(n_370), .Y(n_369) );
AOI221xp5_ASAP7_75t_L g323 ( .A1(n_298), .A2(n_324), .B1(n_327), .B2(n_328), .C(n_332), .Y(n_323) );
INVx1_ASAP7_75t_L g399 ( .A(n_298), .Y(n_399) );
HB1xp67_ASAP7_75t_L g405 ( .A(n_298), .Y(n_405) );
OR2x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
OAI21xp33_ASAP7_75t_L g303 ( .A1(n_304), .A2(n_305), .B(n_308), .Y(n_303) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
NOR2xp33_ASAP7_75t_L g371 ( .A(n_307), .B(n_372), .Y(n_371) );
OAI21xp5_ASAP7_75t_SL g310 ( .A1(n_311), .A2(n_315), .B(n_323), .Y(n_310) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_314), .Y(n_384) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g316 ( .A(n_317), .B(n_320), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_317), .B(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVxp67_ASAP7_75t_SL g318 ( .A(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g336 ( .A(n_319), .Y(n_336) );
INVx1_ASAP7_75t_L g326 ( .A(n_321), .Y(n_326) );
AND2x2_ASAP7_75t_SL g335 ( .A(n_321), .B(n_336), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_321), .B(n_367), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_321), .B(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_SL g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_SL g330 ( .A(n_331), .Y(n_330) );
OR2x2_ASAP7_75t_L g340 ( .A(n_331), .B(n_341), .Y(n_340) );
INVx2_ASAP7_75t_SL g334 ( .A(n_335), .Y(n_334) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_336), .Y(n_401) );
NAND2xp5_ASAP7_75t_SL g337 ( .A(n_338), .B(n_357), .Y(n_337) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g353 ( .A(n_341), .Y(n_353) );
INVx1_ASAP7_75t_SL g343 ( .A(n_344), .Y(n_343) );
OR2x2_ASAP7_75t_L g344 ( .A(n_345), .B(n_346), .Y(n_344) );
INVx1_ASAP7_75t_SL g367 ( .A(n_345), .Y(n_367) );
INVx1_ASAP7_75t_SL g346 ( .A(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_347), .B(n_425), .Y(n_424) );
HB1xp67_ASAP7_75t_L g361 ( .A(n_348), .Y(n_361) );
BUFx2_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
NAND2xp5_ASAP7_75t_SL g358 ( .A(n_359), .B(n_362), .Y(n_358) );
INVxp67_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g372 ( .A(n_364), .Y(n_372) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_SL g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g391 ( .A(n_370), .Y(n_391) );
NOR4xp25_ASAP7_75t_L g373 ( .A(n_374), .B(n_407), .C(n_418), .D(n_431), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_375), .B(n_386), .Y(n_374) );
O2A1O1Ixp33_ASAP7_75t_L g386 ( .A1(n_376), .A2(n_387), .B(n_392), .C(n_395), .Y(n_386) );
INVx1_ASAP7_75t_SL g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx2_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
NAND2xp5_ASAP7_75t_SL g388 ( .A(n_389), .B(n_391), .Y(n_388) );
OAI211xp5_ASAP7_75t_L g398 ( .A1(n_389), .A2(n_399), .B(n_400), .C(n_401), .Y(n_398) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_SL g392 ( .A(n_393), .Y(n_392) );
OAI21xp33_ASAP7_75t_SL g402 ( .A1(n_403), .A2(n_405), .B(n_406), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
AND2x2_ASAP7_75t_SL g437 ( .A(n_406), .B(n_438), .Y(n_437) );
OAI221xp5_ASAP7_75t_SL g407 ( .A1(n_408), .A2(n_410), .B1(n_411), .B2(n_412), .C(n_414), .Y(n_407) );
INVx1_ASAP7_75t_SL g411 ( .A(n_409), .Y(n_411) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
NAND3xp33_ASAP7_75t_SL g418 ( .A(n_419), .B(n_420), .C(n_427), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_421), .B(n_423), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
OAI21xp33_ASAP7_75t_L g431 ( .A1(n_432), .A2(n_434), .B(n_436), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVxp33_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_SL g440 ( .A(n_441), .Y(n_440) );
NOR2xp33_ASAP7_75t_L g448 ( .A(n_449), .B(n_450), .Y(n_448) );
CKINVDCx11_ASAP7_75t_R g450 ( .A(n_451), .Y(n_450) );
CKINVDCx20_ASAP7_75t_R g451 ( .A(n_452), .Y(n_451) );
AND2x2_ASAP7_75t_L g453 ( .A(n_454), .B(n_456), .Y(n_453) );
CKINVDCx5p33_ASAP7_75t_R g454 ( .A(n_455), .Y(n_454) );
OAI21xp5_ASAP7_75t_L g456 ( .A1(n_457), .A2(n_771), .B(n_777), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
OAI22x1_ASAP7_75t_SL g458 ( .A1(n_459), .A2(n_460), .B1(n_462), .B2(n_768), .Y(n_458) );
CKINVDCx5p33_ASAP7_75t_R g460 ( .A(n_461), .Y(n_460) );
CKINVDCx11_ASAP7_75t_R g779 ( .A(n_461), .Y(n_779) );
INVx2_ASAP7_75t_SL g462 ( .A(n_463), .Y(n_462) );
AND2x4_ASAP7_75t_L g463 ( .A(n_464), .B(n_693), .Y(n_463) );
NOR2xp67_ASAP7_75t_L g464 ( .A(n_465), .B(n_612), .Y(n_464) );
NAND5xp2_ASAP7_75t_L g465 ( .A(n_466), .B(n_556), .C(n_566), .D(n_583), .E(n_599), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
OAI22xp5_ASAP7_75t_L g467 ( .A1(n_468), .A2(n_492), .B1(n_534), .B2(n_538), .Y(n_467) );
OR2x2_ASAP7_75t_L g468 ( .A(n_469), .B(n_478), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
AND2x4_ASAP7_75t_L g540 ( .A(n_470), .B(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g558 ( .A(n_470), .B(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g579 ( .A(n_470), .B(n_580), .Y(n_579) );
INVx4_ASAP7_75t_L g593 ( .A(n_470), .Y(n_593) );
AND2x2_ASAP7_75t_L g602 ( .A(n_470), .B(n_603), .Y(n_602) );
AND2x4_ASAP7_75t_SL g624 ( .A(n_470), .B(n_542), .Y(n_624) );
BUFx2_ASAP7_75t_L g667 ( .A(n_470), .Y(n_667) );
AND2x2_ASAP7_75t_L g682 ( .A(n_470), .B(n_479), .Y(n_682) );
OR2x2_ASAP7_75t_L g714 ( .A(n_470), .B(n_715), .Y(n_714) );
NOR4xp25_ASAP7_75t_L g763 ( .A(n_470), .B(n_764), .C(n_765), .D(n_766), .Y(n_763) );
OR2x6_ASAP7_75t_L g470 ( .A(n_471), .B(n_477), .Y(n_470) );
AOI31xp33_ASAP7_75t_L g631 ( .A1(n_478), .A2(n_632), .A3(n_634), .B(n_636), .Y(n_631) );
INVx2_ASAP7_75t_SL g748 ( .A(n_478), .Y(n_748) );
OR2x2_ASAP7_75t_L g478 ( .A(n_479), .B(n_487), .Y(n_478) );
INVx2_ASAP7_75t_L g555 ( .A(n_479), .Y(n_555) );
AND2x2_ASAP7_75t_L g559 ( .A(n_479), .B(n_543), .Y(n_559) );
INVx2_ASAP7_75t_L g582 ( .A(n_479), .Y(n_582) );
AND2x2_ASAP7_75t_L g601 ( .A(n_479), .B(n_542), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_481), .B(n_485), .Y(n_480) );
AND2x2_ASAP7_75t_L g553 ( .A(n_487), .B(n_554), .Y(n_553) );
BUFx3_ASAP7_75t_L g560 ( .A(n_487), .Y(n_560) );
INVx2_ASAP7_75t_L g578 ( .A(n_487), .Y(n_578) );
AND2x2_ASAP7_75t_L g633 ( .A(n_487), .B(n_593), .Y(n_633) );
AND2x4_ASAP7_75t_L g487 ( .A(n_488), .B(n_489), .Y(n_487) );
AND2x4_ASAP7_75t_L g604 ( .A(n_488), .B(n_489), .Y(n_604) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_493), .B(n_524), .Y(n_492) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_494), .B(n_512), .Y(n_493) );
OR2x2_ASAP7_75t_L g534 ( .A(n_494), .B(n_535), .Y(n_534) );
INVx3_ASAP7_75t_L g685 ( .A(n_494), .Y(n_685) );
OR2x2_ASAP7_75t_L g733 ( .A(n_494), .B(n_734), .Y(n_733) );
NAND2x1_ASAP7_75t_L g494 ( .A(n_495), .B(n_503), .Y(n_494) );
OR2x2_ASAP7_75t_SL g525 ( .A(n_495), .B(n_526), .Y(n_525) );
INVx4_ASAP7_75t_L g563 ( .A(n_495), .Y(n_563) );
HB1xp67_ASAP7_75t_L g607 ( .A(n_495), .Y(n_607) );
INVx2_ASAP7_75t_L g615 ( .A(n_495), .Y(n_615) );
OR2x2_ASAP7_75t_L g650 ( .A(n_495), .B(n_514), .Y(n_650) );
AND2x2_ASAP7_75t_L g762 ( .A(n_495), .B(n_617), .Y(n_762) );
AND2x2_ASAP7_75t_L g767 ( .A(n_495), .B(n_527), .Y(n_767) );
OR2x6_ASAP7_75t_L g495 ( .A(n_496), .B(n_497), .Y(n_495) );
OR2x2_ASAP7_75t_L g526 ( .A(n_503), .B(n_527), .Y(n_526) );
AND2x2_ASAP7_75t_L g591 ( .A(n_503), .B(n_513), .Y(n_591) );
OR2x2_ASAP7_75t_L g598 ( .A(n_503), .B(n_563), .Y(n_598) );
NOR2x1_ASAP7_75t_SL g617 ( .A(n_503), .B(n_537), .Y(n_617) );
BUFx2_ASAP7_75t_L g649 ( .A(n_503), .Y(n_649) );
AND2x2_ASAP7_75t_L g658 ( .A(n_503), .B(n_563), .Y(n_658) );
AND2x2_ASAP7_75t_L g691 ( .A(n_503), .B(n_611), .Y(n_691) );
INVx2_ASAP7_75t_SL g700 ( .A(n_503), .Y(n_700) );
AND2x2_ASAP7_75t_L g703 ( .A(n_503), .B(n_514), .Y(n_703) );
OR2x6_ASAP7_75t_L g503 ( .A(n_504), .B(n_511), .Y(n_503) );
NAND3xp33_ASAP7_75t_L g698 ( .A(n_512), .B(n_568), .C(n_653), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_512), .B(n_615), .Y(n_718) );
INVxp67_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_513), .B(n_700), .Y(n_721) );
INVx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
HB1xp67_ASAP7_75t_L g565 ( .A(n_514), .Y(n_565) );
AND2x2_ASAP7_75t_L g609 ( .A(n_514), .B(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g674 ( .A(n_514), .B(n_675), .Y(n_674) );
INVx3_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
AO21x2_ASAP7_75t_L g515 ( .A1(n_516), .A2(n_517), .B(n_523), .Y(n_515) );
AO21x1_ASAP7_75t_SL g537 ( .A1(n_516), .A2(n_517), .B(n_523), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_518), .B(n_522), .Y(n_517) );
AND2x4_ASAP7_75t_L g569 ( .A(n_524), .B(n_570), .Y(n_569) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
OR2x2_ASAP7_75t_L g705 ( .A(n_526), .B(n_650), .Y(n_705) );
AND2x2_ASAP7_75t_L g536 ( .A(n_527), .B(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g573 ( .A(n_527), .Y(n_573) );
HB1xp67_ASAP7_75t_L g590 ( .A(n_527), .Y(n_590) );
INVx2_ASAP7_75t_L g611 ( .A(n_527), .Y(n_611) );
INVx1_ASAP7_75t_L g675 ( .A(n_527), .Y(n_675) );
INVx2_ASAP7_75t_L g757 ( .A(n_534), .Y(n_757) );
OR2x2_ASAP7_75t_L g621 ( .A(n_535), .B(n_598), .Y(n_621) );
INVx2_ASAP7_75t_SL g535 ( .A(n_536), .Y(n_535) );
AND2x2_ASAP7_75t_L g761 ( .A(n_536), .B(n_658), .Y(n_761) );
AND2x2_ASAP7_75t_L g654 ( .A(n_537), .B(n_611), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_539), .B(n_551), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
AOI22xp5_ASAP7_75t_L g745 ( .A1(n_540), .A2(n_668), .B1(n_685), .B2(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx2_ASAP7_75t_L g581 ( .A(n_542), .Y(n_581) );
AND2x2_ASAP7_75t_L g635 ( .A(n_542), .B(n_555), .Y(n_635) );
HB1xp67_ASAP7_75t_L g662 ( .A(n_542), .Y(n_662) );
INVx3_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
HB1xp67_ASAP7_75t_L g630 ( .A(n_543), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_545), .B(n_549), .Y(n_544) );
INVxp67_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_553), .B(n_667), .Y(n_666) );
OAI32xp33_ASAP7_75t_L g683 ( .A1(n_553), .A2(n_684), .A3(n_686), .B1(n_687), .B2(n_689), .Y(n_683) );
BUFx2_ASAP7_75t_L g568 ( .A(n_554), .Y(n_568) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g710 ( .A(n_555), .B(n_604), .Y(n_710) );
OR4x1_ASAP7_75t_L g556 ( .A(n_557), .B(n_560), .C(n_561), .D(n_564), .Y(n_556) );
OAI22xp5_ASAP7_75t_L g741 ( .A1(n_557), .A2(n_648), .B1(n_742), .B2(n_743), .Y(n_741) );
INVx2_ASAP7_75t_SL g557 ( .A(n_558), .Y(n_557) );
HB1xp67_ASAP7_75t_L g750 ( .A(n_558), .Y(n_750) );
AND2x2_ASAP7_75t_L g592 ( .A(n_559), .B(n_593), .Y(n_592) );
BUFx2_ASAP7_75t_L g672 ( .A(n_559), .Y(n_672) );
INVx1_ASAP7_75t_L g688 ( .A(n_559), .Y(n_688) );
INVx1_ASAP7_75t_L g723 ( .A(n_559), .Y(n_723) );
OR2x2_ASAP7_75t_L g680 ( .A(n_560), .B(n_681), .Y(n_680) );
OR2x2_ASAP7_75t_L g724 ( .A(n_560), .B(n_725), .Y(n_724) );
OAI22xp5_ASAP7_75t_L g663 ( .A1(n_561), .A2(n_598), .B1(n_642), .B2(n_661), .Y(n_663) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g707 ( .A(n_562), .B(n_616), .Y(n_707) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
BUFx2_ASAP7_75t_L g574 ( .A(n_563), .Y(n_574) );
NOR2xp67_ASAP7_75t_L g589 ( .A(n_563), .B(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g570 ( .A(n_564), .Y(n_570) );
NAND4xp25_ASAP7_75t_L g697 ( .A(n_564), .B(n_568), .C(n_649), .D(n_661), .Y(n_697) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g734 ( .A(n_565), .Y(n_734) );
AOI22xp5_ASAP7_75t_L g566 ( .A1(n_567), .A2(n_569), .B1(n_571), .B2(n_575), .Y(n_566) );
OAI22xp33_ASAP7_75t_L g717 ( .A1(n_567), .A2(n_568), .B1(n_718), .B2(n_719), .Y(n_717) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVxp67_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_573), .B(n_574), .Y(n_572) );
INVx3_ASAP7_75t_L g596 ( .A(n_573), .Y(n_596) );
AOI32xp33_ASAP7_75t_L g712 ( .A1(n_573), .A2(n_713), .A3(n_717), .B1(n_722), .B2(n_726), .Y(n_712) );
AND2x2_ASAP7_75t_L g575 ( .A(n_576), .B(n_579), .Y(n_575) );
NOR2xp67_ASAP7_75t_L g618 ( .A(n_576), .B(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g671 ( .A(n_576), .B(n_672), .Y(n_671) );
AOI221xp5_ASAP7_75t_L g695 ( .A1(n_576), .A2(n_584), .B1(n_696), .B2(n_701), .C(n_704), .Y(n_695) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
OR2x2_ASAP7_75t_L g628 ( .A(n_577), .B(n_629), .Y(n_628) );
OR2x2_ASAP7_75t_L g743 ( .A(n_577), .B(n_744), .Y(n_743) );
INVx2_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_578), .B(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g585 ( .A(n_580), .Y(n_585) );
AND2x2_ASAP7_75t_L g603 ( .A(n_580), .B(n_604), .Y(n_603) );
AND2x2_ASAP7_75t_L g580 ( .A(n_581), .B(n_582), .Y(n_580) );
INVx1_ASAP7_75t_SL g643 ( .A(n_581), .Y(n_643) );
INVx1_ASAP7_75t_L g627 ( .A(n_582), .Y(n_627) );
AOI22xp5_ASAP7_75t_L g583 ( .A1(n_584), .A2(n_586), .B1(n_592), .B2(n_594), .Y(n_583) );
INVx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
OR2x2_ASAP7_75t_L g729 ( .A(n_585), .B(n_659), .Y(n_729) );
INVx1_ASAP7_75t_SL g586 ( .A(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx2_ASAP7_75t_L g669 ( .A(n_588), .Y(n_669) );
AND2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_591), .Y(n_588) );
AND2x2_ASAP7_75t_L g600 ( .A(n_593), .B(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_593), .B(n_630), .Y(n_629) );
NAND2x1p5_ASAP7_75t_L g642 ( .A(n_593), .B(n_643), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_593), .B(n_635), .Y(n_756) );
AOI22xp33_ASAP7_75t_SL g753 ( .A1(n_594), .A2(n_754), .B1(n_755), .B2(n_757), .Y(n_753) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
OR2x2_ASAP7_75t_L g636 ( .A(n_596), .B(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g646 ( .A(n_596), .B(n_647), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_596), .B(n_658), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_596), .B(n_700), .Y(n_699) );
AND2x4_ASAP7_75t_SL g701 ( .A(n_596), .B(n_702), .Y(n_701) );
INVx2_ASAP7_75t_SL g597 ( .A(n_598), .Y(n_597) );
OR2x2_ASAP7_75t_L g677 ( .A(n_598), .B(n_678), .Y(n_677) );
OAI21xp5_ASAP7_75t_L g599 ( .A1(n_600), .A2(n_602), .B(n_605), .Y(n_599) );
INVx1_ASAP7_75t_L g619 ( .A(n_601), .Y(n_619) );
AOI22xp5_ASAP7_75t_L g638 ( .A1(n_602), .A2(n_639), .B1(n_646), .B2(n_651), .Y(n_638) );
INVx3_ASAP7_75t_L g641 ( .A(n_604), .Y(n_641) );
INVx2_ASAP7_75t_SL g605 ( .A(n_606), .Y(n_605) );
OR2x2_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
OAI32xp33_ASAP7_75t_SL g696 ( .A1(n_607), .A2(n_667), .A3(n_697), .B1(n_698), .B2(n_699), .Y(n_696) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g616 ( .A(n_610), .B(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
NAND4xp25_ASAP7_75t_SL g612 ( .A(n_613), .B(n_638), .C(n_655), .D(n_670), .Y(n_612) );
AOI221xp5_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_618), .B1(n_620), .B2(n_622), .C(n_631), .Y(n_613) );
AND2x2_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
INVx2_ASAP7_75t_L g653 ( .A(n_615), .Y(n_653) );
AND2x2_ASAP7_75t_L g702 ( .A(n_615), .B(n_703), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_615), .B(n_654), .Y(n_740) );
AND2x2_ASAP7_75t_L g751 ( .A(n_615), .B(n_674), .Y(n_751) );
INVx2_ASAP7_75t_L g637 ( .A(n_617), .Y(n_637) );
INVx2_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
OAI21xp5_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_625), .B(n_628), .Y(n_622) );
AND2x2_ASAP7_75t_L g754 ( .A(n_623), .B(n_625), .Y(n_754) );
INVx2_ASAP7_75t_SL g623 ( .A(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_624), .B(n_748), .Y(n_747) );
INVx2_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g731 ( .A(n_629), .Y(n_731) );
INVx1_ASAP7_75t_L g716 ( .A(n_630), .Y(n_716) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_633), .B(n_688), .Y(n_687) );
NOR2x1_ASAP7_75t_L g645 ( .A(n_634), .B(n_641), .Y(n_645) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_SL g744 ( .A(n_635), .Y(n_744) );
INVx1_ASAP7_75t_L g726 ( .A(n_637), .Y(n_726) );
OR2x2_ASAP7_75t_L g742 ( .A(n_637), .B(n_653), .Y(n_742) );
NAND2xp33_ASAP7_75t_SL g639 ( .A(n_640), .B(n_644), .Y(n_639) );
OR2x2_ASAP7_75t_L g640 ( .A(n_641), .B(n_642), .Y(n_640) );
INVx2_ASAP7_75t_L g659 ( .A(n_641), .Y(n_659) );
AND2x2_ASAP7_75t_L g664 ( .A(n_641), .B(n_654), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_641), .B(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g738 ( .A(n_642), .Y(n_738) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
AOI22xp5_ASAP7_75t_L g727 ( .A1(n_647), .A2(n_728), .B1(n_730), .B2(n_732), .Y(n_727) );
INVx1_ASAP7_75t_SL g647 ( .A(n_648), .Y(n_647) );
OR2x2_ASAP7_75t_L g648 ( .A(n_649), .B(n_650), .Y(n_648) );
INVx1_ASAP7_75t_L g692 ( .A(n_650), .Y(n_692) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_653), .B(n_654), .Y(n_652) );
INVx1_ASAP7_75t_L g678 ( .A(n_654), .Y(n_678) );
AOI322xp5_ASAP7_75t_L g655 ( .A1(n_656), .A2(n_659), .A3(n_660), .B1(n_663), .B2(n_664), .C1(n_665), .C2(n_668), .Y(n_655) );
OAI21xp5_ASAP7_75t_SL g706 ( .A1(n_656), .A2(n_707), .B(n_708), .Y(n_706) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
AND2x2_ASAP7_75t_L g673 ( .A(n_658), .B(n_674), .Y(n_673) );
AND2x2_ASAP7_75t_L g730 ( .A(n_659), .B(n_731), .Y(n_730) );
HB1xp67_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx2_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
NOR2xp33_ASAP7_75t_L g704 ( .A(n_666), .B(n_705), .Y(n_704) );
INVx2_ASAP7_75t_L g686 ( .A(n_667), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_667), .B(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
AOI221xp5_ASAP7_75t_L g670 ( .A1(n_671), .A2(n_673), .B1(n_676), .B2(n_679), .C(n_683), .Y(n_670) );
AOI221xp5_ASAP7_75t_L g758 ( .A1(n_672), .A2(n_759), .B1(n_761), .B2(n_762), .C(n_763), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_674), .B(n_685), .Y(n_684) );
BUFx2_ASAP7_75t_L g725 ( .A(n_675), .Y(n_725) );
INVx2_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
OAI21xp5_ASAP7_75t_L g749 ( .A1(n_679), .A2(n_750), .B(n_751), .Y(n_749) );
INVx1_ASAP7_75t_SL g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
NAND2xp33_ASAP7_75t_SL g759 ( .A(n_688), .B(n_760), .Y(n_759) );
INVx3_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
AND2x4_ASAP7_75t_L g690 ( .A(n_691), .B(n_692), .Y(n_690) );
NOR4xp75_ASAP7_75t_L g693 ( .A(n_694), .B(n_711), .C(n_735), .D(n_752), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_695), .B(n_706), .Y(n_694) );
INVx1_ASAP7_75t_L g765 ( .A(n_703), .Y(n_765) );
INVx1_ASAP7_75t_SL g708 ( .A(n_709), .Y(n_708) );
AND2x2_ASAP7_75t_L g737 ( .A(n_710), .B(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g764 ( .A(n_710), .Y(n_764) );
NAND2xp5_ASAP7_75t_SL g711 ( .A(n_712), .B(n_727), .Y(n_711) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
NOR2xp33_ASAP7_75t_L g722 ( .A(n_723), .B(n_724), .Y(n_722) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx2_ASAP7_75t_SL g760 ( .A(n_731), .Y(n_760) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
NAND3x1_ASAP7_75t_L g735 ( .A(n_736), .B(n_745), .C(n_749), .Y(n_735) );
AOI21xp5_ASAP7_75t_L g736 ( .A1(n_737), .A2(n_739), .B(n_741), .Y(n_736) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVxp67_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_753), .B(n_758), .Y(n_752) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
CKINVDCx5p33_ASAP7_75t_R g768 ( .A(n_769), .Y(n_768) );
INVx1_ASAP7_75t_SL g780 ( .A(n_769), .Y(n_780) );
CKINVDCx11_ASAP7_75t_R g769 ( .A(n_770), .Y(n_769) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
INVx1_ASAP7_75t_SL g782 ( .A(n_783), .Y(n_782) );
INVx2_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
endmodule