module fake_netlist_1_10254_n_37 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_37);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_37;
wire n_20;
wire n_36;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVxp33_ASAP7_75t_SL g11 ( .A(n_1), .Y(n_11) );
CKINVDCx20_ASAP7_75t_R g12 ( .A(n_3), .Y(n_12) );
INVx2_ASAP7_75t_L g13 ( .A(n_8), .Y(n_13) );
CKINVDCx20_ASAP7_75t_R g14 ( .A(n_4), .Y(n_14) );
CKINVDCx20_ASAP7_75t_R g15 ( .A(n_1), .Y(n_15) );
INVx2_ASAP7_75t_L g16 ( .A(n_3), .Y(n_16) );
INVx4_ASAP7_75t_L g17 ( .A(n_13), .Y(n_17) );
AND3x1_ASAP7_75t_L g18 ( .A(n_16), .B(n_0), .C(n_2), .Y(n_18) );
INVx4_ASAP7_75t_L g19 ( .A(n_13), .Y(n_19) );
INVx2_ASAP7_75t_L g20 ( .A(n_12), .Y(n_20) );
AOI22xp33_ASAP7_75t_SL g21 ( .A1(n_20), .A2(n_11), .B1(n_15), .B2(n_14), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_17), .Y(n_22) );
CKINVDCx8_ASAP7_75t_R g23 ( .A(n_18), .Y(n_23) );
AOI22xp33_ASAP7_75t_L g24 ( .A1(n_22), .A2(n_17), .B1(n_19), .B2(n_18), .Y(n_24) );
OAI22xp5_ASAP7_75t_L g25 ( .A1(n_23), .A2(n_19), .B1(n_2), .B2(n_4), .Y(n_25) );
NAND2xp5_ASAP7_75t_L g26 ( .A(n_24), .B(n_23), .Y(n_26) );
AND2x2_ASAP7_75t_L g27 ( .A(n_25), .B(n_21), .Y(n_27) );
NOR2x1_ASAP7_75t_L g28 ( .A(n_26), .B(n_0), .Y(n_28) );
INVx1_ASAP7_75t_SL g29 ( .A(n_27), .Y(n_29) );
AOI22xp33_ASAP7_75t_SL g30 ( .A1(n_29), .A2(n_27), .B1(n_6), .B2(n_7), .Y(n_30) );
NOR2xp33_ASAP7_75t_L g31 ( .A(n_28), .B(n_5), .Y(n_31) );
AOI21xp5_ASAP7_75t_L g32 ( .A1(n_28), .A2(n_9), .B(n_10), .Y(n_32) );
NOR2x1p5_ASAP7_75t_L g33 ( .A(n_30), .B(n_5), .Y(n_33) );
BUFx2_ASAP7_75t_L g34 ( .A(n_31), .Y(n_34) );
BUFx2_ASAP7_75t_L g35 ( .A(n_32), .Y(n_35) );
INVx2_ASAP7_75t_L g36 ( .A(n_33), .Y(n_36) );
AOI22xp33_ASAP7_75t_L g37 ( .A1(n_36), .A2(n_35), .B1(n_34), .B2(n_7), .Y(n_37) );
endmodule