module fake_netlist_6_1917_n_901 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_223, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_226, n_228, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_227, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_233, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_234, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_231, n_65, n_230, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_229, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_232, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_901);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_223;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_226;
input n_228;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_227;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_233;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_234;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_231;
input n_65;
input n_230;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_229;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_232;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_901;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_881;
wire n_875;
wire n_465;
wire n_367;
wire n_760;
wire n_741;
wire n_680;
wire n_590;
wire n_625;
wire n_661;
wire n_278;
wire n_362;
wire n_341;
wire n_828;
wire n_462;
wire n_607;
wire n_726;
wire n_671;
wire n_316;
wire n_419;
wire n_304;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_783;
wire n_725;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_628;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_617;
wire n_698;
wire n_898;
wire n_845;
wire n_255;
wire n_807;
wire n_739;
wire n_400;
wire n_284;
wire n_337;
wire n_865;
wire n_893;
wire n_485;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_573;
wire n_769;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_669;
wire n_447;
wire n_872;
wire n_300;
wire n_718;
wire n_248;
wire n_517;
wire n_747;
wire n_852;
wire n_667;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_822;
wire n_693;
wire n_758;
wire n_516;
wire n_631;
wire n_720;
wire n_842;
wire n_525;
wire n_611;
wire n_491;
wire n_878;
wire n_772;
wire n_656;
wire n_843;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_343;
wire n_844;
wire n_448;
wire n_886;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_888;
wire n_454;
wire n_638;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_887;
wire n_752;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_803;
wire n_290;
wire n_809;
wire n_839;
wire n_734;
wire n_708;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_800;
wire n_460;
wire n_854;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_777;
wire n_407;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_650;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_552;
wire n_619;
wire n_885;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_394;
wire n_312;
wire n_519;
wire n_541;
wire n_512;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_792;
wire n_880;
wire n_476;
wire n_714;
wire n_291;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_821;
wire n_325;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_806;
wire n_864;
wire n_879;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_833;
wire n_523;
wire n_322;
wire n_707;
wire n_409;
wire n_345;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_386;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_550;
wire n_487;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_811;
wire n_882;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_299;
wire n_518;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_247;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_285;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_286;
wire n_254;
wire n_834;
wire n_242;
wire n_835;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_816;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_604;
wire n_848;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_722;
wire n_688;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_629;
wire n_388;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_841;
wire n_531;
wire n_827;
wire n_361;
wire n_508;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_664;
wire n_678;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_163),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_154),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_77),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_24),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_177),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_198),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_227),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_233),
.Y(n_242)
);

INVx1_ASAP7_75t_SL g243 ( 
.A(n_221),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_148),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_28),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_145),
.Y(n_246)
);

BUFx10_ASAP7_75t_L g247 ( 
.A(n_116),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_33),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_185),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_135),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_107),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_65),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_42),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_196),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_228),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_195),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_24),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_157),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_100),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_216),
.Y(n_260)
);

BUFx5_ASAP7_75t_L g261 ( 
.A(n_155),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_207),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_210),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_17),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_6),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_66),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_104),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_74),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_170),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_161),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_86),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_43),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_29),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g274 ( 
.A(n_29),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_51),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_92),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_169),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_30),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_87),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_118),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_202),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_225),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_115),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_186),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_125),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_213),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_192),
.Y(n_287)
);

BUFx10_ASAP7_75t_L g288 ( 
.A(n_56),
.Y(n_288)
);

BUFx10_ASAP7_75t_L g289 ( 
.A(n_113),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_212),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_12),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_194),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_62),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_20),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_26),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_139),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_83),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_180),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_165),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_162),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_108),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_72),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_168),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_159),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_201),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_124),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_173),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_226),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_134),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_80),
.Y(n_310)
);

BUFx8_ASAP7_75t_SL g311 ( 
.A(n_175),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_193),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_17),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_91),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_119),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_70),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_90),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_214),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_120),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_122),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_130),
.Y(n_321)
);

BUFx5_ASAP7_75t_L g322 ( 
.A(n_6),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_69),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_7),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_8),
.Y(n_325)
);

BUFx5_ASAP7_75t_L g326 ( 
.A(n_189),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_143),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_85),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_158),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_95),
.Y(n_330)
);

BUFx5_ASAP7_75t_L g331 ( 
.A(n_10),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_99),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_111),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_103),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_82),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_112),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_204),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_47),
.Y(n_338)
);

HB1xp67_ASAP7_75t_L g339 ( 
.A(n_147),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_156),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_136),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_52),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_231),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_41),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_133),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_32),
.Y(n_346)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_73),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_234),
.Y(n_348)
);

BUFx3_ASAP7_75t_L g349 ( 
.A(n_67),
.Y(n_349)
);

INVx1_ASAP7_75t_SL g350 ( 
.A(n_187),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_200),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_224),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_3),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_166),
.Y(n_354)
);

INVx1_ASAP7_75t_SL g355 ( 
.A(n_121),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_3),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_190),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_149),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_76),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_218),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_151),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_146),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_8),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_178),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_176),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_142),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_206),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_102),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_28),
.Y(n_369)
);

BUFx8_ASAP7_75t_SL g370 ( 
.A(n_164),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_229),
.Y(n_371)
);

BUFx3_ASAP7_75t_L g372 ( 
.A(n_39),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_197),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_117),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_50),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_150),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_211),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_30),
.Y(n_378)
);

BUFx10_ASAP7_75t_L g379 ( 
.A(n_128),
.Y(n_379)
);

BUFx2_ASAP7_75t_L g380 ( 
.A(n_54),
.Y(n_380)
);

HB1xp67_ASAP7_75t_L g381 ( 
.A(n_205),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_55),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_172),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_94),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_21),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_220),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_59),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_36),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_10),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_167),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_209),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_98),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_184),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_171),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_0),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_191),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_106),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_105),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_127),
.Y(n_399)
);

INVx4_ASAP7_75t_R g400 ( 
.A(n_137),
.Y(n_400)
);

INVx5_ASAP7_75t_L g401 ( 
.A(n_306),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_380),
.B(n_0),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_274),
.B(n_1),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_306),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_322),
.Y(n_405)
);

NOR2x1_ASAP7_75t_L g406 ( 
.A(n_270),
.B(n_37),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_322),
.Y(n_407)
);

AND2x4_ASAP7_75t_L g408 ( 
.A(n_285),
.B(n_1),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_311),
.Y(n_409)
);

BUFx12f_ASAP7_75t_L g410 ( 
.A(n_247),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_339),
.B(n_2),
.Y(n_411)
);

BUFx12f_ASAP7_75t_L g412 ( 
.A(n_288),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_306),
.Y(n_413)
);

BUFx12f_ASAP7_75t_L g414 ( 
.A(n_288),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_322),
.Y(n_415)
);

AND2x4_ASAP7_75t_L g416 ( 
.A(n_349),
.B(n_2),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_322),
.Y(n_417)
);

OR2x2_ASAP7_75t_L g418 ( 
.A(n_248),
.B(n_4),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_322),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_372),
.B(n_4),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_306),
.Y(n_421)
);

AND2x6_ASAP7_75t_L g422 ( 
.A(n_357),
.B(n_38),
.Y(n_422)
);

BUFx8_ASAP7_75t_SL g423 ( 
.A(n_370),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_300),
.B(n_5),
.Y(n_424)
);

BUFx12f_ASAP7_75t_L g425 ( 
.A(n_289),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_347),
.B(n_5),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_357),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_357),
.Y(n_428)
);

BUFx8_ASAP7_75t_L g429 ( 
.A(n_322),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_296),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_331),
.Y(n_431)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_238),
.Y(n_432)
);

BUFx8_ASAP7_75t_SL g433 ( 
.A(n_369),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_381),
.B(n_7),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_331),
.B(n_9),
.Y(n_435)
);

AND2x4_ASAP7_75t_L g436 ( 
.A(n_305),
.B(n_9),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_331),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_331),
.B(n_11),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_331),
.Y(n_439)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_273),
.Y(n_440)
);

INVx3_ASAP7_75t_L g441 ( 
.A(n_289),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_243),
.B(n_11),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_310),
.Y(n_443)
);

INVx4_ASAP7_75t_L g444 ( 
.A(n_235),
.Y(n_444)
);

BUFx2_ASAP7_75t_L g445 ( 
.A(n_245),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_333),
.B(n_12),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g447 ( 
.A(n_379),
.B(n_388),
.Y(n_447)
);

INVx5_ASAP7_75t_L g448 ( 
.A(n_352),
.Y(n_448)
);

INVx5_ASAP7_75t_L g449 ( 
.A(n_358),
.Y(n_449)
);

OR2x2_ASAP7_75t_L g450 ( 
.A(n_291),
.B(n_13),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_260),
.B(n_13),
.Y(n_451)
);

HB1xp67_ASAP7_75t_L g452 ( 
.A(n_257),
.Y(n_452)
);

BUFx12f_ASAP7_75t_L g453 ( 
.A(n_265),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_261),
.B(n_326),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_295),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_261),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_389),
.B(n_14),
.Y(n_457)
);

BUFx2_ASAP7_75t_L g458 ( 
.A(n_278),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_264),
.B(n_14),
.Y(n_459)
);

AND2x6_ASAP7_75t_L g460 ( 
.A(n_236),
.B(n_40),
.Y(n_460)
);

AND2x4_ASAP7_75t_L g461 ( 
.A(n_239),
.B(n_242),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_313),
.Y(n_462)
);

BUFx2_ASAP7_75t_L g463 ( 
.A(n_294),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_261),
.B(n_15),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_266),
.B(n_15),
.Y(n_465)
);

AND2x4_ASAP7_75t_L g466 ( 
.A(n_246),
.B(n_16),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_261),
.B(n_16),
.Y(n_467)
);

BUFx6f_ASAP7_75t_L g468 ( 
.A(n_249),
.Y(n_468)
);

INVx5_ASAP7_75t_L g469 ( 
.A(n_261),
.Y(n_469)
);

NOR2x1_ASAP7_75t_L g470 ( 
.A(n_251),
.B(n_44),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_346),
.B(n_18),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_268),
.B(n_18),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_350),
.B(n_19),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_261),
.B(n_19),
.Y(n_474)
);

BUFx6f_ASAP7_75t_L g475 ( 
.A(n_253),
.Y(n_475)
);

BUFx8_ASAP7_75t_L g476 ( 
.A(n_324),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_325),
.Y(n_477)
);

NOR2x1_ASAP7_75t_L g478 ( 
.A(n_259),
.B(n_45),
.Y(n_478)
);

AND2x4_ASAP7_75t_L g479 ( 
.A(n_263),
.B(n_20),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_363),
.B(n_21),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_271),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_395),
.B(n_22),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_SL g483 ( 
.A(n_355),
.B(n_23),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_326),
.B(n_23),
.Y(n_484)
);

BUFx2_ASAP7_75t_L g485 ( 
.A(n_353),
.Y(n_485)
);

BUFx8_ASAP7_75t_L g486 ( 
.A(n_356),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_276),
.Y(n_487)
);

INVx4_ASAP7_75t_L g488 ( 
.A(n_237),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_277),
.Y(n_489)
);

INVx5_ASAP7_75t_L g490 ( 
.A(n_326),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_282),
.Y(n_491)
);

AND2x4_ASAP7_75t_L g492 ( 
.A(n_283),
.B(n_25),
.Y(n_492)
);

BUFx12f_ASAP7_75t_L g493 ( 
.A(n_240),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_326),
.B(n_25),
.Y(n_494)
);

BUFx2_ASAP7_75t_L g495 ( 
.A(n_378),
.Y(n_495)
);

HB1xp67_ASAP7_75t_L g496 ( 
.A(n_385),
.Y(n_496)
);

AND2x4_ASAP7_75t_L g497 ( 
.A(n_293),
.B(n_26),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_424),
.A2(n_292),
.B1(n_327),
.B2(n_267),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_427),
.Y(n_499)
);

BUFx10_ASAP7_75t_L g500 ( 
.A(n_409),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_427),
.Y(n_501)
);

AO22x2_ASAP7_75t_L g502 ( 
.A1(n_434),
.A2(n_408),
.B1(n_416),
.B2(n_436),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_402),
.A2(n_361),
.B1(n_391),
.B2(n_337),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_423),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_411),
.A2(n_244),
.B1(n_250),
.B2(n_241),
.Y(n_505)
);

OAI22xp33_ASAP7_75t_L g506 ( 
.A1(n_483),
.A2(n_308),
.B1(n_317),
.B2(n_302),
.Y(n_506)
);

AO22x2_ASAP7_75t_L g507 ( 
.A1(n_408),
.A2(n_321),
.B1(n_330),
.B2(n_318),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_428),
.Y(n_508)
);

INVx4_ASAP7_75t_L g509 ( 
.A(n_493),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_447),
.B(n_252),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_403),
.A2(n_255),
.B1(n_256),
.B2(n_254),
.Y(n_511)
);

OAI22xp33_ASAP7_75t_L g512 ( 
.A1(n_426),
.A2(n_338),
.B1(n_354),
.B2(n_335),
.Y(n_512)
);

AO22x2_ASAP7_75t_L g513 ( 
.A1(n_416),
.A2(n_375),
.B1(n_382),
.B2(n_373),
.Y(n_513)
);

AND2x2_ASAP7_75t_SL g514 ( 
.A(n_459),
.B(n_384),
.Y(n_514)
);

OAI22xp33_ASAP7_75t_SL g515 ( 
.A1(n_441),
.A2(n_387),
.B1(n_390),
.B2(n_386),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_452),
.B(n_258),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_442),
.A2(n_465),
.B1(n_472),
.B2(n_451),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_445),
.B(n_262),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_473),
.A2(n_342),
.B1(n_399),
.B2(n_398),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_SL g520 ( 
.A1(n_418),
.A2(n_345),
.B1(n_272),
.B2(n_275),
.Y(n_520)
);

AND2x4_ASAP7_75t_L g521 ( 
.A(n_420),
.B(n_269),
.Y(n_521)
);

AO22x2_ASAP7_75t_L g522 ( 
.A1(n_436),
.A2(n_400),
.B1(n_31),
.B2(n_32),
.Y(n_522)
);

INVx1_ASAP7_75t_SL g523 ( 
.A(n_433),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_458),
.B(n_279),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_453),
.A2(n_343),
.B1(n_396),
.B2(n_394),
.Y(n_525)
);

OAI22xp33_ASAP7_75t_L g526 ( 
.A1(n_450),
.A2(n_397),
.B1(n_393),
.B2(n_392),
.Y(n_526)
);

INVx3_ASAP7_75t_L g527 ( 
.A(n_430),
.Y(n_527)
);

OR2x2_ASAP7_75t_L g528 ( 
.A(n_463),
.B(n_27),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_L g529 ( 
.A1(n_471),
.A2(n_383),
.B1(n_377),
.B2(n_376),
.Y(n_529)
);

AO22x2_ASAP7_75t_L g530 ( 
.A1(n_466),
.A2(n_27),
.B1(n_33),
.B2(n_34),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g531 ( 
.A1(n_480),
.A2(n_280),
.B1(n_374),
.B2(n_371),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_444),
.B(n_281),
.Y(n_532)
);

AO22x2_ASAP7_75t_L g533 ( 
.A1(n_466),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_533)
);

AO22x2_ASAP7_75t_L g534 ( 
.A1(n_479),
.A2(n_35),
.B1(n_326),
.B2(n_368),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_428),
.Y(n_535)
);

OAI22xp33_ASAP7_75t_SL g536 ( 
.A1(n_464),
.A2(n_367),
.B1(n_366),
.B2(n_365),
.Y(n_536)
);

AOI22xp5_ASAP7_75t_L g537 ( 
.A1(n_482),
.A2(n_364),
.B1(n_362),
.B2(n_360),
.Y(n_537)
);

INVx3_ASAP7_75t_L g538 ( 
.A(n_430),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_404),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_L g540 ( 
.A1(n_457),
.A2(n_315),
.B1(n_351),
.B2(n_348),
.Y(n_540)
);

AO22x2_ASAP7_75t_L g541 ( 
.A1(n_479),
.A2(n_359),
.B1(n_344),
.B2(n_341),
.Y(n_541)
);

AO22x2_ASAP7_75t_L g542 ( 
.A1(n_492),
.A2(n_340),
.B1(n_336),
.B2(n_334),
.Y(n_542)
);

AOI22xp5_ASAP7_75t_L g543 ( 
.A1(n_410),
.A2(n_332),
.B1(n_329),
.B2(n_328),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_488),
.B(n_284),
.Y(n_544)
);

INVx1_ASAP7_75t_SL g545 ( 
.A(n_412),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_430),
.Y(n_546)
);

AOI22xp5_ASAP7_75t_L g547 ( 
.A1(n_414),
.A2(n_323),
.B1(n_320),
.B2(n_319),
.Y(n_547)
);

OAI22xp33_ASAP7_75t_L g548 ( 
.A1(n_435),
.A2(n_316),
.B1(n_314),
.B2(n_312),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_485),
.B(n_286),
.Y(n_549)
);

AOI22xp5_ASAP7_75t_L g550 ( 
.A1(n_425),
.A2(n_309),
.B1(n_307),
.B2(n_304),
.Y(n_550)
);

AOI22xp5_ASAP7_75t_L g551 ( 
.A1(n_492),
.A2(n_301),
.B1(n_299),
.B2(n_298),
.Y(n_551)
);

OR2x2_ASAP7_75t_L g552 ( 
.A(n_495),
.B(n_287),
.Y(n_552)
);

OAI22xp33_ASAP7_75t_L g553 ( 
.A1(n_438),
.A2(n_303),
.B1(n_297),
.B2(n_290),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_413),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_497),
.B(n_46),
.Y(n_555)
);

OAI22xp33_ASAP7_75t_SL g556 ( 
.A1(n_467),
.A2(n_48),
.B1(n_49),
.B2(n_53),
.Y(n_556)
);

OAI22xp33_ASAP7_75t_R g557 ( 
.A1(n_496),
.A2(n_57),
.B1(n_58),
.B2(n_60),
.Y(n_557)
);

AOI22x1_ASAP7_75t_SL g558 ( 
.A1(n_455),
.A2(n_61),
.B1(n_63),
.B2(n_64),
.Y(n_558)
);

OAI22xp33_ASAP7_75t_SL g559 ( 
.A1(n_474),
.A2(n_68),
.B1(n_71),
.B2(n_75),
.Y(n_559)
);

AND2x2_ASAP7_75t_SL g560 ( 
.A(n_497),
.B(n_78),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_461),
.B(n_79),
.Y(n_561)
);

HB1xp67_ASAP7_75t_L g562 ( 
.A(n_552),
.Y(n_562)
);

INVx2_ASAP7_75t_SL g563 ( 
.A(n_549),
.Y(n_563)
);

AOI21xp5_ASAP7_75t_L g564 ( 
.A1(n_502),
.A2(n_514),
.B(n_461),
.Y(n_564)
);

AOI21xp5_ASAP7_75t_L g565 ( 
.A1(n_502),
.A2(n_454),
.B(n_437),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_527),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_555),
.B(n_405),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_538),
.Y(n_568)
);

XNOR2xp5_ASAP7_75t_L g569 ( 
.A(n_503),
.B(n_406),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_546),
.Y(n_570)
);

INVx2_ASAP7_75t_SL g571 ( 
.A(n_518),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_517),
.B(n_446),
.Y(n_572)
);

XNOR2xp5_ASAP7_75t_L g573 ( 
.A(n_498),
.B(n_523),
.Y(n_573)
);

INVx2_ASAP7_75t_SL g574 ( 
.A(n_524),
.Y(n_574)
);

NOR2xp67_ASAP7_75t_L g575 ( 
.A(n_519),
.B(n_401),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_539),
.Y(n_576)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_510),
.B(n_432),
.Y(n_577)
);

INVxp67_ASAP7_75t_SL g578 ( 
.A(n_554),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_516),
.B(n_440),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_526),
.B(n_468),
.Y(n_580)
);

XOR2xp5_ASAP7_75t_L g581 ( 
.A(n_504),
.B(n_470),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_505),
.B(n_468),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_499),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_501),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_508),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_535),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_561),
.Y(n_587)
);

AND2x4_ASAP7_75t_L g588 ( 
.A(n_521),
.B(n_462),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g589 ( 
.A(n_521),
.B(n_477),
.Y(n_589)
);

OAI21xp5_ASAP7_75t_L g590 ( 
.A1(n_560),
.A2(n_460),
.B(n_494),
.Y(n_590)
);

XOR2xp5_ASAP7_75t_L g591 ( 
.A(n_525),
.B(n_478),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_507),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_513),
.Y(n_593)
);

AOI21xp5_ASAP7_75t_L g594 ( 
.A1(n_515),
.A2(n_419),
.B(n_407),
.Y(n_594)
);

AND2x4_ASAP7_75t_L g595 ( 
.A(n_528),
.B(n_460),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_532),
.B(n_415),
.Y(n_596)
);

CKINVDCx20_ASAP7_75t_R g597 ( 
.A(n_500),
.Y(n_597)
);

BUFx2_ASAP7_75t_R g598 ( 
.A(n_530),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_522),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_522),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_530),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_533),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_533),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_544),
.B(n_417),
.Y(n_604)
);

INVx3_ASAP7_75t_L g605 ( 
.A(n_534),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_520),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_511),
.B(n_443),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_534),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_529),
.B(n_475),
.Y(n_609)
);

AND2x6_ASAP7_75t_L g610 ( 
.A(n_551),
.B(n_484),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_559),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_541),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_531),
.B(n_475),
.Y(n_613)
);

INVx2_ASAP7_75t_SL g614 ( 
.A(n_541),
.Y(n_614)
);

AND2x4_ASAP7_75t_L g615 ( 
.A(n_543),
.B(n_460),
.Y(n_615)
);

INVxp33_ASAP7_75t_L g616 ( 
.A(n_542),
.Y(n_616)
);

NOR2xp67_ASAP7_75t_L g617 ( 
.A(n_547),
.B(n_401),
.Y(n_617)
);

INVx3_ASAP7_75t_L g618 ( 
.A(n_542),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_556),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_540),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_537),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_548),
.B(n_431),
.Y(n_622)
);

XNOR2x2_ASAP7_75t_L g623 ( 
.A(n_557),
.B(n_476),
.Y(n_623)
);

CKINVDCx20_ASAP7_75t_R g624 ( 
.A(n_550),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_506),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_512),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_536),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_545),
.Y(n_628)
);

BUFx6f_ASAP7_75t_L g629 ( 
.A(n_576),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_579),
.B(n_509),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_572),
.B(n_460),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_577),
.B(n_481),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_563),
.B(n_481),
.Y(n_633)
);

INVx2_ASAP7_75t_SL g634 ( 
.A(n_571),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_574),
.B(n_481),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_562),
.B(n_487),
.Y(n_636)
);

BUFx6f_ASAP7_75t_L g637 ( 
.A(n_576),
.Y(n_637)
);

INVx3_ASAP7_75t_L g638 ( 
.A(n_576),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_567),
.B(n_553),
.Y(n_639)
);

INVx1_ASAP7_75t_SL g640 ( 
.A(n_628),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_589),
.B(n_487),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_595),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_595),
.Y(n_643)
);

OR2x2_ASAP7_75t_L g644 ( 
.A(n_625),
.B(n_487),
.Y(n_644)
);

INVx1_ASAP7_75t_SL g645 ( 
.A(n_598),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_620),
.B(n_489),
.Y(n_646)
);

NAND2x1p5_ASAP7_75t_L g647 ( 
.A(n_605),
.B(n_615),
.Y(n_647)
);

AND2x4_ASAP7_75t_L g648 ( 
.A(n_588),
.B(n_439),
.Y(n_648)
);

BUFx3_ASAP7_75t_L g649 ( 
.A(n_597),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_567),
.B(n_456),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_596),
.B(n_422),
.Y(n_651)
);

NOR2xp67_ASAP7_75t_R g652 ( 
.A(n_606),
.B(n_558),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_578),
.Y(n_653)
);

BUFx6f_ASAP7_75t_L g654 ( 
.A(n_615),
.Y(n_654)
);

INVx4_ASAP7_75t_L g655 ( 
.A(n_605),
.Y(n_655)
);

BUFx6f_ASAP7_75t_L g656 ( 
.A(n_570),
.Y(n_656)
);

OAI21x1_ASAP7_75t_L g657 ( 
.A1(n_565),
.A2(n_422),
.B(n_429),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_609),
.B(n_489),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_596),
.B(n_422),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_613),
.B(n_491),
.Y(n_660)
);

INVxp67_ASAP7_75t_L g661 ( 
.A(n_580),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_607),
.B(n_582),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_578),
.Y(n_663)
);

INVx2_ASAP7_75t_SL g664 ( 
.A(n_627),
.Y(n_664)
);

INVxp67_ASAP7_75t_L g665 ( 
.A(n_604),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_587),
.B(n_491),
.Y(n_666)
);

INVx1_ASAP7_75t_SL g667 ( 
.A(n_581),
.Y(n_667)
);

BUFx5_ASAP7_75t_L g668 ( 
.A(n_611),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_590),
.B(n_491),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_626),
.B(n_448),
.Y(n_670)
);

AND2x6_ASAP7_75t_L g671 ( 
.A(n_619),
.B(n_421),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_590),
.B(n_421),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_565),
.B(n_421),
.Y(n_673)
);

AND2x2_ASAP7_75t_SL g674 ( 
.A(n_599),
.B(n_81),
.Y(n_674)
);

BUFx4f_ASAP7_75t_L g675 ( 
.A(n_610),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_583),
.Y(n_676)
);

HB1xp67_ASAP7_75t_L g677 ( 
.A(n_592),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_584),
.Y(n_678)
);

AND2x6_ASAP7_75t_L g679 ( 
.A(n_608),
.B(n_84),
.Y(n_679)
);

HB1xp67_ASAP7_75t_L g680 ( 
.A(n_593),
.Y(n_680)
);

OAI21xp5_ASAP7_75t_L g681 ( 
.A1(n_564),
.A2(n_490),
.B(n_469),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_621),
.B(n_476),
.Y(n_682)
);

BUFx2_ASAP7_75t_L g683 ( 
.A(n_610),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_585),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_569),
.B(n_449),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_586),
.Y(n_686)
);

BUFx6f_ASAP7_75t_L g687 ( 
.A(n_622),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_600),
.B(n_469),
.Y(n_688)
);

OR2x2_ASAP7_75t_L g689 ( 
.A(n_640),
.B(n_661),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_636),
.B(n_616),
.Y(n_690)
);

OR2x2_ASAP7_75t_L g691 ( 
.A(n_661),
.B(n_614),
.Y(n_691)
);

NAND2x1p5_ASAP7_75t_L g692 ( 
.A(n_642),
.B(n_618),
.Y(n_692)
);

BUFx5_ASAP7_75t_L g693 ( 
.A(n_679),
.Y(n_693)
);

OR2x6_ASAP7_75t_L g694 ( 
.A(n_683),
.B(n_612),
.Y(n_694)
);

CKINVDCx20_ASAP7_75t_R g695 ( 
.A(n_667),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_642),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_642),
.Y(n_697)
);

OR2x2_ASAP7_75t_L g698 ( 
.A(n_644),
.B(n_601),
.Y(n_698)
);

BUFx8_ASAP7_75t_L g699 ( 
.A(n_649),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_642),
.Y(n_700)
);

AO21x2_ASAP7_75t_L g701 ( 
.A1(n_669),
.A2(n_594),
.B(n_575),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_665),
.B(n_687),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_665),
.B(n_610),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_662),
.B(n_602),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_653),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_643),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_633),
.B(n_618),
.Y(n_707)
);

BUFx6f_ASAP7_75t_L g708 ( 
.A(n_643),
.Y(n_708)
);

BUFx12f_ASAP7_75t_L g709 ( 
.A(n_634),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_635),
.B(n_603),
.Y(n_710)
);

NOR2x1p5_ASAP7_75t_L g711 ( 
.A(n_630),
.B(n_623),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_663),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_685),
.B(n_573),
.Y(n_713)
);

AND2x4_ASAP7_75t_L g714 ( 
.A(n_648),
.B(n_617),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_676),
.Y(n_715)
);

CKINVDCx6p67_ASAP7_75t_R g716 ( 
.A(n_645),
.Y(n_716)
);

AND2x2_ASAP7_75t_SL g717 ( 
.A(n_674),
.B(n_610),
.Y(n_717)
);

OR2x6_ASAP7_75t_L g718 ( 
.A(n_654),
.B(n_594),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_687),
.B(n_591),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_658),
.B(n_566),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_660),
.B(n_568),
.Y(n_721)
);

AND2x4_ASAP7_75t_L g722 ( 
.A(n_648),
.B(n_624),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_655),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_687),
.B(n_650),
.Y(n_724)
);

AND2x4_ASAP7_75t_L g725 ( 
.A(n_654),
.B(n_88),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_675),
.Y(n_726)
);

BUFx2_ASAP7_75t_L g727 ( 
.A(n_654),
.Y(n_727)
);

NAND2x1p5_ASAP7_75t_L g728 ( 
.A(n_654),
.B(n_655),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_678),
.Y(n_729)
);

HB1xp67_ASAP7_75t_L g730 ( 
.A(n_677),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_684),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_SL g732 ( 
.A(n_674),
.B(n_675),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_695),
.Y(n_733)
);

BUFx3_ASAP7_75t_L g734 ( 
.A(n_727),
.Y(n_734)
);

BUFx3_ASAP7_75t_L g735 ( 
.A(n_725),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_723),
.Y(n_736)
);

BUFx2_ASAP7_75t_SL g737 ( 
.A(n_693),
.Y(n_737)
);

INVx1_ASAP7_75t_SL g738 ( 
.A(n_689),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_724),
.Y(n_739)
);

BUFx12f_ASAP7_75t_L g740 ( 
.A(n_699),
.Y(n_740)
);

BUFx3_ASAP7_75t_L g741 ( 
.A(n_725),
.Y(n_741)
);

INVx3_ASAP7_75t_L g742 ( 
.A(n_708),
.Y(n_742)
);

BUFx3_ASAP7_75t_L g743 ( 
.A(n_708),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_705),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_724),
.Y(n_745)
);

INVx3_ASAP7_75t_L g746 ( 
.A(n_708),
.Y(n_746)
);

AND2x2_ASAP7_75t_L g747 ( 
.A(n_702),
.B(n_647),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_712),
.Y(n_748)
);

AND2x4_ASAP7_75t_L g749 ( 
.A(n_696),
.B(n_664),
.Y(n_749)
);

BUFx3_ASAP7_75t_L g750 ( 
.A(n_708),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_702),
.B(n_647),
.Y(n_751)
);

INVx2_ASAP7_75t_SL g752 ( 
.A(n_696),
.Y(n_752)
);

BUFx2_ASAP7_75t_L g753 ( 
.A(n_694),
.Y(n_753)
);

BUFx3_ASAP7_75t_L g754 ( 
.A(n_694),
.Y(n_754)
);

BUFx4f_ASAP7_75t_SL g755 ( 
.A(n_709),
.Y(n_755)
);

INVx3_ASAP7_75t_L g756 ( 
.A(n_728),
.Y(n_756)
);

AOI22xp5_ASAP7_75t_L g757 ( 
.A1(n_717),
.A2(n_639),
.B1(n_668),
.B2(n_646),
.Y(n_757)
);

BUFx12f_ASAP7_75t_L g758 ( 
.A(n_699),
.Y(n_758)
);

INVx8_ASAP7_75t_L g759 ( 
.A(n_718),
.Y(n_759)
);

INVx1_ASAP7_75t_SL g760 ( 
.A(n_690),
.Y(n_760)
);

BUFx3_ASAP7_75t_L g761 ( 
.A(n_694),
.Y(n_761)
);

AOI22xp33_ASAP7_75t_SL g762 ( 
.A1(n_735),
.A2(n_732),
.B1(n_719),
.B2(n_682),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_744),
.Y(n_763)
);

BUFx6f_ASAP7_75t_L g764 ( 
.A(n_743),
.Y(n_764)
);

AOI22xp33_ASAP7_75t_L g765 ( 
.A1(n_757),
.A2(n_703),
.B1(n_719),
.B2(n_704),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_739),
.B(n_707),
.Y(n_766)
);

AOI22xp33_ASAP7_75t_L g767 ( 
.A1(n_739),
.A2(n_679),
.B1(n_711),
.B2(n_646),
.Y(n_767)
);

INVx6_ASAP7_75t_L g768 ( 
.A(n_734),
.Y(n_768)
);

AND2x2_ASAP7_75t_L g769 ( 
.A(n_760),
.B(n_738),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_748),
.Y(n_770)
);

CKINVDCx20_ASAP7_75t_R g771 ( 
.A(n_733),
.Y(n_771)
);

BUFx4f_ASAP7_75t_SL g772 ( 
.A(n_740),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_758),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_748),
.Y(n_774)
);

BUFx8_ASAP7_75t_L g775 ( 
.A(n_758),
.Y(n_775)
);

OAI22xp5_ASAP7_75t_L g776 ( 
.A1(n_735),
.A2(n_726),
.B1(n_631),
.B2(n_728),
.Y(n_776)
);

AOI22xp33_ASAP7_75t_L g777 ( 
.A1(n_745),
.A2(n_679),
.B1(n_731),
.B2(n_729),
.Y(n_777)
);

BUFx3_ASAP7_75t_L g778 ( 
.A(n_755),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_748),
.Y(n_779)
);

INVx3_ASAP7_75t_L g780 ( 
.A(n_759),
.Y(n_780)
);

AOI22xp33_ASAP7_75t_L g781 ( 
.A1(n_745),
.A2(n_679),
.B1(n_715),
.B2(n_718),
.Y(n_781)
);

AOI22xp5_ASAP7_75t_L g782 ( 
.A1(n_735),
.A2(n_713),
.B1(n_722),
.B2(n_682),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_763),
.Y(n_783)
);

AOI22xp33_ASAP7_75t_L g784 ( 
.A1(n_762),
.A2(n_765),
.B1(n_767),
.B2(n_782),
.Y(n_784)
);

BUFx2_ASAP7_75t_L g785 ( 
.A(n_769),
.Y(n_785)
);

BUFx2_ASAP7_75t_L g786 ( 
.A(n_768),
.Y(n_786)
);

HB1xp67_ASAP7_75t_L g787 ( 
.A(n_764),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_766),
.B(n_741),
.Y(n_788)
);

INVx3_ASAP7_75t_L g789 ( 
.A(n_780),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_770),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_771),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_774),
.Y(n_792)
);

OAI22xp5_ASAP7_75t_L g793 ( 
.A1(n_781),
.A2(n_691),
.B1(n_698),
.B2(n_753),
.Y(n_793)
);

BUFx6f_ASAP7_75t_L g794 ( 
.A(n_764),
.Y(n_794)
);

INVx2_ASAP7_75t_SL g795 ( 
.A(n_768),
.Y(n_795)
);

AOI22xp33_ASAP7_75t_L g796 ( 
.A1(n_780),
.A2(n_749),
.B1(n_718),
.B2(n_753),
.Y(n_796)
);

AOI22xp33_ASAP7_75t_L g797 ( 
.A1(n_776),
.A2(n_749),
.B1(n_668),
.B2(n_721),
.Y(n_797)
);

OAI21xp5_ASAP7_75t_SL g798 ( 
.A1(n_777),
.A2(n_714),
.B(n_641),
.Y(n_798)
);

AOI22xp33_ASAP7_75t_L g799 ( 
.A1(n_777),
.A2(n_749),
.B1(n_668),
.B2(n_720),
.Y(n_799)
);

HB1xp67_ASAP7_75t_L g800 ( 
.A(n_764),
.Y(n_800)
);

INVx2_ASAP7_75t_SL g801 ( 
.A(n_768),
.Y(n_801)
);

INVx4_ASAP7_75t_L g802 ( 
.A(n_772),
.Y(n_802)
);

AOI22xp33_ASAP7_75t_L g803 ( 
.A1(n_779),
.A2(n_668),
.B1(n_761),
.B2(n_754),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_783),
.Y(n_804)
);

AOI22xp33_ASAP7_75t_L g805 ( 
.A1(n_784),
.A2(n_486),
.B1(n_666),
.B2(n_747),
.Y(n_805)
);

AND2x2_ASAP7_75t_L g806 ( 
.A(n_785),
.B(n_751),
.Y(n_806)
);

AOI22xp33_ASAP7_75t_L g807 ( 
.A1(n_785),
.A2(n_656),
.B1(n_734),
.B2(n_701),
.Y(n_807)
);

OAI22xp33_ASAP7_75t_L g808 ( 
.A1(n_798),
.A2(n_672),
.B1(n_730),
.B2(n_773),
.Y(n_808)
);

AOI22xp33_ASAP7_75t_L g809 ( 
.A1(n_793),
.A2(n_656),
.B1(n_668),
.B2(n_686),
.Y(n_809)
);

AOI22xp33_ASAP7_75t_L g810 ( 
.A1(n_788),
.A2(n_670),
.B1(n_632),
.B2(n_775),
.Y(n_810)
);

AOI22xp5_ASAP7_75t_L g811 ( 
.A1(n_802),
.A2(n_714),
.B1(n_716),
.B2(n_775),
.Y(n_811)
);

OAI22xp5_ASAP7_75t_L g812 ( 
.A1(n_797),
.A2(n_803),
.B1(n_796),
.B2(n_799),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_786),
.B(n_652),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_787),
.B(n_752),
.Y(n_814)
);

AOI22xp5_ASAP7_75t_L g815 ( 
.A1(n_791),
.A2(n_693),
.B1(n_710),
.B2(n_778),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_790),
.B(n_736),
.Y(n_816)
);

AND2x2_ASAP7_75t_L g817 ( 
.A(n_800),
.B(n_752),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_795),
.B(n_742),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_792),
.Y(n_819)
);

AOI22xp33_ASAP7_75t_L g820 ( 
.A1(n_795),
.A2(n_693),
.B1(n_681),
.B2(n_736),
.Y(n_820)
);

OAI21xp5_ASAP7_75t_SL g821 ( 
.A1(n_801),
.A2(n_681),
.B(n_692),
.Y(n_821)
);

AOI22xp33_ASAP7_75t_SL g822 ( 
.A1(n_789),
.A2(n_693),
.B1(n_737),
.B2(n_756),
.Y(n_822)
);

NAND3xp33_ASAP7_75t_L g823 ( 
.A(n_794),
.B(n_673),
.C(n_651),
.Y(n_823)
);

AOI222xp33_ASAP7_75t_L g824 ( 
.A1(n_794),
.A2(n_680),
.B1(n_677),
.B2(n_688),
.C1(n_671),
.C2(n_659),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_815),
.B(n_810),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_806),
.B(n_794),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_819),
.B(n_794),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_804),
.B(n_742),
.Y(n_828)
);

AOI22xp33_ASAP7_75t_L g829 ( 
.A1(n_805),
.A2(n_671),
.B1(n_680),
.B2(n_697),
.Y(n_829)
);

NOR3xp33_ASAP7_75t_L g830 ( 
.A(n_813),
.B(n_657),
.C(n_746),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_808),
.B(n_746),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_814),
.B(n_817),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_818),
.B(n_743),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_807),
.B(n_750),
.Y(n_834)
);

OA211x2_ASAP7_75t_L g835 ( 
.A1(n_820),
.A2(n_750),
.B(n_89),
.C(n_93),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_816),
.B(n_750),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_824),
.B(n_809),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_812),
.B(n_697),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_821),
.B(n_823),
.Y(n_839)
);

AOI22xp33_ASAP7_75t_L g840 ( 
.A1(n_811),
.A2(n_700),
.B1(n_706),
.B2(n_490),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_SL g841 ( 
.A(n_822),
.B(n_638),
.Y(n_841)
);

OR2x2_ASAP7_75t_L g842 ( 
.A(n_832),
.B(n_96),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_827),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_839),
.B(n_97),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_826),
.B(n_833),
.Y(n_845)
);

INVx2_ASAP7_75t_SL g846 ( 
.A(n_828),
.Y(n_846)
);

AO21x2_ASAP7_75t_L g847 ( 
.A1(n_830),
.A2(n_101),
.B(n_109),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_838),
.B(n_110),
.Y(n_848)
);

HB1xp67_ASAP7_75t_L g849 ( 
.A(n_836),
.Y(n_849)
);

OA211x2_ASAP7_75t_L g850 ( 
.A1(n_825),
.A2(n_114),
.B(n_123),
.C(n_126),
.Y(n_850)
);

AOI22xp33_ASAP7_75t_L g851 ( 
.A1(n_837),
.A2(n_637),
.B1(n_629),
.B2(n_129),
.Y(n_851)
);

OR2x2_ASAP7_75t_L g852 ( 
.A(n_834),
.B(n_831),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_845),
.B(n_849),
.Y(n_853)
);

INVx3_ASAP7_75t_L g854 ( 
.A(n_843),
.Y(n_854)
);

NAND4xp75_ASAP7_75t_L g855 ( 
.A(n_850),
.B(n_835),
.C(n_841),
.D(n_829),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_846),
.B(n_840),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_846),
.B(n_131),
.Y(n_857)
);

INVx2_ASAP7_75t_SL g858 ( 
.A(n_842),
.Y(n_858)
);

XOR2x2_ASAP7_75t_L g859 ( 
.A(n_844),
.B(n_132),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_852),
.Y(n_860)
);

NAND4xp75_ASAP7_75t_L g861 ( 
.A(n_848),
.B(n_138),
.C(n_140),
.D(n_141),
.Y(n_861)
);

AND2x4_ASAP7_75t_L g862 ( 
.A(n_847),
.B(n_232),
.Y(n_862)
);

INVx1_ASAP7_75t_SL g863 ( 
.A(n_853),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_860),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_854),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_854),
.Y(n_866)
);

XNOR2x1_ASAP7_75t_L g867 ( 
.A(n_859),
.B(n_851),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_858),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_856),
.Y(n_869)
);

INVx2_ASAP7_75t_SL g870 ( 
.A(n_857),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_862),
.Y(n_871)
);

INVx1_ASAP7_75t_SL g872 ( 
.A(n_862),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_855),
.B(n_144),
.Y(n_873)
);

NOR2x1_ASAP7_75t_L g874 ( 
.A(n_869),
.B(n_861),
.Y(n_874)
);

INVx1_ASAP7_75t_SL g875 ( 
.A(n_872),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_871),
.Y(n_876)
);

CKINVDCx16_ASAP7_75t_R g877 ( 
.A(n_873),
.Y(n_877)
);

OAI22xp5_ASAP7_75t_L g878 ( 
.A1(n_867),
.A2(n_152),
.B1(n_153),
.B2(n_160),
.Y(n_878)
);

OA22x2_ASAP7_75t_L g879 ( 
.A1(n_863),
.A2(n_870),
.B1(n_868),
.B2(n_865),
.Y(n_879)
);

INVx2_ASAP7_75t_SL g880 ( 
.A(n_864),
.Y(n_880)
);

INVxp67_ASAP7_75t_L g881 ( 
.A(n_866),
.Y(n_881)
);

BUFx2_ASAP7_75t_L g882 ( 
.A(n_879),
.Y(n_882)
);

INVx1_ASAP7_75t_SL g883 ( 
.A(n_875),
.Y(n_883)
);

AOI22xp5_ASAP7_75t_L g884 ( 
.A1(n_882),
.A2(n_877),
.B1(n_874),
.B2(n_878),
.Y(n_884)
);

AO22x1_ASAP7_75t_L g885 ( 
.A1(n_883),
.A2(n_876),
.B1(n_880),
.B2(n_881),
.Y(n_885)
);

HB1xp67_ASAP7_75t_L g886 ( 
.A(n_885),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_884),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_886),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_887),
.Y(n_889)
);

INVx1_ASAP7_75t_SL g890 ( 
.A(n_888),
.Y(n_890)
);

INVxp67_ASAP7_75t_SL g891 ( 
.A(n_889),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_891),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_892),
.B(n_890),
.Y(n_893)
);

AOI22xp33_ASAP7_75t_SL g894 ( 
.A1(n_893),
.A2(n_174),
.B1(n_179),
.B2(n_181),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_894),
.Y(n_895)
);

AOI22xp5_ASAP7_75t_L g896 ( 
.A1(n_895),
.A2(n_182),
.B1(n_183),
.B2(n_188),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_896),
.Y(n_897)
);

OAI22xp5_ASAP7_75t_L g898 ( 
.A1(n_897),
.A2(n_199),
.B1(n_203),
.B2(n_208),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_898),
.Y(n_899)
);

OAI22xp5_ASAP7_75t_L g900 ( 
.A1(n_899),
.A2(n_215),
.B1(n_217),
.B2(n_219),
.Y(n_900)
);

AOI211xp5_ASAP7_75t_L g901 ( 
.A1(n_900),
.A2(n_222),
.B(n_223),
.C(n_230),
.Y(n_901)
);


endmodule