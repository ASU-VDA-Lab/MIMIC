module fake_jpeg_25889_n_136 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_136);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_136;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_14;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

INVx1_ASAP7_75t_SL g15 ( 
.A(n_6),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx6_ASAP7_75t_SL g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

CKINVDCx5p33_ASAP7_75t_R g31 ( 
.A(n_29),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_33),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_36),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_20),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_38),
.Y(n_50)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_15),
.Y(n_53)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_40),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_44),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_18),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_37),
.A2(n_19),
.B1(n_20),
.B2(n_25),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_35),
.B(n_23),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_54),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_36),
.A2(n_19),
.B1(n_15),
.B2(n_23),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_52),
.B(n_30),
.Y(n_57)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_0),
.Y(n_54)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_37),
.A2(n_33),
.B1(n_34),
.B2(n_25),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_56),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_57),
.B(n_0),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_42),
.Y(n_58)
);

OAI21xp33_ASAP7_75t_L g82 ( 
.A1(n_58),
.A2(n_22),
.B(n_21),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_51),
.B(n_54),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_59),
.B(n_73),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_49),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_62),
.B(n_64),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_14),
.Y(n_64)
);

OR2x2_ASAP7_75t_SL g65 ( 
.A(n_41),
.B(n_14),
.Y(n_65)
);

A2O1A1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_65),
.A2(n_68),
.B(n_72),
.C(n_17),
.Y(n_77)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_74),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_53),
.A2(n_50),
.B(n_45),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_42),
.B(n_26),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_24),
.Y(n_78)
);

MAJx2_ASAP7_75t_L g72 ( 
.A(n_45),
.B(n_31),
.C(n_22),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_52),
.B(n_26),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_70),
.A2(n_48),
.B1(n_43),
.B2(n_46),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_76),
.A2(n_80),
.B1(n_74),
.B2(n_60),
.Y(n_98)
);

FAx1_ASAP7_75t_SL g101 ( 
.A(n_77),
.B(n_75),
.CI(n_72),
.CON(n_101),
.SN(n_101)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_78),
.B(n_82),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_70),
.A2(n_48),
.B1(n_43),
.B2(n_46),
.Y(n_80)
);

OAI22x1_ASAP7_75t_SL g81 ( 
.A1(n_61),
.A2(n_22),
.B1(n_29),
.B2(n_38),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_81),
.A2(n_87),
.B1(n_63),
.B2(n_65),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_69),
.B(n_24),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_83),
.B(n_67),
.Y(n_95)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_85),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

INVx13_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_86),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_57),
.A2(n_21),
.B1(n_17),
.B2(n_2),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_88),
.A2(n_64),
.B(n_62),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_90),
.B(n_93),
.Y(n_108)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_89),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_94),
.B(n_98),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_95),
.B(n_101),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_77),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_96),
.B(n_1),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_78),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_97),
.Y(n_109)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_76),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_100),
.B(n_102),
.Y(n_107)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

AOI322xp5_ASAP7_75t_SL g103 ( 
.A1(n_101),
.A2(n_85),
.A3(n_81),
.B1(n_79),
.B2(n_87),
.C1(n_84),
.C2(n_10),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_110),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_99),
.A2(n_88),
.B(n_86),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_106),
.B(n_112),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_60),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_98),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_111),
.B(n_102),
.Y(n_116)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_107),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_113),
.B(n_114),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_110),
.B(n_93),
.C(n_90),
.Y(n_114)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_116),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_111),
.A2(n_100),
.B1(n_91),
.B2(n_101),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_117),
.B(n_118),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_104),
.A2(n_92),
.B1(n_3),
.B2(n_5),
.Y(n_118)
);

OAI322xp33_ASAP7_75t_L g122 ( 
.A1(n_119),
.A2(n_112),
.A3(n_105),
.B1(n_108),
.B2(n_109),
.C1(n_106),
.C2(n_107),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_122),
.B(n_11),
.Y(n_128)
);

NOR3xp33_ASAP7_75t_L g124 ( 
.A(n_114),
.B(n_8),
.C(n_9),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_10),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_125),
.B(n_126),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_123),
.A2(n_118),
.B1(n_115),
.B2(n_12),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_121),
.B(n_115),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_127),
.B(n_128),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_128),
.B(n_120),
.C(n_121),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_130),
.B(n_1),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_13),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_132),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_133),
.C(n_129),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_1),
.Y(n_136)
);


endmodule