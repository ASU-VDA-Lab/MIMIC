module real_aes_853_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_794, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_794;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_791;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_769;
wire n_434;
wire n_527;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_756;
wire n_735;
wire n_728;
wire n_713;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_785;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_335;
wire n_177;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_0), .B(n_152), .Y(n_219) );
AOI21xp5_ASAP7_75t_L g182 ( .A1(n_1), .A2(n_161), .B(n_183), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_2), .B(n_111), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_3), .B(n_152), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_4), .B(n_168), .Y(n_541) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_5), .B(n_168), .Y(n_231) );
INVx1_ASAP7_75t_L g159 ( .A(n_6), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_7), .B(n_168), .Y(n_206) );
CKINVDCx16_ASAP7_75t_R g111 ( .A(n_8), .Y(n_111) );
NAND2xp33_ASAP7_75t_L g169 ( .A(n_9), .B(n_170), .Y(n_169) );
AND2x2_ASAP7_75t_L g483 ( .A(n_10), .B(n_178), .Y(n_483) );
AND2x2_ASAP7_75t_L g543 ( .A(n_11), .B(n_147), .Y(n_543) );
INVx2_ASAP7_75t_L g149 ( .A(n_12), .Y(n_149) );
AOI221x1_ASAP7_75t_L g247 ( .A1(n_13), .A2(n_24), .B1(n_152), .B2(n_161), .C(n_248), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_14), .B(n_168), .Y(n_517) );
CKINVDCx16_ASAP7_75t_R g112 ( .A(n_15), .Y(n_112) );
NAND2xp5_ASAP7_75t_SL g151 ( .A(n_16), .B(n_152), .Y(n_151) );
AO21x2_ASAP7_75t_L g146 ( .A1(n_17), .A2(n_147), .B(n_150), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_18), .B(n_186), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_19), .B(n_168), .Y(n_195) );
AO21x1_ASAP7_75t_L g226 ( .A1(n_20), .A2(n_152), .B(n_227), .Y(n_226) );
NAND2xp5_ASAP7_75t_SL g548 ( .A(n_21), .B(n_152), .Y(n_548) );
INVx1_ASAP7_75t_L g108 ( .A(n_22), .Y(n_108) );
AOI22xp33_ASAP7_75t_L g487 ( .A1(n_23), .A2(n_89), .B1(n_152), .B2(n_488), .Y(n_487) );
NAND2x1_ASAP7_75t_L g217 ( .A(n_25), .B(n_168), .Y(n_217) );
NAND2x1_ASAP7_75t_L g205 ( .A(n_26), .B(n_170), .Y(n_205) );
CKINVDCx20_ASAP7_75t_R g775 ( .A(n_27), .Y(n_775) );
OA21x2_ASAP7_75t_L g148 ( .A1(n_28), .A2(n_86), .B(n_149), .Y(n_148) );
OR2x2_ASAP7_75t_L g173 ( .A(n_28), .B(n_86), .Y(n_173) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_29), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_30), .B(n_170), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_31), .B(n_168), .Y(n_167) );
AO21x2_ASAP7_75t_L g512 ( .A1(n_32), .A2(n_178), .B(n_513), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_33), .B(n_170), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_34), .A2(n_161), .B(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_35), .B(n_168), .Y(n_524) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_36), .A2(n_161), .B(n_237), .Y(n_236) );
AND2x2_ASAP7_75t_L g158 ( .A(n_37), .B(n_159), .Y(n_158) );
AND2x2_ASAP7_75t_L g162 ( .A(n_37), .B(n_163), .Y(n_162) );
INVx1_ASAP7_75t_L g496 ( .A(n_37), .Y(n_496) );
NOR3xp33_ASAP7_75t_L g109 ( .A(n_38), .B(n_110), .C(n_112), .Y(n_109) );
OR2x6_ASAP7_75t_L g126 ( .A(n_38), .B(n_127), .Y(n_126) );
NAND2xp5_ASAP7_75t_SL g240 ( .A(n_39), .B(n_152), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_40), .B(n_152), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_41), .B(n_168), .Y(n_508) );
CKINVDCx20_ASAP7_75t_R g199 ( .A(n_42), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_43), .B(n_170), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_44), .B(n_152), .Y(n_469) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_45), .A2(n_161), .B(n_479), .Y(n_478) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_46), .A2(n_161), .B(n_204), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_47), .B(n_170), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_48), .B(n_170), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_49), .B(n_152), .Y(n_514) );
INVx1_ASAP7_75t_L g155 ( .A(n_50), .Y(n_155) );
INVx1_ASAP7_75t_L g165 ( .A(n_50), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_51), .B(n_168), .Y(n_481) );
AND2x2_ASAP7_75t_L g503 ( .A(n_52), .B(n_186), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_53), .B(n_170), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_54), .B(n_168), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_55), .B(n_170), .Y(n_523) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_56), .A2(n_161), .B(n_216), .Y(n_215) );
NAND2xp5_ASAP7_75t_SL g482 ( .A(n_57), .B(n_152), .Y(n_482) );
NAND2xp5_ASAP7_75t_SL g505 ( .A(n_58), .B(n_152), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_59), .A2(n_161), .B(n_522), .Y(n_521) );
AOI22xp5_ASAP7_75t_L g131 ( .A1(n_60), .A2(n_98), .B1(n_132), .B2(n_133), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g133 ( .A(n_60), .Y(n_133) );
AO21x1_ASAP7_75t_L g228 ( .A1(n_61), .A2(n_161), .B(n_229), .Y(n_228) );
AND2x2_ASAP7_75t_L g554 ( .A(n_62), .B(n_187), .Y(n_554) );
NAND2xp5_ASAP7_75t_SL g181 ( .A(n_63), .B(n_152), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_64), .B(n_170), .Y(n_509) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_65), .B(n_152), .Y(n_207) );
AOI22xp5_ASAP7_75t_L g784 ( .A1(n_66), .A2(n_78), .B1(n_785), .B2(n_786), .Y(n_784) );
CKINVDCx20_ASAP7_75t_R g786 ( .A(n_66), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_67), .B(n_170), .Y(n_518) );
AOI22xp5_ASAP7_75t_L g493 ( .A1(n_68), .A2(n_93), .B1(n_161), .B2(n_494), .Y(n_493) );
AND2x2_ASAP7_75t_L g241 ( .A(n_69), .B(n_187), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_70), .B(n_168), .Y(n_551) );
INVx1_ASAP7_75t_L g157 ( .A(n_71), .Y(n_157) );
INVx1_ASAP7_75t_L g163 ( .A(n_71), .Y(n_163) );
AND2x2_ASAP7_75t_L g209 ( .A(n_72), .B(n_178), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_73), .B(n_170), .Y(n_540) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_74), .A2(n_161), .B(n_507), .Y(n_506) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_75), .A2(n_161), .B(n_471), .Y(n_470) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_76), .A2(n_161), .B(n_516), .Y(n_515) );
AND2x2_ASAP7_75t_L g526 ( .A(n_77), .B(n_187), .Y(n_526) );
CKINVDCx20_ASAP7_75t_R g785 ( .A(n_78), .Y(n_785) );
NAND2xp5_ASAP7_75t_SL g485 ( .A(n_79), .B(n_186), .Y(n_485) );
NOR2xp33_ASAP7_75t_L g107 ( .A(n_80), .B(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g128 ( .A(n_80), .Y(n_128) );
AND2x2_ASAP7_75t_L g177 ( .A(n_81), .B(n_178), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_82), .B(n_152), .Y(n_197) );
AND2x2_ASAP7_75t_L g474 ( .A(n_83), .B(n_147), .Y(n_474) );
INVxp33_ASAP7_75t_L g792 ( .A(n_84), .Y(n_792) );
AND2x2_ASAP7_75t_L g227 ( .A(n_85), .B(n_172), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_87), .B(n_170), .Y(n_196) );
AND2x2_ASAP7_75t_L g221 ( .A(n_88), .B(n_178), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_90), .B(n_168), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g193 ( .A1(n_91), .A2(n_161), .B(n_194), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_92), .B(n_170), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_94), .A2(n_161), .B(n_550), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_95), .B(n_168), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_96), .B(n_168), .Y(n_184) );
BUFx2_ASAP7_75t_L g553 ( .A(n_97), .Y(n_553) );
CKINVDCx20_ASAP7_75t_R g132 ( .A(n_98), .Y(n_132) );
BUFx2_ASAP7_75t_L g117 ( .A(n_99), .Y(n_117) );
BUFx2_ASAP7_75t_SL g781 ( .A(n_99), .Y(n_781) );
AOI21xp5_ASAP7_75t_L g160 ( .A1(n_100), .A2(n_161), .B(n_166), .Y(n_160) );
AOI21xp33_ASAP7_75t_SL g101 ( .A1(n_102), .A2(n_113), .B(n_791), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
NOR2xp33_ASAP7_75t_L g791 ( .A(n_104), .B(n_792), .Y(n_791) );
INVx1_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
INVx3_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
AND2x2_ASAP7_75t_SL g106 ( .A(n_107), .B(n_109), .Y(n_106) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_108), .B(n_128), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_112), .B(n_125), .Y(n_124) );
OR2x6_ASAP7_75t_SL g139 ( .A(n_112), .B(n_125), .Y(n_139) );
AND2x6_ASAP7_75t_SL g768 ( .A(n_112), .B(n_126), .Y(n_768) );
OR2x2_ASAP7_75t_L g778 ( .A(n_112), .B(n_126), .Y(n_778) );
OA21x2_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_130), .B(n_779), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_115), .B(n_118), .Y(n_114) );
HB1xp67_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
HB1xp67_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVxp67_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
AOI21xp5_ASAP7_75t_L g782 ( .A1(n_119), .A2(n_783), .B(n_788), .Y(n_782) );
NOR2xp33_ASAP7_75t_SL g119 ( .A(n_120), .B(n_129), .Y(n_119) );
INVx1_ASAP7_75t_SL g120 ( .A(n_121), .Y(n_120) );
BUFx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_123), .Y(n_122) );
BUFx3_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
BUFx2_ASAP7_75t_L g790 ( .A(n_124), .Y(n_790) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_126), .Y(n_125) );
OAI21xp5_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_134), .B(n_769), .Y(n_130) );
AOI21xp5_ASAP7_75t_L g769 ( .A1(n_131), .A2(n_770), .B(n_774), .Y(n_769) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
OAI22xp5_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_140), .B1(n_462), .B2(n_765), .Y(n_135) );
BUFx4f_ASAP7_75t_SL g136 ( .A(n_137), .Y(n_136) );
OAI22x1_ASAP7_75t_L g770 ( .A1(n_137), .A2(n_771), .B1(n_772), .B2(n_773), .Y(n_770) );
CKINVDCx20_ASAP7_75t_R g137 ( .A(n_138), .Y(n_137) );
CKINVDCx11_ASAP7_75t_R g138 ( .A(n_139), .Y(n_138) );
INVx1_ASAP7_75t_L g771 ( .A(n_140), .Y(n_771) );
AND2x4_ASAP7_75t_L g140 ( .A(n_141), .B(n_383), .Y(n_140) );
NOR3xp33_ASAP7_75t_SL g141 ( .A(n_142), .B(n_295), .C(n_335), .Y(n_141) );
OAI221xp5_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_210), .B1(n_259), .B2(n_274), .C(n_277), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
AND2x2_ASAP7_75t_L g144 ( .A(n_145), .B(n_174), .Y(n_144) );
INVx2_ASAP7_75t_L g292 ( .A(n_145), .Y(n_292) );
AND2x2_ASAP7_75t_L g322 ( .A(n_145), .B(n_323), .Y(n_322) );
BUFx3_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AND2x2_ASAP7_75t_L g260 ( .A(n_146), .B(n_261), .Y(n_260) );
OR2x2_ASAP7_75t_L g267 ( .A(n_146), .B(n_200), .Y(n_267) );
INVx2_ASAP7_75t_L g273 ( .A(n_146), .Y(n_273) );
AND2x2_ASAP7_75t_L g282 ( .A(n_146), .B(n_176), .Y(n_282) );
INVx1_ASAP7_75t_L g298 ( .A(n_146), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_146), .B(n_344), .Y(n_343) );
AOI21xp5_ASAP7_75t_L g547 ( .A1(n_147), .A2(n_548), .B(n_549), .Y(n_547) );
BUFx4f_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx3_ASAP7_75t_L g179 ( .A(n_148), .Y(n_179) );
AND2x4_ASAP7_75t_L g172 ( .A(n_149), .B(n_173), .Y(n_172) );
AND2x2_ASAP7_75t_SL g187 ( .A(n_149), .B(n_173), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_160), .B(n_172), .Y(n_150) );
AND2x4_ASAP7_75t_L g152 ( .A(n_153), .B(n_158), .Y(n_152) );
AND2x4_ASAP7_75t_L g153 ( .A(n_154), .B(n_156), .Y(n_153) );
AND2x6_ASAP7_75t_L g170 ( .A(n_154), .B(n_163), .Y(n_170) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
AND2x4_ASAP7_75t_L g168 ( .A(n_156), .B(n_165), .Y(n_168) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx5_ASAP7_75t_L g171 ( .A(n_158), .Y(n_171) );
AND2x2_ASAP7_75t_L g164 ( .A(n_159), .B(n_165), .Y(n_164) );
HB1xp67_ASAP7_75t_L g491 ( .A(n_159), .Y(n_491) );
AND2x6_ASAP7_75t_L g161 ( .A(n_162), .B(n_164), .Y(n_161) );
BUFx3_ASAP7_75t_L g492 ( .A(n_162), .Y(n_492) );
INVx2_ASAP7_75t_L g498 ( .A(n_163), .Y(n_498) );
AND2x4_ASAP7_75t_L g494 ( .A(n_164), .B(n_495), .Y(n_494) );
INVx2_ASAP7_75t_L g490 ( .A(n_165), .Y(n_490) );
AOI21xp5_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_169), .B(n_171), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_170), .B(n_553), .Y(n_552) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_171), .A2(n_184), .B(n_185), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_171), .A2(n_195), .B(n_196), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_171), .A2(n_205), .B(n_206), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_171), .A2(n_217), .B(n_218), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_171), .A2(n_230), .B(n_231), .Y(n_229) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_171), .A2(n_238), .B(n_239), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_171), .A2(n_249), .B(n_250), .Y(n_248) );
AOI21xp5_ASAP7_75t_L g471 ( .A1(n_171), .A2(n_472), .B(n_473), .Y(n_471) );
AOI21xp5_ASAP7_75t_L g479 ( .A1(n_171), .A2(n_480), .B(n_481), .Y(n_479) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_171), .A2(n_508), .B(n_509), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_171), .A2(n_517), .B(n_518), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_171), .A2(n_523), .B(n_524), .Y(n_522) );
AOI21xp5_ASAP7_75t_L g539 ( .A1(n_171), .A2(n_540), .B(n_541), .Y(n_539) );
AOI21xp5_ASAP7_75t_L g550 ( .A1(n_171), .A2(n_551), .B(n_552), .Y(n_550) );
INVx1_ASAP7_75t_SL g191 ( .A(n_172), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_172), .B(n_233), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g504 ( .A1(n_172), .A2(n_505), .B(n_506), .Y(n_504) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_172), .A2(n_514), .B(n_515), .Y(n_513) );
AND2x2_ASAP7_75t_SL g174 ( .A(n_175), .B(n_188), .Y(n_174) );
INVx4_ASAP7_75t_L g263 ( .A(n_175), .Y(n_263) );
AND2x2_ASAP7_75t_L g294 ( .A(n_175), .B(n_201), .Y(n_294) );
AND2x2_ASAP7_75t_L g370 ( .A(n_175), .B(n_344), .Y(n_370) );
NAND2x1p5_ASAP7_75t_L g412 ( .A(n_175), .B(n_200), .Y(n_412) );
INVx5_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_176), .B(n_200), .Y(n_299) );
AND2x2_ASAP7_75t_L g323 ( .A(n_176), .B(n_201), .Y(n_323) );
BUFx2_ASAP7_75t_L g339 ( .A(n_176), .Y(n_339) );
NOR2x1_ASAP7_75t_SL g442 ( .A(n_176), .B(n_344), .Y(n_442) );
OR2x6_ASAP7_75t_L g176 ( .A(n_177), .B(n_180), .Y(n_176) );
INVx3_ASAP7_75t_L g220 ( .A(n_178), .Y(n_220) );
INVx4_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
AO21x2_ASAP7_75t_L g476 ( .A1(n_179), .A2(n_477), .B(n_483), .Y(n_476) );
AOI21xp5_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_182), .B(n_186), .Y(n_180) );
CKINVDCx5p33_ASAP7_75t_R g208 ( .A(n_186), .Y(n_208) );
OA21x2_ASAP7_75t_L g246 ( .A1(n_186), .A2(n_247), .B(n_251), .Y(n_246) );
OA21x2_ASAP7_75t_L g309 ( .A1(n_186), .A2(n_247), .B(n_251), .Y(n_309) );
AOI21xp5_ASAP7_75t_L g468 ( .A1(n_186), .A2(n_469), .B(n_470), .Y(n_468) );
AO21x2_ASAP7_75t_L g486 ( .A1(n_186), .A2(n_487), .B(n_493), .Y(n_486) );
BUFx6f_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
INVx2_ASAP7_75t_L g319 ( .A(n_188), .Y(n_319) );
AOI221xp5_ASAP7_75t_L g385 ( .A1(n_188), .A2(n_386), .B1(n_388), .B2(n_390), .C(n_395), .Y(n_385) );
AND2x2_ASAP7_75t_L g405 ( .A(n_188), .B(n_298), .Y(n_405) );
AND2x4_ASAP7_75t_L g188 ( .A(n_189), .B(n_200), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVx2_ASAP7_75t_L g261 ( .A(n_190), .Y(n_261) );
INVx1_ASAP7_75t_L g314 ( .A(n_190), .Y(n_314) );
AO21x2_ASAP7_75t_L g190 ( .A1(n_191), .A2(n_192), .B(n_198), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_191), .B(n_199), .Y(n_198) );
AO21x2_ASAP7_75t_L g344 ( .A1(n_191), .A2(n_192), .B(n_198), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_193), .B(n_197), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_200), .B(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g283 ( .A(n_200), .B(n_271), .Y(n_283) );
INVx2_ASAP7_75t_L g325 ( .A(n_200), .Y(n_325) );
AND2x2_ASAP7_75t_L g458 ( .A(n_200), .B(n_273), .Y(n_458) );
INVx4_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
HB1xp67_ASAP7_75t_L g315 ( .A(n_201), .Y(n_315) );
AO21x2_ASAP7_75t_L g201 ( .A1(n_202), .A2(n_208), .B(n_209), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_203), .B(n_207), .Y(n_202) );
AOI21x1_ASAP7_75t_L g536 ( .A1(n_208), .A2(n_537), .B(n_543), .Y(n_536) );
NOR3xp33_ASAP7_75t_L g210 ( .A(n_211), .B(n_242), .C(n_257), .Y(n_210) );
AND2x2_ASAP7_75t_L g211 ( .A(n_212), .B(n_222), .Y(n_211) );
INVx2_ASAP7_75t_L g372 ( .A(n_212), .Y(n_372) );
AND2x2_ASAP7_75t_L g417 ( .A(n_212), .B(n_294), .Y(n_417) );
BUFx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
INVx1_ASAP7_75t_L g362 ( .A(n_213), .Y(n_362) );
AND2x4_ASAP7_75t_SL g377 ( .A(n_213), .B(n_289), .Y(n_377) );
AO21x2_ASAP7_75t_L g213 ( .A1(n_214), .A2(n_220), .B(n_221), .Y(n_213) );
AO21x2_ASAP7_75t_L g256 ( .A1(n_214), .A2(n_220), .B(n_221), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_215), .B(n_219), .Y(n_214) );
AO21x2_ASAP7_75t_L g234 ( .A1(n_220), .A2(n_235), .B(n_241), .Y(n_234) );
AO21x2_ASAP7_75t_L g254 ( .A1(n_220), .A2(n_235), .B(n_241), .Y(n_254) );
AO21x1_ASAP7_75t_SL g519 ( .A1(n_220), .A2(n_520), .B(n_526), .Y(n_519) );
AO21x2_ASAP7_75t_L g577 ( .A1(n_220), .A2(n_520), .B(n_526), .Y(n_577) );
INVx2_ASAP7_75t_L g331 ( .A(n_222), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_222), .B(n_361), .Y(n_387) );
AND2x4_ASAP7_75t_L g420 ( .A(n_222), .B(n_367), .Y(n_420) );
AND2x4_ASAP7_75t_L g222 ( .A(n_223), .B(n_234), .Y(n_222) );
AND2x2_ASAP7_75t_L g258 ( .A(n_223), .B(n_253), .Y(n_258) );
OR2x2_ASAP7_75t_L g288 ( .A(n_223), .B(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_SL g357 ( .A(n_223), .B(n_309), .Y(n_357) );
INVx2_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
BUFx2_ASAP7_75t_L g302 ( .A(n_224), .Y(n_302) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
INVx2_ASAP7_75t_L g276 ( .A(n_225), .Y(n_276) );
OAI21x1_ASAP7_75t_SL g225 ( .A1(n_226), .A2(n_228), .B(n_232), .Y(n_225) );
INVx1_ASAP7_75t_L g233 ( .A(n_227), .Y(n_233) );
INVx2_ASAP7_75t_L g289 ( .A(n_234), .Y(n_289) );
NAND2xp5_ASAP7_75t_SL g235 ( .A(n_236), .B(n_240), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g451 ( .A(n_242), .B(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_244), .B(n_252), .Y(n_243) );
AND2x2_ASAP7_75t_L g257 ( .A(n_244), .B(n_258), .Y(n_257) );
OR2x2_ASAP7_75t_L g330 ( .A(n_244), .B(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g415 ( .A(n_244), .Y(n_415) );
BUFx2_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
AND2x4_ASAP7_75t_L g275 ( .A(n_245), .B(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g394 ( .A(n_245), .B(n_254), .Y(n_394) );
AND2x2_ASAP7_75t_L g398 ( .A(n_245), .B(n_264), .Y(n_398) );
INVx2_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
INVx2_ASAP7_75t_L g367 ( .A(n_246), .Y(n_367) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_246), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_252), .B(n_275), .Y(n_351) );
AND2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_255), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_253), .B(n_276), .Y(n_461) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g265 ( .A(n_254), .B(n_256), .Y(n_265) );
AND2x2_ASAP7_75t_L g347 ( .A(n_254), .B(n_309), .Y(n_347) );
AND2x2_ASAP7_75t_L g366 ( .A(n_254), .B(n_255), .Y(n_366) );
BUFx2_ASAP7_75t_L g287 ( .A(n_255), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_255), .B(n_347), .Y(n_346) );
INVx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
BUFx3_ASAP7_75t_L g264 ( .A(n_256), .Y(n_264) );
INVxp67_ASAP7_75t_L g307 ( .A(n_256), .Y(n_307) );
INVx1_ASAP7_75t_L g280 ( .A(n_258), .Y(n_280) );
AND2x2_ASAP7_75t_L g316 ( .A(n_258), .B(n_287), .Y(n_316) );
NAND2xp33_ASAP7_75t_L g397 ( .A(n_258), .B(n_398), .Y(n_397) );
AND2x2_ASAP7_75t_L g434 ( .A(n_258), .B(n_435), .Y(n_434) );
AOI221xp5_ASAP7_75t_L g259 ( .A1(n_260), .A2(n_262), .B1(n_265), .B2(n_266), .C(n_268), .Y(n_259) );
AND2x2_ASAP7_75t_L g363 ( .A(n_260), .B(n_263), .Y(n_363) );
AND2x2_ASAP7_75t_SL g382 ( .A(n_260), .B(n_323), .Y(n_382) );
AND2x2_ASAP7_75t_L g400 ( .A(n_260), .B(n_325), .Y(n_400) );
AND2x2_ASAP7_75t_L g455 ( .A(n_260), .B(n_294), .Y(n_455) );
INVx1_ASAP7_75t_L g271 ( .A(n_261), .Y(n_271) );
HB1xp67_ASAP7_75t_L g327 ( .A(n_261), .Y(n_327) );
CKINVDCx16_ASAP7_75t_R g407 ( .A(n_262), .Y(n_407) );
AND2x4_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_263), .B(n_273), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_263), .B(n_314), .Y(n_389) );
AND2x2_ASAP7_75t_L g356 ( .A(n_264), .B(n_357), .Y(n_356) );
INVx1_ASAP7_75t_SL g392 ( .A(n_264), .Y(n_392) );
AND2x2_ASAP7_75t_L g301 ( .A(n_265), .B(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_265), .B(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g443 ( .A(n_265), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_265), .B(n_367), .Y(n_453) );
AND2x4_ASAP7_75t_L g369 ( .A(n_266), .B(n_370), .Y(n_369) );
INVx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
OR2x2_ASAP7_75t_L g440 ( .A(n_267), .B(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
OR2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_272), .Y(n_269) );
OR2x2_ASAP7_75t_L g311 ( .A(n_272), .B(n_312), .Y(n_311) );
OR2x2_ASAP7_75t_L g318 ( .A(n_273), .B(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g349 ( .A(n_273), .B(n_323), .Y(n_349) );
AND2x2_ASAP7_75t_L g423 ( .A(n_273), .B(n_344), .Y(n_423) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g371 ( .A(n_275), .B(n_372), .Y(n_371) );
OAI32xp33_ASAP7_75t_L g436 ( .A1(n_275), .A2(n_437), .A3(n_439), .B1(n_440), .B2(n_443), .Y(n_436) );
AND2x4_ASAP7_75t_L g308 ( .A(n_276), .B(n_309), .Y(n_308) );
OR2x2_ASAP7_75t_L g406 ( .A(n_276), .B(n_309), .Y(n_406) );
AOI22xp5_ASAP7_75t_L g277 ( .A1(n_278), .A2(n_281), .B1(n_284), .B2(n_290), .Y(n_277) );
INVxp67_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
O2A1O1Ixp33_ASAP7_75t_SL g395 ( .A1(n_279), .A2(n_293), .B(n_396), .C(n_397), .Y(n_395) );
HB1xp67_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
OR2x2_ASAP7_75t_L g379 ( .A(n_280), .B(n_307), .Y(n_379) );
INVx1_ASAP7_75t_SL g450 ( .A(n_281), .Y(n_450) );
AND2x4_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
AND2x4_ASAP7_75t_L g353 ( .A(n_283), .B(n_292), .Y(n_353) );
AOI221xp5_ASAP7_75t_L g431 ( .A1(n_283), .A2(n_432), .B1(n_433), .B2(n_434), .C(n_436), .Y(n_431) );
INVx1_ASAP7_75t_SL g284 ( .A(n_285), .Y(n_284) );
OR2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_288), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
NOR2xp33_ASAP7_75t_L g359 ( .A(n_288), .B(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
OAI22xp33_ASAP7_75t_L g373 ( .A1(n_291), .A2(n_321), .B1(n_374), .B2(n_375), .Y(n_373) );
OR2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
OAI211xp5_ASAP7_75t_SL g409 ( .A1(n_292), .A2(n_410), .B(n_418), .C(n_431), .Y(n_409) );
INVx2_ASAP7_75t_SL g293 ( .A(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g329 ( .A(n_294), .B(n_298), .Y(n_329) );
OAI211xp5_ASAP7_75t_SL g295 ( .A1(n_296), .A2(n_300), .B(n_303), .C(n_332), .Y(n_295) );
OR2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_299), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g326 ( .A(n_298), .B(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g446 ( .A(n_298), .B(n_442), .Y(n_446) );
OAI32xp33_ASAP7_75t_L g403 ( .A1(n_299), .A2(n_404), .A3(n_406), .B1(n_407), .B2(n_408), .Y(n_403) );
INVx1_ASAP7_75t_SL g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_SL g393 ( .A(n_302), .B(n_394), .Y(n_393) );
AOI221xp5_ASAP7_75t_L g303 ( .A1(n_304), .A2(n_310), .B1(n_316), .B2(n_317), .C(n_320), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_SL g305 ( .A(n_306), .B(n_308), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
OR2x2_ASAP7_75t_L g460 ( .A(n_307), .B(n_461), .Y(n_460) );
NAND2xp5_ASAP7_75t_SL g374 ( .A(n_308), .B(n_372), .Y(n_374) );
A2O1A1O1Ixp25_ASAP7_75t_L g445 ( .A1(n_308), .A2(n_377), .B(n_393), .C(n_439), .D(n_446), .Y(n_445) );
AOI31xp33_ASAP7_75t_L g447 ( .A1(n_308), .A2(n_329), .A3(n_439), .B(n_446), .Y(n_447) );
AND2x2_ASAP7_75t_L g361 ( .A(n_309), .B(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_SL g449 ( .A(n_311), .B(n_450), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_313), .B(n_315), .Y(n_312) );
INVx2_ASAP7_75t_L g438 ( .A(n_313), .Y(n_438) );
INVx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g433 ( .A(n_314), .B(n_325), .Y(n_433) );
INVx1_ASAP7_75t_L g348 ( .A(n_316), .Y(n_348) );
AND2x2_ASAP7_75t_L g333 ( .A(n_317), .B(n_334), .Y(n_333) );
INVx2_ASAP7_75t_SL g317 ( .A(n_318), .Y(n_317) );
AOI31xp33_ASAP7_75t_L g320 ( .A1(n_321), .A2(n_324), .A3(n_328), .B(n_330), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_323), .B(n_438), .Y(n_437) );
AND2x2_ASAP7_75t_L g456 ( .A(n_323), .B(n_402), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
AND2x2_ASAP7_75t_L g401 ( .A(n_325), .B(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g427 ( .A(n_325), .Y(n_427) );
INVxp67_ASAP7_75t_L g396 ( .A(n_326), .Y(n_396) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx2_ASAP7_75t_L g334 ( .A(n_330), .Y(n_334) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
NAND3xp33_ASAP7_75t_SL g335 ( .A(n_336), .B(n_352), .C(n_368), .Y(n_335) );
AOI22xp5_ASAP7_75t_L g336 ( .A1(n_337), .A2(n_345), .B1(n_349), .B2(n_350), .Y(n_336) );
INVxp67_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
INVx2_ASAP7_75t_L g422 ( .A(n_339), .Y(n_422) );
INVx1_ASAP7_75t_SL g340 ( .A(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVxp67_ASAP7_75t_SL g402 ( .A(n_343), .Y(n_402) );
INVxp67_ASAP7_75t_SL g428 ( .A(n_343), .Y(n_428) );
OR2x2_ASAP7_75t_L g429 ( .A(n_343), .B(n_412), .Y(n_429) );
NAND2xp33_ASAP7_75t_L g345 ( .A(n_346), .B(n_348), .Y(n_345) );
INVx1_ASAP7_75t_L g380 ( .A(n_347), .Y(n_380) );
INVx1_ASAP7_75t_SL g350 ( .A(n_351), .Y(n_350) );
AOI22xp33_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_354), .B1(n_363), .B2(n_364), .Y(n_352) );
NAND2xp5_ASAP7_75t_SL g354 ( .A(n_355), .B(n_358), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_SL g360 ( .A(n_361), .Y(n_360) );
AOI221xp5_ASAP7_75t_L g399 ( .A1(n_361), .A2(n_366), .B1(n_400), .B2(n_401), .C(n_403), .Y(n_399) );
INVx2_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
NAND2x1_ASAP7_75t_L g365 ( .A(n_366), .B(n_367), .Y(n_365) );
INVx1_ASAP7_75t_L g439 ( .A(n_366), .Y(n_439) );
AND2x2_ASAP7_75t_L g376 ( .A(n_367), .B(n_377), .Y(n_376) );
O2A1O1Ixp33_ASAP7_75t_SL g424 ( .A1(n_367), .A2(n_425), .B(n_429), .C(n_430), .Y(n_424) );
AOI211xp5_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_371), .B(n_373), .C(n_378), .Y(n_368) );
AND2x2_ASAP7_75t_L g419 ( .A(n_372), .B(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g430 ( .A(n_377), .Y(n_430) );
AOI21xp33_ASAP7_75t_SL g378 ( .A1(n_379), .A2(n_380), .B(n_381), .Y(n_378) );
INVx2_ASAP7_75t_SL g381 ( .A(n_382), .Y(n_381) );
NOR3xp33_ASAP7_75t_L g383 ( .A(n_384), .B(n_409), .C(n_444), .Y(n_383) );
NAND2xp5_ASAP7_75t_SL g384 ( .A(n_385), .B(n_399), .Y(n_384) );
INVx1_ASAP7_75t_SL g386 ( .A(n_387), .Y(n_386) );
INVxp67_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
NAND2xp5_ASAP7_75t_SL g391 ( .A(n_392), .B(n_393), .Y(n_391) );
INVx1_ASAP7_75t_L g408 ( .A(n_393), .Y(n_408) );
INVxp67_ASAP7_75t_L g432 ( .A(n_397), .Y(n_432) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_SL g416 ( .A(n_406), .Y(n_416) );
AOI22xp5_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_413), .B1(n_416), .B2(n_417), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
AOI21xp5_ASAP7_75t_L g418 ( .A1(n_419), .A2(n_421), .B(n_424), .Y(n_418) );
AND2x2_ASAP7_75t_L g421 ( .A(n_422), .B(n_423), .Y(n_421) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_427), .B(n_428), .Y(n_426) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
AND2x2_ASAP7_75t_L g457 ( .A(n_442), .B(n_458), .Y(n_457) );
OAI221xp5_ASAP7_75t_L g444 ( .A1(n_445), .A2(n_447), .B1(n_448), .B2(n_451), .C(n_454), .Y(n_444) );
INVxp67_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
OAI31xp33_ASAP7_75t_SL g454 ( .A1(n_455), .A2(n_456), .A3(n_457), .B(n_459), .Y(n_454) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx3_ASAP7_75t_SL g772 ( .A(n_462), .Y(n_772) );
OAI22xp5_ASAP7_75t_SL g783 ( .A1(n_462), .A2(n_772), .B1(n_784), .B2(n_787), .Y(n_783) );
AND2x4_ASAP7_75t_SL g462 ( .A(n_463), .B(n_661), .Y(n_462) );
NOR3xp33_ASAP7_75t_SL g463 ( .A(n_464), .B(n_570), .C(n_602), .Y(n_463) );
OAI221xp5_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_499), .B1(n_527), .B2(n_544), .C(n_555), .Y(n_464) );
OR2x2_ASAP7_75t_L g465 ( .A(n_466), .B(n_475), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
AND2x2_ASAP7_75t_L g533 ( .A(n_467), .B(n_476), .Y(n_533) );
INVx4_ASAP7_75t_L g561 ( .A(n_467), .Y(n_561) );
AND2x4_ASAP7_75t_SL g601 ( .A(n_467), .B(n_535), .Y(n_601) );
BUFx2_ASAP7_75t_L g611 ( .A(n_467), .Y(n_611) );
NOR2x1_ASAP7_75t_L g677 ( .A(n_467), .B(n_616), .Y(n_677) );
AND2x2_ASAP7_75t_L g686 ( .A(n_467), .B(n_614), .Y(n_686) );
OR2x2_ASAP7_75t_L g694 ( .A(n_467), .B(n_695), .Y(n_694) );
AND2x2_ASAP7_75t_L g720 ( .A(n_467), .B(n_559), .Y(n_720) );
AND2x4_ASAP7_75t_L g739 ( .A(n_467), .B(n_740), .Y(n_739) );
OR2x6_ASAP7_75t_L g467 ( .A(n_468), .B(n_474), .Y(n_467) );
INVx2_ASAP7_75t_SL g652 ( .A(n_475), .Y(n_652) );
OR2x2_ASAP7_75t_L g475 ( .A(n_476), .B(n_484), .Y(n_475) );
AND2x2_ASAP7_75t_L g559 ( .A(n_476), .B(n_536), .Y(n_559) );
INVx2_ASAP7_75t_L g586 ( .A(n_476), .Y(n_586) );
INVx2_ASAP7_75t_L g616 ( .A(n_476), .Y(n_616) );
AND2x2_ASAP7_75t_L g630 ( .A(n_476), .B(n_535), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_478), .B(n_482), .Y(n_477) );
AND2x2_ASAP7_75t_L g560 ( .A(n_484), .B(n_561), .Y(n_560) );
INVx2_ASAP7_75t_L g583 ( .A(n_484), .Y(n_583) );
BUFx3_ASAP7_75t_L g597 ( .A(n_484), .Y(n_597) );
AND2x2_ASAP7_75t_L g626 ( .A(n_484), .B(n_627), .Y(n_626) );
AND2x4_ASAP7_75t_L g484 ( .A(n_485), .B(n_486), .Y(n_484) );
AND2x4_ASAP7_75t_L g531 ( .A(n_485), .B(n_486), .Y(n_531) );
AND2x4_ASAP7_75t_L g488 ( .A(n_489), .B(n_492), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_490), .B(n_491), .Y(n_489) );
NOR2x1p5_ASAP7_75t_L g495 ( .A(n_496), .B(n_497), .Y(n_495) );
INVx3_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g632 ( .A(n_499), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_500), .B(n_510), .Y(n_499) );
OR2x2_ASAP7_75t_L g743 ( .A(n_500), .B(n_544), .Y(n_743) );
INVx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
AND2x2_ASAP7_75t_L g599 ( .A(n_501), .B(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_501), .B(n_510), .Y(n_660) );
OR2x2_ASAP7_75t_L g758 ( .A(n_501), .B(n_680), .Y(n_758) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
AND2x2_ASAP7_75t_L g569 ( .A(n_502), .B(n_545), .Y(n_569) );
OR2x2_ASAP7_75t_SL g579 ( .A(n_502), .B(n_580), .Y(n_579) );
INVx4_ASAP7_75t_L g590 ( .A(n_502), .Y(n_590) );
HB1xp67_ASAP7_75t_L g641 ( .A(n_502), .Y(n_641) );
NAND2x1_ASAP7_75t_L g647 ( .A(n_502), .B(n_546), .Y(n_647) );
AND2x2_ASAP7_75t_L g672 ( .A(n_502), .B(n_512), .Y(n_672) );
OR2x2_ASAP7_75t_L g693 ( .A(n_502), .B(n_576), .Y(n_693) );
OR2x6_ASAP7_75t_L g502 ( .A(n_503), .B(n_504), .Y(n_502) );
INVx1_ASAP7_75t_L g588 ( .A(n_510), .Y(n_588) );
O2A1O1Ixp33_ASAP7_75t_L g681 ( .A1(n_510), .A2(n_682), .B(n_685), .C(n_687), .Y(n_681) );
AND2x2_ASAP7_75t_L g754 ( .A(n_510), .B(n_530), .Y(n_754) );
AND2x2_ASAP7_75t_L g510 ( .A(n_511), .B(n_519), .Y(n_510) );
INVx1_ASAP7_75t_L g621 ( .A(n_511), .Y(n_621) );
AND2x2_ASAP7_75t_L g691 ( .A(n_511), .B(n_546), .Y(n_691) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g565 ( .A(n_512), .Y(n_565) );
OR2x2_ASAP7_75t_L g580 ( .A(n_512), .B(n_546), .Y(n_580) );
INVx1_ASAP7_75t_L g596 ( .A(n_512), .Y(n_596) );
AND2x2_ASAP7_75t_L g608 ( .A(n_512), .B(n_519), .Y(n_608) );
HB1xp67_ASAP7_75t_L g714 ( .A(n_512), .Y(n_714) );
NOR2x1_ASAP7_75t_SL g545 ( .A(n_519), .B(n_546), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_521), .B(n_525), .Y(n_520) );
INVxp67_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_529), .B(n_532), .Y(n_528) );
OR2x2_ASAP7_75t_L g678 ( .A(n_529), .B(n_613), .Y(n_678) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_530), .B(n_696), .Y(n_695) );
OR2x2_ASAP7_75t_L g760 ( .A(n_530), .B(n_657), .Y(n_760) );
INVx3_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
AND2x2_ASAP7_75t_L g605 ( .A(n_531), .B(n_586), .Y(n_605) );
AND2x2_ASAP7_75t_L g701 ( .A(n_531), .B(n_614), .Y(n_701) );
INVx1_ASAP7_75t_L g618 ( .A(n_532), .Y(n_618) );
AND2x2_ASAP7_75t_L g532 ( .A(n_533), .B(n_534), .Y(n_532) );
INVx1_ASAP7_75t_L g668 ( .A(n_533), .Y(n_668) );
INVx2_ASAP7_75t_L g635 ( .A(n_534), .Y(n_635) );
HB1xp67_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
AND2x2_ASAP7_75t_L g585 ( .A(n_535), .B(n_586), .Y(n_585) );
INVx2_ASAP7_75t_L g615 ( .A(n_535), .Y(n_615) );
INVx1_ASAP7_75t_L g740 ( .A(n_535), .Y(n_740) );
INVx3_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
HB1xp67_ASAP7_75t_L g697 ( .A(n_536), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_538), .B(n_542), .Y(n_537) );
OR2x2_ASAP7_75t_L g711 ( .A(n_544), .B(n_712), .Y(n_711) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx2_ASAP7_75t_SL g566 ( .A(n_546), .Y(n_566) );
OR2x2_ASAP7_75t_L g589 ( .A(n_546), .B(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g600 ( .A(n_546), .B(n_576), .Y(n_600) );
AND2x2_ASAP7_75t_L g674 ( .A(n_546), .B(n_590), .Y(n_674) );
BUFx2_ASAP7_75t_L g757 ( .A(n_546), .Y(n_757) );
OR2x6_ASAP7_75t_L g546 ( .A(n_547), .B(n_554), .Y(n_546) );
AOI21xp5_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_562), .B(n_567), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_558), .B(n_560), .Y(n_557) );
AND2x2_ASAP7_75t_L g709 ( .A(n_558), .B(n_631), .Y(n_709) );
BUFx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g568 ( .A(n_559), .B(n_561), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_560), .B(n_630), .Y(n_731) );
INVx1_ASAP7_75t_L g761 ( .A(n_560), .Y(n_761) );
NAND2x1p5_ASAP7_75t_L g657 ( .A(n_561), .B(n_658), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_561), .B(n_697), .Y(n_734) );
INVxp67_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_564), .B(n_566), .Y(n_563) );
AND2x4_ASAP7_75t_SL g598 ( .A(n_564), .B(n_599), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_564), .B(n_592), .Y(n_745) );
INVx3_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
NOR2xp33_ASAP7_75t_L g703 ( .A(n_565), .B(n_647), .Y(n_703) );
AND2x2_ASAP7_75t_L g721 ( .A(n_565), .B(n_674), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_566), .B(n_608), .Y(n_624) );
A2O1A1Ixp33_ASAP7_75t_L g653 ( .A1(n_566), .A2(n_612), .B(n_654), .C(n_659), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_566), .B(n_684), .Y(n_683) );
AND2x2_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
AOI221xp5_ASAP7_75t_L g748 ( .A1(n_568), .A2(n_641), .B1(n_749), .B2(n_755), .C(n_759), .Y(n_748) );
INVx1_ASAP7_75t_SL g736 ( .A(n_569), .Y(n_736) );
OAI221xp5_ASAP7_75t_L g570 ( .A1(n_571), .A2(n_581), .B1(n_587), .B2(n_591), .C(n_794), .Y(n_570) );
INVx2_ASAP7_75t_SL g571 ( .A(n_572), .Y(n_571) );
AND2x4_ASAP7_75t_L g572 ( .A(n_573), .B(n_578), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g646 ( .A(n_575), .Y(n_646) );
HB1xp67_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g620 ( .A(n_576), .B(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g651 ( .A(n_576), .B(n_596), .Y(n_651) );
INVx2_ASAP7_75t_L g684 ( .A(n_576), .Y(n_684) );
INVx3_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
OAI32xp33_ASAP7_75t_L g735 ( .A1(n_579), .A2(n_626), .A3(n_657), .B1(n_736), .B2(n_737), .Y(n_735) );
OR2x2_ASAP7_75t_L g706 ( .A(n_580), .B(n_693), .Y(n_706) );
INVx1_ASAP7_75t_L g716 ( .A(n_581), .Y(n_716) );
OR2x2_ASAP7_75t_L g581 ( .A(n_582), .B(n_584), .Y(n_581) );
INVx2_ASAP7_75t_L g631 ( .A(n_582), .Y(n_631) );
AND2x2_ASAP7_75t_L g702 ( .A(n_582), .B(n_677), .Y(n_702) );
OR2x2_ASAP7_75t_L g733 ( .A(n_582), .B(n_734), .Y(n_733) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_583), .B(n_638), .Y(n_637) );
INVx1_ASAP7_75t_SL g584 ( .A(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g627 ( .A(n_586), .Y(n_627) );
OR2x2_ASAP7_75t_L g587 ( .A(n_588), .B(n_589), .Y(n_587) );
INVx2_ASAP7_75t_SL g592 ( .A(n_589), .Y(n_592) );
OR2x2_ASAP7_75t_L g679 ( .A(n_589), .B(n_680), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_590), .B(n_608), .Y(n_607) );
NOR2xp67_ASAP7_75t_L g713 ( .A(n_590), .B(n_714), .Y(n_713) );
BUFx2_ASAP7_75t_L g726 ( .A(n_590), .Y(n_726) );
A2O1A1Ixp33_ASAP7_75t_L g591 ( .A1(n_592), .A2(n_593), .B(n_598), .C(n_601), .Y(n_591) );
AND2x2_ASAP7_75t_L g741 ( .A(n_593), .B(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
OR2x2_ASAP7_75t_L g594 ( .A(n_595), .B(n_597), .Y(n_594) );
BUFx2_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
OR2x2_ASAP7_75t_L g667 ( .A(n_597), .B(n_668), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_597), .B(n_601), .Y(n_688) );
AND2x2_ASAP7_75t_L g719 ( .A(n_597), .B(n_720), .Y(n_719) );
O2A1O1Ixp33_ASAP7_75t_L g729 ( .A1(n_599), .A2(n_730), .B(n_732), .C(n_735), .Y(n_729) );
AOI222xp33_ASAP7_75t_L g603 ( .A1(n_600), .A2(n_604), .B1(n_606), .B2(n_609), .C1(n_617), .C2(n_619), .Y(n_603) );
AND2x2_ASAP7_75t_L g671 ( .A(n_600), .B(n_672), .Y(n_671) );
AND2x2_ASAP7_75t_L g604 ( .A(n_601), .B(n_605), .Y(n_604) );
INVx2_ASAP7_75t_SL g625 ( .A(n_601), .Y(n_625) );
NAND4xp25_ASAP7_75t_L g602 ( .A(n_603), .B(n_622), .C(n_643), .D(n_653), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_605), .B(n_611), .Y(n_665) );
INVx1_ASAP7_75t_SL g606 ( .A(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g673 ( .A(n_608), .B(n_674), .Y(n_673) );
INVx2_ASAP7_75t_SL g680 ( .A(n_608), .Y(n_680) );
AND2x2_ASAP7_75t_L g609 ( .A(n_610), .B(n_612), .Y(n_609) );
A2O1A1Ixp33_ASAP7_75t_L g643 ( .A1(n_610), .A2(n_644), .B(n_648), .C(n_652), .Y(n_643) );
INVx2_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_611), .B(n_626), .Y(n_747) );
OR2x2_ASAP7_75t_L g751 ( .A(n_611), .B(n_637), .Y(n_751) );
INVx1_ASAP7_75t_L g724 ( .A(n_612), .Y(n_724) );
INVx2_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
AND2x2_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
INVx1_ASAP7_75t_SL g658 ( .A(n_615), .Y(n_658) );
INVx1_ASAP7_75t_L g638 ( .A(n_616), .Y(n_638) );
INVx2_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_618), .B(n_655), .Y(n_654) );
BUFx2_ASAP7_75t_SL g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g642 ( .A(n_620), .Y(n_642) );
AOI322xp5_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_625), .A3(n_626), .B1(n_628), .B2(n_632), .C1(n_633), .C2(n_639), .Y(n_622) );
INVxp67_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
O2A1O1Ixp33_ASAP7_75t_SL g704 ( .A1(n_625), .A2(n_705), .B(n_706), .C(n_707), .Y(n_704) );
INVx1_ASAP7_75t_L g727 ( .A(n_626), .Y(n_727) );
NOR2xp67_ASAP7_75t_L g628 ( .A(n_629), .B(n_631), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g685 ( .A(n_631), .B(n_686), .Y(n_685) );
AND2x2_ASAP7_75t_L g633 ( .A(n_634), .B(n_636), .Y(n_633) );
INVx2_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx2_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
HB1xp67_ASAP7_75t_L g707 ( .A(n_637), .Y(n_707) );
INVx2_ASAP7_75t_SL g639 ( .A(n_640), .Y(n_639) );
OR2x2_ASAP7_75t_L g640 ( .A(n_641), .B(n_642), .Y(n_640) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
OR2x2_ASAP7_75t_L g645 ( .A(n_646), .B(n_647), .Y(n_645) );
INVx3_ASAP7_75t_L g650 ( .A(n_647), .Y(n_650) );
OR2x2_ASAP7_75t_L g718 ( .A(n_647), .B(n_680), .Y(n_718) );
NOR2xp33_ASAP7_75t_L g763 ( .A(n_647), .B(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_650), .B(n_651), .Y(n_649) );
INVx1_ASAP7_75t_SL g750 ( .A(n_651), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_652), .B(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
NAND3xp33_ASAP7_75t_SL g755 ( .A(n_660), .B(n_756), .C(n_758), .Y(n_755) );
NOR3xp33_ASAP7_75t_SL g661 ( .A(n_662), .B(n_699), .C(n_728), .Y(n_661) );
NAND2xp5_ASAP7_75t_SL g662 ( .A(n_663), .B(n_681), .Y(n_662) );
O2A1O1Ixp33_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_666), .B(n_669), .C(n_675), .Y(n_663) );
OAI31xp33_ASAP7_75t_L g708 ( .A1(n_664), .A2(n_686), .A3(n_709), .B(n_710), .Y(n_708) );
INVx1_ASAP7_75t_SL g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_SL g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
NOR2xp33_ASAP7_75t_L g670 ( .A(n_671), .B(n_673), .Y(n_670) );
INVx2_ASAP7_75t_L g723 ( .A(n_671), .Y(n_723) );
INVx1_ASAP7_75t_L g698 ( .A(n_673), .Y(n_698) );
AOI21xp5_ASAP7_75t_L g675 ( .A1(n_676), .A2(n_678), .B(n_679), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
OR2x2_ASAP7_75t_L g725 ( .A(n_683), .B(n_726), .Y(n_725) );
INVxp67_ASAP7_75t_L g764 ( .A(n_684), .Y(n_764) );
OAI22xp33_ASAP7_75t_SL g687 ( .A1(n_688), .A2(n_689), .B1(n_694), .B2(n_698), .Y(n_687) );
INVx3_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
AND2x4_ASAP7_75t_L g690 ( .A(n_691), .B(n_692), .Y(n_690) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
HB1xp67_ASAP7_75t_L g705 ( .A(n_693), .Y(n_705) );
OR2x2_ASAP7_75t_L g756 ( .A(n_693), .B(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
NAND3xp33_ASAP7_75t_SL g699 ( .A(n_700), .B(n_708), .C(n_715), .Y(n_699) );
O2A1O1Ixp33_ASAP7_75t_L g700 ( .A1(n_701), .A2(n_702), .B(n_703), .C(n_704), .Y(n_700) );
INVx2_ASAP7_75t_L g737 ( .A(n_701), .Y(n_737) );
INVx1_ASAP7_75t_SL g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
AOI221xp5_ASAP7_75t_L g715 ( .A1(n_716), .A2(n_717), .B1(n_719), .B2(n_721), .C(n_722), .Y(n_715) );
INVx2_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
OAI22xp33_ASAP7_75t_L g722 ( .A1(n_723), .A2(n_724), .B1(n_725), .B2(n_727), .Y(n_722) );
NAND3xp33_ASAP7_75t_SL g728 ( .A(n_729), .B(n_738), .C(n_748), .Y(n_728) );
INVxp33_ASAP7_75t_SL g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_SL g732 ( .A(n_733), .Y(n_732) );
AOI22xp5_ASAP7_75t_L g738 ( .A1(n_739), .A2(n_741), .B1(n_744), .B2(n_746), .Y(n_738) );
INVx2_ASAP7_75t_L g752 ( .A(n_739), .Y(n_752) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
OAI22xp5_ASAP7_75t_L g749 ( .A1(n_750), .A2(n_751), .B1(n_752), .B2(n_753), .Y(n_749) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
OAI22xp33_ASAP7_75t_SL g759 ( .A1(n_758), .A2(n_760), .B1(n_761), .B2(n_762), .Y(n_759) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
INVx4_ASAP7_75t_SL g765 ( .A(n_766), .Y(n_765) );
CKINVDCx6p67_ASAP7_75t_R g773 ( .A(n_766), .Y(n_773) );
INVx3_ASAP7_75t_SL g766 ( .A(n_767), .Y(n_766) );
CKINVDCx5p33_ASAP7_75t_R g767 ( .A(n_768), .Y(n_767) );
NOR2xp33_ASAP7_75t_L g774 ( .A(n_775), .B(n_776), .Y(n_774) );
INVx1_ASAP7_75t_SL g776 ( .A(n_777), .Y(n_776) );
INVx2_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_780), .B(n_782), .Y(n_779) );
INVx1_ASAP7_75t_SL g780 ( .A(n_781), .Y(n_780) );
CKINVDCx16_ASAP7_75t_R g787 ( .A(n_784), .Y(n_787) );
INVx1_ASAP7_75t_SL g788 ( .A(n_789), .Y(n_788) );
INVx1_ASAP7_75t_SL g789 ( .A(n_790), .Y(n_789) );
endmodule