module real_jpeg_32573_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_83;
wire n_78;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_292;
wire n_221;
wire n_249;
wire n_288;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_276;
wire n_163;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_105;
wire n_173;
wire n_40;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_184;
wire n_56;
wire n_48;
wire n_164;
wire n_200;
wire n_293;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_267;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_285;
wire n_268;
wire n_42;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_148;
wire n_19;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_137;
wire n_31;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_195;
wire n_61;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_278;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_240;
wire n_185;
wire n_209;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_210;
wire n_53;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_283;
wire n_85;
wire n_102;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

HB1xp67_ASAP7_75t_L g59 ( 
.A(n_0),
.Y(n_59)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_0),
.Y(n_171)
);

BUFx12f_ASAP7_75t_L g270 ( 
.A(n_0),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_0),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_1),
.A2(n_144),
.B1(n_148),
.B2(n_152),
.Y(n_143)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_1),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_1),
.A2(n_152),
.B1(n_210),
.B2(n_212),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_1),
.A2(n_152),
.B1(n_240),
.B2(n_242),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_2),
.A2(n_105),
.B1(n_106),
.B2(n_110),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_2),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_2),
.A2(n_105),
.B1(n_265),
.B2(n_267),
.Y(n_264)
);

OAI32xp33_ASAP7_75t_L g20 ( 
.A1(n_3),
.A2(n_21),
.A3(n_25),
.B1(n_29),
.B2(n_36),
.Y(n_20)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_3),
.A2(n_37),
.B1(n_133),
.B2(n_137),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_3),
.A2(n_43),
.B1(n_209),
.B2(n_215),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_3),
.B(n_281),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_5),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_5),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_6),
.A2(n_49),
.B1(n_53),
.B2(n_54),
.Y(n_48)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_6),
.A2(n_53),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

OAI22x1_ASAP7_75t_SL g60 ( 
.A1(n_7),
.A2(n_61),
.B1(n_65),
.B2(n_66),
.Y(n_60)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_7),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_8),
.A2(n_77),
.B1(n_82),
.B2(n_83),
.Y(n_76)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_8),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_8),
.A2(n_82),
.B1(n_158),
.B2(n_162),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_8),
.A2(n_82),
.B1(n_227),
.B2(n_229),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_9),
.A2(n_173),
.B1(n_174),
.B2(n_178),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_9),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_10),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_10),
.Y(n_85)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_11),
.Y(n_187)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_12),
.Y(n_91)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_12),
.Y(n_95)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_12),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_13),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_13),
.Y(n_147)
);

HAxp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_202),
.CON(n_14),
.SN(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_201),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

NOR2xp67_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_153),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_18),
.B(n_153),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_74),
.C(n_116),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_19),
.B(n_290),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_41),
.B1(n_72),
.B2(n_73),
.Y(n_19)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_20),
.B(n_73),
.Y(n_200)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_24),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_24),
.Y(n_151)
);

OAI21xp33_ASAP7_75t_SL g245 ( 
.A1(n_25),
.A2(n_37),
.B(n_246),
.Y(n_245)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_28),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_28),
.Y(n_244)
);

AO21x2_ASAP7_75t_L g118 ( 
.A1(n_29),
.A2(n_119),
.B(n_123),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_33),
.Y(n_29)
);

AOI22x1_ASAP7_75t_L g183 ( 
.A1(n_30),
.A2(n_184),
.B1(n_188),
.B2(n_189),
.Y(n_183)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_32),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_32),
.Y(n_161)
);

BUFx5_ASAP7_75t_L g165 ( 
.A(n_32),
.Y(n_165)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_33),
.Y(n_120)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_34),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_35),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_38),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_37),
.B(n_182),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_37),
.B(n_215),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_37),
.B(n_114),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_37),
.B(n_247),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_39),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_40),
.Y(n_89)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_40),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_40),
.Y(n_128)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_48),
.B1(n_58),
.B2(n_60),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_42),
.A2(n_60),
.B1(n_168),
.B2(n_172),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_42),
.A2(n_262),
.B1(n_263),
.B2(n_268),
.Y(n_261)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_43),
.A2(n_209),
.B1(n_226),
.B2(n_233),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_43),
.A2(n_264),
.B1(n_276),
.B2(n_278),
.Y(n_275)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_46),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_45),
.Y(n_218)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_46),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_47),
.Y(n_102)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_47),
.Y(n_177)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_47),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_48),
.Y(n_278)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx4f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_63),
.Y(n_103)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_63),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_63),
.Y(n_232)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_64),
.Y(n_223)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_71),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_71),
.Y(n_228)
);

BUFx2_ASAP7_75t_L g267 ( 
.A(n_71),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_74),
.A2(n_116),
.B1(n_117),
.B2(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_74),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_86),
.B1(n_104),
.B2(n_113),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_76),
.A2(n_87),
.B1(n_114),
.B2(n_283),
.Y(n_282)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_77),
.Y(n_195)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_81),
.Y(n_130)
);

INVx3_ASAP7_75t_SL g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_85),
.Y(n_241)
);

AO22x1_ASAP7_75t_SL g238 ( 
.A1(n_86),
.A2(n_113),
.B1(n_239),
.B2(n_245),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_87),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_87),
.A2(n_114),
.B1(n_194),
.B2(n_199),
.Y(n_193)
);

AO21x2_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_92),
.B(n_97),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_88),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_90),
.Y(n_88)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_89),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_90),
.A2(n_98),
.B1(n_101),
.B2(n_103),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_96),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_97),
.Y(n_115)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_100),
.Y(n_255)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_104),
.Y(n_199)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_SL g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx4f_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_132),
.B1(n_141),
.B2(n_143),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_118),
.A2(n_143),
.B1(n_156),
.B2(n_157),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_121),
.Y(n_119)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_122),
.Y(n_188)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_124),
.Y(n_142)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_124),
.Y(n_281)
);

OA22x2_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_127),
.B1(n_129),
.B2(n_131),
.Y(n_124)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_142),
.Y(n_156)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx8_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_192),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_166),
.Y(n_154)
);

BUFx2_ASAP7_75t_SL g158 ( 
.A(n_159),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_181),
.B1(n_190),
.B2(n_191),
.Y(n_166)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_167),
.Y(n_190)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_181),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx4_ASAP7_75t_SL g189 ( 
.A(n_186),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_200),
.Y(n_192)
);

INVx2_ASAP7_75t_SL g196 ( 
.A(n_197),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

OAI31xp67_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_286),
.A3(n_292),
.B(n_293),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_271),
.B(n_272),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_236),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_224),
.B(n_235),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_208),
.B(n_219),
.Y(n_207)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx3_ASAP7_75t_SL g215 ( 
.A(n_216),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_217),
.Y(n_233)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_223),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_234),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_225),
.B(n_234),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_226),
.Y(n_262)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_232),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_237),
.B(n_261),
.Y(n_236)
);

OR2x2_ASAP7_75t_L g271 ( 
.A(n_237),
.B(n_261),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_249),
.Y(n_237)
);

NAND2xp33_ASAP7_75t_R g273 ( 
.A(n_238),
.B(n_249),
.Y(n_273)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_239),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx5_ASAP7_75t_L g248 ( 
.A(n_241),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_246),
.Y(n_256)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

AO22x1_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_256),
.B1(n_257),
.B2(n_260),
.Y(n_249)
);

NAND2xp33_ASAP7_75t_SL g250 ( 
.A(n_251),
.B(n_253),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

BUFx2_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

BUFx2_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx5_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx8_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_273),
.B(n_274),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_279),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_275),
.B(n_284),
.C(n_288),
.Y(n_287)
);

INVx5_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_282),
.B1(n_284),
.B2(n_285),
.Y(n_279)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_280),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_282),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_282),
.Y(n_288)
);

NOR2xp67_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_289),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_287),
.B(n_289),
.Y(n_293)
);


endmodule