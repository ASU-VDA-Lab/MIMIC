module fake_jpeg_11881_n_157 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_157);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_157;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_93;
wire n_54;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_33),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_30),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_0),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_6),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_23),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_39),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_17),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_19),
.B(n_10),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_5),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_8),
.Y(n_62)
);

BUFx12_ASAP7_75t_L g63 ( 
.A(n_9),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_12),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_65),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_0),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_66),
.B(n_67),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_52),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_45),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_68),
.A2(n_70),
.B1(n_72),
.B2(n_73),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_1),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_69),
.B(n_60),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_57),
.A2(n_26),
.B1(n_43),
.B2(n_42),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_45),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_55),
.A2(n_27),
.B1(n_41),
.B2(n_40),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_66),
.B(n_59),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_77),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_59),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_78),
.B(n_81),
.Y(n_104)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_67),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_82),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_73),
.B(n_47),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_56),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_71),
.B(n_64),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_79),
.Y(n_100)
);

BUFx12_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_84),
.Y(n_92)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_77),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_93),
.B(n_95),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_75),
.A2(n_55),
.B1(n_48),
.B2(n_62),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_94),
.A2(n_103),
.B1(n_63),
.B2(n_8),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_64),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_51),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_96),
.B(n_98),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_51),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_86),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_99),
.B(n_58),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_106),
.Y(n_111)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_102),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_75),
.A2(n_48),
.B1(n_62),
.B2(n_61),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_87),
.A2(n_61),
.B1(n_54),
.B2(n_53),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_105),
.A2(n_84),
.B1(n_63),
.B2(n_52),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_49),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_102),
.B(n_85),
.Y(n_107)
);

OAI21xp33_ASAP7_75t_L g139 ( 
.A1(n_107),
.A2(n_25),
.B(n_31),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_100),
.B(n_28),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_108),
.B(n_109),
.Y(n_134)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_101),
.A2(n_84),
.B(n_58),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_110),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_94),
.A2(n_103),
.B1(n_101),
.B2(n_90),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_112),
.A2(n_121),
.B1(n_15),
.B2(n_20),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_114),
.B(n_116),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_104),
.A2(n_63),
.B(n_52),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_115),
.A2(n_122),
.B(n_125),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_89),
.B(n_4),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_6),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_120),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_118),
.A2(n_126),
.B1(n_127),
.B2(n_14),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_91),
.B(n_7),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_92),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_90),
.B(n_44),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_123),
.B(n_13),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_7),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_97),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_100),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_128),
.B(n_129),
.Y(n_146)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_113),
.Y(n_129)
);

AO22x1_ASAP7_75t_L g131 ( 
.A1(n_115),
.A2(n_121),
.B1(n_111),
.B2(n_110),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_131),
.B(n_109),
.Y(n_143)
);

AO21x1_ASAP7_75t_L g148 ( 
.A1(n_132),
.A2(n_139),
.B(n_134),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_135),
.A2(n_137),
.B1(n_140),
.B2(n_35),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_108),
.A2(n_15),
.B1(n_21),
.B2(n_22),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_124),
.A2(n_119),
.B1(n_123),
.B2(n_118),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_107),
.Y(n_141)
);

NAND3xp33_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_127),
.C(n_107),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_142),
.B(n_147),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_143),
.A2(n_144),
.B(n_148),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_130),
.A2(n_32),
.B(n_34),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_145),
.A2(n_128),
.B1(n_139),
.B2(n_138),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_136),
.A2(n_36),
.B(n_37),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_150),
.B(n_133),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_149),
.A2(n_143),
.B(n_146),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_152),
.B(n_153),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_154),
.A2(n_131),
.B(n_130),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_151),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_133),
.Y(n_157)
);


endmodule