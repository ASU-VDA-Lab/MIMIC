module real_aes_7117_n_350 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_323, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_346, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_350);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_323;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_346;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_350;
wire n_480;
wire n_1073;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_1066;
wire n_684;
wire n_390;
wire n_1096;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_1092;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_905;
wire n_1067;
wire n_878;
wire n_665;
wire n_991;
wire n_667;
wire n_580;
wire n_577;
wire n_1004;
wire n_469;
wire n_987;
wire n_362;
wire n_759;
wire n_979;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_540;
wire n_1064;
wire n_1075;
wire n_657;
wire n_900;
wire n_841;
wire n_718;
wire n_355;
wire n_669;
wire n_1091;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_364;
wire n_555;
wire n_421;
wire n_766;
wire n_852;
wire n_974;
wire n_857;
wire n_919;
wire n_1089;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_491;
wire n_894;
wire n_923;
wire n_1034;
wire n_952;
wire n_429;
wire n_752;
wire n_448;
wire n_556;
wire n_545;
wire n_593;
wire n_460;
wire n_937;
wire n_989;
wire n_773;
wire n_401;
wire n_538;
wire n_353;
wire n_431;
wire n_1044;
wire n_963;
wire n_865;
wire n_551;
wire n_666;
wire n_537;
wire n_884;
wire n_560;
wire n_660;
wire n_1094;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_983;
wire n_767;
wire n_889;
wire n_696;
wire n_955;
wire n_975;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_1046;
wire n_677;
wire n_958;
wire n_1021;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_1093;
wire n_870;
wire n_961;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_415;
wire n_572;
wire n_815;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_816;
wire n_539;
wire n_400;
wire n_626;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_990;
wire n_550;
wire n_966;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_356;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_994;
wire n_892;
wire n_1078;
wire n_495;
wire n_528;
wire n_578;
wire n_370;
wire n_1072;
wire n_384;
wire n_938;
wire n_744;
wire n_352;
wire n_935;
wire n_824;
wire n_951;
wire n_467;
wire n_875;
wire n_774;
wire n_992;
wire n_813;
wire n_791;
wire n_981;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_976;
wire n_1049;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_1086;
wire n_1070;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_962;
wire n_1082;
wire n_468;
wire n_755;
wire n_532;
wire n_746;
wire n_656;
wire n_1025;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_523;
wire n_909;
wire n_996;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_801;
wire n_383;
wire n_529;
wire n_504;
wire n_455;
wire n_725;
wire n_973;
wire n_1081;
wire n_671;
wire n_960;
wire n_1084;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_885;
wire n_1059;
wire n_950;
wire n_381;
wire n_993;
wire n_493;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_1013;
wire n_1017;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_641;
wire n_1063;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_745;
wire n_722;
wire n_867;
wire n_398;
wire n_688;
wire n_425;
wire n_609;
wire n_1042;
wire n_879;
wire n_1006;
wire n_363;
wire n_417;
wire n_607;
wire n_449;
wire n_754;
wire n_690;
wire n_629;
wire n_1053;
wire n_499;
wire n_508;
wire n_706;
wire n_901;
wire n_561;
wire n_970;
wire n_947;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_1012;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_986;
wire n_1083;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1031;
wire n_1037;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_999;
wire n_490;
wire n_913;
wire n_619;
wire n_391;
wire n_1095;
wire n_360;
wire n_1060;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_1080;
wire n_361;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_985;
wire n_777;
wire n_1077;
wire n_488;
wire n_501;
wire n_1041;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_957;
wire n_995;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_351;
wire n_945;
wire n_898;
wire n_604;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_997;
wire n_569;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_1079;
wire n_579;
wire n_1033;
wire n_699;
wire n_533;
wire n_1028;
wire n_1000;
wire n_1003;
wire n_366;
wire n_727;
wire n_1014;
wire n_649;
wire n_358;
wire n_397;
wire n_385;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_851;
wire n_470;
wire n_915;
wire n_1002;
wire n_934;
wire n_1001;
wire n_494;
wire n_711;
wire n_864;
wire n_1027;
wire n_377;
wire n_1058;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_1085;
wire n_382;
wire n_845;
wire n_1043;
wire n_850;
wire n_354;
wire n_720;
wire n_972;
wire n_968;
wire n_435;
wire n_1026;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_1068;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_1005;
wire n_939;
wire n_487;
wire n_831;
wire n_653;
wire n_365;
wire n_526;
wire n_928;
wire n_637;
wire n_899;
wire n_692;
wire n_544;
wire n_789;
wire n_1087;
wire n_1051;
wire n_389;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_922;
wire n_926;
wire n_942;
wire n_1048;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_1052;
wire n_787;
wire n_1071;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_959;
wire n_715;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_741;
wire n_753;
wire n_623;
wire n_1032;
wire n_721;
wire n_446;
wire n_681;
wire n_1090;
wire n_359;
wire n_982;
wire n_456;
wire n_717;
wire n_712;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_762;
wire n_575;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_1074;
wire n_674;
wire n_644;
wire n_836;
wire n_888;
wire n_793;
wire n_1056;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_1045;
wire n_465;
wire n_473;
wire n_566;
wire n_719;
wire n_837;
wire n_967;
wire n_871;
wire n_474;
wire n_829;
wire n_1030;
wire n_988;
wire n_1055;
wire n_1088;
wire n_921;
wire n_375;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_1036;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_1040;
wire n_393;
wire n_703;
wire n_652;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_1076;
wire n_804;
wire n_396;
wire n_447;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_1039;
wire n_574;
wire n_1069;
wire n_1024;
wire n_842;
wire n_1061;
wire n_849;
wire n_554;
wire n_475;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_SL g757 ( .A1(n_0), .A2(n_262), .B1(n_450), .B2(n_585), .Y(n_757) );
CKINVDCx20_ASAP7_75t_R g808 ( .A(n_1), .Y(n_808) );
CKINVDCx20_ASAP7_75t_R g659 ( .A(n_2), .Y(n_659) );
CKINVDCx20_ASAP7_75t_R g534 ( .A(n_3), .Y(n_534) );
AOI211xp5_ASAP7_75t_L g350 ( .A1(n_4), .A2(n_351), .B(n_359), .C(n_1043), .Y(n_350) );
AOI22xp33_ASAP7_75t_L g1077 ( .A1(n_5), .A2(n_82), .B1(n_512), .B2(n_1078), .Y(n_1077) );
CKINVDCx20_ASAP7_75t_R g743 ( .A(n_6), .Y(n_743) );
AOI22xp33_ASAP7_75t_L g925 ( .A1(n_7), .A2(n_47), .B1(n_607), .B2(n_895), .Y(n_925) );
AOI22x1_ASAP7_75t_L g977 ( .A1(n_8), .A2(n_978), .B1(n_1005), .B2(n_1006), .Y(n_977) );
INVx1_ASAP7_75t_L g1005 ( .A(n_8), .Y(n_1005) );
CKINVDCx20_ASAP7_75t_R g477 ( .A(n_9), .Y(n_477) );
AO22x2_ASAP7_75t_L g371 ( .A1(n_10), .A2(n_204), .B1(n_372), .B2(n_373), .Y(n_371) );
INVx1_ASAP7_75t_L g1041 ( .A(n_10), .Y(n_1041) );
AOI22xp33_ASAP7_75t_L g794 ( .A1(n_11), .A2(n_144), .B1(n_587), .B2(n_795), .Y(n_794) );
CKINVDCx20_ASAP7_75t_R g937 ( .A(n_12), .Y(n_937) );
CKINVDCx20_ASAP7_75t_R g1003 ( .A(n_13), .Y(n_1003) );
CKINVDCx20_ASAP7_75t_R g884 ( .A(n_14), .Y(n_884) );
CKINVDCx20_ASAP7_75t_R g811 ( .A(n_15), .Y(n_811) );
AOI22xp33_ASAP7_75t_L g758 ( .A1(n_16), .A2(n_267), .B1(n_553), .B2(n_723), .Y(n_758) );
CKINVDCx20_ASAP7_75t_R g869 ( .A(n_17), .Y(n_869) );
AOI22xp33_ASAP7_75t_L g1083 ( .A1(n_18), .A2(n_293), .B1(n_502), .B2(n_795), .Y(n_1083) );
CKINVDCx20_ASAP7_75t_R g734 ( .A(n_19), .Y(n_734) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_20), .A2(n_141), .B1(n_648), .B2(n_649), .Y(n_647) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_21), .Y(n_750) );
CKINVDCx20_ASAP7_75t_R g714 ( .A(n_22), .Y(n_714) );
CKINVDCx20_ASAP7_75t_R g916 ( .A(n_23), .Y(n_916) );
AOI22xp33_ASAP7_75t_L g949 ( .A1(n_24), .A2(n_332), .B1(n_438), .B2(n_517), .Y(n_949) );
CKINVDCx20_ASAP7_75t_R g837 ( .A(n_25), .Y(n_837) );
CKINVDCx20_ASAP7_75t_R g728 ( .A(n_26), .Y(n_728) );
AOI222xp33_ASAP7_75t_L g969 ( .A1(n_27), .A2(n_48), .B1(n_320), .B2(n_567), .C1(n_601), .C2(n_970), .Y(n_969) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_28), .A2(n_110), .B1(n_502), .B2(n_504), .Y(n_501) );
CKINVDCx20_ASAP7_75t_R g1061 ( .A(n_29), .Y(n_1061) );
AO22x2_ASAP7_75t_L g375 ( .A1(n_30), .A2(n_95), .B1(n_372), .B2(n_376), .Y(n_375) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_31), .A2(n_345), .B1(n_512), .B2(n_513), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g967 ( .A1(n_32), .A2(n_225), .B1(n_504), .B2(n_732), .Y(n_967) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_33), .A2(n_100), .B1(n_430), .B2(n_582), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g909 ( .A1(n_34), .A2(n_146), .B1(n_779), .B2(n_910), .Y(n_909) );
AOI22xp5_ASAP7_75t_L g826 ( .A1(n_35), .A2(n_252), .B1(n_507), .B2(n_827), .Y(n_826) );
CKINVDCx20_ASAP7_75t_R g453 ( .A(n_36), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_37), .B(n_572), .Y(n_571) );
AOI22xp5_ASAP7_75t_SL g760 ( .A1(n_38), .A2(n_761), .B1(n_762), .B2(n_784), .Y(n_760) );
INVx1_ASAP7_75t_L g784 ( .A(n_38), .Y(n_784) );
AOI22xp33_ASAP7_75t_L g712 ( .A1(n_39), .A2(n_271), .B1(n_422), .B2(n_642), .Y(n_712) );
AOI22xp5_ASAP7_75t_L g838 ( .A1(n_40), .A2(n_198), .B1(n_413), .B2(n_422), .Y(n_838) );
AOI22xp33_ASAP7_75t_L g777 ( .A1(n_41), .A2(n_223), .B1(n_778), .B2(n_779), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_42), .B(n_392), .Y(n_644) );
CKINVDCx20_ASAP7_75t_R g999 ( .A(n_43), .Y(n_999) );
AOI222xp33_ASAP7_75t_L g1089 ( .A1(n_44), .A2(n_272), .B1(n_291), .B2(n_368), .C1(n_575), .C2(n_970), .Y(n_1089) );
CKINVDCx20_ASAP7_75t_R g807 ( .A(n_45), .Y(n_807) );
CKINVDCx20_ASAP7_75t_R g877 ( .A(n_46), .Y(n_877) );
AOI22xp33_ASAP7_75t_L g798 ( .A1(n_49), .A2(n_221), .B1(n_690), .B2(n_799), .Y(n_798) );
AOI22xp33_ASAP7_75t_L g990 ( .A1(n_50), .A2(n_116), .B1(n_801), .B2(n_991), .Y(n_990) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_51), .B(n_674), .Y(n_673) );
AOI22xp33_ASAP7_75t_L g911 ( .A1(n_52), .A2(n_297), .B1(n_618), .B2(n_912), .Y(n_911) );
AOI22xp33_ASAP7_75t_SL g856 ( .A1(n_53), .A2(n_251), .B1(n_440), .B2(n_658), .Y(n_856) );
CKINVDCx20_ASAP7_75t_R g538 ( .A(n_54), .Y(n_538) );
CKINVDCx20_ASAP7_75t_R g893 ( .A(n_55), .Y(n_893) );
INVx1_ASAP7_75t_L g605 ( .A(n_56), .Y(n_605) );
CKINVDCx20_ASAP7_75t_R g448 ( .A(n_57), .Y(n_448) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_58), .A2(n_90), .B1(n_476), .B2(n_504), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g617 ( .A1(n_59), .A2(n_317), .B1(n_618), .B2(n_619), .Y(n_617) );
CKINVDCx20_ASAP7_75t_R g383 ( .A(n_60), .Y(n_383) );
AOI22xp33_ASAP7_75t_L g1065 ( .A1(n_61), .A2(n_84), .B1(n_438), .B2(n_1066), .Y(n_1065) );
CKINVDCx20_ASAP7_75t_R g933 ( .A(n_62), .Y(n_933) );
AOI22xp33_ASAP7_75t_L g397 ( .A1(n_63), .A2(n_228), .B1(n_398), .B2(n_403), .Y(n_397) );
AOI222xp33_ASAP7_75t_L g894 ( .A1(n_64), .A2(n_257), .B1(n_316), .B2(n_601), .C1(n_674), .C2(n_895), .Y(n_894) );
AOI22xp5_ASAP7_75t_L g641 ( .A1(n_65), .A2(n_235), .B1(n_422), .B2(n_642), .Y(n_641) );
AOI22xp33_ASAP7_75t_L g968 ( .A1(n_66), .A2(n_270), .B1(n_551), .B2(n_554), .Y(n_968) );
AOI22xp5_ASAP7_75t_L g565 ( .A1(n_67), .A2(n_194), .B1(n_566), .B2(n_567), .Y(n_565) );
INVx1_ASAP7_75t_L g823 ( .A(n_68), .Y(n_823) );
CKINVDCx20_ASAP7_75t_R g938 ( .A(n_69), .Y(n_938) );
CKINVDCx20_ASAP7_75t_R g994 ( .A(n_70), .Y(n_994) );
AOI22xp33_ASAP7_75t_L g930 ( .A1(n_71), .A2(n_119), .B1(n_646), .B2(n_770), .Y(n_930) );
AO22x2_ASAP7_75t_L g381 ( .A1(n_72), .A2(n_229), .B1(n_372), .B2(n_373), .Y(n_381) );
INVx1_ASAP7_75t_L g1038 ( .A(n_72), .Y(n_1038) );
CKINVDCx20_ASAP7_75t_R g1013 ( .A(n_73), .Y(n_1013) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_74), .A2(n_75), .B1(n_553), .B2(n_554), .Y(n_552) );
CKINVDCx20_ASAP7_75t_R g725 ( .A(n_76), .Y(n_725) );
AOI22xp5_ASAP7_75t_L g830 ( .A1(n_77), .A2(n_93), .B1(n_547), .B2(n_653), .Y(n_830) );
AOI22xp5_ASAP7_75t_L g746 ( .A1(n_78), .A2(n_210), .B1(n_423), .B2(n_642), .Y(n_746) );
OA22x2_ASAP7_75t_L g701 ( .A1(n_79), .A2(n_702), .B1(n_703), .B2(n_704), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_79), .Y(n_702) );
OA22x2_ASAP7_75t_L g1073 ( .A1(n_80), .A2(n_1074), .B1(n_1075), .B2(n_1090), .Y(n_1073) );
INVx1_ASAP7_75t_L g1074 ( .A(n_80), .Y(n_1074) );
AOI22xp33_ASAP7_75t_L g437 ( .A1(n_81), .A2(n_134), .B1(n_438), .B2(n_444), .Y(n_437) );
CKINVDCx20_ASAP7_75t_R g489 ( .A(n_83), .Y(n_489) );
INVx1_ASAP7_75t_L g813 ( .A(n_85), .Y(n_813) );
AOI221xp5_ASAP7_75t_L g888 ( .A1(n_86), .A2(n_307), .B1(n_889), .B2(n_890), .C(n_891), .Y(n_888) );
AOI22xp33_ASAP7_75t_L g766 ( .A1(n_87), .A2(n_128), .B1(n_403), .B2(n_420), .Y(n_766) );
CKINVDCx20_ASAP7_75t_R g539 ( .A(n_88), .Y(n_539) );
CKINVDCx20_ASAP7_75t_R g530 ( .A(n_89), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g965 ( .A1(n_91), .A2(n_168), .B1(n_649), .B2(n_716), .Y(n_965) );
AOI22xp33_ASAP7_75t_SL g773 ( .A1(n_92), .A2(n_334), .B1(n_774), .B2(n_775), .Y(n_773) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_94), .A2(n_135), .B1(n_460), .B2(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g1042 ( .A(n_95), .Y(n_1042) );
AOI22xp33_ASAP7_75t_SL g768 ( .A1(n_96), .A2(n_153), .B1(n_536), .B2(n_716), .Y(n_768) );
CKINVDCx20_ASAP7_75t_R g924 ( .A(n_97), .Y(n_924) );
CKINVDCx20_ASAP7_75t_R g834 ( .A(n_98), .Y(n_834) );
CKINVDCx20_ASAP7_75t_R g493 ( .A(n_99), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_101), .A2(n_200), .B1(n_513), .B2(n_658), .Y(n_691) );
CKINVDCx20_ASAP7_75t_R g871 ( .A(n_102), .Y(n_871) );
CKINVDCx20_ASAP7_75t_R g745 ( .A(n_103), .Y(n_745) );
CKINVDCx20_ASAP7_75t_R g844 ( .A(n_104), .Y(n_844) );
CKINVDCx20_ASAP7_75t_R g988 ( .A(n_105), .Y(n_988) );
AOI22xp33_ASAP7_75t_L g654 ( .A1(n_106), .A2(n_266), .B1(n_464), .B2(n_551), .Y(n_654) );
CKINVDCx20_ASAP7_75t_R g995 ( .A(n_107), .Y(n_995) );
AOI22xp33_ASAP7_75t_L g427 ( .A1(n_108), .A2(n_288), .B1(n_428), .B2(n_433), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g685 ( .A1(n_109), .A2(n_120), .B1(n_686), .B2(n_687), .Y(n_685) );
AOI22xp5_ASAP7_75t_L g753 ( .A1(n_111), .A2(n_284), .B1(n_436), .B2(n_504), .Y(n_753) );
CKINVDCx20_ASAP7_75t_R g480 ( .A(n_112), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_113), .B(n_391), .Y(n_390) );
AOI22xp33_ASAP7_75t_SL g1018 ( .A1(n_114), .A2(n_163), .B1(n_536), .B2(n_648), .Y(n_1018) );
AOI22xp33_ASAP7_75t_SL g1021 ( .A1(n_115), .A2(n_279), .B1(n_517), .B2(n_553), .Y(n_1021) );
AOI22xp33_ASAP7_75t_L g1084 ( .A1(n_117), .A2(n_311), .B1(n_755), .B2(n_1085), .Y(n_1084) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_118), .A2(n_310), .B1(n_423), .B2(n_536), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g942 ( .A1(n_121), .A2(n_289), .B1(n_398), .B2(n_413), .Y(n_942) );
AOI22xp33_ASAP7_75t_SL g852 ( .A1(n_122), .A2(n_303), .B1(n_642), .B2(n_649), .Y(n_852) );
AOI22xp33_ASAP7_75t_L g958 ( .A1(n_123), .A2(n_308), .B1(n_782), .B2(n_959), .Y(n_958) );
AOI22xp33_ASAP7_75t_L g985 ( .A1(n_124), .A2(n_287), .B1(n_579), .B2(n_986), .Y(n_985) );
AOI22xp33_ASAP7_75t_L g948 ( .A1(n_125), .A2(n_179), .B1(n_580), .B2(n_859), .Y(n_948) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_126), .A2(n_185), .B1(n_587), .B2(n_588), .Y(n_586) );
CKINVDCx20_ASAP7_75t_R g833 ( .A(n_127), .Y(n_833) );
NAND2xp5_ASAP7_75t_L g847 ( .A(n_129), .B(n_848), .Y(n_847) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_130), .A2(n_183), .B1(n_507), .B2(n_509), .Y(n_506) );
CKINVDCx20_ASAP7_75t_R g365 ( .A(n_131), .Y(n_365) );
AOI22xp33_ASAP7_75t_L g1088 ( .A1(n_132), .A2(n_249), .B1(n_398), .B2(n_406), .Y(n_1088) );
AND2x6_ASAP7_75t_L g353 ( .A(n_133), .B(n_354), .Y(n_353) );
HB1xp67_ASAP7_75t_L g1035 ( .A(n_133), .Y(n_1035) );
AOI22xp33_ASAP7_75t_L g683 ( .A1(n_136), .A2(n_216), .B1(n_616), .B2(n_684), .Y(n_683) );
AOI22xp33_ASAP7_75t_SL g927 ( .A1(n_137), .A2(n_253), .B1(n_403), .B2(n_928), .Y(n_927) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_138), .A2(n_161), .B1(n_514), .B2(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g679 ( .A(n_139), .Y(n_679) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_140), .A2(n_238), .B1(n_547), .B2(n_548), .Y(n_546) );
CKINVDCx20_ASAP7_75t_R g1050 ( .A(n_142), .Y(n_1050) );
AOI22xp5_ASAP7_75t_L g720 ( .A1(n_143), .A2(n_236), .B1(n_452), .B2(n_721), .Y(n_720) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_145), .A2(n_169), .B1(n_579), .B2(n_580), .Y(n_578) );
AOI22xp5_ASAP7_75t_SL g590 ( .A1(n_147), .A2(n_591), .B1(n_630), .B2(n_631), .Y(n_590) );
INVx1_ASAP7_75t_L g631 ( .A(n_147), .Y(n_631) );
AOI22xp33_ASAP7_75t_SL g845 ( .A1(n_148), .A2(n_256), .B1(n_422), .B2(n_575), .Y(n_845) );
CKINVDCx20_ASAP7_75t_R g946 ( .A(n_149), .Y(n_946) );
AOI22xp5_ASAP7_75t_L g828 ( .A1(n_150), .A2(n_283), .B1(n_514), .B2(n_588), .Y(n_828) );
NAND2xp5_ASAP7_75t_SL g1017 ( .A(n_151), .B(n_889), .Y(n_1017) );
INVx1_ASAP7_75t_L g594 ( .A(n_152), .Y(n_594) );
AO22x2_ASAP7_75t_L g379 ( .A1(n_154), .A2(n_219), .B1(n_372), .B2(n_376), .Y(n_379) );
NOR2xp33_ASAP7_75t_L g1039 ( .A(n_154), .B(n_1040), .Y(n_1039) );
CKINVDCx20_ASAP7_75t_R g1001 ( .A(n_155), .Y(n_1001) );
AOI22xp33_ASAP7_75t_SL g1024 ( .A1(n_156), .A2(n_234), .B1(n_727), .B2(n_779), .Y(n_1024) );
CKINVDCx20_ASAP7_75t_R g461 ( .A(n_157), .Y(n_461) );
AOI211xp5_ASAP7_75t_L g367 ( .A1(n_158), .A2(n_368), .B(n_382), .C(n_409), .Y(n_367) );
CKINVDCx20_ASAP7_75t_R g881 ( .A(n_159), .Y(n_881) );
AOI22xp5_ASAP7_75t_L g950 ( .A1(n_160), .A2(n_331), .B1(n_951), .B2(n_952), .Y(n_950) );
AOI22xp33_ASAP7_75t_SL g1014 ( .A1(n_162), .A2(n_244), .B1(n_566), .B2(n_642), .Y(n_1014) );
CKINVDCx20_ASAP7_75t_R g640 ( .A(n_164), .Y(n_640) );
CKINVDCx20_ASAP7_75t_R g1052 ( .A(n_165), .Y(n_1052) );
CKINVDCx20_ASAP7_75t_R g1054 ( .A(n_166), .Y(n_1054) );
CKINVDCx20_ASAP7_75t_R g418 ( .A(n_167), .Y(n_418) );
CKINVDCx20_ASAP7_75t_R g742 ( .A(n_170), .Y(n_742) );
AOI22xp33_ASAP7_75t_SL g652 ( .A1(n_171), .A2(n_207), .B1(n_434), .B2(n_653), .Y(n_652) );
AOI22xp33_ASAP7_75t_SL g1023 ( .A1(n_172), .A2(n_182), .B1(n_653), .B2(n_686), .Y(n_1023) );
AOI22xp5_ASAP7_75t_L g831 ( .A1(n_173), .A2(n_212), .B1(n_553), .B2(n_755), .Y(n_831) );
AOI22xp33_ASAP7_75t_L g769 ( .A1(n_174), .A2(n_208), .B1(n_646), .B2(n_770), .Y(n_769) );
AOI22xp33_ASAP7_75t_SL g781 ( .A1(n_175), .A2(n_336), .B1(n_721), .B2(n_782), .Y(n_781) );
INVx1_ASAP7_75t_L g765 ( .A(n_176), .Y(n_765) );
AOI22xp33_ASAP7_75t_L g800 ( .A1(n_177), .A2(n_295), .B1(n_513), .B2(n_801), .Y(n_800) );
CKINVDCx20_ASAP7_75t_R g495 ( .A(n_178), .Y(n_495) );
CKINVDCx20_ASAP7_75t_R g971 ( .A(n_180), .Y(n_971) );
AOI22xp33_ASAP7_75t_L g961 ( .A1(n_181), .A2(n_341), .B1(n_553), .B2(n_723), .Y(n_961) );
AOI22xp33_ASAP7_75t_L g722 ( .A1(n_184), .A2(n_269), .B1(n_623), .B2(n_723), .Y(n_722) );
AOI22xp33_ASAP7_75t_SL g656 ( .A1(n_186), .A2(n_278), .B1(n_440), .B2(n_452), .Y(n_656) );
AOI22xp33_ASAP7_75t_SL g1020 ( .A1(n_187), .A2(n_329), .B1(n_512), .B2(n_959), .Y(n_1020) );
CKINVDCx20_ASAP7_75t_R g963 ( .A(n_188), .Y(n_963) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_189), .B(n_674), .Y(n_809) );
CKINVDCx20_ASAP7_75t_R g483 ( .A(n_190), .Y(n_483) );
AOI22xp33_ASAP7_75t_SL g855 ( .A1(n_191), .A2(n_233), .B1(n_504), .B2(n_551), .Y(n_855) );
CKINVDCx20_ASAP7_75t_R g805 ( .A(n_192), .Y(n_805) );
CKINVDCx20_ASAP7_75t_R g984 ( .A(n_193), .Y(n_984) );
CKINVDCx20_ASAP7_75t_R g668 ( .A(n_195), .Y(n_668) );
AOI22xp33_ASAP7_75t_L g1056 ( .A1(n_196), .A2(n_203), .B1(n_566), .B2(n_1057), .Y(n_1056) );
AOI22xp33_ASAP7_75t_L g953 ( .A1(n_197), .A2(n_309), .B1(n_436), .B2(n_778), .Y(n_953) );
CKINVDCx20_ASAP7_75t_R g882 ( .A(n_199), .Y(n_882) );
AOI22xp33_ASAP7_75t_L g796 ( .A1(n_201), .A2(n_232), .B1(n_554), .B2(n_686), .Y(n_796) );
CKINVDCx20_ASAP7_75t_R g892 ( .A(n_202), .Y(n_892) );
CKINVDCx20_ASAP7_75t_R g945 ( .A(n_205), .Y(n_945) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_206), .A2(n_323), .B1(n_622), .B2(n_623), .Y(n_621) );
AOI22xp33_ASAP7_75t_L g783 ( .A1(n_209), .A2(n_302), .B1(n_553), .B2(n_723), .Y(n_783) );
AOI22xp33_ASAP7_75t_L g624 ( .A1(n_211), .A2(n_250), .B1(n_625), .B2(n_628), .Y(n_624) );
OA22x2_ASAP7_75t_L g523 ( .A1(n_213), .A2(n_524), .B1(n_525), .B2(n_555), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_213), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g1016 ( .A(n_214), .B(n_890), .Y(n_1016) );
XNOR2x2_ASAP7_75t_L g905 ( .A(n_215), .B(n_906), .Y(n_905) );
AND2x2_ASAP7_75t_L g357 ( .A(n_217), .B(n_358), .Y(n_357) );
AOI22xp5_ASAP7_75t_L g790 ( .A1(n_218), .A2(n_791), .B1(n_815), .B2(n_816), .Y(n_790) );
INVx1_ASAP7_75t_L g815 ( .A(n_218), .Y(n_815) );
AOI22xp5_ASAP7_75t_L g1068 ( .A1(n_220), .A2(n_231), .B1(n_502), .B2(n_951), .Y(n_1068) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_222), .B(n_646), .Y(n_645) );
AOI22xp33_ASAP7_75t_SL g860 ( .A1(n_224), .A2(n_347), .B1(n_460), .B2(n_755), .Y(n_860) );
CKINVDCx20_ASAP7_75t_R g914 ( .A(n_226), .Y(n_914) );
AOI22xp33_ASAP7_75t_SL g858 ( .A1(n_227), .A2(n_343), .B1(n_827), .B2(n_859), .Y(n_858) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_230), .A2(n_324), .B1(n_399), .B2(n_575), .Y(n_574) );
CKINVDCx20_ASAP7_75t_R g676 ( .A(n_237), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g1080 ( .A1(n_239), .A2(n_349), .B1(n_912), .B2(n_1081), .Y(n_1080) );
AOI22xp33_ASAP7_75t_L g689 ( .A1(n_240), .A2(n_281), .B1(n_452), .B2(n_690), .Y(n_689) );
CKINVDCx20_ASAP7_75t_R g708 ( .A(n_241), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_242), .B(n_570), .Y(n_569) );
AOI22xp5_ASAP7_75t_L g865 ( .A1(n_243), .A2(n_866), .B1(n_897), .B2(n_898), .Y(n_865) );
CKINVDCx20_ASAP7_75t_R g897 ( .A(n_243), .Y(n_897) );
AOI22xp33_ASAP7_75t_L g1064 ( .A1(n_245), .A2(n_344), .B1(n_509), .B2(n_727), .Y(n_1064) );
CKINVDCx20_ASAP7_75t_R g733 ( .A(n_246), .Y(n_733) );
AOI22xp33_ASAP7_75t_L g1087 ( .A1(n_247), .A2(n_290), .B1(n_889), .B2(n_890), .Y(n_1087) );
CKINVDCx20_ASAP7_75t_R g528 ( .A(n_248), .Y(n_528) );
INVx1_ASAP7_75t_L g603 ( .A(n_254), .Y(n_603) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_255), .A2(n_280), .B1(n_516), .B2(n_517), .Y(n_515) );
INVx1_ASAP7_75t_L g609 ( .A(n_258), .Y(n_609) );
INVx1_ASAP7_75t_L g372 ( .A(n_259), .Y(n_372) );
INVx1_ASAP7_75t_L g374 ( .A(n_259), .Y(n_374) );
AOI22xp33_ASAP7_75t_L g1069 ( .A1(n_260), .A2(n_342), .B1(n_504), .B2(n_547), .Y(n_1069) );
CKINVDCx20_ASAP7_75t_R g717 ( .A(n_261), .Y(n_717) );
CKINVDCx20_ASAP7_75t_R g748 ( .A(n_263), .Y(n_748) );
CKINVDCx20_ASAP7_75t_R g1004 ( .A(n_264), .Y(n_1004) );
AOI22xp5_ASAP7_75t_L g1044 ( .A1(n_265), .A2(n_1045), .B1(n_1046), .B2(n_1070), .Y(n_1044) );
CKINVDCx20_ASAP7_75t_R g1070 ( .A(n_265), .Y(n_1070) );
CKINVDCx20_ASAP7_75t_R g458 ( .A(n_268), .Y(n_458) );
CKINVDCx20_ASAP7_75t_R g666 ( .A(n_273), .Y(n_666) );
CKINVDCx20_ASAP7_75t_R g886 ( .A(n_274), .Y(n_886) );
CKINVDCx20_ASAP7_75t_R g519 ( .A(n_275), .Y(n_519) );
CKINVDCx20_ASAP7_75t_R g997 ( .A(n_276), .Y(n_997) );
INVx1_ASAP7_75t_L g804 ( .A(n_277), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g964 ( .A(n_282), .B(n_570), .Y(n_964) );
CKINVDCx20_ASAP7_75t_R g707 ( .A(n_285), .Y(n_707) );
AOI22xp33_ASAP7_75t_SL g584 ( .A1(n_286), .A2(n_338), .B1(n_450), .B2(n_585), .Y(n_584) );
AOI22xp33_ASAP7_75t_L g754 ( .A1(n_292), .A2(n_328), .B1(n_551), .B2(n_755), .Y(n_754) );
AOI22xp33_ASAP7_75t_L g835 ( .A1(n_294), .A2(n_315), .B1(n_399), .B2(n_405), .Y(n_835) );
INVx1_ASAP7_75t_L g358 ( .A(n_296), .Y(n_358) );
CKINVDCx20_ASAP7_75t_R g670 ( .A(n_298), .Y(n_670) );
CKINVDCx20_ASAP7_75t_R g1025 ( .A(n_299), .Y(n_1025) );
INVx1_ASAP7_75t_L g354 ( .A(n_300), .Y(n_354) );
CKINVDCx20_ASAP7_75t_R g920 ( .A(n_301), .Y(n_920) );
OA22x2_ASAP7_75t_L g839 ( .A1(n_304), .A2(n_840), .B1(n_841), .B2(n_861), .Y(n_839) );
INVx1_ASAP7_75t_L g840 ( .A(n_304), .Y(n_840) );
AOI22xp33_ASAP7_75t_L g615 ( .A1(n_305), .A2(n_335), .B1(n_554), .B2(n_616), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g850 ( .A(n_306), .B(n_851), .Y(n_850) );
CKINVDCx20_ASAP7_75t_R g941 ( .A(n_312), .Y(n_941) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_313), .B(n_607), .Y(n_606) );
CKINVDCx20_ASAP7_75t_R g921 ( .A(n_314), .Y(n_921) );
CKINVDCx20_ASAP7_75t_R g981 ( .A(n_318), .Y(n_981) );
CKINVDCx20_ASAP7_75t_R g410 ( .A(n_319), .Y(n_410) );
CKINVDCx20_ASAP7_75t_R g564 ( .A(n_321), .Y(n_564) );
CKINVDCx20_ASAP7_75t_R g672 ( .A(n_322), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_325), .B(n_403), .Y(n_481) );
INVx1_ASAP7_75t_L g597 ( .A(n_326), .Y(n_597) );
CKINVDCx20_ASAP7_75t_R g1059 ( .A(n_327), .Y(n_1059) );
CKINVDCx20_ASAP7_75t_R g710 ( .A(n_330), .Y(n_710) );
CKINVDCx20_ASAP7_75t_R g989 ( .A(n_333), .Y(n_989) );
CKINVDCx20_ASAP7_75t_R g874 ( .A(n_337), .Y(n_874) );
INVx1_ASAP7_75t_L g759 ( .A(n_339), .Y(n_759) );
CKINVDCx20_ASAP7_75t_R g589 ( .A(n_340), .Y(n_589) );
OA22x2_ASAP7_75t_SL g661 ( .A1(n_346), .A2(n_662), .B1(n_663), .B2(n_692), .Y(n_661) );
INVx1_ASAP7_75t_L g692 ( .A(n_346), .Y(n_692) );
INVx1_ASAP7_75t_L g610 ( .A(n_348), .Y(n_610) );
INVx1_ASAP7_75t_SL g351 ( .A(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_353), .B(n_355), .Y(n_352) );
HB1xp67_ASAP7_75t_L g1034 ( .A(n_354), .Y(n_1034) );
OAI21xp5_ASAP7_75t_L g1095 ( .A1(n_355), .A2(n_1033), .B(n_1096), .Y(n_1095) );
CKINVDCx20_ASAP7_75t_R g355 ( .A(n_356), .Y(n_355) );
INVxp67_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AOI221xp5_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_903), .B1(n_1028), .B2(n_1029), .C(n_1030), .Y(n_359) );
INVx1_ASAP7_75t_L g1028 ( .A(n_360), .Y(n_1028) );
AOI22xp5_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_696), .B1(n_901), .B2(n_902), .Y(n_360) );
INVx1_ASAP7_75t_L g901 ( .A(n_361), .Y(n_901) );
AOI22xp5_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_556), .B1(n_694), .B2(n_695), .Y(n_361) );
INVx1_ASAP7_75t_L g694 ( .A(n_362), .Y(n_694) );
AOI22xp5_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_364), .B1(n_467), .B2(n_468), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
XNOR2x1_ASAP7_75t_L g364 ( .A(n_365), .B(n_366), .Y(n_364) );
AND2x2_ASAP7_75t_L g366 ( .A(n_367), .B(n_425), .Y(n_366) );
INVx3_ASAP7_75t_L g711 ( .A(n_368), .Y(n_711) );
BUFx3_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
BUFx6f_ASAP7_75t_L g476 ( .A(n_369), .Y(n_476) );
INVx4_ASAP7_75t_L g602 ( .A(n_369), .Y(n_602) );
INVx2_ASAP7_75t_L g639 ( .A(n_369), .Y(n_639) );
INVx2_ASAP7_75t_L g1012 ( .A(n_369), .Y(n_1012) );
AND2x6_ASAP7_75t_L g369 ( .A(n_370), .B(n_377), .Y(n_369) );
AND2x4_ASAP7_75t_L g406 ( .A(n_370), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g541 ( .A(n_370), .Y(n_541) );
AND2x2_ASAP7_75t_L g370 ( .A(n_371), .B(n_375), .Y(n_370) );
INVx2_ASAP7_75t_L g388 ( .A(n_371), .Y(n_388) );
AND2x2_ASAP7_75t_L g402 ( .A(n_371), .B(n_379), .Y(n_402) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g376 ( .A(n_374), .Y(n_376) );
AND2x2_ASAP7_75t_L g387 ( .A(n_375), .B(n_388), .Y(n_387) );
OR2x2_ASAP7_75t_L g396 ( .A(n_375), .B(n_388), .Y(n_396) );
INVx1_ASAP7_75t_L g401 ( .A(n_375), .Y(n_401) );
INVx2_ASAP7_75t_L g417 ( .A(n_375), .Y(n_417) );
AND2x2_ASAP7_75t_L g431 ( .A(n_377), .B(n_432), .Y(n_431) );
AND2x6_ASAP7_75t_L g436 ( .A(n_377), .B(n_395), .Y(n_436) );
AND2x4_ASAP7_75t_L g452 ( .A(n_377), .B(n_387), .Y(n_452) );
AND2x2_ASAP7_75t_L g377 ( .A(n_378), .B(n_380), .Y(n_377) );
AND2x2_ASAP7_75t_L g389 ( .A(n_378), .B(n_381), .Y(n_389) );
INVx2_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
AND2x2_ASAP7_75t_L g443 ( .A(n_379), .B(n_408), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_379), .B(n_381), .Y(n_446) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g408 ( .A(n_381), .Y(n_408) );
INVx1_ASAP7_75t_L g416 ( .A(n_381), .Y(n_416) );
OAI211xp5_ASAP7_75t_L g382 ( .A1(n_383), .A2(n_384), .B(n_390), .C(n_397), .Y(n_382) );
BUFx3_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx2_ASAP7_75t_L g491 ( .A(n_385), .Y(n_491) );
OAI22xp5_ASAP7_75t_L g803 ( .A1(n_385), .A2(n_486), .B1(n_804), .B2(n_805), .Y(n_803) );
OAI221xp5_ASAP7_75t_L g832 ( .A1(n_385), .A2(n_487), .B1(n_833), .B2(n_834), .C(n_835), .Y(n_832) );
BUFx3_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g532 ( .A(n_386), .Y(n_532) );
NAND2x1p5_ASAP7_75t_L g386 ( .A(n_387), .B(n_389), .Y(n_386) );
AND2x2_ASAP7_75t_L g442 ( .A(n_387), .B(n_443), .Y(n_442) );
AND2x6_ASAP7_75t_L g573 ( .A(n_387), .B(n_389), .Y(n_573) );
NAND2xp5_ASAP7_75t_SL g876 ( .A(n_387), .B(n_443), .Y(n_876) );
AND2x2_ASAP7_75t_L g432 ( .A(n_388), .B(n_417), .Y(n_432) );
AND2x4_ASAP7_75t_L g394 ( .A(n_389), .B(n_395), .Y(n_394) );
AND2x4_ASAP7_75t_L g460 ( .A(n_389), .B(n_432), .Y(n_460) );
INVx1_ASAP7_75t_L g488 ( .A(n_389), .Y(n_488) );
BUFx2_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx2_ASAP7_75t_L g570 ( .A(n_393), .Y(n_570) );
INVx2_ASAP7_75t_L g770 ( .A(n_393), .Y(n_770) );
INVx5_ASAP7_75t_L g851 ( .A(n_393), .Y(n_851) );
INVx4_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
OR2x2_ASAP7_75t_L g487 ( .A(n_396), .B(n_488), .Y(n_487) );
BUFx2_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
BUFx2_ASAP7_75t_L g536 ( .A(n_399), .Y(n_536) );
BUFx3_ASAP7_75t_L g649 ( .A(n_399), .Y(n_649) );
INVx1_ASAP7_75t_L g929 ( .A(n_399), .Y(n_929) );
AND2x4_ASAP7_75t_L g399 ( .A(n_400), .B(n_402), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
OR2x6_ASAP7_75t_L g445 ( .A(n_401), .B(n_446), .Y(n_445) );
AND2x4_ASAP7_75t_L g414 ( .A(n_402), .B(n_415), .Y(n_414) );
AND2x4_ASAP7_75t_L g423 ( .A(n_402), .B(n_424), .Y(n_423) );
NAND2x1p5_ASAP7_75t_L g497 ( .A(n_402), .B(n_498), .Y(n_497) );
INVx2_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_SL g404 ( .A(n_405), .Y(n_404) );
BUFx6f_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
BUFx2_ASAP7_75t_SL g567 ( .A(n_406), .Y(n_567) );
BUFx2_ASAP7_75t_SL g642 ( .A(n_406), .Y(n_642) );
INVx1_ASAP7_75t_L g542 ( .A(n_407), .Y(n_542) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
OAI22xp5_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_411), .B1(n_418), .B2(n_419), .Y(n_409) );
OAI222xp33_ASAP7_75t_L g996 ( .A1(n_411), .A2(n_997), .B1(n_998), .B2(n_999), .C1(n_1000), .C2(n_1001), .Y(n_996) );
INVx2_ASAP7_75t_SL g411 ( .A(n_412), .Y(n_411) );
INVx2_ASAP7_75t_SL g749 ( .A(n_412), .Y(n_749) );
BUFx6f_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g494 ( .A(n_413), .Y(n_494) );
BUFx6f_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
BUFx2_ASAP7_75t_L g548 ( .A(n_414), .Y(n_548) );
BUFx4f_ASAP7_75t_SL g575 ( .A(n_414), .Y(n_575) );
BUFx6f_ASAP7_75t_L g648 ( .A(n_414), .Y(n_648) );
BUFx6f_ASAP7_75t_L g716 ( .A(n_414), .Y(n_716) );
AND2x2_ASAP7_75t_L g415 ( .A(n_416), .B(n_417), .Y(n_415) );
INVx1_ASAP7_75t_L g424 ( .A(n_416), .Y(n_424) );
INVx1_ASAP7_75t_L g498 ( .A(n_417), .Y(n_498) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx3_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
BUFx4f_ASAP7_75t_SL g970 ( .A(n_422), .Y(n_970) );
BUFx12f_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
BUFx6f_ASAP7_75t_L g479 ( .A(n_423), .Y(n_479) );
BUFx6f_ASAP7_75t_L g566 ( .A(n_423), .Y(n_566) );
NOR3xp33_ASAP7_75t_L g425 ( .A(n_426), .B(n_447), .C(n_457), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_427), .B(n_437), .Y(n_426) );
INVx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
OAI221xp5_ASAP7_75t_SL g980 ( .A1(n_429), .A2(n_981), .B1(n_982), .B2(n_984), .C(n_985), .Y(n_980) );
INVx3_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
BUFx3_ASAP7_75t_L g616 ( .A(n_430), .Y(n_616) );
BUFx3_ASAP7_75t_L g795 ( .A(n_430), .Y(n_795) );
BUFx6f_ASAP7_75t_L g910 ( .A(n_430), .Y(n_910) );
BUFx6f_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g508 ( .A(n_431), .Y(n_508) );
BUFx2_ASAP7_75t_SL g727 ( .A(n_431), .Y(n_727) );
BUFx2_ASAP7_75t_SL g778 ( .A(n_431), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_432), .B(n_443), .Y(n_456) );
AND2x4_ASAP7_75t_L g465 ( .A(n_432), .B(n_466), .Y(n_465) );
AND2x2_ASAP7_75t_L g505 ( .A(n_432), .B(n_443), .Y(n_505) );
INVx1_ASAP7_75t_L g885 ( .A(n_433), .Y(n_885) );
HB1xp67_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g915 ( .A(n_434), .Y(n_915) );
INVx5_ASAP7_75t_SL g434 ( .A(n_435), .Y(n_434) );
INVx4_ASAP7_75t_L g579 ( .A(n_435), .Y(n_579) );
INVx2_ASAP7_75t_L g622 ( .A(n_435), .Y(n_622) );
INVx1_ASAP7_75t_L g732 ( .A(n_435), .Y(n_732) );
INVx11_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx11_ASAP7_75t_L g503 ( .A(n_436), .Y(n_503) );
INVx3_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
BUFx6f_ASAP7_75t_L g618 ( .A(n_440), .Y(n_618) );
BUFx2_ASAP7_75t_L g1081 ( .A(n_440), .Y(n_1081) );
INVx4_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx5_ASAP7_75t_L g514 ( .A(n_441), .Y(n_514) );
INVx3_ASAP7_75t_L g585 ( .A(n_441), .Y(n_585) );
INVx1_ASAP7_75t_L g721 ( .A(n_441), .Y(n_721) );
BUFx3_ASAP7_75t_L g960 ( .A(n_441), .Y(n_960) );
INVx8_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_SL g444 ( .A(n_445), .Y(n_444) );
INVx6_ASAP7_75t_SL g518 ( .A(n_445), .Y(n_518) );
OAI22xp5_ASAP7_75t_L g537 ( .A1(n_445), .A2(n_538), .B1(n_539), .B2(n_540), .Y(n_537) );
INVx1_ASAP7_75t_SL g658 ( .A(n_445), .Y(n_658) );
INVx1_ASAP7_75t_L g1066 ( .A(n_445), .Y(n_1066) );
INVx1_ASAP7_75t_L g466 ( .A(n_446), .Y(n_466) );
OAI22xp5_ASAP7_75t_L g447 ( .A1(n_448), .A2(n_449), .B1(n_453), .B2(n_454), .Y(n_447) );
OAI22xp5_ASAP7_75t_L g880 ( .A1(n_449), .A2(n_454), .B1(n_881), .B2(n_882), .Y(n_880) );
INVxp67_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx2_ASAP7_75t_L g512 ( .A(n_451), .Y(n_512) );
INVx2_ASAP7_75t_L g782 ( .A(n_451), .Y(n_782) );
INVx3_ASAP7_75t_L g859 ( .A(n_451), .Y(n_859) );
OAI22xp5_ASAP7_75t_L g919 ( .A1(n_451), .A2(n_735), .B1(n_920), .B2(n_921), .Y(n_919) );
INVx6_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
BUFx3_ASAP7_75t_L g547 ( .A(n_452), .Y(n_547) );
BUFx3_ASAP7_75t_L g627 ( .A(n_452), .Y(n_627) );
BUFx3_ASAP7_75t_L g799 ( .A(n_452), .Y(n_799) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g735 ( .A(n_455), .Y(n_735) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
OAI22xp5_ASAP7_75t_L g457 ( .A1(n_458), .A2(n_459), .B1(n_461), .B2(n_462), .Y(n_457) );
INVx2_ASAP7_75t_L g587 ( .A(n_459), .Y(n_587) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
BUFx3_ASAP7_75t_L g516 ( .A(n_460), .Y(n_516) );
BUFx3_ASAP7_75t_L g553 ( .A(n_460), .Y(n_553) );
BUFx3_ASAP7_75t_L g623 ( .A(n_460), .Y(n_623) );
BUFx6f_ASAP7_75t_L g918 ( .A(n_460), .Y(n_918) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
BUFx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
BUFx3_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
BUFx2_ASAP7_75t_SL g509 ( .A(n_465), .Y(n_509) );
BUFx3_ASAP7_75t_L g554 ( .A(n_465), .Y(n_554) );
BUFx3_ASAP7_75t_L g582 ( .A(n_465), .Y(n_582) );
BUFx3_ASAP7_75t_L g687 ( .A(n_465), .Y(n_687) );
BUFx2_ASAP7_75t_L g755 ( .A(n_465), .Y(n_755) );
BUFx2_ASAP7_75t_SL g779 ( .A(n_465), .Y(n_779) );
AND2x2_ASAP7_75t_L g588 ( .A(n_466), .B(n_498), .Y(n_588) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
OAI22xp5_ASAP7_75t_L g468 ( .A1(n_469), .A2(n_470), .B1(n_520), .B2(n_521), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
XOR2x2_ASAP7_75t_L g471 ( .A(n_472), .B(n_519), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_473), .B(n_499), .Y(n_472) );
NOR3xp33_ASAP7_75t_L g473 ( .A(n_474), .B(n_482), .C(n_492), .Y(n_473) );
OAI221xp5_ASAP7_75t_L g474 ( .A1(n_475), .A2(n_477), .B1(n_478), .B2(n_480), .C(n_481), .Y(n_474) );
OAI21xp5_ASAP7_75t_L g563 ( .A1(n_475), .A2(n_564), .B(n_565), .Y(n_563) );
INVx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx2_ASAP7_75t_SL g998 ( .A(n_476), .Y(n_998) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
BUFx4f_ASAP7_75t_L g607 ( .A(n_479), .Y(n_607) );
OAI22xp5_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_484), .B1(n_489), .B2(n_490), .Y(n_482) );
OAI22xp5_ASAP7_75t_L g936 ( .A1(n_484), .A2(n_937), .B1(n_938), .B2(n_939), .Y(n_936) );
OAI22xp5_ASAP7_75t_L g993 ( .A1(n_484), .A2(n_490), .B1(n_994), .B2(n_995), .Y(n_993) );
INVx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
BUFx6f_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
BUFx3_ASAP7_75t_L g529 ( .A(n_487), .Y(n_529) );
INVx2_ASAP7_75t_L g596 ( .A(n_487), .Y(n_596) );
OAI22xp5_ASAP7_75t_L g665 ( .A1(n_490), .A2(n_666), .B1(n_667), .B2(n_668), .Y(n_665) );
OAI22xp5_ASAP7_75t_SL g706 ( .A1(n_490), .A2(n_595), .B1(n_707), .B2(n_708), .Y(n_706) );
OAI22xp5_ASAP7_75t_L g1049 ( .A1(n_490), .A2(n_1050), .B1(n_1051), .B2(n_1052), .Y(n_1049) );
INVx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
OAI22xp5_ASAP7_75t_L g492 ( .A1(n_493), .A2(n_494), .B1(n_495), .B2(n_496), .Y(n_492) );
OAI22xp33_ASAP7_75t_L g713 ( .A1(n_496), .A2(n_714), .B1(n_715), .B2(n_717), .Y(n_713) );
BUFx3_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
OAI22xp5_ASAP7_75t_L g608 ( .A1(n_497), .A2(n_609), .B1(n_610), .B2(n_611), .Y(n_608) );
INVx4_ASAP7_75t_L g678 ( .A(n_497), .Y(n_678) );
OAI22xp5_ASAP7_75t_L g747 ( .A1(n_497), .A2(n_748), .B1(n_749), .B2(n_750), .Y(n_747) );
HB1xp67_ASAP7_75t_L g812 ( .A(n_497), .Y(n_812) );
OAI22xp5_ASAP7_75t_L g891 ( .A1(n_497), .A2(n_540), .B1(n_892), .B2(n_893), .Y(n_891) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_500), .B(n_510), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_501), .B(n_506), .Y(n_500) );
INVx2_ASAP7_75t_SL g502 ( .A(n_503), .Y(n_502) );
OAI21xp33_ASAP7_75t_SL g533 ( .A1(n_503), .A2(n_534), .B(n_535), .Y(n_533) );
INVx4_ASAP7_75t_L g686 ( .A(n_503), .Y(n_686) );
INVx3_ASAP7_75t_L g774 ( .A(n_503), .Y(n_774) );
INVx4_ASAP7_75t_L g827 ( .A(n_503), .Y(n_827) );
INVx1_ASAP7_75t_L g1079 ( .A(n_504), .Y(n_1079) );
BUFx3_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
BUFx3_ASAP7_75t_L g580 ( .A(n_505), .Y(n_580) );
BUFx3_ASAP7_75t_L g653 ( .A(n_505), .Y(n_653) );
BUFx3_ASAP7_75t_L g776 ( .A(n_505), .Y(n_776) );
INVxp67_ASAP7_75t_L g870 ( .A(n_507), .Y(n_870) );
INVx3_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx3_ASAP7_75t_L g551 ( .A(n_508), .Y(n_551) );
INVx1_ASAP7_75t_SL g729 ( .A(n_509), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_511), .B(n_515), .Y(n_510) );
BUFx6f_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
BUFx2_ASAP7_75t_L g991 ( .A(n_514), .Y(n_991) );
BUFx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
BUFx2_ASAP7_75t_L g619 ( .A(n_518), .Y(n_619) );
BUFx2_ASAP7_75t_L g723 ( .A(n_518), .Y(n_723) );
BUFx4f_ASAP7_75t_SL g801 ( .A(n_518), .Y(n_801) );
BUFx2_ASAP7_75t_L g912 ( .A(n_518), .Y(n_912) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx2_ASAP7_75t_L g555 ( .A(n_525), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_526), .B(n_543), .Y(n_525) );
NOR3xp33_ASAP7_75t_L g526 ( .A(n_527), .B(n_533), .C(n_537), .Y(n_526) );
OAI22xp5_ASAP7_75t_L g527 ( .A1(n_528), .A2(n_529), .B1(n_530), .B2(n_531), .Y(n_527) );
OAI22xp5_ASAP7_75t_L g741 ( .A1(n_529), .A2(n_598), .B1(n_742), .B2(n_743), .Y(n_741) );
OA211x2_ASAP7_75t_L g962 ( .A1(n_531), .A2(n_963), .B(n_964), .C(n_965), .Y(n_962) );
INVx1_ASAP7_75t_SL g531 ( .A(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g598 ( .A(n_532), .Y(n_598) );
INVx2_ASAP7_75t_L g939 ( .A(n_532), .Y(n_939) );
CKINVDCx16_ASAP7_75t_R g612 ( .A(n_540), .Y(n_612) );
BUFx2_ASAP7_75t_L g680 ( .A(n_540), .Y(n_680) );
OR2x6_ASAP7_75t_L g540 ( .A(n_541), .B(n_542), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g543 ( .A(n_544), .B(n_549), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_545), .B(n_546), .Y(n_544) );
INVx1_ASAP7_75t_L g604 ( .A(n_548), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_550), .B(n_552), .Y(n_549) );
HB1xp67_ASAP7_75t_L g983 ( .A(n_553), .Y(n_983) );
INVx1_ASAP7_75t_L g695 ( .A(n_556), .Y(n_695) );
AOI22xp5_ASAP7_75t_L g556 ( .A1(n_557), .A2(n_632), .B1(n_633), .B2(n_693), .Y(n_556) );
INVx4_ASAP7_75t_L g693 ( .A(n_557), .Y(n_693) );
XOR2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_590), .Y(n_557) );
INVx2_ASAP7_75t_SL g558 ( .A(n_559), .Y(n_558) );
OAI22x1_ASAP7_75t_L g634 ( .A1(n_559), .A2(n_560), .B1(n_635), .B2(n_660), .Y(n_634) );
INVx3_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
XOR2x2_ASAP7_75t_L g560 ( .A(n_561), .B(n_589), .Y(n_560) );
NAND2xp5_ASAP7_75t_SL g561 ( .A(n_562), .B(n_576), .Y(n_561) );
NOR2xp33_ASAP7_75t_L g562 ( .A(n_563), .B(n_568), .Y(n_562) );
BUFx3_ASAP7_75t_L g674 ( .A(n_566), .Y(n_674) );
INVx2_ASAP7_75t_L g944 ( .A(n_566), .Y(n_944) );
NAND3xp33_ASAP7_75t_L g568 ( .A(n_569), .B(n_571), .C(n_574), .Y(n_568) );
BUFx4f_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
BUFx2_ASAP7_75t_L g646 ( .A(n_573), .Y(n_646) );
INVx1_ASAP7_75t_SL g849 ( .A(n_573), .Y(n_849) );
BUFx2_ASAP7_75t_L g890 ( .A(n_573), .Y(n_890) );
NOR2x1_ASAP7_75t_L g576 ( .A(n_577), .B(n_583), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_578), .B(n_581), .Y(n_577) );
INVx1_ASAP7_75t_L g629 ( .A(n_580), .Y(n_629) );
INVx2_ASAP7_75t_L g872 ( .A(n_582), .Y(n_872) );
HB1xp67_ASAP7_75t_L g986 ( .A(n_582), .Y(n_986) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_584), .B(n_586), .Y(n_583) );
INVx1_ASAP7_75t_SL g630 ( .A(n_591), .Y(n_630) );
AND2x2_ASAP7_75t_SL g591 ( .A(n_592), .B(n_613), .Y(n_591) );
NOR3xp33_ASAP7_75t_L g592 ( .A(n_593), .B(n_599), .C(n_608), .Y(n_592) );
OAI22xp5_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_595), .B1(n_597), .B2(n_598), .Y(n_593) );
INVx2_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVx2_ASAP7_75t_L g667 ( .A(n_596), .Y(n_667) );
INVx1_ASAP7_75t_SL g1051 ( .A(n_596), .Y(n_1051) );
OAI221xp5_ASAP7_75t_SL g599 ( .A1(n_600), .A2(n_603), .B1(n_604), .B2(n_605), .C(n_606), .Y(n_599) );
OAI221xp5_ASAP7_75t_L g669 ( .A1(n_600), .A2(n_670), .B1(n_671), .B2(n_672), .C(n_673), .Y(n_669) );
OAI21xp5_ASAP7_75t_SL g764 ( .A1(n_600), .A2(n_765), .B(n_766), .Y(n_764) );
OAI221xp5_ASAP7_75t_SL g806 ( .A1(n_600), .A2(n_604), .B1(n_807), .B2(n_808), .C(n_809), .Y(n_806) );
OAI21xp33_ASAP7_75t_SL g940 ( .A1(n_600), .A2(n_941), .B(n_942), .Y(n_940) );
INVx2_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx4_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
OAI21xp5_ASAP7_75t_SL g744 ( .A1(n_602), .A2(n_745), .B(n_746), .Y(n_744) );
BUFx2_ASAP7_75t_L g1055 ( .A(n_602), .Y(n_1055) );
OAI22xp5_ASAP7_75t_L g1058 ( .A1(n_611), .A2(n_1059), .B1(n_1060), .B2(n_1061), .Y(n_1058) );
INVx2_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx2_ASAP7_75t_L g814 ( .A(n_612), .Y(n_814) );
NOR2xp33_ASAP7_75t_L g613 ( .A(n_614), .B(n_620), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_615), .B(n_617), .Y(n_614) );
INVxp67_ASAP7_75t_L g878 ( .A(n_619), .Y(n_878) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_621), .B(n_624), .Y(n_620) );
BUFx2_ASAP7_75t_L g684 ( .A(n_623), .Y(n_684) );
INVx1_ASAP7_75t_L g887 ( .A(n_623), .Y(n_887) );
INVx2_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
OAI221xp5_ASAP7_75t_SL g987 ( .A1(n_626), .A2(n_735), .B1(n_988), .B2(n_989), .C(n_990), .Y(n_987) );
INVx3_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx2_ASAP7_75t_SL g632 ( .A(n_633), .Y(n_632) );
XNOR2x2_ASAP7_75t_L g633 ( .A(n_634), .B(n_661), .Y(n_633) );
INVx3_ASAP7_75t_L g660 ( .A(n_635), .Y(n_660) );
XOR2x2_ASAP7_75t_L g635 ( .A(n_636), .B(n_659), .Y(n_635) );
NAND2x1_ASAP7_75t_SL g636 ( .A(n_637), .B(n_650), .Y(n_636) );
NOR2xp33_ASAP7_75t_L g637 ( .A(n_638), .B(n_643), .Y(n_637) );
OAI21xp5_ASAP7_75t_SL g638 ( .A1(n_639), .A2(n_640), .B(n_641), .Y(n_638) );
OAI21xp5_ASAP7_75t_SL g923 ( .A1(n_639), .A2(n_924), .B(n_925), .Y(n_923) );
NAND3xp33_ASAP7_75t_L g643 ( .A(n_644), .B(n_645), .C(n_647), .Y(n_643) );
INVx2_ASAP7_75t_L g671 ( .A(n_648), .Y(n_671) );
INVx4_ASAP7_75t_L g896 ( .A(n_648), .Y(n_896) );
BUFx2_ASAP7_75t_L g1057 ( .A(n_648), .Y(n_1057) );
NOR2x1_ASAP7_75t_L g650 ( .A(n_651), .B(n_655), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_652), .B(n_654), .Y(n_651) );
BUFx3_ASAP7_75t_L g690 ( .A(n_653), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_656), .B(n_657), .Y(n_655) );
INVx2_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
AND2x2_ASAP7_75t_SL g663 ( .A(n_664), .B(n_681), .Y(n_663) );
NOR3xp33_ASAP7_75t_L g664 ( .A(n_665), .B(n_669), .C(n_675), .Y(n_664) );
INVx2_ASAP7_75t_L g1000 ( .A(n_674), .Y(n_1000) );
OAI22xp5_ASAP7_75t_L g675 ( .A1(n_676), .A2(n_677), .B1(n_679), .B2(n_680), .Y(n_675) );
OAI22xp5_ASAP7_75t_L g1002 ( .A1(n_677), .A2(n_814), .B1(n_1003), .B2(n_1004), .Y(n_1002) );
INVx2_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx3_ASAP7_75t_SL g1060 ( .A(n_678), .Y(n_1060) );
OAI22xp5_ASAP7_75t_SL g943 ( .A1(n_680), .A2(n_944), .B1(n_945), .B2(n_946), .Y(n_943) );
NOR2xp33_ASAP7_75t_L g681 ( .A(n_682), .B(n_688), .Y(n_681) );
NAND2xp5_ASAP7_75t_SL g682 ( .A(n_683), .B(n_685), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_689), .B(n_691), .Y(n_688) );
INVx1_ASAP7_75t_L g902 ( .A(n_696), .Y(n_902) );
AOI22xp5_ASAP7_75t_L g696 ( .A1(n_697), .A2(n_698), .B1(n_787), .B2(n_900), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
HB1xp67_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
AOI22xp5_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_701), .B1(n_736), .B2(n_786), .Y(n_699) );
INVx2_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx2_ASAP7_75t_SL g703 ( .A(n_704), .Y(n_703) );
AND2x2_ASAP7_75t_L g704 ( .A(n_705), .B(n_718), .Y(n_704) );
NOR3xp33_ASAP7_75t_L g705 ( .A(n_706), .B(n_709), .C(n_713), .Y(n_705) );
OAI21xp33_ASAP7_75t_L g709 ( .A1(n_710), .A2(n_711), .B(n_712), .Y(n_709) );
OAI21xp5_ASAP7_75t_SL g836 ( .A1(n_711), .A2(n_837), .B(n_838), .Y(n_836) );
OAI21xp5_ASAP7_75t_SL g843 ( .A1(n_711), .A2(n_844), .B(n_845), .Y(n_843) );
CKINVDCx20_ASAP7_75t_R g715 ( .A(n_716), .Y(n_715) );
NOR3xp33_ASAP7_75t_L g718 ( .A(n_719), .B(n_724), .C(n_730), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_720), .B(n_722), .Y(n_719) );
OAI22xp5_ASAP7_75t_L g724 ( .A1(n_725), .A2(n_726), .B1(n_728), .B2(n_729), .Y(n_724) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
OAI22xp5_ASAP7_75t_L g730 ( .A1(n_731), .A2(n_733), .B1(n_734), .B2(n_735), .Y(n_730) );
INVx2_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g786 ( .A(n_736), .Y(n_786) );
OA22x2_ASAP7_75t_L g736 ( .A1(n_737), .A2(n_738), .B1(n_760), .B2(n_785), .Y(n_736) );
INVx2_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
OAI22xp5_ASAP7_75t_L g788 ( .A1(n_738), .A2(n_789), .B1(n_790), .B2(n_817), .Y(n_788) );
INVx1_ASAP7_75t_L g817 ( .A(n_738), .Y(n_817) );
XOR2x2_ASAP7_75t_L g738 ( .A(n_739), .B(n_759), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_740), .B(n_751), .Y(n_739) );
NOR3xp33_ASAP7_75t_L g740 ( .A(n_741), .B(n_744), .C(n_747), .Y(n_740) );
NOR2xp33_ASAP7_75t_L g751 ( .A(n_752), .B(n_756), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_753), .B(n_754), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_757), .B(n_758), .Y(n_756) );
INVx1_ASAP7_75t_L g785 ( .A(n_760), .Y(n_785) );
INVx1_ASAP7_75t_SL g761 ( .A(n_762), .Y(n_761) );
NAND2xp5_ASAP7_75t_SL g762 ( .A(n_763), .B(n_771), .Y(n_762) );
NOR2xp33_ASAP7_75t_L g763 ( .A(n_764), .B(n_767), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_768), .B(n_769), .Y(n_767) );
NOR2xp33_ASAP7_75t_L g771 ( .A(n_772), .B(n_780), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_773), .B(n_777), .Y(n_772) );
BUFx4f_ASAP7_75t_SL g775 ( .A(n_776), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_781), .B(n_783), .Y(n_780) );
INVx1_ASAP7_75t_L g900 ( .A(n_787), .Y(n_900) );
AOI22xp33_ASAP7_75t_L g787 ( .A1(n_788), .A2(n_818), .B1(n_819), .B2(n_899), .Y(n_787) );
INVx1_ASAP7_75t_L g899 ( .A(n_788), .Y(n_899) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
INVx1_ASAP7_75t_L g816 ( .A(n_791), .Y(n_816) );
AND2x2_ASAP7_75t_SL g791 ( .A(n_792), .B(n_802), .Y(n_791) );
NOR2xp33_ASAP7_75t_L g792 ( .A(n_793), .B(n_797), .Y(n_792) );
NAND2xp33_ASAP7_75t_SL g793 ( .A(n_794), .B(n_796), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g797 ( .A(n_798), .B(n_800), .Y(n_797) );
NOR3xp33_ASAP7_75t_L g802 ( .A(n_803), .B(n_806), .C(n_810), .Y(n_802) );
OAI22xp5_ASAP7_75t_L g810 ( .A1(n_811), .A2(n_812), .B1(n_813), .B2(n_814), .Y(n_810) );
INVx1_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
OAI22xp5_ASAP7_75t_SL g819 ( .A1(n_820), .A2(n_821), .B1(n_864), .B2(n_865), .Y(n_819) );
INVx1_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
AOI22xp5_ASAP7_75t_L g821 ( .A1(n_822), .A2(n_839), .B1(n_862), .B2(n_863), .Y(n_821) );
INVx2_ASAP7_75t_SL g862 ( .A(n_822), .Y(n_862) );
XNOR2x2_ASAP7_75t_L g822 ( .A(n_823), .B(n_824), .Y(n_822) );
NOR4xp75_ASAP7_75t_L g824 ( .A(n_825), .B(n_829), .C(n_832), .D(n_836), .Y(n_824) );
NAND2xp5_ASAP7_75t_SL g825 ( .A(n_826), .B(n_828), .Y(n_825) );
NAND2xp5_ASAP7_75t_SL g829 ( .A(n_830), .B(n_831), .Y(n_829) );
INVx1_ASAP7_75t_L g863 ( .A(n_839), .Y(n_863) );
INVx1_ASAP7_75t_L g861 ( .A(n_841), .Y(n_861) );
NAND2xp5_ASAP7_75t_L g841 ( .A(n_842), .B(n_853), .Y(n_841) );
NOR2xp67_ASAP7_75t_L g842 ( .A(n_843), .B(n_846), .Y(n_842) );
NAND3xp33_ASAP7_75t_L g846 ( .A(n_847), .B(n_850), .C(n_852), .Y(n_846) );
INVx1_ASAP7_75t_SL g848 ( .A(n_849), .Y(n_848) );
BUFx6f_ASAP7_75t_L g889 ( .A(n_851), .Y(n_889) );
NOR2x1_ASAP7_75t_L g853 ( .A(n_854), .B(n_857), .Y(n_853) );
NAND2xp5_ASAP7_75t_L g854 ( .A(n_855), .B(n_856), .Y(n_854) );
NAND2xp5_ASAP7_75t_L g857 ( .A(n_858), .B(n_860), .Y(n_857) );
INVx1_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
INVx1_ASAP7_75t_L g898 ( .A(n_866), .Y(n_898) );
AND4x1_ASAP7_75t_L g866 ( .A(n_867), .B(n_879), .C(n_888), .D(n_894), .Y(n_866) );
NOR2xp33_ASAP7_75t_SL g867 ( .A(n_868), .B(n_873), .Y(n_867) );
OAI22xp5_ASAP7_75t_L g868 ( .A1(n_869), .A2(n_870), .B1(n_871), .B2(n_872), .Y(n_868) );
INVx2_ASAP7_75t_L g952 ( .A(n_872), .Y(n_952) );
OAI22xp5_ASAP7_75t_L g873 ( .A1(n_874), .A2(n_875), .B1(n_877), .B2(n_878), .Y(n_873) );
BUFx2_ASAP7_75t_R g875 ( .A(n_876), .Y(n_875) );
NOR2xp33_ASAP7_75t_L g879 ( .A(n_880), .B(n_883), .Y(n_879) );
OAI22xp5_ASAP7_75t_L g883 ( .A1(n_884), .A2(n_885), .B1(n_886), .B2(n_887), .Y(n_883) );
INVx3_ASAP7_75t_L g895 ( .A(n_896), .Y(n_895) );
INVx1_ASAP7_75t_L g1029 ( .A(n_903), .Y(n_1029) );
AOI22xp5_ASAP7_75t_SL g903 ( .A1(n_904), .A2(n_974), .B1(n_975), .B2(n_1027), .Y(n_903) );
INVx1_ASAP7_75t_L g1027 ( .A(n_904), .Y(n_1027) );
AOI22xp5_ASAP7_75t_L g904 ( .A1(n_905), .A2(n_931), .B1(n_972), .B2(n_973), .Y(n_904) );
INVx2_ASAP7_75t_L g972 ( .A(n_905), .Y(n_972) );
NAND2xp5_ASAP7_75t_SL g906 ( .A(n_907), .B(n_922), .Y(n_906) );
NOR3xp33_ASAP7_75t_L g907 ( .A(n_908), .B(n_913), .C(n_919), .Y(n_907) );
NAND2xp5_ASAP7_75t_L g908 ( .A(n_909), .B(n_911), .Y(n_908) );
OAI22xp5_ASAP7_75t_L g913 ( .A1(n_914), .A2(n_915), .B1(n_916), .B2(n_917), .Y(n_913) );
INVx4_ASAP7_75t_L g951 ( .A(n_917), .Y(n_951) );
INVx3_ASAP7_75t_L g1085 ( .A(n_917), .Y(n_1085) );
INVx4_ASAP7_75t_L g917 ( .A(n_918), .Y(n_917) );
NOR2xp33_ASAP7_75t_L g922 ( .A(n_923), .B(n_926), .Y(n_922) );
NAND2xp5_ASAP7_75t_L g926 ( .A(n_927), .B(n_930), .Y(n_926) );
INVx1_ASAP7_75t_L g928 ( .A(n_929), .Y(n_928) );
INVx1_ASAP7_75t_L g973 ( .A(n_931), .Y(n_973) );
XNOR2xp5_ASAP7_75t_L g931 ( .A(n_932), .B(n_954), .Y(n_931) );
XNOR2x1_ASAP7_75t_L g932 ( .A(n_933), .B(n_934), .Y(n_932) );
AND2x2_ASAP7_75t_L g934 ( .A(n_935), .B(n_947), .Y(n_934) );
NOR3xp33_ASAP7_75t_L g935 ( .A(n_936), .B(n_940), .C(n_943), .Y(n_935) );
AND4x1_ASAP7_75t_L g947 ( .A(n_948), .B(n_949), .C(n_950), .D(n_953), .Y(n_947) );
INVx2_ASAP7_75t_L g954 ( .A(n_955), .Y(n_954) );
XOR2x2_ASAP7_75t_L g955 ( .A(n_956), .B(n_971), .Y(n_955) );
NAND4xp75_ASAP7_75t_L g956 ( .A(n_957), .B(n_962), .C(n_966), .D(n_969), .Y(n_956) );
AND2x2_ASAP7_75t_L g957 ( .A(n_958), .B(n_961), .Y(n_957) );
INVx3_ASAP7_75t_L g959 ( .A(n_960), .Y(n_959) );
AND2x2_ASAP7_75t_L g966 ( .A(n_967), .B(n_968), .Y(n_966) );
INVx1_ASAP7_75t_L g974 ( .A(n_975), .Y(n_974) );
OAI22xp5_ASAP7_75t_SL g975 ( .A1(n_976), .A2(n_977), .B1(n_1007), .B2(n_1026), .Y(n_975) );
INVx2_ASAP7_75t_L g976 ( .A(n_977), .Y(n_976) );
INVx1_ASAP7_75t_SL g1006 ( .A(n_978), .Y(n_1006) );
AND2x2_ASAP7_75t_SL g978 ( .A(n_979), .B(n_992), .Y(n_978) );
NOR2xp33_ASAP7_75t_L g979 ( .A(n_980), .B(n_987), .Y(n_979) );
INVx1_ASAP7_75t_L g982 ( .A(n_983), .Y(n_982) );
NOR3xp33_ASAP7_75t_L g992 ( .A(n_993), .B(n_996), .C(n_1002), .Y(n_992) );
INVx1_ASAP7_75t_L g1026 ( .A(n_1007), .Y(n_1026) );
INVx1_ASAP7_75t_L g1007 ( .A(n_1008), .Y(n_1007) );
XOR2x2_ASAP7_75t_L g1008 ( .A(n_1009), .B(n_1025), .Y(n_1008) );
NAND3x1_ASAP7_75t_L g1009 ( .A(n_1010), .B(n_1019), .C(n_1022), .Y(n_1009) );
NOR2xp33_ASAP7_75t_L g1010 ( .A(n_1011), .B(n_1015), .Y(n_1010) );
OAI21xp5_ASAP7_75t_SL g1011 ( .A1(n_1012), .A2(n_1013), .B(n_1014), .Y(n_1011) );
NAND3xp33_ASAP7_75t_L g1015 ( .A(n_1016), .B(n_1017), .C(n_1018), .Y(n_1015) );
AND2x2_ASAP7_75t_L g1019 ( .A(n_1020), .B(n_1021), .Y(n_1019) );
AND2x2_ASAP7_75t_L g1022 ( .A(n_1023), .B(n_1024), .Y(n_1022) );
INVx1_ASAP7_75t_SL g1030 ( .A(n_1031), .Y(n_1030) );
NOR2x1_ASAP7_75t_L g1031 ( .A(n_1032), .B(n_1036), .Y(n_1031) );
OR2x2_ASAP7_75t_SL g1093 ( .A(n_1032), .B(n_1037), .Y(n_1093) );
NAND2xp5_ASAP7_75t_L g1032 ( .A(n_1033), .B(n_1035), .Y(n_1032) );
NAND2xp5_ASAP7_75t_L g1071 ( .A(n_1033), .B(n_1072), .Y(n_1071) );
INVx1_ASAP7_75t_L g1033 ( .A(n_1034), .Y(n_1033) );
NAND2xp5_ASAP7_75t_L g1096 ( .A(n_1034), .B(n_1072), .Y(n_1096) );
CKINVDCx16_ASAP7_75t_R g1072 ( .A(n_1035), .Y(n_1072) );
CKINVDCx20_ASAP7_75t_R g1036 ( .A(n_1037), .Y(n_1036) );
NAND2xp5_ASAP7_75t_L g1037 ( .A(n_1038), .B(n_1039), .Y(n_1037) );
NAND2xp5_ASAP7_75t_L g1040 ( .A(n_1041), .B(n_1042), .Y(n_1040) );
OAI222xp33_ASAP7_75t_L g1043 ( .A1(n_1044), .A2(n_1071), .B1(n_1073), .B2(n_1074), .C1(n_1091), .C2(n_1094), .Y(n_1043) );
CKINVDCx20_ASAP7_75t_R g1045 ( .A(n_1046), .Y(n_1045) );
HB1xp67_ASAP7_75t_L g1046 ( .A(n_1047), .Y(n_1046) );
NAND2xp5_ASAP7_75t_L g1047 ( .A(n_1048), .B(n_1062), .Y(n_1047) );
NOR3xp33_ASAP7_75t_L g1048 ( .A(n_1049), .B(n_1053), .C(n_1058), .Y(n_1048) );
OAI21xp33_ASAP7_75t_L g1053 ( .A1(n_1054), .A2(n_1055), .B(n_1056), .Y(n_1053) );
NOR2xp33_ASAP7_75t_L g1062 ( .A(n_1063), .B(n_1067), .Y(n_1062) );
NAND2xp5_ASAP7_75t_L g1063 ( .A(n_1064), .B(n_1065), .Y(n_1063) );
NAND2xp5_ASAP7_75t_L g1067 ( .A(n_1068), .B(n_1069), .Y(n_1067) );
INVx1_ASAP7_75t_SL g1090 ( .A(n_1075), .Y(n_1090) );
NAND4xp75_ASAP7_75t_L g1075 ( .A(n_1076), .B(n_1082), .C(n_1086), .D(n_1089), .Y(n_1075) );
AND2x2_ASAP7_75t_L g1076 ( .A(n_1077), .B(n_1080), .Y(n_1076) );
INVx2_ASAP7_75t_L g1078 ( .A(n_1079), .Y(n_1078) );
AND2x2_ASAP7_75t_L g1082 ( .A(n_1083), .B(n_1084), .Y(n_1082) );
AND2x2_ASAP7_75t_SL g1086 ( .A(n_1087), .B(n_1088), .Y(n_1086) );
CKINVDCx20_ASAP7_75t_R g1091 ( .A(n_1092), .Y(n_1091) );
CKINVDCx20_ASAP7_75t_R g1092 ( .A(n_1093), .Y(n_1092) );
CKINVDCx16_ASAP7_75t_R g1094 ( .A(n_1095), .Y(n_1094) );
endmodule