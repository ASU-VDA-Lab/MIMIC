module fake_jpeg_27460_n_323 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_323);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_323;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

OR2x2_ASAP7_75t_L g16 ( 
.A(n_11),
.B(n_2),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_18),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_34),
.B(n_38),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_16),
.B(n_7),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_42),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_20),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_18),
.Y(n_42)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

OA22x2_ASAP7_75t_L g49 ( 
.A1(n_39),
.A2(n_19),
.B1(n_20),
.B2(n_22),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_49),
.A2(n_40),
.B1(n_22),
.B2(n_42),
.Y(n_62)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_39),
.A2(n_19),
.B1(n_24),
.B2(n_31),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_52),
.A2(n_28),
.B1(n_29),
.B2(n_27),
.Y(n_75)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_54),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_38),
.C(n_40),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_57),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_35),
.B(n_21),
.Y(n_57)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_42),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_61),
.B(n_69),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_62),
.A2(n_75),
.B1(n_29),
.B2(n_27),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_49),
.A2(n_26),
.B1(n_30),
.B2(n_33),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_64),
.A2(n_51),
.B1(n_58),
.B2(n_25),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_44),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_67),
.B(n_77),
.Y(n_96)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_68),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_34),
.Y(n_69)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

BUFx12_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_72),
.Y(n_110)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_54),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_73),
.B(n_53),
.Y(n_95)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_74),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_35),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_78),
.Y(n_101)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_80),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_34),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

BUFx4f_ASAP7_75t_SL g111 ( 
.A(n_81),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_56),
.B(n_38),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_84),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_53),
.B(n_31),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_85),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_86),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g87 ( 
.A(n_49),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_87),
.Y(n_92)
);

AO22x1_ASAP7_75t_SL g88 ( 
.A1(n_68),
.A2(n_50),
.B1(n_48),
.B2(n_46),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_88),
.B(n_108),
.Y(n_130)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_66),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_89),
.B(n_104),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_71),
.A2(n_58),
.B1(n_24),
.B2(n_25),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_94),
.A2(n_103),
.B1(n_113),
.B2(n_75),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_95),
.A2(n_72),
.B(n_70),
.Y(n_141)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_86),
.A2(n_50),
.B1(n_59),
.B2(n_47),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_99),
.A2(n_100),
.B1(n_102),
.B2(n_81),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_62),
.A2(n_59),
.B1(n_47),
.B2(n_54),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_63),
.A2(n_51),
.B1(n_48),
.B2(n_46),
.Y(n_103)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_66),
.Y(n_104)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_60),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_106),
.B(n_112),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_67),
.B(n_53),
.Y(n_108)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_60),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_65),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_114),
.B(n_115),
.Y(n_132)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_65),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_116),
.B(n_76),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_103),
.B(n_63),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_117),
.A2(n_138),
.B(n_141),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_109),
.B(n_77),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_118),
.B(n_123),
.Y(n_148)
);

BUFx2_ASAP7_75t_L g119 ( 
.A(n_111),
.Y(n_119)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_119),
.Y(n_150)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_120),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_90),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_122),
.B(n_135),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_96),
.B(n_77),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_125),
.A2(n_95),
.B1(n_79),
.B2(n_74),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_96),
.B(n_37),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_126),
.B(n_131),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_37),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_127),
.B(n_105),
.Y(n_161)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_101),
.Y(n_128)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_128),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_98),
.B(n_26),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_129),
.B(n_134),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_91),
.B(n_72),
.C(n_53),
.Y(n_131)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_110),
.Y(n_133)
);

INVxp33_ASAP7_75t_L g155 ( 
.A(n_133),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_100),
.B(n_73),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_88),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_91),
.B(n_72),
.C(n_53),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_136),
.B(n_111),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_110),
.B(n_78),
.Y(n_137)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_137),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_107),
.A2(n_0),
.B(n_1),
.Y(n_138)
);

AND2x6_ASAP7_75t_L g139 ( 
.A(n_93),
.B(n_15),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_139),
.B(n_10),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_114),
.B(n_115),
.Y(n_140)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_140),
.Y(n_166)
);

AO22x2_ASAP7_75t_L g142 ( 
.A1(n_93),
.A2(n_85),
.B1(n_83),
.B2(n_76),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_142),
.A2(n_112),
.B1(n_106),
.B2(n_88),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_92),
.B(n_70),
.Y(n_143)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_143),
.Y(n_171)
);

NAND2xp33_ASAP7_75t_SL g144 ( 
.A(n_142),
.B(n_92),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_144),
.A2(n_152),
.B(n_157),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_119),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_145),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_121),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_151),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_130),
.A2(n_117),
.B(n_135),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_153),
.A2(n_168),
.B1(n_172),
.B2(n_32),
.Y(n_205)
);

OAI32xp33_ASAP7_75t_L g154 ( 
.A1(n_130),
.A2(n_105),
.A3(n_95),
.B1(n_97),
.B2(n_33),
.Y(n_154)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_154),
.Y(n_194)
);

OAI21xp33_ASAP7_75t_L g180 ( 
.A1(n_156),
.A2(n_11),
.B(n_15),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_124),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_158),
.B(n_175),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_117),
.A2(n_138),
.B(n_123),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_159),
.A2(n_169),
.B(n_174),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_161),
.B(n_165),
.C(n_170),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_162),
.A2(n_141),
.B1(n_128),
.B2(n_120),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_127),
.B(n_89),
.Y(n_165)
);

CKINVDCx11_ASAP7_75t_R g167 ( 
.A(n_142),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_167),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_116),
.A2(n_142),
.B1(n_131),
.B2(n_136),
.Y(n_168)
);

OA21x2_ASAP7_75t_L g169 ( 
.A1(n_142),
.A2(n_111),
.B(n_104),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_143),
.A2(n_97),
.B1(n_83),
.B2(n_76),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_118),
.A2(n_23),
.B(n_1),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_132),
.Y(n_175)
);

AND2x2_ASAP7_75t_SL g176 ( 
.A(n_126),
.B(n_83),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_176),
.A2(n_0),
.B(n_1),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_146),
.B(n_129),
.Y(n_178)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_178),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_SL g221 ( 
.A(n_179),
.B(n_180),
.C(n_185),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_152),
.A2(n_139),
.B1(n_133),
.B2(n_33),
.Y(n_181)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_181),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_171),
.B(n_23),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_182),
.B(n_189),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_183),
.A2(n_204),
.B(n_205),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_155),
.B(n_23),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_184),
.B(n_188),
.Y(n_210)
);

AND2x6_ASAP7_75t_L g185 ( 
.A(n_156),
.B(n_9),
.Y(n_185)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_150),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_187),
.B(n_198),
.Y(n_229)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_172),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_148),
.B(n_23),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_153),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_190),
.B(n_201),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_176),
.B(n_32),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_193),
.B(n_207),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_161),
.B(n_32),
.C(n_30),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_197),
.B(n_164),
.C(n_157),
.Y(n_230)
);

INVx2_ASAP7_75t_SL g198 ( 
.A(n_169),
.Y(n_198)
);

AND2x6_ASAP7_75t_L g199 ( 
.A(n_159),
.B(n_9),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_199),
.B(n_203),
.Y(n_231)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_169),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_154),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_202),
.B(n_208),
.Y(n_216)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_150),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_168),
.B(n_170),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_149),
.A2(n_0),
.B(n_1),
.Y(n_206)
);

AOI21xp33_ASAP7_75t_L g232 ( 
.A1(n_206),
.A2(n_0),
.B(n_2),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_176),
.B(n_30),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_166),
.B(n_26),
.Y(n_208)
);

AND2x6_ASAP7_75t_L g214 ( 
.A(n_204),
.B(n_149),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_214),
.B(n_231),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_191),
.Y(n_215)
);

OR2x2_ASAP7_75t_L g248 ( 
.A(n_215),
.B(n_218),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_196),
.B(n_163),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_217),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_177),
.Y(n_218)
);

BUFx2_ASAP7_75t_L g220 ( 
.A(n_187),
.Y(n_220)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_220),
.Y(n_236)
);

OAI21xp33_ASAP7_75t_L g222 ( 
.A1(n_178),
.A2(n_173),
.B(n_162),
.Y(n_222)
);

NOR2xp67_ASAP7_75t_SL g243 ( 
.A(n_222),
.B(n_227),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_195),
.B(n_165),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_224),
.B(n_197),
.Y(n_235)
);

NOR2x1_ASAP7_75t_L g225 ( 
.A(n_205),
.B(n_144),
.Y(n_225)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_225),
.Y(n_240)
);

BUFx2_ASAP7_75t_L g226 ( 
.A(n_203),
.Y(n_226)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_226),
.Y(n_245)
);

NAND3xp33_ASAP7_75t_L g227 ( 
.A(n_189),
.B(n_174),
.C(n_11),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_181),
.B(n_160),
.Y(n_228)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_228),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_230),
.B(n_233),
.C(n_193),
.Y(n_247)
);

AO21x1_ASAP7_75t_L g241 ( 
.A1(n_232),
.A2(n_206),
.B(n_192),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_195),
.B(n_164),
.C(n_157),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_234),
.B(n_210),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_235),
.B(n_239),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_215),
.B(n_155),
.Y(n_238)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_238),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_224),
.B(n_192),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_241),
.B(n_242),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_218),
.B(n_182),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_233),
.B(n_207),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_244),
.B(n_246),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_230),
.B(n_204),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_247),
.B(n_253),
.C(n_211),
.Y(n_258)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_220),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_251),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_212),
.B(n_200),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_212),
.B(n_183),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_252),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_211),
.B(n_186),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_223),
.A2(n_194),
.B1(n_198),
.B2(n_199),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_254),
.A2(n_225),
.B1(n_221),
.B2(n_185),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_240),
.A2(n_223),
.B1(n_194),
.B2(n_179),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_255),
.A2(n_265),
.B1(n_232),
.B2(n_8),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_237),
.B(n_209),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_257),
.B(n_264),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_258),
.B(n_236),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_247),
.B(n_209),
.C(n_219),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_259),
.B(n_267),
.C(n_270),
.Y(n_273)
);

O2A1O1Ixp33_ASAP7_75t_L g260 ( 
.A1(n_251),
.A2(n_229),
.B(n_213),
.C(n_198),
.Y(n_260)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_260),
.Y(n_275)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_263),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_243),
.A2(n_216),
.B1(n_221),
.B2(n_219),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_235),
.B(n_214),
.C(n_186),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_248),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_268),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_244),
.B(n_147),
.C(n_226),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_261),
.B(n_248),
.Y(n_272)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_272),
.Y(n_288)
);

FAx1_ASAP7_75t_L g274 ( 
.A(n_269),
.B(n_253),
.CI(n_241),
.CON(n_274),
.SN(n_274)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_274),
.B(n_283),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_270),
.B(n_246),
.C(n_239),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_276),
.B(n_281),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_259),
.B(n_249),
.Y(n_278)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_278),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_262),
.B(n_252),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_280),
.B(n_266),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_266),
.B(n_250),
.C(n_245),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_282),
.B(n_4),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_256),
.A2(n_267),
.B1(n_258),
.B2(n_262),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_284),
.A2(n_6),
.B1(n_13),
.B2(n_4),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_271),
.A2(n_7),
.B(n_14),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_285),
.B(n_255),
.C(n_17),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_287),
.B(n_298),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_SL g289 ( 
.A(n_276),
.B(n_260),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_289),
.B(n_297),
.Y(n_307)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_290),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_294),
.A2(n_296),
.B(n_13),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_279),
.B(n_17),
.Y(n_295)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_295),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_286),
.A2(n_6),
.B(n_10),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_273),
.B(n_5),
.C(n_9),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_295),
.B(n_277),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_299),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_291),
.A2(n_275),
.B1(n_274),
.B2(n_282),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_303),
.A2(n_2),
.B1(n_3),
.B2(n_302),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_297),
.B(n_281),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_304),
.B(n_305),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_288),
.B(n_273),
.Y(n_305)
);

OAI321xp33_ASAP7_75t_L g308 ( 
.A1(n_306),
.A2(n_291),
.A3(n_274),
.B1(n_289),
.B2(n_292),
.C(n_293),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_308),
.A2(n_309),
.B(n_301),
.Y(n_316)
);

INVxp33_ASAP7_75t_L g309 ( 
.A(n_299),
.Y(n_309)
);

NOR2x1_ASAP7_75t_L g310 ( 
.A(n_304),
.B(n_284),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_310),
.B(n_311),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_313),
.B(n_307),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_315),
.B(n_316),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_317),
.B(n_312),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_314),
.C(n_300),
.Y(n_319)
);

BUFx24_ASAP7_75t_SL g320 ( 
.A(n_319),
.Y(n_320)
);

BUFx24_ASAP7_75t_SL g321 ( 
.A(n_320),
.Y(n_321)
);

BUFx24_ASAP7_75t_SL g322 ( 
.A(n_321),
.Y(n_322)
);

MAJx2_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_3),
.C(n_319),
.Y(n_323)
);


endmodule