module fake_jpeg_4173_n_180 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_180);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_180;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_14),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_29),
.B(n_31),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_35),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_15),
.B(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_14),
.B(n_1),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_32),
.B(n_36),
.Y(n_48)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_26),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_41),
.B(n_44),
.Y(n_68)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_35),
.A2(n_24),
.B1(n_28),
.B2(n_16),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_43),
.A2(n_20),
.B1(n_24),
.B2(n_26),
.Y(n_65)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_29),
.B(n_22),
.Y(n_45)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_32),
.B(n_22),
.Y(n_49)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_31),
.B(n_28),
.C(n_18),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_18),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_53),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_58),
.B(n_13),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_15),
.Y(n_60)
);

NAND3xp33_ASAP7_75t_L g86 ( 
.A(n_60),
.B(n_64),
.C(n_21),
.Y(n_86)
);

AO21x1_ASAP7_75t_L g62 ( 
.A1(n_38),
.A2(n_16),
.B(n_20),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_66),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_36),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_64),
.Y(n_76)
);

AND2x2_ASAP7_75t_SL g64 ( 
.A(n_48),
.B(n_36),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_65),
.A2(n_67),
.B1(n_47),
.B2(n_46),
.Y(n_84)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

OA22x2_ASAP7_75t_L g67 ( 
.A1(n_47),
.A2(n_36),
.B1(n_24),
.B2(n_21),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_41),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_70),
.B(n_59),
.Y(n_73)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_71),
.Y(n_99)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_75),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_63),
.B(n_39),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_76),
.B(n_85),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_48),
.C(n_50),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_77),
.B(n_89),
.C(n_58),
.Y(n_92)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_55),
.B(n_44),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_88),
.Y(n_94)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_67),
.Y(n_82)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_83),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_84),
.A2(n_46),
.B1(n_54),
.B2(n_61),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_56),
.B(n_53),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_86),
.B(n_87),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_55),
.B(n_21),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_76),
.A2(n_60),
.B(n_66),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_90),
.A2(n_79),
.B(n_89),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_91),
.A2(n_95),
.B1(n_97),
.B2(n_106),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_77),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_82),
.A2(n_62),
.B1(n_61),
.B2(n_57),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_78),
.A2(n_57),
.B1(n_56),
.B2(n_40),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_81),
.A2(n_51),
.B1(n_40),
.B2(n_26),
.Y(n_106)
);

OA21x2_ASAP7_75t_L g107 ( 
.A1(n_103),
.A2(n_72),
.B(n_88),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_107),
.A2(n_109),
.B(n_117),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_108),
.B(n_112),
.C(n_114),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_94),
.B(n_74),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_110),
.B(n_111),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_93),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_84),
.C(n_83),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_97),
.Y(n_113)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_113),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_90),
.B(n_87),
.C(n_80),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_100),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_115),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_94),
.B(n_21),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_116),
.B(n_101),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_105),
.A2(n_17),
.B(n_21),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_106),
.Y(n_118)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_118),
.Y(n_132)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_95),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_119),
.Y(n_130)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_91),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_121),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_96),
.B(n_2),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_122),
.B(n_99),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_127),
.B(n_17),
.C(n_27),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_131),
.B(n_116),
.Y(n_140)
);

NAND2xp67_ASAP7_75t_SL g133 ( 
.A(n_107),
.B(n_105),
.Y(n_133)
);

AOI321xp33_ASAP7_75t_L g146 ( 
.A1(n_133),
.A2(n_130),
.A3(n_125),
.B1(n_124),
.B2(n_134),
.C(n_129),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_113),
.A2(n_101),
.B1(n_102),
.B2(n_98),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_134),
.A2(n_120),
.B1(n_118),
.B2(n_114),
.Y(n_137)
);

AOI221xp5_ASAP7_75t_L g135 ( 
.A1(n_107),
.A2(n_27),
.B1(n_17),
.B2(n_104),
.C(n_13),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_109),
.Y(n_136)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_136),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_137),
.B(n_138),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_128),
.A2(n_112),
.B1(n_120),
.B2(n_108),
.Y(n_138)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_132),
.Y(n_139)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_139),
.Y(n_155)
);

AOI31xp67_ASAP7_75t_L g150 ( 
.A1(n_140),
.A2(n_146),
.A3(n_127),
.B(n_141),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_141),
.B(n_142),
.C(n_143),
.Y(n_151)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_131),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_126),
.B(n_51),
.C(n_71),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_126),
.B(n_27),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_144),
.B(n_145),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_125),
.A2(n_25),
.B1(n_23),
.B2(n_69),
.Y(n_145)
);

XNOR2x1_ASAP7_75t_L g149 ( 
.A(n_136),
.B(n_133),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_149),
.A2(n_150),
.B(n_9),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_143),
.B(n_144),
.C(n_123),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_152),
.B(n_154),
.C(n_25),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_143),
.B(n_128),
.C(n_130),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_148),
.A2(n_132),
.B(n_25),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_156),
.A2(n_158),
.B(n_159),
.Y(n_165)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_155),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_157),
.B(n_160),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_151),
.B(n_12),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_155),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_147),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_161),
.B(n_153),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_162),
.B(n_23),
.C(n_3),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_163),
.B(n_166),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_156),
.B(n_149),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_164),
.B(n_168),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_162),
.B(n_10),
.Y(n_166)
);

AOI31xp33_ASAP7_75t_L g171 ( 
.A1(n_165),
.A2(n_2),
.A3(n_3),
.B(n_5),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_171),
.A2(n_172),
.B(n_5),
.Y(n_173)
);

AOI21x1_ASAP7_75t_SL g172 ( 
.A1(n_163),
.A2(n_167),
.B(n_6),
.Y(n_172)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_173),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_170),
.A2(n_69),
.B1(n_23),
.B2(n_7),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_174),
.B(n_175),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_169),
.A2(n_5),
.B(n_6),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_177),
.A2(n_7),
.B(n_8),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_176),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_179),
.B(n_7),
.Y(n_180)
);


endmodule