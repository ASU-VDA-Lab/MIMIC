module fake_jpeg_13029_n_104 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_29, n_12, n_8, n_15, n_7, n_104);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_104;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx5_ASAP7_75t_L g30 ( 
.A(n_29),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_18),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

BUFx16f_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_4),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_28),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_39),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_43),
.B(n_49),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_42),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_48),
.C(n_33),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_50),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_42),
.A2(n_14),
.B1(n_27),
.B2(n_23),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_1),
.Y(n_49)
);

BUFx4f_ASAP7_75t_SL g50 ( 
.A(n_30),
.Y(n_50)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_55),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_50),
.B(n_41),
.Y(n_55)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_36),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_SL g69 ( 
.A(n_59),
.B(n_60),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_32),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_54),
.A2(n_51),
.B1(n_56),
.B2(n_32),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_63),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_57),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_SL g64 ( 
.A(n_60),
.B(n_38),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_64),
.B(n_67),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_53),
.A2(n_35),
.B(n_34),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_56),
.A2(n_39),
.B(n_37),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_71),
.Y(n_79)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_58),
.Y(n_70)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g71 ( 
.A1(n_60),
.A2(n_39),
.B(n_37),
.Y(n_71)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

CKINVDCx14_ASAP7_75t_R g83 ( 
.A(n_72),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_57),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_4),
.Y(n_86)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_78),
.Y(n_88)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_2),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_72),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_65),
.B(n_3),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_84),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_86),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_84),
.A2(n_69),
.B1(n_16),
.B2(n_17),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_87),
.A2(n_79),
.B(n_75),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_89),
.B(n_92),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_80),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_90),
.B(n_85),
.C(n_77),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_95),
.A2(n_96),
.B(n_97),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_88),
.A2(n_82),
.B(n_83),
.Y(n_97)
);

AO221x1_ASAP7_75t_L g99 ( 
.A1(n_94),
.A2(n_91),
.B1(n_93),
.B2(n_11),
.C(n_13),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_9),
.C(n_10),
.Y(n_100)
);

AOI21x1_ASAP7_75t_L g101 ( 
.A1(n_100),
.A2(n_98),
.B(n_19),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_15),
.Y(n_102)
);

BUFx24_ASAP7_75t_SL g103 ( 
.A(n_102),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_103),
.Y(n_104)
);


endmodule