module fake_ariane_2098_n_192 (n_8, n_24, n_7, n_22, n_1, n_6, n_13, n_20, n_27, n_29, n_17, n_4, n_2, n_18, n_28, n_9, n_11, n_26, n_3, n_14, n_0, n_19, n_30, n_31, n_16, n_5, n_12, n_15, n_21, n_23, n_10, n_25, n_192);

input n_8;
input n_24;
input n_7;
input n_22;
input n_1;
input n_6;
input n_13;
input n_20;
input n_27;
input n_29;
input n_17;
input n_4;
input n_2;
input n_18;
input n_28;
input n_9;
input n_11;
input n_26;
input n_3;
input n_14;
input n_0;
input n_19;
input n_30;
input n_31;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_23;
input n_10;
input n_25;

output n_192;

wire n_83;
wire n_56;
wire n_60;
wire n_170;
wire n_190;
wire n_160;
wire n_64;
wire n_179;
wire n_180;
wire n_119;
wire n_124;
wire n_167;
wire n_90;
wire n_38;
wire n_47;
wire n_110;
wire n_153;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_176;
wire n_149;
wire n_34;
wire n_158;
wire n_172;
wire n_69;
wire n_95;
wire n_175;
wire n_92;
wire n_143;
wire n_183;
wire n_150;
wire n_98;
wire n_74;
wire n_113;
wire n_114;
wire n_33;
wire n_40;
wire n_181;
wire n_152;
wire n_120;
wire n_169;
wire n_106;
wire n_53;
wire n_173;
wire n_111;
wire n_115;
wire n_133;
wire n_66;
wire n_71;
wire n_109;
wire n_96;
wire n_156;
wire n_49;
wire n_174;
wire n_100;
wire n_50;
wire n_187;
wire n_132;
wire n_62;
wire n_147;
wire n_51;
wire n_166;
wire n_76;
wire n_103;
wire n_79;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_159;
wire n_107;
wire n_189;
wire n_72;
wire n_105;
wire n_128;
wire n_44;
wire n_82;
wire n_178;
wire n_42;
wire n_57;
wire n_131;
wire n_70;
wire n_117;
wire n_139;
wire n_165;
wire n_85;
wire n_130;
wire n_144;
wire n_48;
wire n_94;
wire n_101;
wire n_134;
wire n_188;
wire n_185;
wire n_32;
wire n_37;
wire n_58;
wire n_65;
wire n_123;
wire n_138;
wire n_112;
wire n_45;
wire n_162;
wire n_129;
wire n_126;
wire n_137;
wire n_122;
wire n_148;
wire n_164;
wire n_52;
wire n_157;
wire n_184;
wire n_177;
wire n_135;
wire n_73;
wire n_77;
wire n_171;
wire n_118;
wire n_93;
wire n_121;
wire n_61;
wire n_108;
wire n_102;
wire n_182;
wire n_125;
wire n_168;
wire n_43;
wire n_87;
wire n_81;
wire n_41;
wire n_140;
wire n_55;
wire n_191;
wire n_151;
wire n_136;
wire n_146;
wire n_80;
wire n_97;
wire n_154;
wire n_142;
wire n_161;
wire n_163;
wire n_88;
wire n_186;
wire n_141;
wire n_68;
wire n_116;
wire n_104;
wire n_145;
wire n_78;
wire n_39;
wire n_59;
wire n_63;
wire n_99;
wire n_155;
wire n_127;
wire n_35;
wire n_54;

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_16),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_15),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

CKINVDCx5p33_ASAP7_75t_R g43 ( 
.A(n_6),
.Y(n_43)
);

INVxp67_ASAP7_75t_SL g44 ( 
.A(n_17),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_2),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

INVxp67_ASAP7_75t_SL g48 ( 
.A(n_3),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_20),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

INVxp67_ASAP7_75t_SL g51 ( 
.A(n_15),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_13),
.Y(n_53)
);

INVxp67_ASAP7_75t_SL g54 ( 
.A(n_7),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_9),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_33),
.B(n_0),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_49),
.A2(n_46),
.B1(n_41),
.B2(n_53),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

AND2x4_ASAP7_75t_L g64 ( 
.A(n_33),
.B(n_1),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_35),
.B(n_4),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_38),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_44),
.B(n_5),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

OR2x2_ASAP7_75t_SL g77 ( 
.A(n_74),
.B(n_52),
.Y(n_77)
);

OAI221xp5_ASAP7_75t_L g78 ( 
.A1(n_58),
.A2(n_50),
.B1(n_54),
.B2(n_51),
.C(n_48),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

OAI221xp5_ASAP7_75t_L g80 ( 
.A1(n_58),
.A2(n_55),
.B1(n_42),
.B2(n_32),
.C(n_43),
.Y(n_80)
);

NOR2x1p5_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_43),
.Y(n_81)
);

AO22x2_ASAP7_75t_L g82 ( 
.A1(n_64),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_82)
);

OAI221xp5_ASAP7_75t_L g83 ( 
.A1(n_60),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.C(n_12),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_14),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

AO22x2_ASAP7_75t_L g86 ( 
.A1(n_64),
.A2(n_16),
.B1(n_19),
.B2(n_21),
.Y(n_86)
);

NAND3xp33_ASAP7_75t_L g87 ( 
.A(n_59),
.B(n_22),
.C(n_24),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_60),
.B(n_26),
.Y(n_88)
);

AND3x1_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_28),
.C(n_29),
.Y(n_89)
);

AO22x2_ASAP7_75t_L g90 ( 
.A1(n_64),
.A2(n_30),
.B1(n_31),
.B2(n_67),
.Y(n_90)
);

NAND2x1p5_ASAP7_75t_L g91 ( 
.A(n_61),
.B(n_64),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_61),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g93 ( 
.A(n_59),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

AND2x2_ASAP7_75t_SL g95 ( 
.A(n_89),
.B(n_67),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_91),
.B(n_65),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_82),
.A2(n_62),
.B1(n_57),
.B2(n_68),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_90),
.A2(n_65),
.B1(n_63),
.B2(n_56),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_63),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_72),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_77),
.B(n_93),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_103),
.B(n_92),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_95),
.B(n_87),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_103),
.B(n_90),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_103),
.B(n_88),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_94),
.A2(n_84),
.B(n_88),
.Y(n_111)
);

O2A1O1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_99),
.A2(n_83),
.B(n_98),
.C(n_102),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_R g113 ( 
.A(n_96),
.B(n_79),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_106),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_110),
.B(n_96),
.Y(n_115)
);

OA21x2_ASAP7_75t_L g116 ( 
.A1(n_111),
.A2(n_105),
.B(n_100),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_107),
.A2(n_95),
.B1(n_110),
.B2(n_90),
.Y(n_117)
);

HB1xp67_ASAP7_75t_L g118 ( 
.A(n_113),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_104),
.Y(n_119)
);

AO32x1_ASAP7_75t_L g120 ( 
.A1(n_109),
.A2(n_99),
.A3(n_105),
.B1(n_90),
.B2(n_86),
.Y(n_120)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_115),
.B(n_104),
.Y(n_121)
);

OA21x2_ASAP7_75t_L g122 ( 
.A1(n_117),
.A2(n_87),
.B(n_108),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_116),
.Y(n_123)
);

CKINVDCx5p33_ASAP7_75t_R g124 ( 
.A(n_118),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_114),
.B(n_101),
.Y(n_125)
);

NAND3xp33_ASAP7_75t_L g126 ( 
.A(n_125),
.B(n_107),
.C(n_118),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_123),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_123),
.Y(n_128)
);

AND2x4_ASAP7_75t_L g129 ( 
.A(n_121),
.B(n_119),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_123),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_123),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_123),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_124),
.B(n_114),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_123),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_123),
.Y(n_135)
);

INVxp67_ASAP7_75t_SL g136 ( 
.A(n_125),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_129),
.B(n_82),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_127),
.Y(n_138)
);

NAND2xp33_ASAP7_75t_SL g139 ( 
.A(n_129),
.B(n_121),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_127),
.Y(n_140)
);

INVx1_ASAP7_75t_SL g141 ( 
.A(n_133),
.Y(n_141)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_129),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_126),
.A2(n_95),
.B1(n_89),
.B2(n_86),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_138),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_142),
.B(n_136),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_141),
.B(n_121),
.Y(n_146)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_138),
.B(n_135),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_137),
.B(n_135),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_137),
.B(n_130),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_139),
.B(n_130),
.Y(n_150)
);

OR2x2_ASAP7_75t_L g151 ( 
.A(n_140),
.B(n_132),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_140),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_146),
.B(n_112),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_145),
.B(n_132),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_148),
.B(n_128),
.Y(n_155)
);

OAI221xp5_ASAP7_75t_L g156 ( 
.A1(n_150),
.A2(n_143),
.B1(n_80),
.B2(n_78),
.C(n_70),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_144),
.B(n_134),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_149),
.B(n_66),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_152),
.A2(n_82),
.B1(n_86),
.B2(n_122),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_147),
.Y(n_160)
);

OAI32xp33_ASAP7_75t_L g161 ( 
.A1(n_151),
.A2(n_57),
.A3(n_75),
.B1(n_72),
.B2(n_73),
.Y(n_161)
);

AND2x2_ASAP7_75t_SL g162 ( 
.A(n_160),
.B(n_149),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_160),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_160),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_159),
.B(n_82),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_155),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_154),
.B(n_134),
.Y(n_167)
);

NOR2x1_ASAP7_75t_L g168 ( 
.A(n_158),
.B(n_70),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_157),
.Y(n_169)
);

AOI322xp5_ASAP7_75t_L g170 ( 
.A1(n_162),
.A2(n_153),
.A3(n_73),
.B1(n_75),
.B2(n_120),
.C1(n_76),
.C2(n_66),
.Y(n_170)
);

OAI221xp5_ASAP7_75t_L g171 ( 
.A1(n_165),
.A2(n_156),
.B1(n_71),
.B2(n_76),
.C(n_66),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_169),
.B(n_66),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_165),
.A2(n_86),
.B1(n_122),
.B2(n_81),
.Y(n_173)
);

NAND3x1_ASAP7_75t_L g174 ( 
.A(n_163),
.B(n_120),
.C(n_161),
.Y(n_174)
);

A2O1A1Ixp33_ASAP7_75t_L g175 ( 
.A1(n_162),
.A2(n_66),
.B(n_71),
.C(n_76),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_169),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_175),
.A2(n_164),
.B(n_166),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_173),
.B(n_167),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_171),
.A2(n_122),
.B1(n_167),
.B2(n_168),
.Y(n_179)
);

OAI211xp5_ASAP7_75t_L g180 ( 
.A1(n_170),
.A2(n_66),
.B(n_71),
.C(n_76),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_176),
.B(n_71),
.Y(n_181)
);

AOI221xp5_ASAP7_75t_L g182 ( 
.A1(n_172),
.A2(n_71),
.B1(n_76),
.B2(n_77),
.C(n_120),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_181),
.Y(n_183)
);

AOI322xp5_ASAP7_75t_L g184 ( 
.A1(n_179),
.A2(n_173),
.A3(n_71),
.B1(n_76),
.B2(n_174),
.C1(n_122),
.C2(n_81),
.Y(n_184)
);

AOI322xp5_ASAP7_75t_L g185 ( 
.A1(n_182),
.A2(n_122),
.A3(n_96),
.B1(n_128),
.B2(n_131),
.C1(n_101),
.C2(n_105),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_178),
.A2(n_131),
.B1(n_104),
.B2(n_116),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_177),
.A2(n_94),
.B1(n_98),
.B2(n_102),
.Y(n_187)
);

AOI211xp5_ASAP7_75t_L g188 ( 
.A1(n_187),
.A2(n_180),
.B(n_101),
.C(n_97),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_183),
.Y(n_189)
);

AOI21xp33_ASAP7_75t_L g190 ( 
.A1(n_189),
.A2(n_186),
.B(n_184),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_188),
.B(n_185),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_191),
.A2(n_97),
.B1(n_108),
.B2(n_190),
.Y(n_192)
);


endmodule