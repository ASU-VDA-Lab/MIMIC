module real_jpeg_29354_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_330, n_12, n_6, n_11, n_14, n_7, n_329, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_330;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_329;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_0),
.Y(n_77)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_0),
.Y(n_83)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_0),
.Y(n_178)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_1),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_L g38 ( 
.A1(n_2),
.A2(n_29),
.B1(n_30),
.B2(n_39),
.Y(n_38)
);

CKINVDCx14_ASAP7_75t_R g39 ( 
.A(n_2),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_2),
.A2(n_39),
.B1(n_61),
.B2(n_62),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_2),
.A2(n_35),
.B1(n_36),
.B2(n_39),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_2),
.A2(n_39),
.B1(n_52),
.B2(n_54),
.Y(n_168)
);

BUFx8_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

OAI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_4),
.A2(n_61),
.B1(n_62),
.B2(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_4),
.Y(n_69)
);

AOI21xp33_ASAP7_75t_SL g74 ( 
.A1(n_4),
.A2(n_30),
.B(n_64),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_4),
.B(n_66),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_4),
.A2(n_35),
.B(n_148),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_4),
.B(n_35),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_4),
.B(n_92),
.Y(n_157)
);

OAI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_4),
.A2(n_103),
.B1(n_174),
.B2(n_178),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_4),
.A2(n_29),
.B(n_190),
.Y(n_189)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_5),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_6),
.A2(n_52),
.B1(n_54),
.B2(n_79),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_6),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_6),
.A2(n_35),
.B1(n_36),
.B2(n_79),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_79),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_6),
.A2(n_61),
.B1(n_62),
.B2(n_79),
.Y(n_282)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_7),
.A2(n_61),
.B1(n_62),
.B2(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_7),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_7),
.A2(n_29),
.B1(n_30),
.B2(n_71),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_7),
.A2(n_35),
.B1(n_36),
.B2(n_71),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_7),
.A2(n_52),
.B1(n_54),
.B2(n_71),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_8),
.A2(n_52),
.B1(n_54),
.B2(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_8),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_8),
.A2(n_35),
.B1(n_36),
.B2(n_106),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_8),
.A2(n_29),
.B1(n_30),
.B2(n_106),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_SL g321 ( 
.A1(n_8),
.A2(n_61),
.B1(n_62),
.B2(n_106),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_9),
.A2(n_35),
.B1(n_36),
.B2(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_9),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_9),
.A2(n_29),
.B1(n_30),
.B2(n_46),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_9),
.A2(n_46),
.B1(n_52),
.B2(n_54),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_9),
.A2(n_46),
.B1(n_61),
.B2(n_62),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_41),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_10),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_10),
.A2(n_41),
.B1(n_61),
.B2(n_62),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_10),
.A2(n_41),
.B1(n_52),
.B2(n_54),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_10),
.A2(n_35),
.B1(n_36),
.B2(n_41),
.Y(n_194)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_12),
.A2(n_52),
.B1(n_54),
.B2(n_128),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_12),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_12),
.A2(n_35),
.B1(n_36),
.B2(n_128),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_12),
.A2(n_29),
.B1(n_30),
.B2(n_128),
.Y(n_300)
);

BUFx24_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

A2O1A1Ixp33_ASAP7_75t_L g28 ( 
.A1(n_14),
.A2(n_29),
.B(n_31),
.C(n_34),
.Y(n_28)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_14),
.A2(n_33),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_14),
.Y(n_200)
);

OAI22xp33_ASAP7_75t_L g56 ( 
.A1(n_15),
.A2(n_35),
.B1(n_36),
.B2(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_15),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_15),
.A2(n_52),
.B1(n_54),
.B2(n_57),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_15),
.A2(n_29),
.B1(n_30),
.B2(n_57),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_15),
.A2(n_57),
.B1(n_61),
.B2(n_62),
.Y(n_260)
);

INVx11_ASAP7_75t_SL g53 ( 
.A(n_16),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_17),
.A2(n_52),
.B1(n_54),
.B2(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_17),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_17),
.A2(n_35),
.B1(n_36),
.B2(n_85),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_17),
.A2(n_29),
.B1(n_30),
.B2(n_85),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_17),
.A2(n_61),
.B1(n_62),
.B2(n_85),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_309),
.Y(n_18)
);

OAI321xp33_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_277),
.A3(n_304),
.B1(n_307),
.B2(n_308),
.C(n_329),
.Y(n_19)
);

AOI321xp33_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_228),
.A3(n_266),
.B1(n_271),
.B2(n_276),
.C(n_330),
.Y(n_20)
);

NOR3xp33_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_120),
.C(n_139),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_96),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_23),
.B(n_96),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_72),
.C(n_86),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_24),
.B(n_225),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_59),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_42),
.B2(n_43),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_26),
.B(n_43),
.C(n_59),
.Y(n_107)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_28),
.A2(n_34),
.B1(n_37),
.B2(n_40),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_28),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_28),
.A2(n_34),
.B1(n_40),
.B2(n_117),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_28),
.A2(n_34),
.B1(n_90),
.B2(n_189),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_28),
.A2(n_34),
.B1(n_250),
.B2(n_251),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_28),
.A2(n_34),
.B(n_317),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_29),
.B(n_32),
.Y(n_31)
);

AO22x1_ASAP7_75t_L g66 ( 
.A1(n_29),
.A2(n_30),
.B1(n_64),
.B2(n_67),
.Y(n_66)
);

OAI32xp33_ASAP7_75t_L g198 ( 
.A1(n_29),
.A2(n_36),
.A3(n_191),
.B1(n_199),
.B2(n_201),
.Y(n_198)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_30),
.B(n_69),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_34),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_L g55 ( 
.A1(n_35),
.A2(n_36),
.B1(n_50),
.B2(n_51),
.Y(n_55)
);

OAI32xp33_ASAP7_75t_L g151 ( 
.A1(n_35),
.A2(n_50),
.A3(n_54),
.B1(n_152),
.B2(n_153),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_35),
.B(n_202),
.Y(n_201)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_38),
.A2(n_89),
.B1(n_91),
.B2(n_92),
.Y(n_88)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_47),
.B1(n_56),
.B2(n_58),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_45),
.A2(n_48),
.B1(n_49),
.B2(n_218),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_47),
.A2(n_58),
.B1(n_193),
.B2(n_194),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_47),
.A2(n_58),
.B1(n_239),
.B2(n_240),
.Y(n_238)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_48),
.A2(n_49),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_48),
.A2(n_49),
.B1(n_101),
.B2(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_48),
.A2(n_49),
.B1(n_147),
.B2(n_149),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_48),
.A2(n_49),
.B1(n_149),
.B2(n_160),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_48),
.A2(n_49),
.B1(n_241),
.B2(n_253),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_48),
.A2(n_49),
.B(n_253),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_49),
.B(n_55),
.Y(n_48)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_49),
.B(n_69),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_51),
.B1(n_52),
.B2(n_54),
.Y(n_49)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_51),
.B(n_52),
.Y(n_153)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_52),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_52),
.B(n_77),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_52),
.B(n_180),
.Y(n_179)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_56),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_66),
.B1(n_68),
.B2(n_70),
.Y(n_59)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_60),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_60),
.A2(n_66),
.B1(n_115),
.B2(n_135),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_60),
.A2(n_66),
.B1(n_135),
.B2(n_232),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_60),
.A2(n_66),
.B1(n_296),
.B2(n_297),
.Y(n_295)
);

O2A1O1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_64),
.B(n_65),
.C(n_66),
.Y(n_60)
);

NAND2xp33_ASAP7_75t_SL g65 ( 
.A(n_61),
.B(n_64),
.Y(n_65)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

A2O1A1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_62),
.A2(n_67),
.B(n_69),
.C(n_74),
.Y(n_73)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_64),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_66),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_69),
.B(n_83),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_70),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_72),
.A2(n_86),
.B1(n_87),
.B2(n_226),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_72),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_75),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_73),
.B(n_75),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_78),
.B1(n_80),
.B2(n_84),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_76),
.A2(n_78),
.B1(n_82),
.B2(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_76),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_76),
.A2(n_80),
.B1(n_167),
.B2(n_169),
.Y(n_166)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_81),
.A2(n_103),
.B1(n_104),
.B2(n_105),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_81),
.A2(n_103),
.B1(n_105),
.B2(n_127),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_81),
.A2(n_103),
.B1(n_162),
.B2(n_163),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_81),
.A2(n_103),
.B1(n_168),
.B2(n_174),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_81),
.A2(n_103),
.B1(n_163),
.B2(n_204),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_81),
.A2(n_103),
.B(n_127),
.Y(n_243)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_84),
.Y(n_104)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_93),
.C(n_95),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_88),
.B(n_213),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_91),
.A2(n_92),
.B1(n_118),
.B2(n_137),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_91),
.A2(n_92),
.B1(n_137),
.B2(n_234),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_91),
.A2(n_92),
.B1(n_285),
.B2(n_286),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_91),
.A2(n_92),
.B1(n_286),
.B2(n_300),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_93),
.B(n_95),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_94),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_108),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_107),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_98),
.B(n_107),
.C(n_108),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_102),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_99),
.B(n_102),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g108 ( 
.A(n_109),
.B(n_119),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_116),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_110),
.B(n_116),
.C(n_119),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_111),
.A2(n_112),
.B1(n_113),
.B2(n_114),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_111),
.A2(n_113),
.B1(n_259),
.B2(n_260),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_111),
.A2(n_113),
.B1(n_260),
.B2(n_282),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_111),
.A2(n_113),
.B1(n_320),
.B2(n_321),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

AOI21xp33_ASAP7_75t_L g272 ( 
.A1(n_121),
.A2(n_273),
.B(n_274),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_123),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_122),
.B(n_123),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_138),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_131),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_125),
.B(n_131),
.C(n_138),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_129),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_126),
.B(n_129),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_130),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_133),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_132),
.B(n_134),
.C(n_136),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_136),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_222),
.B(n_227),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_208),
.B(n_221),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_184),
.B(n_207),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_164),
.B(n_183),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_154),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_144),
.B(n_154),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_145),
.B(n_150),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_145),
.A2(n_146),
.B1(n_150),
.B2(n_151),
.Y(n_170)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_148),
.Y(n_152)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_161),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_157),
.B1(n_158),
.B2(n_159),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_156),
.B(n_159),
.C(n_161),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_160),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_162),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_171),
.B(n_182),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_170),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_166),
.B(n_170),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_176),
.B(n_181),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_175),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_173),
.B(n_175),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_177),
.B(n_179),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_185),
.B(n_186),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_187),
.A2(n_197),
.B1(n_205),
.B2(n_206),
.Y(n_186)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_187),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_192),
.B1(n_195),
.B2(n_196),
.Y(n_187)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_188),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_192),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_192),
.B(n_196),
.C(n_206),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_194),
.Y(n_218)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_197),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_203),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_198),
.B(n_203),
.Y(n_216)
);

INVx6_ASAP7_75t_L g202 ( 
.A(n_199),
.Y(n_202)
);

INVx8_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_209),
.B(n_210),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_211),
.A2(n_212),
.B1(n_214),
.B2(n_215),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_211),
.B(n_217),
.C(n_219),
.Y(n_223)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_216),
.A2(n_217),
.B1(n_219),
.B2(n_220),
.Y(n_215)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_216),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_217),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_223),
.B(n_224),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_245),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_229),
.B(n_245),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_236),
.C(n_244),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_230),
.B(n_236),
.Y(n_270)
);

BUFx24_ASAP7_75t_SL g327 ( 
.A(n_230),
.Y(n_327)
);

FAx1_ASAP7_75t_SL g230 ( 
.A(n_231),
.B(n_233),
.CI(n_235),
.CON(n_230),
.SN(n_230)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_231),
.B(n_233),
.C(n_235),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_232),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_234),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_237),
.A2(n_238),
.B1(n_242),
.B2(n_243),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_237),
.B(n_243),
.Y(n_262)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_241),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_242),
.A2(n_243),
.B1(n_257),
.B2(n_258),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_242),
.A2(n_258),
.B(n_261),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_243),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_244),
.B(n_270),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_246),
.A2(n_247),
.B1(n_264),
.B2(n_265),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_255),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_248),
.B(n_255),
.C(n_265),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_252),
.B(n_254),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_249),
.B(n_252),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_251),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_254),
.B(n_279),
.C(n_291),
.Y(n_278)
);

FAx1_ASAP7_75t_SL g306 ( 
.A(n_254),
.B(n_279),
.CI(n_291),
.CON(n_306),
.SN(n_306)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_261),
.B1(n_262),
.B2(n_263),
.Y(n_255)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_256),
.Y(n_263)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_264),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_267),
.A2(n_272),
.B(n_275),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_268),
.B(n_269),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_292),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_278),
.B(n_292),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_281),
.B1(n_283),
.B2(n_290),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_280),
.A2(n_281),
.B1(n_294),
.B2(n_302),
.Y(n_293)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_281),
.B(n_284),
.C(n_289),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_281),
.B(n_302),
.C(n_303),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_282),
.Y(n_296)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_283),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_287),
.B1(n_288),
.B2(n_289),
.Y(n_283)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_284),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_287),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_287),
.A2(n_289),
.B1(n_299),
.B2(n_301),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_287),
.B(n_295),
.C(n_299),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_303),
.Y(n_292)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_294),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_SL g294 ( 
.A(n_295),
.B(n_298),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_297),
.Y(n_320)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_299),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_300),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_305),
.B(n_306),
.Y(n_307)
);

BUFx24_ASAP7_75t_SL g328 ( 
.A(n_306),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_324),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_311),
.B(n_312),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_314),
.B1(n_322),
.B2(n_323),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_315),
.A2(n_316),
.B1(n_318),
.B2(n_319),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_316),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_319),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_323),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);


endmodule