module fake_jpeg_18081_n_78 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_78);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_78;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

INVx1_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_6),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

BUFx3_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_18),
.B(n_20),
.Y(n_24)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_10),
.B(n_0),
.Y(n_21)
);

AOI21xp33_ASAP7_75t_L g28 ( 
.A1(n_21),
.A2(n_22),
.B(n_13),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_23),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_19),
.A2(n_15),
.B1(n_10),
.B2(n_13),
.Y(n_26)
);

CKINVDCx14_ASAP7_75t_R g35 ( 
.A(n_26),
.Y(n_35)
);

A2O1A1Ixp33_ASAP7_75t_L g36 ( 
.A1(n_28),
.A2(n_26),
.B(n_20),
.C(n_11),
.Y(n_36)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

HB1xp67_ASAP7_75t_L g30 ( 
.A(n_29),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_24),
.B(n_21),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_32),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_24),
.B(n_18),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_28),
.A2(n_23),
.B1(n_18),
.B2(n_20),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_33),
.A2(n_36),
.B(n_0),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_25),
.B(n_19),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_38),
.B(n_27),
.C(n_19),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_27),
.C(n_22),
.Y(n_50)
);

NAND2xp33_ASAP7_75t_SL g42 ( 
.A(n_36),
.B(n_29),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_SL g49 ( 
.A1(n_42),
.A2(n_44),
.B(n_33),
.Y(n_49)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_46),
.Y(n_53)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

AO21x2_ASAP7_75t_L g47 ( 
.A1(n_35),
.A2(n_29),
.B(n_25),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_47),
.A2(n_25),
.B1(n_37),
.B2(n_17),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_39),
.B(n_16),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_48),
.B(n_55),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g58 ( 
.A1(n_49),
.A2(n_51),
.B(n_52),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_44),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_12),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g59 ( 
.A1(n_54),
.A2(n_43),
.B(n_16),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_17),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_57),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_59),
.B(n_60),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_54),
.Y(n_60)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_64),
.Y(n_67)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_61),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_57),
.B(n_5),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_66),
.B(n_8),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_68),
.B(n_3),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g69 ( 
.A1(n_63),
.A2(n_52),
.B(n_47),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_69),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_67),
.A2(n_47),
.B1(n_65),
.B2(n_62),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_71),
.A2(n_47),
.B(n_2),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_4),
.Y(n_73)
);

AOI322xp5_ASAP7_75t_L g75 ( 
.A1(n_73),
.A2(n_74),
.A3(n_70),
.B1(n_8),
.B2(n_2),
.C1(n_1),
.C2(n_12),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_75),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_1),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_1),
.Y(n_78)
);


endmodule