module fake_aes_7437_n_677 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_677);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_677;
wire n_117;
wire n_663;
wire n_513;
wire n_361;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_624;
wire n_426;
wire n_255;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_415;
wire n_482;
wire n_394;
wire n_235;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_428;
wire n_364;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_515;
wire n_253;
wire n_670;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVxp67_ASAP7_75t_SL g79 ( .A(n_25), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_54), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_75), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_8), .Y(n_82) );
INVxp67_ASAP7_75t_SL g83 ( .A(n_22), .Y(n_83) );
CKINVDCx20_ASAP7_75t_R g84 ( .A(n_69), .Y(n_84) );
INVxp67_ASAP7_75t_SL g85 ( .A(n_62), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_15), .Y(n_86) );
INVx2_ASAP7_75t_L g87 ( .A(n_65), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_13), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_31), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_43), .Y(n_90) );
CKINVDCx16_ASAP7_75t_R g91 ( .A(n_34), .Y(n_91) );
INVxp67_ASAP7_75t_SL g92 ( .A(n_42), .Y(n_92) );
INVxp67_ASAP7_75t_SL g93 ( .A(n_52), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_33), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_77), .Y(n_95) );
INVx2_ASAP7_75t_L g96 ( .A(n_24), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_41), .Y(n_97) );
INVx2_ASAP7_75t_L g98 ( .A(n_32), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_63), .Y(n_99) );
INVxp33_ASAP7_75t_L g100 ( .A(n_58), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_48), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_78), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_56), .Y(n_103) );
BUFx3_ASAP7_75t_L g104 ( .A(n_38), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_2), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_12), .B(n_7), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_76), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g108 ( .A(n_70), .B(n_71), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_44), .Y(n_109) );
INVxp33_ASAP7_75t_SL g110 ( .A(n_37), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g111 ( .A(n_49), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_59), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_64), .Y(n_113) );
HB1xp67_ASAP7_75t_L g114 ( .A(n_26), .Y(n_114) );
CKINVDCx16_ASAP7_75t_R g115 ( .A(n_36), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_27), .Y(n_116) );
INVxp67_ASAP7_75t_SL g117 ( .A(n_3), .Y(n_117) );
INVx2_ASAP7_75t_L g118 ( .A(n_30), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_11), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_29), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_18), .Y(n_121) );
BUFx3_ASAP7_75t_L g122 ( .A(n_19), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_74), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_23), .Y(n_124) );
INVxp33_ASAP7_75t_L g125 ( .A(n_6), .Y(n_125) );
INVxp67_ASAP7_75t_L g126 ( .A(n_20), .Y(n_126) );
INVxp67_ASAP7_75t_SL g127 ( .A(n_20), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_66), .Y(n_128) );
NAND2xp33_ASAP7_75t_R g129 ( .A(n_110), .B(n_0), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_87), .Y(n_130) );
INVx3_ASAP7_75t_L g131 ( .A(n_122), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g132 ( .A(n_91), .Y(n_132) );
INVx3_ASAP7_75t_L g133 ( .A(n_122), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_114), .B(n_0), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_122), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_82), .B(n_1), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_80), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_80), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_81), .Y(n_139) );
INVx6_ASAP7_75t_L g140 ( .A(n_104), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_81), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_87), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_87), .Y(n_143) );
OR2x6_ASAP7_75t_L g144 ( .A(n_106), .B(n_28), .Y(n_144) );
HB1xp67_ASAP7_75t_L g145 ( .A(n_126), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_82), .B(n_1), .Y(n_146) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_104), .Y(n_147) );
NAND2xp5_ASAP7_75t_SL g148 ( .A(n_91), .B(n_2), .Y(n_148) );
AND2x2_ASAP7_75t_L g149 ( .A(n_125), .B(n_3), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g150 ( .A(n_115), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_89), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_89), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_96), .Y(n_153) );
CKINVDCx5p33_ASAP7_75t_R g154 ( .A(n_115), .Y(n_154) );
HB1xp67_ASAP7_75t_L g155 ( .A(n_126), .Y(n_155) );
CKINVDCx20_ASAP7_75t_R g156 ( .A(n_84), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_86), .B(n_4), .Y(n_157) );
AND2x4_ASAP7_75t_L g158 ( .A(n_104), .B(n_4), .Y(n_158) );
BUFx2_ASAP7_75t_L g159 ( .A(n_86), .Y(n_159) );
CKINVDCx5p33_ASAP7_75t_R g160 ( .A(n_107), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_96), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_90), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_90), .Y(n_163) );
CKINVDCx5p33_ASAP7_75t_R g164 ( .A(n_111), .Y(n_164) );
INVx3_ASAP7_75t_L g165 ( .A(n_96), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_98), .Y(n_166) );
CKINVDCx5p33_ASAP7_75t_R g167 ( .A(n_99), .Y(n_167) );
HB1xp67_ASAP7_75t_L g168 ( .A(n_88), .Y(n_168) );
CKINVDCx20_ASAP7_75t_R g169 ( .A(n_106), .Y(n_169) );
INVxp67_ASAP7_75t_SL g170 ( .A(n_88), .Y(n_170) );
INVx3_ASAP7_75t_L g171 ( .A(n_98), .Y(n_171) );
INVx3_ASAP7_75t_L g172 ( .A(n_98), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_94), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_137), .B(n_100), .Y(n_174) );
AND2x4_ASAP7_75t_L g175 ( .A(n_170), .B(n_105), .Y(n_175) );
NAND2xp5_ASAP7_75t_SL g176 ( .A(n_158), .B(n_118), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_147), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_158), .Y(n_178) );
NAND2x1p5_ASAP7_75t_L g179 ( .A(n_149), .B(n_105), .Y(n_179) );
NAND2xp5_ASAP7_75t_SL g180 ( .A(n_158), .B(n_118), .Y(n_180) );
AND2x4_ASAP7_75t_L g181 ( .A(n_170), .B(n_119), .Y(n_181) );
AND2x2_ASAP7_75t_L g182 ( .A(n_145), .B(n_121), .Y(n_182) );
INVx2_ASAP7_75t_SL g183 ( .A(n_158), .Y(n_183) );
CKINVDCx5p33_ASAP7_75t_R g184 ( .A(n_150), .Y(n_184) );
AND2x4_ASAP7_75t_L g185 ( .A(n_159), .B(n_119), .Y(n_185) );
INVx1_ASAP7_75t_SL g186 ( .A(n_154), .Y(n_186) );
HB1xp67_ASAP7_75t_L g187 ( .A(n_145), .Y(n_187) );
INVx3_ASAP7_75t_L g188 ( .A(n_165), .Y(n_188) );
INVx4_ASAP7_75t_L g189 ( .A(n_144), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_168), .Y(n_190) );
INVxp67_ASAP7_75t_L g191 ( .A(n_155), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_168), .Y(n_192) );
INVx3_ASAP7_75t_L g193 ( .A(n_165), .Y(n_193) );
BUFx3_ASAP7_75t_L g194 ( .A(n_140), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_155), .B(n_116), .Y(n_195) );
INVx4_ASAP7_75t_L g196 ( .A(n_144), .Y(n_196) );
OAI22xp33_ASAP7_75t_L g197 ( .A1(n_129), .A2(n_121), .B1(n_117), .B2(n_127), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_137), .Y(n_198) );
BUFx6f_ASAP7_75t_L g199 ( .A(n_147), .Y(n_199) );
INVx5_ASAP7_75t_L g200 ( .A(n_140), .Y(n_200) );
NAND2xp5_ASAP7_75t_SL g201 ( .A(n_138), .B(n_118), .Y(n_201) );
OAI22xp5_ASAP7_75t_L g202 ( .A1(n_169), .A2(n_128), .B1(n_124), .B2(n_123), .Y(n_202) );
AND2x2_ASAP7_75t_L g203 ( .A(n_159), .B(n_101), .Y(n_203) );
INVx4_ASAP7_75t_L g204 ( .A(n_144), .Y(n_204) );
INVx4_ASAP7_75t_L g205 ( .A(n_144), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g206 ( .A(n_138), .B(n_128), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_147), .Y(n_207) );
AND2x4_ASAP7_75t_L g208 ( .A(n_139), .B(n_124), .Y(n_208) );
BUFx3_ASAP7_75t_L g209 ( .A(n_140), .Y(n_209) );
INVx4_ASAP7_75t_L g210 ( .A(n_144), .Y(n_210) );
OR2x2_ASAP7_75t_SL g211 ( .A(n_156), .B(n_123), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_139), .Y(n_212) );
OAI22xp33_ASAP7_75t_L g213 ( .A1(n_129), .A2(n_120), .B1(n_113), .B2(n_112), .Y(n_213) );
BUFx2_ASAP7_75t_L g214 ( .A(n_167), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_141), .Y(n_215) );
AOI22xp5_ASAP7_75t_L g216 ( .A1(n_149), .A2(n_79), .B1(n_83), .B2(n_85), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_141), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_151), .B(n_120), .Y(n_218) );
AND2x4_ASAP7_75t_L g219 ( .A(n_173), .B(n_113), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_151), .Y(n_220) );
INVx6_ASAP7_75t_L g221 ( .A(n_140), .Y(n_221) );
HB1xp67_ASAP7_75t_L g222 ( .A(n_149), .Y(n_222) );
AND2x4_ASAP7_75t_L g223 ( .A(n_173), .B(n_112), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_152), .B(n_109), .Y(n_224) );
INVx3_ASAP7_75t_L g225 ( .A(n_165), .Y(n_225) );
AOI22x1_ASAP7_75t_L g226 ( .A1(n_135), .A2(n_109), .B1(n_94), .B2(n_95), .Y(n_226) );
BUFx6f_ASAP7_75t_L g227 ( .A(n_147), .Y(n_227) );
OAI22xp33_ASAP7_75t_L g228 ( .A1(n_132), .A2(n_102), .B1(n_97), .B2(n_95), .Y(n_228) );
INVx1_ASAP7_75t_SL g229 ( .A(n_160), .Y(n_229) );
BUFx2_ASAP7_75t_L g230 ( .A(n_164), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_152), .B(n_102), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_162), .Y(n_232) );
NAND2x1p5_ASAP7_75t_L g233 ( .A(n_148), .B(n_97), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_162), .Y(n_234) );
BUFx3_ASAP7_75t_L g235 ( .A(n_140), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_163), .Y(n_236) );
AND2x2_ASAP7_75t_L g237 ( .A(n_131), .B(n_103), .Y(n_237) );
AND2x2_ASAP7_75t_L g238 ( .A(n_163), .B(n_92), .Y(n_238) );
INVx1_ASAP7_75t_SL g239 ( .A(n_134), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_165), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_171), .Y(n_241) );
BUFx2_ASAP7_75t_L g242 ( .A(n_187), .Y(n_242) );
CKINVDCx5p33_ASAP7_75t_R g243 ( .A(n_229), .Y(n_243) );
CKINVDCx5p33_ASAP7_75t_R g244 ( .A(n_214), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_240), .Y(n_245) );
INVxp67_ASAP7_75t_SL g246 ( .A(n_191), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_239), .B(n_134), .Y(n_247) );
NAND3xp33_ASAP7_75t_SL g248 ( .A(n_186), .B(n_157), .C(n_146), .Y(n_248) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_195), .B(n_157), .Y(n_249) );
INVx2_ASAP7_75t_L g250 ( .A(n_177), .Y(n_250) );
OR2x6_ASAP7_75t_L g251 ( .A(n_179), .B(n_144), .Y(n_251) );
NOR2xp33_ASAP7_75t_R g252 ( .A(n_184), .B(n_133), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_177), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_207), .Y(n_254) );
INVx2_ASAP7_75t_L g255 ( .A(n_207), .Y(n_255) );
AND2x2_ASAP7_75t_L g256 ( .A(n_222), .B(n_136), .Y(n_256) );
NOR3xp33_ASAP7_75t_SL g257 ( .A(n_184), .B(n_136), .C(n_146), .Y(n_257) );
CKINVDCx5p33_ASAP7_75t_R g258 ( .A(n_230), .Y(n_258) );
INVx2_ASAP7_75t_L g259 ( .A(n_199), .Y(n_259) );
INVx2_ASAP7_75t_SL g260 ( .A(n_185), .Y(n_260) );
BUFx5_ASAP7_75t_L g261 ( .A(n_178), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_174), .B(n_131), .Y(n_262) );
AND2x2_ASAP7_75t_L g263 ( .A(n_185), .B(n_131), .Y(n_263) );
INVx3_ASAP7_75t_L g264 ( .A(n_188), .Y(n_264) );
NAND2xp5_ASAP7_75t_SL g265 ( .A(n_185), .B(n_135), .Y(n_265) );
NOR2xp33_ASAP7_75t_L g266 ( .A(n_190), .B(n_93), .Y(n_266) );
INVx2_ASAP7_75t_L g267 ( .A(n_199), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_241), .Y(n_268) );
HB1xp67_ASAP7_75t_L g269 ( .A(n_203), .Y(n_269) );
INVx3_ASAP7_75t_L g270 ( .A(n_188), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_199), .Y(n_271) );
AND3x1_ASAP7_75t_SL g272 ( .A(n_192), .B(n_5), .C(n_6), .Y(n_272) );
BUFx2_ASAP7_75t_L g273 ( .A(n_179), .Y(n_273) );
BUFx6f_ASAP7_75t_L g274 ( .A(n_199), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_174), .B(n_131), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_238), .B(n_133), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_238), .B(n_133), .Y(n_277) );
BUFx3_ASAP7_75t_L g278 ( .A(n_194), .Y(n_278) );
NOR2xp33_ASAP7_75t_R g279 ( .A(n_189), .B(n_133), .Y(n_279) );
OR2x6_ASAP7_75t_L g280 ( .A(n_189), .B(n_172), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_188), .Y(n_281) );
INVx4_ASAP7_75t_L g282 ( .A(n_189), .Y(n_282) );
BUFx2_ASAP7_75t_L g283 ( .A(n_196), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_193), .Y(n_284) );
AOI22xp5_ASAP7_75t_L g285 ( .A1(n_197), .A2(n_172), .B1(n_171), .B2(n_166), .Y(n_285) );
INVxp33_ASAP7_75t_L g286 ( .A(n_182), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_227), .Y(n_287) );
NOR2xp33_ASAP7_75t_R g288 ( .A(n_196), .B(n_172), .Y(n_288) );
AOI21xp5_ASAP7_75t_L g289 ( .A1(n_176), .A2(n_130), .B(n_166), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_193), .Y(n_290) );
AO22x1_ASAP7_75t_L g291 ( .A1(n_196), .A2(n_153), .B1(n_143), .B2(n_166), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_193), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_227), .Y(n_293) );
NOR2xp33_ASAP7_75t_L g294 ( .A(n_216), .B(n_175), .Y(n_294) );
INVx3_ASAP7_75t_L g295 ( .A(n_225), .Y(n_295) );
AND2x4_ASAP7_75t_L g296 ( .A(n_175), .B(n_172), .Y(n_296) );
HB1xp67_ASAP7_75t_L g297 ( .A(n_175), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_181), .B(n_171), .Y(n_298) );
INVxp67_ASAP7_75t_L g299 ( .A(n_202), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_225), .Y(n_300) );
INVx3_ASAP7_75t_L g301 ( .A(n_225), .Y(n_301) );
OR2x2_ASAP7_75t_L g302 ( .A(n_211), .B(n_171), .Y(n_302) );
INVx2_ASAP7_75t_SL g303 ( .A(n_208), .Y(n_303) );
INVxp67_ASAP7_75t_SL g304 ( .A(n_183), .Y(n_304) );
NOR3xp33_ASAP7_75t_SL g305 ( .A(n_228), .B(n_108), .C(n_7), .Y(n_305) );
BUFx4_ASAP7_75t_SL g306 ( .A(n_198), .Y(n_306) );
NOR2xp67_ASAP7_75t_L g307 ( .A(n_181), .B(n_161), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_183), .Y(n_308) );
NAND2xp5_ASAP7_75t_SL g309 ( .A(n_181), .B(n_153), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_208), .Y(n_310) );
AND2x2_ASAP7_75t_L g311 ( .A(n_208), .B(n_161), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_212), .Y(n_312) );
OR2x6_ASAP7_75t_L g313 ( .A(n_251), .B(n_204), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_245), .Y(n_314) );
INVx5_ASAP7_75t_L g315 ( .A(n_280), .Y(n_315) );
NAND2xp33_ASAP7_75t_L g316 ( .A(n_279), .B(n_215), .Y(n_316) );
OAI22xp33_ASAP7_75t_L g317 ( .A1(n_243), .A2(n_210), .B1(n_204), .B2(n_205), .Y(n_317) );
BUFx2_ASAP7_75t_L g318 ( .A(n_242), .Y(n_318) );
AND2x4_ASAP7_75t_L g319 ( .A(n_260), .B(n_204), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_312), .Y(n_320) );
NOR2x1p5_ASAP7_75t_L g321 ( .A(n_243), .B(n_244), .Y(n_321) );
AOI22xp33_ASAP7_75t_L g322 ( .A1(n_251), .A2(n_210), .B1(n_205), .B2(n_213), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_312), .Y(n_323) );
BUFx12f_ASAP7_75t_L g324 ( .A(n_244), .Y(n_324) );
INVx5_ASAP7_75t_L g325 ( .A(n_280), .Y(n_325) );
BUFx4_ASAP7_75t_SL g326 ( .A(n_258), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_256), .B(n_219), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_245), .Y(n_328) );
CKINVDCx16_ASAP7_75t_R g329 ( .A(n_252), .Y(n_329) );
BUFx2_ASAP7_75t_L g330 ( .A(n_242), .Y(n_330) );
AND2x2_ASAP7_75t_L g331 ( .A(n_256), .B(n_219), .Y(n_331) );
AOI22xp33_ASAP7_75t_L g332 ( .A1(n_251), .A2(n_210), .B1(n_205), .B2(n_219), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_268), .Y(n_333) );
INVxp67_ASAP7_75t_L g334 ( .A(n_247), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_249), .B(n_223), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g336 ( .A(n_286), .B(n_233), .Y(n_336) );
INVx2_ASAP7_75t_SL g337 ( .A(n_303), .Y(n_337) );
BUFx3_ASAP7_75t_L g338 ( .A(n_278), .Y(n_338) );
BUFx3_ASAP7_75t_L g339 ( .A(n_278), .Y(n_339) );
INVx2_ASAP7_75t_SL g340 ( .A(n_303), .Y(n_340) );
NOR2xp33_ASAP7_75t_L g341 ( .A(n_246), .B(n_294), .Y(n_341) );
AOI22xp33_ASAP7_75t_L g342 ( .A1(n_251), .A2(n_223), .B1(n_180), .B2(n_176), .Y(n_342) );
BUFx3_ASAP7_75t_L g343 ( .A(n_280), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_260), .B(n_223), .Y(n_344) );
AOI21xp5_ASAP7_75t_L g345 ( .A1(n_304), .A2(n_180), .B(n_237), .Y(n_345) );
BUFx6f_ASAP7_75t_L g346 ( .A(n_280), .Y(n_346) );
AND2x4_ASAP7_75t_L g347 ( .A(n_273), .B(n_236), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_268), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_273), .B(n_220), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_310), .Y(n_350) );
BUFx3_ASAP7_75t_L g351 ( .A(n_283), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_281), .Y(n_352) );
BUFx6f_ASAP7_75t_L g353 ( .A(n_282), .Y(n_353) );
INVxp67_ASAP7_75t_SL g354 ( .A(n_297), .Y(n_354) );
BUFx3_ASAP7_75t_L g355 ( .A(n_283), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_296), .B(n_217), .Y(n_356) );
BUFx2_ASAP7_75t_L g357 ( .A(n_288), .Y(n_357) );
BUFx6f_ASAP7_75t_L g358 ( .A(n_282), .Y(n_358) );
NOR2x1_ASAP7_75t_L g359 ( .A(n_282), .B(n_231), .Y(n_359) );
AOI21xp33_ASAP7_75t_SL g360 ( .A1(n_258), .A2(n_233), .B(n_206), .Y(n_360) );
BUFx6f_ASAP7_75t_L g361 ( .A(n_274), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_296), .B(n_234), .Y(n_362) );
BUFx2_ASAP7_75t_L g363 ( .A(n_261), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_281), .Y(n_364) );
BUFx2_ASAP7_75t_L g365 ( .A(n_261), .Y(n_365) );
CKINVDCx5p33_ASAP7_75t_R g366 ( .A(n_306), .Y(n_366) );
INVx3_ASAP7_75t_L g367 ( .A(n_264), .Y(n_367) );
INVx3_ASAP7_75t_L g368 ( .A(n_264), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_320), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_334), .B(n_299), .Y(n_370) );
OAI22xp5_ASAP7_75t_L g371 ( .A1(n_313), .A2(n_307), .B1(n_296), .B2(n_311), .Y(n_371) );
AND2x4_ASAP7_75t_L g372 ( .A(n_315), .B(n_257), .Y(n_372) );
OAI22xp33_ASAP7_75t_L g373 ( .A1(n_313), .A2(n_302), .B1(n_285), .B2(n_248), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_327), .B(n_269), .Y(n_374) );
AOI22xp33_ASAP7_75t_L g375 ( .A1(n_341), .A2(n_263), .B1(n_266), .B2(n_265), .Y(n_375) );
OAI22xp5_ASAP7_75t_L g376 ( .A1(n_313), .A2(n_311), .B1(n_298), .B2(n_263), .Y(n_376) );
OR2x6_ASAP7_75t_L g377 ( .A(n_313), .B(n_291), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_327), .B(n_309), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_320), .Y(n_379) );
INVx4_ASAP7_75t_L g380 ( .A(n_315), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_320), .Y(n_381) );
AOI21xp5_ASAP7_75t_L g382 ( .A1(n_345), .A2(n_262), .B(n_275), .Y(n_382) );
BUFx2_ASAP7_75t_L g383 ( .A(n_318), .Y(n_383) );
AO221x2_ASAP7_75t_L g384 ( .A1(n_317), .A2(n_291), .B1(n_272), .B2(n_305), .C(n_153), .Y(n_384) );
AND2x4_ASAP7_75t_L g385 ( .A(n_315), .B(n_325), .Y(n_385) );
OAI22xp5_ASAP7_75t_L g386 ( .A1(n_313), .A2(n_308), .B1(n_302), .B2(n_276), .Y(n_386) );
AOI22xp5_ASAP7_75t_L g387 ( .A1(n_318), .A2(n_261), .B1(n_301), .B2(n_270), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_349), .Y(n_388) );
INVx4_ASAP7_75t_L g389 ( .A(n_315), .Y(n_389) );
NOR2xp33_ASAP7_75t_L g390 ( .A(n_331), .B(n_264), .Y(n_390) );
OR2x6_ASAP7_75t_L g391 ( .A(n_324), .B(n_277), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_323), .Y(n_392) );
AOI22xp33_ASAP7_75t_L g393 ( .A1(n_335), .A2(n_226), .B1(n_231), .B2(n_224), .Y(n_393) );
OAI22xp5_ASAP7_75t_L g394 ( .A1(n_322), .A2(n_308), .B1(n_232), .B2(n_301), .Y(n_394) );
OAI22xp5_ASAP7_75t_L g395 ( .A1(n_332), .A2(n_301), .B1(n_270), .B2(n_295), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_349), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_331), .Y(n_397) );
CKINVDCx8_ASAP7_75t_R g398 ( .A(n_366), .Y(n_398) );
OAI22xp33_ASAP7_75t_SL g399 ( .A1(n_329), .A2(n_330), .B1(n_325), .B2(n_315), .Y(n_399) );
CKINVDCx6p67_ASAP7_75t_R g400 ( .A(n_324), .Y(n_400) );
OA21x2_ASAP7_75t_L g401 ( .A1(n_314), .A2(n_289), .B(n_142), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g402 ( .A1(n_335), .A2(n_224), .B1(n_206), .B2(n_218), .Y(n_402) );
NOR2x1p5_ASAP7_75t_L g403 ( .A(n_400), .B(n_343), .Y(n_403) );
BUFx2_ASAP7_75t_L g404 ( .A(n_377), .Y(n_404) );
OAI211xp5_ASAP7_75t_L g405 ( .A1(n_370), .A2(n_360), .B(n_330), .C(n_336), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_369), .B(n_323), .Y(n_406) );
OA21x2_ASAP7_75t_L g407 ( .A1(n_382), .A2(n_314), .B(n_328), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_388), .B(n_347), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_369), .Y(n_409) );
AND2x4_ASAP7_75t_L g410 ( .A(n_385), .B(n_315), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g411 ( .A1(n_384), .A2(n_321), .B1(n_347), .B2(n_343), .Y(n_411) );
AOI22xp33_ASAP7_75t_SL g412 ( .A1(n_384), .A2(n_329), .B1(n_343), .B2(n_325), .Y(n_412) );
OAI22xp5_ASAP7_75t_SL g413 ( .A1(n_391), .A2(n_342), .B1(n_325), .B2(n_347), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_396), .B(n_347), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_379), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_384), .A2(n_321), .B1(n_328), .B2(n_348), .Y(n_416) );
AO31x2_ASAP7_75t_L g417 ( .A1(n_379), .A2(n_348), .A3(n_333), .B(n_323), .Y(n_417) );
OAI22xp5_ASAP7_75t_L g418 ( .A1(n_377), .A2(n_325), .B1(n_351), .B2(n_355), .Y(n_418) );
OAI221xp5_ASAP7_75t_L g419 ( .A1(n_375), .A2(n_360), .B1(n_354), .B2(n_344), .C(n_218), .Y(n_419) );
AOI21xp33_ASAP7_75t_L g420 ( .A1(n_373), .A2(n_316), .B(n_357), .Y(n_420) );
AOI22xp33_ASAP7_75t_L g421 ( .A1(n_373), .A2(n_333), .B1(n_357), .B2(n_356), .Y(n_421) );
AOI22xp33_ASAP7_75t_L g422 ( .A1(n_386), .A2(n_362), .B1(n_356), .B2(n_346), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_381), .Y(n_423) );
OAI221xp5_ASAP7_75t_L g424 ( .A1(n_375), .A2(n_350), .B1(n_362), .B2(n_337), .C(n_340), .Y(n_424) );
OAI22xp5_ASAP7_75t_L g425 ( .A1(n_377), .A2(n_325), .B1(n_346), .B2(n_355), .Y(n_425) );
OAI22xp33_ASAP7_75t_L g426 ( .A1(n_391), .A2(n_346), .B1(n_351), .B2(n_355), .Y(n_426) );
AND2x4_ASAP7_75t_L g427 ( .A(n_385), .B(n_363), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_397), .B(n_350), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_381), .Y(n_429) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_372), .A2(n_346), .B1(n_351), .B2(n_319), .Y(n_430) );
AOI22xp33_ASAP7_75t_L g431 ( .A1(n_372), .A2(n_346), .B1(n_319), .B2(n_340), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_417), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_406), .B(n_392), .Y(n_433) );
NOR2xp33_ASAP7_75t_SL g434 ( .A(n_425), .B(n_380), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_417), .Y(n_435) );
AND2x6_ASAP7_75t_SL g436 ( .A(n_410), .B(n_391), .Y(n_436) );
INVx1_ASAP7_75t_SL g437 ( .A(n_406), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_409), .B(n_392), .Y(n_438) );
OR2x2_ASAP7_75t_L g439 ( .A(n_417), .B(n_409), .Y(n_439) );
AO21x2_ASAP7_75t_L g440 ( .A1(n_420), .A2(n_394), .B(n_371), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_417), .Y(n_441) );
AOI221xp5_ASAP7_75t_L g442 ( .A1(n_419), .A2(n_374), .B1(n_383), .B2(n_402), .C(n_378), .Y(n_442) );
NOR2x2_ASAP7_75t_L g443 ( .A(n_403), .B(n_326), .Y(n_443) );
AO21x2_ASAP7_75t_L g444 ( .A1(n_425), .A2(n_376), .B(n_130), .Y(n_444) );
AND2x4_ASAP7_75t_L g445 ( .A(n_417), .B(n_380), .Y(n_445) );
OR2x2_ASAP7_75t_L g446 ( .A(n_417), .B(n_389), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_423), .Y(n_447) );
AOI221xp5_ASAP7_75t_L g448 ( .A1(n_405), .A2(n_402), .B1(n_390), .B2(n_399), .C(n_372), .Y(n_448) );
AOI33xp33_ASAP7_75t_L g449 ( .A1(n_416), .A2(n_161), .A3(n_143), .B1(n_142), .B2(n_130), .B3(n_393), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_415), .Y(n_450) );
INVx4_ASAP7_75t_SL g451 ( .A(n_413), .Y(n_451) );
OAI21xp5_ASAP7_75t_L g452 ( .A1(n_421), .A2(n_393), .B(n_390), .Y(n_452) );
AO221x2_ASAP7_75t_L g453 ( .A1(n_413), .A2(n_395), .B1(n_8), .B2(n_9), .C(n_10), .Y(n_453) );
CKINVDCx5p33_ASAP7_75t_R g454 ( .A(n_403), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_415), .B(n_389), .Y(n_455) );
HB1xp67_ASAP7_75t_L g456 ( .A(n_415), .Y(n_456) );
AO21x2_ASAP7_75t_L g457 ( .A1(n_429), .A2(n_143), .B(n_142), .Y(n_457) );
NAND2xp33_ASAP7_75t_R g458 ( .A(n_404), .B(n_401), .Y(n_458) );
AOI22xp33_ASAP7_75t_L g459 ( .A1(n_404), .A2(n_346), .B1(n_319), .B2(n_368), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_424), .A2(n_319), .B1(n_368), .B2(n_367), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_429), .B(n_401), .Y(n_461) );
AOI211xp5_ASAP7_75t_L g462 ( .A1(n_426), .A2(n_387), .B(n_201), .C(n_353), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_429), .B(n_401), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_427), .B(n_352), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_408), .B(n_352), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_428), .B(n_364), .Y(n_466) );
BUFx2_ASAP7_75t_L g467 ( .A(n_418), .Y(n_467) );
OAI221xp5_ASAP7_75t_L g468 ( .A1(n_411), .A2(n_398), .B1(n_337), .B2(n_359), .C(n_367), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_447), .Y(n_469) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_454), .B(n_414), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_437), .B(n_407), .Y(n_471) );
AOI22xp33_ASAP7_75t_L g472 ( .A1(n_453), .A2(n_422), .B1(n_412), .B2(n_427), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_450), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_433), .B(n_427), .Y(n_474) );
OR2x2_ASAP7_75t_L g475 ( .A(n_439), .B(n_407), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_447), .Y(n_476) );
INVxp67_ASAP7_75t_SL g477 ( .A(n_456), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_437), .B(n_407), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_433), .B(n_427), .Y(n_479) );
OR2x2_ASAP7_75t_L g480 ( .A(n_439), .B(n_407), .Y(n_480) );
OR2x2_ASAP7_75t_L g481 ( .A(n_446), .B(n_410), .Y(n_481) );
AND2x4_ASAP7_75t_L g482 ( .A(n_445), .B(n_410), .Y(n_482) );
BUFx3_ASAP7_75t_L g483 ( .A(n_455), .Y(n_483) );
NAND3xp33_ASAP7_75t_L g484 ( .A(n_453), .B(n_147), .C(n_431), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_445), .B(n_430), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_445), .B(n_5), .Y(n_486) );
INVx4_ASAP7_75t_L g487 ( .A(n_436), .Y(n_487) );
INVx2_ASAP7_75t_SL g488 ( .A(n_445), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_438), .B(n_364), .Y(n_489) );
OR2x2_ASAP7_75t_L g490 ( .A(n_432), .B(n_201), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_450), .Y(n_491) );
INVxp67_ASAP7_75t_SL g492 ( .A(n_450), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_435), .Y(n_493) );
OAI221xp5_ASAP7_75t_L g494 ( .A1(n_448), .A2(n_359), .B1(n_290), .B2(n_292), .C(n_284), .Y(n_494) );
OR2x2_ASAP7_75t_L g495 ( .A(n_441), .B(n_10), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_461), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_441), .B(n_11), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_455), .B(n_12), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_464), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_461), .B(n_13), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_464), .Y(n_501) );
OR2x2_ASAP7_75t_L g502 ( .A(n_467), .B(n_14), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_463), .B(n_14), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_463), .B(n_15), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_466), .Y(n_505) );
INVx1_ASAP7_75t_SL g506 ( .A(n_443), .Y(n_506) );
OR2x2_ASAP7_75t_L g507 ( .A(n_467), .B(n_16), .Y(n_507) );
OR2x2_ASAP7_75t_L g508 ( .A(n_444), .B(n_453), .Y(n_508) );
OAI33xp33_ASAP7_75t_L g509 ( .A1(n_466), .A2(n_16), .A3(n_17), .B1(n_18), .B2(n_19), .B3(n_284), .Y(n_509) );
INVx4_ASAP7_75t_L g510 ( .A(n_436), .Y(n_510) );
AND2x4_ASAP7_75t_L g511 ( .A(n_451), .B(n_68), .Y(n_511) );
INVx2_ASAP7_75t_SL g512 ( .A(n_453), .Y(n_512) );
INVxp67_ASAP7_75t_L g513 ( .A(n_458), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_457), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_451), .B(n_17), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_457), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_452), .A2(n_338), .B1(n_339), .B2(n_368), .Y(n_517) );
OR2x6_ASAP7_75t_L g518 ( .A(n_487), .B(n_451), .Y(n_518) );
INVxp67_ASAP7_75t_SL g519 ( .A(n_492), .Y(n_519) );
NOR3xp33_ASAP7_75t_L g520 ( .A(n_509), .B(n_468), .C(n_442), .Y(n_520) );
INVxp67_ASAP7_75t_L g521 ( .A(n_477), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_505), .B(n_452), .Y(n_522) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_502), .B(n_444), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_469), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_483), .B(n_451), .Y(n_525) );
OR2x2_ASAP7_75t_L g526 ( .A(n_481), .B(n_444), .Y(n_526) );
NAND2xp33_ASAP7_75t_R g527 ( .A(n_511), .B(n_451), .Y(n_527) );
NOR2xp33_ASAP7_75t_R g528 ( .A(n_506), .B(n_434), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_500), .B(n_444), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_476), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_500), .B(n_462), .Y(n_531) );
INVx1_ASAP7_75t_SL g532 ( .A(n_483), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_503), .B(n_462), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_473), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_503), .B(n_449), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_486), .B(n_434), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_486), .B(n_440), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_493), .Y(n_538) );
HB1xp67_ASAP7_75t_L g539 ( .A(n_473), .Y(n_539) );
INVxp67_ASAP7_75t_L g540 ( .A(n_475), .Y(n_540) );
INVx2_ASAP7_75t_L g541 ( .A(n_491), .Y(n_541) );
NOR4xp75_ASAP7_75t_L g542 ( .A(n_512), .B(n_465), .C(n_368), .D(n_367), .Y(n_542) );
OAI22xp5_ASAP7_75t_SL g543 ( .A1(n_487), .A2(n_460), .B1(n_459), .B2(n_353), .Y(n_543) );
AND2x4_ASAP7_75t_L g544 ( .A(n_488), .B(n_457), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_495), .Y(n_545) );
AND2x4_ASAP7_75t_SL g546 ( .A(n_487), .B(n_353), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_499), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_504), .B(n_440), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_504), .B(n_440), .Y(n_549) );
NOR2xp67_ASAP7_75t_L g550 ( .A(n_510), .B(n_147), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_501), .Y(n_551) );
NAND4xp75_ASAP7_75t_L g552 ( .A(n_515), .B(n_292), .C(n_300), .D(n_39), .Y(n_552) );
OR2x2_ASAP7_75t_L g553 ( .A(n_496), .B(n_457), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_498), .B(n_147), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_482), .B(n_353), .Y(n_555) );
NAND2xp33_ASAP7_75t_SL g556 ( .A(n_510), .B(n_353), .Y(n_556) );
AND2x4_ASAP7_75t_L g557 ( .A(n_488), .B(n_21), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_497), .Y(n_558) );
NAND4xp25_ASAP7_75t_L g559 ( .A(n_472), .B(n_300), .C(n_270), .D(n_295), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g560 ( .A(n_502), .B(n_35), .Y(n_560) );
INVx2_ASAP7_75t_L g561 ( .A(n_491), .Y(n_561) );
HB1xp67_ASAP7_75t_L g562 ( .A(n_475), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_507), .B(n_358), .Y(n_563) );
NOR2x1_ASAP7_75t_L g564 ( .A(n_510), .B(n_339), .Y(n_564) );
AOI32xp33_ASAP7_75t_L g565 ( .A1(n_515), .A2(n_365), .A3(n_363), .B1(n_295), .B2(n_338), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_482), .B(n_358), .Y(n_566) );
INVx1_ASAP7_75t_SL g567 ( .A(n_482), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_507), .Y(n_568) );
AOI221xp5_ASAP7_75t_L g569 ( .A1(n_568), .A2(n_512), .B1(n_484), .B2(n_513), .C(n_470), .Y(n_569) );
INVx2_ASAP7_75t_L g570 ( .A(n_539), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_547), .B(n_471), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_551), .B(n_471), .Y(n_572) );
AOI22xp33_ASAP7_75t_SL g573 ( .A1(n_528), .A2(n_511), .B1(n_508), .B2(n_485), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_524), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_530), .Y(n_575) );
INVx2_ASAP7_75t_SL g576 ( .A(n_532), .Y(n_576) );
OAI31xp33_ASAP7_75t_L g577 ( .A1(n_559), .A2(n_508), .A3(n_485), .B(n_480), .Y(n_577) );
AOI21xp5_ASAP7_75t_L g578 ( .A1(n_556), .A2(n_516), .B(n_514), .Y(n_578) );
NOR2xp67_ASAP7_75t_L g579 ( .A(n_562), .B(n_480), .Y(n_579) );
OAI22xp5_ASAP7_75t_L g580 ( .A1(n_518), .A2(n_474), .B1(n_479), .B2(n_489), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_538), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_540), .B(n_478), .Y(n_582) );
AOI22xp33_ASAP7_75t_SL g583 ( .A1(n_528), .A2(n_478), .B1(n_490), .B2(n_494), .Y(n_583) );
OAI32xp33_ASAP7_75t_L g584 ( .A1(n_527), .A2(n_490), .A3(n_517), .B1(n_339), .B2(n_338), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_567), .B(n_40), .Y(n_585) );
OR4x1_ASAP7_75t_L g586 ( .A(n_558), .B(n_45), .C(n_46), .D(n_47), .Y(n_586) );
AOI21xp33_ASAP7_75t_SL g587 ( .A1(n_527), .A2(n_50), .B(n_51), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_540), .B(n_53), .Y(n_588) );
INVxp67_ASAP7_75t_SL g589 ( .A(n_519), .Y(n_589) );
NAND3xp33_ASAP7_75t_L g590 ( .A(n_520), .B(n_358), .C(n_274), .Y(n_590) );
OAI22xp5_ASAP7_75t_L g591 ( .A1(n_531), .A2(n_358), .B1(n_221), .B2(n_361), .Y(n_591) );
OAI22xp33_ASAP7_75t_L g592 ( .A1(n_518), .A2(n_358), .B1(n_361), .B2(n_221), .Y(n_592) );
AOI22xp5_ASAP7_75t_L g593 ( .A1(n_533), .A2(n_261), .B1(n_221), .B2(n_361), .Y(n_593) );
INVx3_ASAP7_75t_SL g594 ( .A(n_546), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_562), .B(n_55), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_521), .Y(n_596) );
OAI22xp5_ASAP7_75t_L g597 ( .A1(n_560), .A2(n_361), .B1(n_200), .B2(n_274), .Y(n_597) );
INVx2_ASAP7_75t_L g598 ( .A(n_521), .Y(n_598) );
AND2x4_ASAP7_75t_L g599 ( .A(n_525), .B(n_57), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_519), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_536), .B(n_60), .Y(n_601) );
NAND2x1p5_ASAP7_75t_L g602 ( .A(n_557), .B(n_361), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_545), .Y(n_603) );
NAND2x1_ASAP7_75t_L g604 ( .A(n_557), .B(n_361), .Y(n_604) );
INVx2_ASAP7_75t_L g605 ( .A(n_534), .Y(n_605) );
AND2x4_ASAP7_75t_L g606 ( .A(n_546), .B(n_61), .Y(n_606) );
AOI32xp33_ASAP7_75t_L g607 ( .A1(n_560), .A2(n_209), .A3(n_235), .B1(n_194), .B2(n_73), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_526), .Y(n_608) );
A2O1A1Ixp33_ASAP7_75t_L g609 ( .A1(n_550), .A2(n_209), .B(n_235), .C(n_72), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_534), .Y(n_610) );
OAI21xp33_ASAP7_75t_L g611 ( .A1(n_523), .A2(n_259), .B(n_293), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_574), .Y(n_612) );
INVx1_ASAP7_75t_SL g613 ( .A(n_594), .Y(n_613) );
NOR2xp33_ASAP7_75t_L g614 ( .A(n_596), .B(n_522), .Y(n_614) );
OR2x2_ASAP7_75t_L g615 ( .A(n_582), .B(n_529), .Y(n_615) );
AOI22xp5_ASAP7_75t_L g616 ( .A1(n_580), .A2(n_523), .B1(n_543), .B2(n_537), .Y(n_616) );
NOR3xp33_ASAP7_75t_SL g617 ( .A(n_590), .B(n_552), .C(n_535), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_575), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_581), .Y(n_619) );
NAND4xp75_ASAP7_75t_L g620 ( .A(n_577), .B(n_564), .C(n_548), .D(n_549), .Y(n_620) );
NOR2xp33_ASAP7_75t_L g621 ( .A(n_603), .B(n_554), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_608), .B(n_563), .Y(n_622) );
INVxp67_ASAP7_75t_L g623 ( .A(n_589), .Y(n_623) );
AND2x2_ASAP7_75t_L g624 ( .A(n_576), .B(n_544), .Y(n_624) );
XNOR2x2_ASAP7_75t_L g625 ( .A(n_569), .B(n_542), .Y(n_625) );
INVx2_ASAP7_75t_L g626 ( .A(n_605), .Y(n_626) );
INVx2_ASAP7_75t_L g627 ( .A(n_610), .Y(n_627) );
BUFx2_ASAP7_75t_L g628 ( .A(n_598), .Y(n_628) );
AND2x4_ASAP7_75t_L g629 ( .A(n_579), .B(n_561), .Y(n_629) );
AND2x2_ASAP7_75t_SL g630 ( .A(n_606), .B(n_541), .Y(n_630) );
XNOR2xp5_ASAP7_75t_L g631 ( .A(n_573), .B(n_566), .Y(n_631) );
XNOR2x1_ASAP7_75t_SL g632 ( .A(n_602), .B(n_555), .Y(n_632) );
AND2x2_ASAP7_75t_L g633 ( .A(n_571), .B(n_553), .Y(n_633) );
OAI211xp5_ASAP7_75t_L g634 ( .A1(n_577), .A2(n_565), .B(n_200), .C(n_293), .Y(n_634) );
INVx1_ASAP7_75t_SL g635 ( .A(n_606), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_572), .B(n_67), .Y(n_636) );
INVx2_ASAP7_75t_SL g637 ( .A(n_570), .Y(n_637) );
NAND2xp5_ASAP7_75t_SL g638 ( .A(n_613), .B(n_587), .Y(n_638) );
AOI221x1_ASAP7_75t_SL g639 ( .A1(n_612), .A2(n_600), .B1(n_611), .B2(n_599), .C(n_591), .Y(n_639) );
OAI21x1_ASAP7_75t_SL g640 ( .A1(n_632), .A2(n_625), .B(n_631), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_618), .Y(n_641) );
AOI221x1_ASAP7_75t_L g642 ( .A1(n_619), .A2(n_611), .B1(n_591), .B2(n_595), .C(n_588), .Y(n_642) );
OAI22xp33_ASAP7_75t_L g643 ( .A1(n_616), .A2(n_604), .B1(n_602), .B2(n_592), .Y(n_643) );
AOI22xp5_ASAP7_75t_L g644 ( .A1(n_620), .A2(n_583), .B1(n_601), .B2(n_599), .Y(n_644) );
AOI211x1_ASAP7_75t_L g645 ( .A1(n_634), .A2(n_584), .B(n_578), .C(n_585), .Y(n_645) );
XNOR2xp5_ASAP7_75t_L g646 ( .A(n_625), .B(n_593), .Y(n_646) );
AOI22xp5_ASAP7_75t_L g647 ( .A1(n_635), .A2(n_614), .B1(n_621), .B2(n_624), .Y(n_647) );
OAI211xp5_ASAP7_75t_L g648 ( .A1(n_623), .A2(n_607), .B(n_593), .C(n_609), .Y(n_648) );
INVxp67_ASAP7_75t_L g649 ( .A(n_628), .Y(n_649) );
INVxp67_ASAP7_75t_L g650 ( .A(n_614), .Y(n_650) );
OAI21xp5_ASAP7_75t_L g651 ( .A1(n_623), .A2(n_597), .B(n_586), .Y(n_651) );
OAI22xp33_ASAP7_75t_L g652 ( .A1(n_615), .A2(n_200), .B1(n_274), .B2(n_287), .Y(n_652) );
AOI321xp33_ASAP7_75t_SL g653 ( .A1(n_621), .A2(n_261), .A3(n_200), .B1(n_253), .B2(n_254), .C(n_255), .Y(n_653) );
INVxp67_ASAP7_75t_L g654 ( .A(n_640), .Y(n_654) );
AOI221xp5_ASAP7_75t_L g655 ( .A1(n_639), .A2(n_637), .B1(n_622), .B2(n_633), .C(n_629), .Y(n_655) );
OA22x2_ASAP7_75t_L g656 ( .A1(n_644), .A2(n_627), .B1(n_636), .B2(n_626), .Y(n_656) );
CKINVDCx16_ASAP7_75t_R g657 ( .A(n_647), .Y(n_657) );
NOR2x1p5_ASAP7_75t_L g658 ( .A(n_645), .B(n_630), .Y(n_658) );
AOI22xp5_ASAP7_75t_L g659 ( .A1(n_638), .A2(n_617), .B1(n_261), .B2(n_267), .Y(n_659) );
AOI211xp5_ASAP7_75t_L g660 ( .A1(n_648), .A2(n_271), .B(n_267), .C(n_253), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_641), .B(n_250), .Y(n_661) );
XNOR2x1_ASAP7_75t_L g662 ( .A(n_653), .B(n_652), .Y(n_662) );
AOI22xp5_ASAP7_75t_L g663 ( .A1(n_642), .A2(n_646), .B1(n_643), .B2(n_650), .Y(n_663) );
NOR5xp2_ASAP7_75t_L g664 ( .A(n_649), .B(n_640), .C(n_623), .D(n_634), .E(n_651), .Y(n_664) );
AOI21xp5_ASAP7_75t_L g665 ( .A1(n_640), .A2(n_638), .B(n_634), .Y(n_665) );
CKINVDCx5p33_ASAP7_75t_R g666 ( .A(n_654), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_663), .B(n_657), .Y(n_667) );
INVxp67_ASAP7_75t_SL g668 ( .A(n_664), .Y(n_668) );
AOI32xp33_ASAP7_75t_L g669 ( .A1(n_667), .A2(n_662), .A3(n_660), .B1(n_655), .B2(n_665), .Y(n_669) );
NOR3xp33_ASAP7_75t_L g670 ( .A(n_668), .B(n_659), .C(n_661), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_666), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_671), .Y(n_672) );
INVx2_ASAP7_75t_L g673 ( .A(n_670), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_672), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_673), .B(n_666), .Y(n_675) );
AOI22xp5_ASAP7_75t_L g676 ( .A1(n_675), .A2(n_673), .B1(n_658), .B2(n_656), .Y(n_676) );
AOI21xp5_ASAP7_75t_L g677 ( .A1(n_676), .A2(n_674), .B(n_669), .Y(n_677) );
endmodule