module fake_jpeg_7627_n_94 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_94);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_94;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_82;

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_28),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_19),
.B(n_26),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_30),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_7),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_13),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_33),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

NOR3xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_0),
.C(n_1),
.Y(n_49)
);

OA22x2_ASAP7_75t_L g60 ( 
.A1(n_49),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_47),
.B(n_2),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_50),
.B(n_56),
.Y(n_66)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_34),
.B(n_2),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_56),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_65),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_60),
.B(n_61),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_56),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_52),
.A2(n_40),
.B1(n_36),
.B2(n_35),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_63),
.A2(n_64),
.B1(n_67),
.B2(n_6),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_52),
.A2(n_43),
.B1(n_41),
.B2(n_38),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_52),
.A2(n_45),
.B1(n_9),
.B2(n_11),
.Y(n_67)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_71),
.Y(n_77)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_74),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_69),
.A2(n_12),
.B(n_14),
.Y(n_74)
);

A2O1A1Ixp33_ASAP7_75t_SL g76 ( 
.A1(n_60),
.A2(n_16),
.B(n_17),
.C(n_20),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_76),
.A2(n_79),
.B1(n_80),
.B2(n_58),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_66),
.B(n_21),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_82),
.B(n_75),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_83),
.B(n_73),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_84),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_85),
.A2(n_81),
.B1(n_78),
.B2(n_62),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_86),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_87),
.Y(n_88)
);

MAJx2_ASAP7_75t_L g89 ( 
.A(n_88),
.B(n_76),
.C(n_77),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_89),
.B(n_22),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_90),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_91),
.A2(n_23),
.B(n_24),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_92),
.B(n_25),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_27),
.Y(n_94)
);


endmodule