module real_jpeg_25610_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_126;
wire n_13;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_110;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_206;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_0),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_1),
.A2(n_38),
.B1(n_42),
.B2(n_45),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_1),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_1),
.A2(n_45),
.B1(n_59),
.B2(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_1),
.A2(n_45),
.B1(n_53),
.B2(n_54),
.Y(n_95)
);

O2A1O1Ixp33_ASAP7_75t_L g105 ( 
.A1(n_1),
.A2(n_57),
.B(n_106),
.C(n_107),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_1),
.B(n_52),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_1),
.A2(n_21),
.B1(n_23),
.B2(n_45),
.Y(n_127)
);

O2A1O1Ixp33_ASAP7_75t_L g135 ( 
.A1(n_1),
.A2(n_54),
.B(n_77),
.C(n_136),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_1),
.B(n_23),
.C(n_40),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_1),
.B(n_84),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_1),
.B(n_11),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_1),
.B(n_43),
.Y(n_184)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_4),
.A2(n_21),
.B1(n_23),
.B2(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_4),
.A2(n_33),
.B1(n_38),
.B2(n_42),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_4),
.A2(n_33),
.B1(n_53),
.B2(n_54),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_4),
.A2(n_33),
.B1(n_99),
.B2(n_100),
.Y(n_98)
);

BUFx10_ASAP7_75t_L g57 ( 
.A(n_5),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_6),
.A2(n_59),
.B1(n_60),
.B2(n_61),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_6),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_6),
.A2(n_53),
.B1(n_54),
.B2(n_61),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_6),
.A2(n_38),
.B1(n_42),
.B2(n_61),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_6),
.A2(n_21),
.B1(n_23),
.B2(n_61),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_7),
.A2(n_21),
.B1(n_23),
.B2(n_24),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_8),
.Y(n_78)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_9),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_11),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_129),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_128),
.Y(n_13)
);

OR2x2_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_114),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_15),
.B(n_114),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g15 ( 
.A1(n_16),
.A2(n_17),
.B1(n_88),
.B2(n_113),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_48),
.B1(n_86),
.B2(n_87),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_18),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_34),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_25),
.B(n_27),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_20),
.A2(n_109),
.B(n_112),
.Y(n_108)
);

CKINVDCx5p33_ASAP7_75t_R g23 ( 
.A(n_21),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_21),
.A2(n_23),
.B1(n_39),
.B2(n_40),
.Y(n_43)
);

INVx6_ASAP7_75t_SL g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_23),
.B(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_23),
.B(n_180),
.Y(n_179)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_25),
.B(n_32),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_25),
.B(n_127),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_25),
.A2(n_31),
.B(n_127),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_25),
.B(n_168),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_28),
.B(n_126),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_28),
.B(n_167),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_32),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_30),
.B(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_30),
.B(n_169),
.Y(n_174)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_46),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_35),
.B(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_36),
.B(n_44),
.Y(n_35)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_36),
.B(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_36),
.B(n_47),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_43),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_39),
.B1(n_40),
.B2(n_42),
.Y(n_37)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_38),
.A2(n_42),
.B1(n_77),
.B2(n_79),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_38),
.B(n_155),
.Y(n_154)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx24_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI21xp33_ASAP7_75t_L g136 ( 
.A1(n_42),
.A2(n_45),
.B(n_79),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_43),
.B(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_43),
.B(n_142),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_44),
.Y(n_72)
);

OAI21xp33_ASAP7_75t_L g106 ( 
.A1(n_45),
.A2(n_54),
.B(n_56),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_46),
.B(n_141),
.Y(n_160)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_68),
.C(n_73),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_49),
.A2(n_50),
.B1(n_117),
.B2(n_118),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_62),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_58),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_52),
.B(n_98),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_54),
.B1(n_56),
.B2(n_57),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_53),
.A2(n_54),
.B1(n_77),
.B2(n_79),
.Y(n_76)
);

INVx3_ASAP7_75t_SL g53 ( 
.A(n_54),
.Y(n_53)
);

CKINVDCx6p67_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_56),
.A2(n_57),
.B1(n_59),
.B2(n_60),
.Y(n_67)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_58),
.B(n_66),
.Y(n_101)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_59),
.Y(n_107)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_60),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_66),
.Y(n_62)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_68),
.A2(n_69),
.B1(n_73),
.B2(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_SL g69 ( 
.A1(n_70),
.A2(n_71),
.B(n_72),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_71),
.B(n_72),
.Y(n_139)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_73),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_74),
.B(n_82),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_81),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_75),
.B(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_75),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_80),
.Y(n_75)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_77),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_80),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_94),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_80),
.B(n_81),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_83),
.B(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_85),
.Y(n_83)
);

INVxp67_ASAP7_75t_SL g92 ( 
.A(n_85),
.Y(n_92)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_88),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_104),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_96),
.B1(n_102),
.B2(n_103),
.Y(n_89)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_90),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_91),
.B(n_93),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_91),
.B(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_95),
.B(n_195),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_96),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_101),
.Y(n_96)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_99),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_108),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_105),
.B(n_108),
.Y(n_120)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_112),
.B(n_174),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_120),
.C(n_121),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_115),
.A2(n_116),
.B1(n_144),
.B2(n_145),
.Y(n_143)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_120),
.B(n_121),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_124),
.C(n_125),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_122),
.B(n_133),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_124),
.B(n_125),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_126),
.B(n_182),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_127),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_146),
.B(n_207),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_143),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_131),
.B(n_143),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_134),
.C(n_138),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_132),
.B(n_205),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_134),
.B(n_138),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_137),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_135),
.A2(n_137),
.B1(n_199),
.B2(n_200),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_135),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_137),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

INVxp33_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_202),
.B(n_206),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_148),
.A2(n_189),
.B(n_201),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_171),
.B(n_188),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_156),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_150),
.B(n_156),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_153),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_151),
.A2(n_153),
.B1(n_154),
.B2(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_151),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_152),
.B(n_197),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_158),
.B1(n_163),
.B2(n_170),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_160),
.B1(n_161),
.B2(n_162),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_159),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_159),
.B(n_162),
.C(n_170),
.Y(n_190)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_160),
.Y(n_162)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_163),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_166),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_177),
.B(n_187),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_175),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_173),
.B(n_175),
.Y(n_187)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_174),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_183),
.B(n_186),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_181),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_184),
.B(n_185),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_190),
.B(n_191),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_198),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_196),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_193),
.B(n_196),
.C(n_198),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_203),
.B(n_204),
.Y(n_206)
);


endmodule