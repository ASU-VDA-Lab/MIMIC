module fake_jpeg_19157_n_212 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_212);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_212;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_3),
.B(n_11),
.Y(n_26)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx6_ASAP7_75t_SL g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_1),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_26),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_19),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_31),
.Y(n_50)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_37),
.Y(n_61)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_38),
.Y(n_57)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

BUFx24_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_35),
.A2(n_19),
.B1(n_15),
.B2(n_18),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_43),
.A2(n_56),
.B1(n_24),
.B2(n_22),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_30),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_46),
.B(n_60),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_47),
.B(n_28),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g48 ( 
.A(n_33),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_48),
.B(n_50),
.Y(n_72)
);

AOI22x1_ASAP7_75t_SL g51 ( 
.A1(n_33),
.A2(n_17),
.B1(n_27),
.B2(n_29),
.Y(n_51)
);

OA22x2_ASAP7_75t_L g85 ( 
.A1(n_51),
.A2(n_37),
.B1(n_29),
.B2(n_42),
.Y(n_85)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_36),
.A2(n_16),
.B1(n_31),
.B2(n_18),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_54),
.A2(n_64),
.B1(n_42),
.B2(n_41),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_20),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_59),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_38),
.A2(n_15),
.B1(n_23),
.B2(n_25),
.Y(n_56)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_30),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_30),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_62),
.B(n_21),
.Y(n_91)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_66),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_36),
.A2(n_16),
.B1(n_23),
.B2(n_25),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_36),
.B(n_20),
.Y(n_66)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_68),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_51),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_69),
.A2(n_84),
.B1(n_88),
.B2(n_89),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_53),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_70),
.B(n_79),
.Y(n_103)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_71),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_39),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_73),
.B(n_75),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_74),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_16),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_76),
.Y(n_113)
);

AND2x2_ASAP7_75t_SL g77 ( 
.A(n_60),
.B(n_32),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_77),
.B(n_82),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_39),
.C(n_32),
.Y(n_82)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_83),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_57),
.A2(n_42),
.B1(n_41),
.B2(n_29),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_85),
.B(n_86),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_61),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_52),
.B(n_24),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_92),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_59),
.A2(n_32),
.B1(n_22),
.B2(n_17),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_63),
.A2(n_32),
.B1(n_27),
.B2(n_21),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_96),
.Y(n_117)
);

BUFx4f_ASAP7_75t_SL g92 ( 
.A(n_61),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_67),
.A2(n_27),
.B1(n_21),
.B2(n_28),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_93),
.A2(n_49),
.B1(n_58),
.B2(n_5),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_65),
.A2(n_27),
.B1(n_2),
.B2(n_3),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_94),
.A2(n_53),
.B1(n_65),
.B2(n_67),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_53),
.B(n_13),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_12),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_45),
.B(n_37),
.C(n_2),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_97),
.A2(n_122),
.B1(n_95),
.B2(n_86),
.Y(n_131)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_71),
.Y(n_100)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_100),
.Y(n_136)
);

NOR3xp33_ASAP7_75t_SL g102 ( 
.A(n_72),
.B(n_37),
.C(n_4),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_102),
.B(n_116),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_80),
.A2(n_49),
.B1(n_44),
.B2(n_45),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_106),
.A2(n_108),
.B1(n_110),
.B2(n_115),
.Y(n_140)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_107),
.B(n_120),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_80),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_68),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_115)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_90),
.Y(n_118)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_118),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_69),
.A2(n_6),
.B(n_7),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_119),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_78),
.B(n_6),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_77),
.Y(n_121)
);

INVx13_ASAP7_75t_L g125 ( 
.A(n_121),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_82),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_105),
.A2(n_73),
.B1(n_96),
.B2(n_85),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_123),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_77),
.C(n_91),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_124),
.B(n_129),
.Y(n_150)
);

AND2x6_ASAP7_75t_L g126 ( 
.A(n_99),
.B(n_73),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_126),
.B(n_127),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_104),
.Y(n_127)
);

INVx13_ASAP7_75t_L g128 ( 
.A(n_114),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_128),
.B(n_138),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_117),
.B(n_77),
.C(n_75),
.Y(n_129)
);

NAND2xp33_ASAP7_75t_SL g130 ( 
.A(n_114),
.B(n_85),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_130),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_131),
.A2(n_132),
.B1(n_144),
.B2(n_115),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_121),
.A2(n_79),
.B1(n_88),
.B2(n_86),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_78),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_133),
.B(n_135),
.Y(n_159)
);

AO22x2_ASAP7_75t_L g135 ( 
.A1(n_98),
.A2(n_85),
.B1(n_83),
.B2(n_81),
.Y(n_135)
);

AOI32xp33_ASAP7_75t_L g138 ( 
.A1(n_103),
.A2(n_72),
.A3(n_81),
.B1(n_70),
.B2(n_83),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_107),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_142),
.B(n_143),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_118),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_119),
.A2(n_92),
.B1(n_10),
.B2(n_11),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_SL g145 ( 
.A(n_126),
.B(n_101),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_145),
.B(n_133),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_137),
.A2(n_140),
.B1(n_127),
.B2(n_109),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_147),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_148),
.A2(n_135),
.B1(n_132),
.B2(n_130),
.Y(n_164)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_141),
.Y(n_149)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_149),
.Y(n_168)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_141),
.Y(n_151)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_151),
.Y(n_175)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_136),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_152),
.Y(n_173)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_136),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_154),
.B(n_161),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_134),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_155),
.B(n_102),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_135),
.A2(n_98),
.B1(n_108),
.B2(n_109),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_160),
.B(n_148),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_140),
.A2(n_101),
.B1(n_113),
.B2(n_106),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_162),
.B(n_172),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_153),
.A2(n_123),
.B(n_128),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_163),
.A2(n_153),
.B(n_146),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_164),
.A2(n_165),
.B1(n_169),
.B2(n_135),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_159),
.A2(n_135),
.B1(n_124),
.B2(n_129),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_159),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_166),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_170),
.B(n_171),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_150),
.B(n_125),
.C(n_122),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_150),
.B(n_110),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_176),
.A2(n_181),
.B1(n_185),
.B2(n_186),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_167),
.A2(n_146),
.B(n_157),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_177),
.A2(n_179),
.B(n_183),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_174),
.B(n_158),
.Y(n_178)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_178),
.Y(n_189)
);

XNOR2x1_ASAP7_75t_L g179 ( 
.A(n_165),
.B(n_145),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_168),
.A2(n_111),
.B1(n_151),
.B2(n_149),
.Y(n_181)
);

XOR2x2_ASAP7_75t_L g183 ( 
.A(n_163),
.B(n_156),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_167),
.A2(n_154),
.B1(n_152),
.B2(n_125),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_180),
.B(n_171),
.C(n_179),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_187),
.B(n_182),
.C(n_176),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_183),
.A2(n_164),
.B1(n_174),
.B2(n_172),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_188),
.A2(n_191),
.B1(n_185),
.B2(n_111),
.Y(n_198)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_186),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_190),
.B(n_193),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_184),
.A2(n_175),
.B1(n_173),
.B2(n_162),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_177),
.B(n_142),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_187),
.B(n_180),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_195),
.B(n_196),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_198),
.B(n_199),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_194),
.B(n_139),
.Y(n_199)
);

OR2x2_ASAP7_75t_L g200 ( 
.A(n_193),
.B(n_188),
.Y(n_200)
);

AOI21x1_ASAP7_75t_L g203 ( 
.A1(n_200),
.A2(n_192),
.B(n_191),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_197),
.A2(n_194),
.B(n_189),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_202),
.B(n_203),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_204),
.A2(n_200),
.B1(n_197),
.B2(n_100),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_205),
.Y(n_208)
);

OAI21xp33_ASAP7_75t_L g206 ( 
.A1(n_201),
.A2(n_9),
.B(n_92),
.Y(n_206)
);

OAI21x1_ASAP7_75t_L g209 ( 
.A1(n_206),
.A2(n_9),
.B(n_92),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_209),
.A2(n_207),
.B(n_112),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_210),
.A2(n_208),
.B(n_112),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_211),
.B(n_201),
.Y(n_212)
);


endmodule