module fake_jpeg_13264_n_517 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_517);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_517;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_13),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_8),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_2),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_8),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_5),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_3),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_52),
.Y(n_106)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_53),
.Y(n_125)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

INVx11_ASAP7_75t_L g121 ( 
.A(n_54),
.Y(n_121)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_55),
.Y(n_112)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g114 ( 
.A(n_56),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_58),
.Y(n_131)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_59),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_60),
.Y(n_135)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_61),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_62),
.Y(n_140)
);

BUFx4f_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_63),
.Y(n_108)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_64),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_65),
.Y(n_148)
);

BUFx4f_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_66),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_67),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_19),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_68),
.B(n_74),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_69),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_70),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g151 ( 
.A(n_71),
.Y(n_151)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_72),
.Y(n_157)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_73),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_19),
.B(n_14),
.Y(n_74)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_26),
.Y(n_75)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_75),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_26),
.Y(n_76)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_76),
.Y(n_130)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_77),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_38),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_78),
.B(n_84),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_26),
.Y(n_79)
);

INVx3_ASAP7_75t_SL g105 ( 
.A(n_79),
.Y(n_105)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_37),
.Y(n_80)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_80),
.Y(n_122)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_41),
.Y(n_81)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_81),
.Y(n_133)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_82),
.Y(n_147)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_32),
.Y(n_83)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_83),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_38),
.B(n_14),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_85),
.Y(n_149)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_16),
.Y(n_86)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_86),
.Y(n_153)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_32),
.Y(n_87)
);

INVx2_ASAP7_75t_SL g129 ( 
.A(n_87),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_26),
.Y(n_88)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_88),
.Y(n_127)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_33),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_89),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_39),
.Y(n_90)
);

INVx3_ASAP7_75t_SL g136 ( 
.A(n_90),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_36),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_91),
.B(n_94),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_39),
.Y(n_92)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_92),
.Y(n_144)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_36),
.Y(n_93)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_93),
.Y(n_158)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_16),
.Y(n_94)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_39),
.Y(n_95)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_95),
.Y(n_134)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_39),
.Y(n_96)
);

BUFx24_ASAP7_75t_L g101 ( 
.A(n_96),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_44),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_97),
.B(n_98),
.Y(n_146)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_32),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_36),
.B(n_14),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_99),
.B(n_100),
.Y(n_155)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_33),
.Y(n_100)
);

BUFx12_ASAP7_75t_L g102 ( 
.A(n_70),
.Y(n_102)
);

BUFx16f_ASAP7_75t_L g178 ( 
.A(n_102),
.Y(n_178)
);

OA22x2_ASAP7_75t_L g104 ( 
.A1(n_51),
.A2(n_33),
.B1(n_46),
.B2(n_44),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_104),
.A2(n_59),
.B1(n_56),
.B2(n_71),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_29),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_107),
.B(n_113),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_75),
.B(n_29),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_96),
.A2(n_50),
.B1(n_49),
.B2(n_48),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_115),
.A2(n_30),
.B1(n_47),
.B2(n_21),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_57),
.B(n_45),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_117),
.B(n_137),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_70),
.B(n_50),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_128),
.B(n_150),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_58),
.B(n_45),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_60),
.B(n_31),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_138),
.B(n_142),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_62),
.B(n_31),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_65),
.B(n_49),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_143),
.B(n_152),
.Y(n_197)
);

NOR3xp33_ASAP7_75t_L g150 ( 
.A(n_67),
.B(n_32),
.C(n_27),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_69),
.B(n_47),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_160),
.A2(n_175),
.B1(n_23),
.B2(n_105),
.Y(n_245)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_103),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_161),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_145),
.B(n_32),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_162),
.B(n_166),
.Y(n_242)
);

CKINVDCx12_ASAP7_75t_R g163 ( 
.A(n_129),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_163),
.Y(n_209)
);

INVxp67_ASAP7_75t_SL g164 ( 
.A(n_124),
.Y(n_164)
);

BUFx24_ASAP7_75t_L g235 ( 
.A(n_164),
.Y(n_235)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_139),
.Y(n_165)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_165),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_145),
.B(n_34),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_125),
.Y(n_167)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_167),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_111),
.B(n_34),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_168),
.B(n_179),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_114),
.A2(n_40),
.B1(n_42),
.B2(n_28),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_169),
.Y(n_244)
);

BUFx12f_ASAP7_75t_L g170 ( 
.A(n_139),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_170),
.Y(n_215)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_118),
.Y(n_171)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_171),
.Y(n_217)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_126),
.Y(n_172)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_172),
.Y(n_222)
);

INVx4_ASAP7_75t_SL g173 ( 
.A(n_129),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_173),
.B(n_202),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_114),
.A2(n_42),
.B1(n_17),
.B2(n_28),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_174),
.A2(n_177),
.B1(n_180),
.B2(n_193),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_146),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_176),
.B(n_194),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_153),
.A2(n_17),
.B1(n_40),
.B2(n_27),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_111),
.B(n_30),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_119),
.A2(n_27),
.B1(n_48),
.B2(n_21),
.Y(n_180)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_133),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_181),
.Y(n_241)
);

INVx5_ASAP7_75t_SL g182 ( 
.A(n_102),
.Y(n_182)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_182),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_141),
.B(n_13),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_184),
.B(n_186),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_103),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_185),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_141),
.B(n_112),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_151),
.Y(n_187)
);

BUFx12f_ASAP7_75t_L g212 ( 
.A(n_187),
.Y(n_212)
);

CKINVDCx12_ASAP7_75t_R g188 ( 
.A(n_123),
.Y(n_188)
);

BUFx8_ASAP7_75t_L g210 ( 
.A(n_188),
.Y(n_210)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_151),
.Y(n_189)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_189),
.Y(n_231)
);

INVx6_ASAP7_75t_L g190 ( 
.A(n_109),
.Y(n_190)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_190),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_104),
.A2(n_79),
.B1(n_92),
.B2(n_90),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_192),
.A2(n_105),
.B1(n_136),
.B2(n_140),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_156),
.A2(n_46),
.B1(n_44),
.B2(n_88),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_106),
.B(n_97),
.Y(n_194)
);

INVx6_ASAP7_75t_L g196 ( 
.A(n_109),
.Y(n_196)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_196),
.Y(n_238)
);

INVx5_ASAP7_75t_SL g198 ( 
.A(n_121),
.Y(n_198)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_198),
.Y(n_243)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_127),
.Y(n_199)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_199),
.Y(n_247)
);

CKINVDCx12_ASAP7_75t_R g200 ( 
.A(n_101),
.Y(n_200)
);

OR2x2_ASAP7_75t_L g240 ( 
.A(n_200),
.B(n_134),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_151),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_201),
.B(n_204),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_108),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_158),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_203),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_146),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_154),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_205),
.B(n_208),
.Y(n_227)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_147),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_206),
.Y(n_224)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_122),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_207),
.B(n_136),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_149),
.B(n_97),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_183),
.A2(n_104),
.B1(n_132),
.B2(n_157),
.Y(n_218)
);

OAI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_218),
.A2(n_232),
.B1(n_175),
.B2(n_131),
.Y(n_283)
);

FAx1_ASAP7_75t_SL g225 ( 
.A(n_183),
.B(n_155),
.CI(n_101),
.CON(n_225),
.SN(n_225)
);

MAJIxp5_ASAP7_75t_SL g268 ( 
.A(n_225),
.B(n_195),
.C(n_197),
.Y(n_268)
);

NAND2x1_ASAP7_75t_L g229 ( 
.A(n_176),
.B(n_150),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_229),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_192),
.A2(n_132),
.B1(n_110),
.B2(n_120),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_233),
.A2(n_163),
.B1(n_200),
.B2(n_144),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_234),
.Y(n_254)
);

AND2x2_ASAP7_75t_SL g236 ( 
.A(n_207),
.B(n_155),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_236),
.B(n_173),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_195),
.B(n_130),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_239),
.B(n_167),
.Y(n_280)
);

INVxp33_ASAP7_75t_L g281 ( 
.A(n_240),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_245),
.A2(n_244),
.B1(n_236),
.B2(n_233),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_L g248 ( 
.A1(n_204),
.A2(n_130),
.B1(n_110),
.B2(n_120),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g277 ( 
.A1(n_248),
.A2(n_198),
.B1(n_196),
.B2(n_190),
.Y(n_277)
);

INVx13_ASAP7_75t_L g249 ( 
.A(n_209),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_249),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_209),
.A2(n_159),
.B(n_191),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_250),
.A2(n_265),
.B(n_268),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_246),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_251),
.B(n_258),
.Y(n_290)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_217),
.Y(n_252)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_252),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_253),
.A2(n_269),
.B1(n_277),
.B2(n_240),
.Y(n_289)
);

INVx13_ASAP7_75t_L g255 ( 
.A(n_235),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_255),
.Y(n_316)
);

INVx8_ASAP7_75t_L g256 ( 
.A(n_213),
.Y(n_256)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_256),
.Y(n_303)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_217),
.Y(n_257)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_257),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_246),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_242),
.B(n_191),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_259),
.B(n_267),
.Y(n_286)
);

INVx8_ASAP7_75t_L g260 ( 
.A(n_213),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_260),
.B(n_266),
.Y(n_295)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_234),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_261),
.Y(n_312)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_243),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_263),
.B(n_264),
.Y(n_296)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_243),
.Y(n_264)
);

INVx8_ASAP7_75t_L g266 ( 
.A(n_219),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_239),
.B(n_197),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_236),
.B(n_171),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_270),
.B(n_272),
.Y(n_297)
);

CKINVDCx12_ASAP7_75t_R g271 ( 
.A(n_235),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_271),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_216),
.B(n_205),
.Y(n_272)
);

AND2x6_ASAP7_75t_L g273 ( 
.A(n_225),
.B(n_182),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_273),
.B(n_274),
.Y(n_299)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_246),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_222),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_275),
.B(n_280),
.Y(n_302)
);

AND2x2_ASAP7_75t_SL g276 ( 
.A(n_225),
.B(n_172),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_276),
.B(n_247),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_223),
.B(n_178),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_278),
.B(n_224),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_218),
.B(n_173),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_279),
.A2(n_23),
.B(n_210),
.Y(n_315)
);

INVx13_ASAP7_75t_L g282 ( 
.A(n_235),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_282),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_283),
.A2(n_220),
.B1(n_238),
.B2(n_230),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_227),
.B(n_202),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_284),
.B(n_285),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_221),
.B(n_188),
.Y(n_285)
);

FAx1_ASAP7_75t_SL g287 ( 
.A(n_268),
.B(n_229),
.CI(n_226),
.CON(n_287),
.SN(n_287)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_287),
.B(n_294),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_269),
.A2(n_232),
.B1(n_211),
.B2(n_244),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_288),
.A2(n_289),
.B1(n_293),
.B2(n_258),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_254),
.A2(n_229),
.B1(n_238),
.B2(n_230),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_298),
.B(n_310),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_SL g334 ( 
.A(n_300),
.B(n_308),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_249),
.Y(n_301)
);

BUFx12f_ASAP7_75t_L g333 ( 
.A(n_301),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_281),
.B(n_228),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_304),
.B(n_284),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_262),
.B(n_228),
.C(n_247),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_306),
.B(n_309),
.C(n_311),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_267),
.B(n_222),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_276),
.B(n_237),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_279),
.A2(n_161),
.B1(n_219),
.B2(n_214),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_262),
.B(n_241),
.C(n_237),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_279),
.A2(n_214),
.B1(n_185),
.B2(n_148),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_314),
.B(n_317),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_315),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_276),
.A2(n_185),
.B1(n_135),
.B2(n_148),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_265),
.A2(n_210),
.B(n_178),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_319),
.A2(n_274),
.B(n_265),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_308),
.B(n_270),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_322),
.B(n_320),
.C(n_297),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_296),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_323),
.B(n_324),
.Y(n_355)
);

INVx8_ASAP7_75t_L g324 ( 
.A(n_301),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_325),
.A2(n_338),
.B(n_290),
.Y(n_358)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_291),
.Y(n_327)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_327),
.Y(n_370)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_291),
.Y(n_330)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_330),
.Y(n_384)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_307),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_331),
.B(n_332),
.Y(n_381)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_307),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_335),
.A2(n_345),
.B1(n_314),
.B2(n_253),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_299),
.A2(n_273),
.B(n_250),
.Y(n_336)
);

AO21x1_ASAP7_75t_L g378 ( 
.A1(n_336),
.A2(n_352),
.B(n_210),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_337),
.B(n_340),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_299),
.A2(n_285),
.B(n_251),
.Y(n_338)
);

BUFx3_ASAP7_75t_L g339 ( 
.A(n_303),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_339),
.B(n_342),
.Y(n_367)
);

CKINVDCx16_ASAP7_75t_R g340 ( 
.A(n_296),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_319),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_SL g382 ( 
.A1(n_341),
.A2(n_348),
.B1(n_351),
.B2(n_354),
.Y(n_382)
);

AND2x6_ASAP7_75t_L g342 ( 
.A(n_287),
.B(n_254),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_312),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_343),
.B(n_344),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_302),
.Y(n_344)
);

AOI22xp33_ASAP7_75t_SL g345 ( 
.A1(n_288),
.A2(n_263),
.B1(n_264),
.B2(n_271),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_302),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_346),
.B(n_350),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_286),
.B(n_272),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_SL g357 ( 
.A(n_347),
.B(n_320),
.Y(n_357)
);

INVx4_ASAP7_75t_L g348 ( 
.A(n_313),
.Y(n_348)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_304),
.Y(n_350)
);

INVx1_ASAP7_75t_SL g351 ( 
.A(n_306),
.Y(n_351)
);

AND2x6_ASAP7_75t_L g352 ( 
.A(n_287),
.B(n_292),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_294),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_353),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_311),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_356),
.B(n_331),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_357),
.B(n_260),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_358),
.A2(n_366),
.B(n_379),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_324),
.B(n_310),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_359),
.Y(n_388)
);

O2A1O1Ixp33_ASAP7_75t_L g360 ( 
.A1(n_349),
.A2(n_305),
.B(n_292),
.C(n_316),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_360),
.B(n_231),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_321),
.A2(n_261),
.B1(n_280),
.B2(n_298),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_361),
.A2(n_369),
.B1(n_378),
.B2(n_326),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_333),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_362),
.B(n_170),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_351),
.B(n_300),
.C(n_309),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_365),
.B(n_374),
.C(n_376),
.Y(n_396)
);

NAND2x1p5_ASAP7_75t_L g366 ( 
.A(n_338),
.B(n_315),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_321),
.A2(n_305),
.B1(n_303),
.B2(n_317),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_SL g371 ( 
.A(n_334),
.B(n_257),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_SL g394 ( 
.A(n_371),
.B(n_375),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_372),
.A2(n_328),
.B1(n_326),
.B2(n_332),
.Y(n_393)
);

NOR2xp67_ASAP7_75t_L g373 ( 
.A(n_342),
.B(n_252),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_373),
.B(n_170),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_354),
.B(n_275),
.C(n_316),
.Y(n_374)
);

XNOR2x1_ASAP7_75t_L g375 ( 
.A(n_329),
.B(n_318),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_329),
.B(n_295),
.C(n_199),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_335),
.A2(n_328),
.B1(n_336),
.B2(n_352),
.Y(n_377)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_377),
.Y(n_392)
);

A2O1A1Ixp33_ASAP7_75t_SL g379 ( 
.A1(n_325),
.A2(n_282),
.B(n_255),
.C(n_212),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_334),
.B(n_165),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_380),
.B(n_385),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g383 ( 
.A1(n_341),
.A2(n_215),
.B(n_187),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_383),
.A2(n_386),
.B(n_189),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_322),
.B(n_178),
.Y(n_385)
);

A2O1A1Ixp33_ASAP7_75t_SL g386 ( 
.A1(n_333),
.A2(n_212),
.B(n_266),
.C(n_215),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_387),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_389),
.B(n_407),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_364),
.B(n_333),
.Y(n_390)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_390),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_393),
.A2(n_410),
.B1(n_382),
.B2(n_383),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_395),
.A2(n_366),
.B1(n_379),
.B2(n_386),
.Y(n_439)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_368),
.Y(n_397)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_397),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_398),
.B(n_380),
.Y(n_431)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_381),
.Y(n_399)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_399),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_364),
.B(n_327),
.Y(n_400)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_400),
.Y(n_434)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_370),
.Y(n_401)
);

INVx1_ASAP7_75t_SL g420 ( 
.A(n_401),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_375),
.B(n_348),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_403),
.B(n_385),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_404),
.B(n_413),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_363),
.B(n_339),
.Y(n_405)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_405),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_SL g432 ( 
.A1(n_406),
.A2(n_379),
.B(n_386),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_355),
.B(n_256),
.Y(n_408)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_408),
.Y(n_437)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_384),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_409),
.B(n_411),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_360),
.A2(n_231),
.B1(n_135),
.B2(n_131),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_361),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_369),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_412),
.B(n_414),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_359),
.B(n_212),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_367),
.B(n_212),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_415),
.B(n_201),
.Y(n_433)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_416),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_396),
.B(n_376),
.C(n_374),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_419),
.B(n_430),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_SL g426 ( 
.A(n_394),
.B(n_371),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_426),
.B(n_427),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_428),
.B(n_438),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_396),
.B(n_365),
.C(n_378),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_431),
.B(n_438),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_432),
.A2(n_435),
.B(n_391),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_L g446 ( 
.A1(n_433),
.A2(n_439),
.B1(n_404),
.B2(n_410),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_391),
.A2(n_366),
.B(n_379),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_398),
.B(n_356),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_420),
.B(n_390),
.Y(n_440)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_440),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_441),
.B(n_443),
.Y(n_462)
);

BUFx2_ASAP7_75t_L g442 ( 
.A(n_422),
.Y(n_442)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_442),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_419),
.B(n_430),
.C(n_431),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_444),
.B(n_448),
.Y(n_465)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_425),
.Y(n_445)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_445),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_446),
.A2(n_427),
.B1(n_417),
.B2(n_437),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_SL g447 ( 
.A(n_418),
.B(n_405),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_447),
.B(n_442),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_424),
.B(n_414),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_420),
.B(n_400),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_449),
.B(n_454),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_L g450 ( 
.A1(n_439),
.A2(n_392),
.B1(n_393),
.B2(n_388),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_450),
.A2(n_457),
.B1(n_413),
.B2(n_402),
.Y(n_473)
);

AOI21xp5_ASAP7_75t_L g452 ( 
.A1(n_435),
.A2(n_406),
.B(n_388),
.Y(n_452)
);

AOI21xp5_ASAP7_75t_L g464 ( 
.A1(n_452),
.A2(n_432),
.B(n_406),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_423),
.B(n_408),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_429),
.B(n_403),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_455),
.B(n_458),
.Y(n_471)
);

CKINVDCx14_ASAP7_75t_R g457 ( 
.A(n_417),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_434),
.Y(n_458)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_459),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_SL g463 ( 
.A(n_451),
.B(n_428),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_463),
.B(n_467),
.Y(n_477)
);

AOI21x1_ASAP7_75t_L g487 ( 
.A1(n_464),
.A2(n_386),
.B(n_426),
.Y(n_487)
);

A2O1A1Ixp33_ASAP7_75t_L g466 ( 
.A1(n_441),
.A2(n_421),
.B(n_417),
.C(n_436),
.Y(n_466)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_466),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_456),
.B(n_401),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_469),
.B(n_470),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_444),
.B(n_453),
.C(n_443),
.Y(n_470)
);

HB1xp67_ASAP7_75t_L g481 ( 
.A(n_473),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_455),
.B(n_402),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_474),
.B(n_475),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_451),
.B(n_394),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_465),
.B(n_440),
.Y(n_476)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_476),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_SL g480 ( 
.A(n_470),
.B(n_468),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_SL g498 ( 
.A(n_480),
.B(n_483),
.Y(n_498)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_462),
.B(n_453),
.Y(n_482)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_482),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_SL g483 ( 
.A(n_462),
.B(n_449),
.Y(n_483)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_466),
.A2(n_452),
.B(n_413),
.Y(n_485)
);

AOI21xp5_ASAP7_75t_SL g495 ( 
.A1(n_485),
.A2(n_488),
.B(n_475),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_487),
.B(n_116),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_472),
.B(n_170),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_474),
.B(n_140),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_489),
.B(n_76),
.Y(n_497)
);

AOI22xp33_ASAP7_75t_L g491 ( 
.A1(n_484),
.A2(n_461),
.B1(n_460),
.B2(n_467),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_491),
.B(n_493),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_486),
.B(n_471),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_L g502 ( 
.A1(n_492),
.A2(n_499),
.B(n_488),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_479),
.B(n_463),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_495),
.B(n_477),
.C(n_478),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_496),
.B(n_497),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_476),
.B(n_46),
.Y(n_499)
);

HB1xp67_ASAP7_75t_L g507 ( 
.A(n_502),
.Y(n_507)
);

AOI21xp5_ASAP7_75t_L g503 ( 
.A1(n_494),
.A2(n_477),
.B(n_481),
.Y(n_503)
);

NAND3xp33_ASAP7_75t_L g509 ( 
.A(n_503),
.B(n_500),
.C(n_501),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_504),
.B(n_505),
.Y(n_510)
);

AOI322xp5_ASAP7_75t_L g505 ( 
.A1(n_490),
.A2(n_46),
.A3(n_44),
.B1(n_66),
.B2(n_63),
.C1(n_6),
.C2(n_7),
.Y(n_505)
);

AOI322xp5_ASAP7_75t_L g506 ( 
.A1(n_498),
.A2(n_1),
.A3(n_2),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_7),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_506),
.B(n_492),
.C(n_2),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_508),
.B(n_509),
.Y(n_512)
);

AOI322xp5_ASAP7_75t_L g511 ( 
.A1(n_510),
.A2(n_1),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C1(n_10),
.C2(n_11),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_511),
.B(n_507),
.C(n_512),
.Y(n_513)
);

OAI22xp33_ASAP7_75t_R g514 ( 
.A1(n_513),
.A2(n_1),
.B1(n_5),
.B2(n_6),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_514),
.B(n_1),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_515),
.B(n_10),
.Y(n_516)
);

AO21x1_ASAP7_75t_L g517 ( 
.A1(n_516),
.A2(n_10),
.B(n_11),
.Y(n_517)
);


endmodule