module real_aes_14655_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_673;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_89;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_502;
wire n_434;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_85;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_87;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_288;
wire n_147;
wire n_150;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_691;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_623;
wire n_249;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
wire n_91;
INVx2_ASAP7_75t_SL g146 ( .A(n_0), .Y(n_146) );
CKINVDCx5p33_ASAP7_75t_R g215 ( .A(n_1), .Y(n_215) );
OA21x2_ASAP7_75t_L g94 ( .A1(n_2), .A2(n_41), .B(n_95), .Y(n_94) );
INVx1_ASAP7_75t_L g154 ( .A(n_2), .Y(n_154) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_3), .B(n_143), .Y(n_237) );
NAND2xp5_ASAP7_75t_SL g164 ( .A(n_4), .B(n_165), .Y(n_164) );
AOI22xp5_ASAP7_75t_L g689 ( .A1(n_4), .A2(n_690), .B1(n_691), .B2(n_692), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_4), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_5), .A2(n_31), .B1(n_572), .B2(n_573), .Y(n_571) );
INVxp33_ASAP7_75t_SL g662 ( .A(n_5), .Y(n_662) );
AOI221xp5_ASAP7_75t_L g575 ( .A1(n_6), .A2(n_19), .B1(n_576), .B2(n_577), .C(n_578), .Y(n_575) );
INVxp33_ASAP7_75t_SL g610 ( .A(n_6), .Y(n_610) );
AND2x2_ASAP7_75t_L g287 ( .A(n_7), .B(n_92), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g103 ( .A(n_8), .B(n_104), .Y(n_103) );
BUFx3_ASAP7_75t_L g604 ( .A(n_9), .Y(n_604) );
INVx3_ASAP7_75t_L g521 ( .A(n_10), .Y(n_521) );
INVx1_ASAP7_75t_L g609 ( .A(n_11), .Y(n_609) );
INVx2_ASAP7_75t_L g621 ( .A(n_11), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_12), .B(n_191), .Y(n_230) );
AOI22xp33_ASAP7_75t_SL g551 ( .A1(n_13), .A2(n_16), .B1(n_552), .B2(n_555), .Y(n_551) );
INVx1_ASAP7_75t_L g674 ( .A(n_13), .Y(n_674) );
BUFx3_ASAP7_75t_L g102 ( .A(n_14), .Y(n_102) );
INVx1_ASAP7_75t_L g107 ( .A(n_14), .Y(n_107) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_15), .B(n_91), .Y(n_241) );
AOI22xp33_ASAP7_75t_SL g629 ( .A1(n_16), .A2(n_65), .B1(n_630), .B2(n_634), .Y(n_629) );
CKINVDCx5p33_ASAP7_75t_R g696 ( .A(n_17), .Y(n_696) );
BUFx10_ASAP7_75t_L g715 ( .A(n_18), .Y(n_715) );
INVxp33_ASAP7_75t_SL g657 ( .A(n_19), .Y(n_657) );
HB1xp67_ASAP7_75t_L g699 ( .A(n_20), .Y(n_699) );
CKINVDCx5p33_ASAP7_75t_R g204 ( .A(n_21), .Y(n_204) );
NAND3xp33_ASAP7_75t_L g173 ( .A(n_22), .B(n_168), .C(n_174), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_23), .B(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g528 ( .A(n_24), .B(n_529), .Y(n_528) );
AND2x2_ASAP7_75t_L g545 ( .A(n_24), .B(n_33), .Y(n_545) );
INVx1_ASAP7_75t_L g570 ( .A(n_24), .Y(n_570) );
INVx1_ASAP7_75t_L g125 ( .A(n_25), .Y(n_125) );
INVx2_ASAP7_75t_L g533 ( .A(n_26), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_27), .Y(n_534) );
AOI221xp5_ASAP7_75t_L g669 ( .A1(n_27), .A2(n_55), .B1(n_631), .B2(n_670), .C(n_673), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_28), .B(n_135), .Y(n_134) );
INVx1_ASAP7_75t_L g541 ( .A(n_29), .Y(n_541) );
INVx1_ASAP7_75t_L g546 ( .A(n_30), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g617 ( .A1(n_30), .A2(n_46), .B1(n_618), .B2(n_623), .Y(n_617) );
INVxp67_ASAP7_75t_SL g676 ( .A(n_31), .Y(n_676) );
HB1xp67_ASAP7_75t_L g698 ( .A(n_32), .Y(n_698) );
INVx2_ASAP7_75t_L g529 ( .A(n_33), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_33), .B(n_570), .Y(n_579) );
NAND2xp5_ASAP7_75t_SL g252 ( .A(n_34), .B(n_253), .Y(n_252) );
INVx1_ASAP7_75t_L g744 ( .A(n_34), .Y(n_744) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_35), .B(n_219), .Y(n_218) );
INVx1_ASAP7_75t_L g691 ( .A(n_35), .Y(n_691) );
AND2x4_ASAP7_75t_L g124 ( .A(n_36), .B(n_125), .Y(n_124) );
HB1xp67_ASAP7_75t_L g709 ( .A(n_36), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_37), .B(n_91), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_38), .B(n_120), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g90 ( .A(n_39), .B(n_91), .Y(n_90) );
INVx1_ASAP7_75t_L g615 ( .A(n_40), .Y(n_615) );
INVx1_ASAP7_75t_L g622 ( .A(n_40), .Y(n_622) );
INVx1_ASAP7_75t_L g153 ( .A(n_41), .Y(n_153) );
CKINVDCx5p33_ASAP7_75t_R g284 ( .A(n_42), .Y(n_284) );
A2O1A1Ixp33_ASAP7_75t_L g141 ( .A1(n_43), .A2(n_142), .B(n_144), .C(n_147), .Y(n_141) );
INVx1_ASAP7_75t_L g95 ( .A(n_44), .Y(n_95) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_45), .B(n_91), .Y(n_221) );
AOI221xp5_ASAP7_75t_L g558 ( .A1(n_46), .A2(n_55), .B1(n_559), .B2(n_563), .C(n_568), .Y(n_558) );
INVx3_ASAP7_75t_L g201 ( .A(n_47), .Y(n_201) );
INVx1_ASAP7_75t_L g589 ( .A(n_48), .Y(n_589) );
NAND2xp5_ASAP7_75t_SL g115 ( .A(n_49), .B(n_99), .Y(n_115) );
INVx1_ASAP7_75t_L g233 ( .A(n_50), .Y(n_233) );
HB1xp67_ASAP7_75t_L g687 ( .A(n_51), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_52), .B(n_163), .Y(n_162) );
CKINVDCx5p33_ASAP7_75t_R g279 ( .A(n_53), .Y(n_279) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_54), .B(n_174), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_56), .B(n_171), .Y(n_257) );
HB1xp67_ASAP7_75t_L g745 ( .A(n_56), .Y(n_745) );
BUFx2_ASAP7_75t_L g685 ( .A(n_57), .Y(n_685) );
INVx1_ASAP7_75t_L g133 ( .A(n_58), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_59), .B(n_239), .Y(n_238) );
CKINVDCx5p33_ASAP7_75t_R g285 ( .A(n_60), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_61), .B(n_168), .Y(n_167) );
INVx1_ASAP7_75t_L g110 ( .A(n_62), .Y(n_110) );
INVx1_ASAP7_75t_L g149 ( .A(n_62), .Y(n_149) );
BUFx3_ASAP7_75t_L g191 ( .A(n_62), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_63), .B(n_163), .Y(n_212) );
INVx1_ASAP7_75t_L g199 ( .A(n_64), .Y(n_199) );
INVx1_ASAP7_75t_L g524 ( .A(n_65), .Y(n_524) );
INVx1_ASAP7_75t_L g581 ( .A(n_66), .Y(n_581) );
INVx2_ASAP7_75t_L g532 ( .A(n_67), .Y(n_532) );
AND2x2_ASAP7_75t_L g549 ( .A(n_67), .B(n_533), .Y(n_549) );
INVxp67_ASAP7_75t_SL g566 ( .A(n_67), .Y(n_566) );
AOI22xp5_ASAP7_75t_L g727 ( .A1(n_68), .A2(n_514), .B1(n_703), .B2(n_728), .Y(n_727) );
CKINVDCx5p33_ASAP7_75t_R g728 ( .A(n_68), .Y(n_728) );
NAND2xp5_ASAP7_75t_SL g255 ( .A(n_69), .B(n_256), .Y(n_255) );
INVx1_ASAP7_75t_L g593 ( .A(n_70), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_71), .B(n_92), .Y(n_258) );
INVx2_ASAP7_75t_L g606 ( .A(n_72), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_73), .B(n_113), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g194 ( .A(n_74), .Y(n_194) );
INVx1_ASAP7_75t_L g189 ( .A(n_75), .Y(n_189) );
CKINVDCx5p33_ASAP7_75t_R g281 ( .A(n_76), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g98 ( .A(n_77), .B(n_99), .Y(n_98) );
AOI21xp33_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_505), .B(n_512), .Y(n_78) );
INVx3_ASAP7_75t_L g79 ( .A(n_80), .Y(n_79) );
AND2x4_ASAP7_75t_L g80 ( .A(n_81), .B(n_410), .Y(n_80) );
NOR3xp33_ASAP7_75t_L g81 ( .A(n_82), .B(n_346), .C(n_381), .Y(n_81) );
NAND3xp33_ASAP7_75t_SL g82 ( .A(n_83), .B(n_288), .C(n_318), .Y(n_82) );
AOI22xp5_ASAP7_75t_L g83 ( .A1(n_84), .A2(n_178), .B1(n_242), .B2(n_264), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_85), .Y(n_84) );
NOR2xp33_ASAP7_75t_L g452 ( .A(n_85), .B(n_453), .Y(n_452) );
OR2x2_ASAP7_75t_L g85 ( .A(n_86), .B(n_126), .Y(n_85) );
AND2x2_ASAP7_75t_L g426 ( .A(n_86), .B(n_427), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_86), .B(n_373), .Y(n_439) );
INVx2_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
NAND3xp33_ASAP7_75t_L g405 ( .A(n_87), .B(n_223), .C(n_327), .Y(n_405) );
INVx1_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
AND2x2_ASAP7_75t_L g291 ( .A(n_88), .B(n_244), .Y(n_291) );
INVx2_ASAP7_75t_L g322 ( .A(n_88), .Y(n_322) );
OR2x2_ASAP7_75t_L g345 ( .A(n_88), .B(n_321), .Y(n_345) );
AND2x2_ASAP7_75t_L g361 ( .A(n_88), .B(n_157), .Y(n_361) );
BUFx2_ASAP7_75t_L g415 ( .A(n_88), .Y(n_415) );
AND2x4_ASAP7_75t_L g423 ( .A(n_88), .B(n_380), .Y(n_423) );
INVx2_ASAP7_75t_L g433 ( .A(n_88), .Y(n_433) );
BUFx6f_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
NAND2x1_ASAP7_75t_L g89 ( .A(n_90), .B(n_96), .Y(n_89) );
HB1xp67_ASAP7_75t_L g263 ( .A(n_91), .Y(n_263) );
BUFx6f_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
INVx2_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_94), .Y(n_93) );
BUFx6f_ASAP7_75t_L g120 ( .A(n_94), .Y(n_120) );
BUFx2_ASAP7_75t_L g208 ( .A(n_94), .Y(n_208) );
INVx1_ASAP7_75t_L g155 ( .A(n_95), .Y(n_155) );
OAI21x1_ASAP7_75t_SL g96 ( .A1(n_97), .A2(n_111), .B(n_118), .Y(n_96) );
AOI21xp5_ASAP7_75t_L g97 ( .A1(n_98), .A2(n_103), .B(n_108), .Y(n_97) );
AOI22xp33_ASAP7_75t_L g197 ( .A1(n_99), .A2(n_198), .B1(n_200), .B2(n_202), .Y(n_197) );
INVx2_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_100), .B(n_194), .Y(n_193) );
INVx2_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
INVx2_ASAP7_75t_L g145 ( .A(n_101), .Y(n_145) );
INVx1_ASAP7_75t_L g239 ( .A(n_101), .Y(n_239) );
BUFx6f_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_102), .Y(n_132) );
INVx2_ASAP7_75t_L g175 ( .A(n_102), .Y(n_175) );
INVx2_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx2_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g114 ( .A(n_106), .Y(n_114) );
INVx2_ASAP7_75t_L g143 ( .A(n_106), .Y(n_143) );
INVx2_ASAP7_75t_L g219 ( .A(n_106), .Y(n_219) );
BUFx6f_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx2_ASAP7_75t_L g137 ( .A(n_107), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_108), .Y(n_138) );
INVx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx2_ASAP7_75t_L g196 ( .A(n_109), .Y(n_196) );
INVx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
BUFx3_ASAP7_75t_L g117 ( .A(n_110), .Y(n_117) );
AOI21xp5_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_115), .B(n_116), .Y(n_111) );
INVx1_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_117), .A2(n_250), .B(n_252), .Y(n_249) );
NOR2x1_ASAP7_75t_SL g118 ( .A(n_119), .B(n_121), .Y(n_118) );
BUFx6f_ASAP7_75t_L g247 ( .A(n_119), .Y(n_247) );
BUFx6f_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_L g159 ( .A(n_120), .Y(n_159) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx2_ASAP7_75t_SL g122 ( .A(n_123), .Y(n_122) );
INVx1_ASAP7_75t_L g176 ( .A(n_123), .Y(n_176) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx1_ASAP7_75t_L g156 ( .A(n_124), .Y(n_156) );
INVx3_ASAP7_75t_L g192 ( .A(n_124), .Y(n_192) );
BUFx6f_ASAP7_75t_SL g240 ( .A(n_124), .Y(n_240) );
HB1xp67_ASAP7_75t_L g711 ( .A(n_125), .Y(n_711) );
OR2x2_ASAP7_75t_L g418 ( .A(n_126), .B(n_297), .Y(n_418) );
INVx2_ASAP7_75t_L g476 ( .A(n_126), .Y(n_476) );
OR2x2_ASAP7_75t_SL g126 ( .A(n_127), .B(n_157), .Y(n_126) );
OR2x6_ASAP7_75t_L g259 ( .A(n_127), .B(n_260), .Y(n_259) );
INVx2_ASAP7_75t_L g298 ( .A(n_127), .Y(n_298) );
INVx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx2_ASAP7_75t_L g294 ( .A(n_128), .Y(n_294) );
OAI21x1_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_139), .B(n_150), .Y(n_128) );
AOI21x1_ASAP7_75t_SL g129 ( .A1(n_130), .A2(n_134), .B(n_138), .Y(n_129) );
OR2x2_ASAP7_75t_L g130 ( .A(n_131), .B(n_133), .Y(n_130) );
INVx3_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx2_ASAP7_75t_L g163 ( .A(n_132), .Y(n_163) );
INVx2_ASAP7_75t_L g217 ( .A(n_132), .Y(n_217) );
INVx2_ASAP7_75t_L g229 ( .A(n_132), .Y(n_229) );
INVx2_ASAP7_75t_L g251 ( .A(n_132), .Y(n_251) );
INVx3_ASAP7_75t_L g278 ( .A(n_132), .Y(n_278) );
HB1xp67_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx2_ASAP7_75t_L g165 ( .A(n_136), .Y(n_165) );
INVx2_ASAP7_75t_L g253 ( .A(n_136), .Y(n_253) );
INVx2_ASAP7_75t_L g256 ( .A(n_136), .Y(n_256) );
INVx3_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_137), .Y(n_172) );
AOI22x1_ASAP7_75t_L g275 ( .A1(n_138), .A2(n_148), .B1(n_276), .B2(n_282), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_140), .B(n_141), .Y(n_139) );
OAI21xp33_ASAP7_75t_L g150 ( .A1(n_140), .A2(n_151), .B(n_156), .Y(n_150) );
OAI22xp5_ASAP7_75t_L g282 ( .A1(n_142), .A2(n_283), .B1(n_284), .B2(n_285), .Y(n_282) );
INVx1_ASAP7_75t_L g511 ( .A(n_142), .Y(n_511) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
NOR2xp33_ASAP7_75t_L g144 ( .A(n_145), .B(n_146), .Y(n_144) );
INVx1_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
AOI21x1_ASAP7_75t_L g161 ( .A1(n_148), .A2(n_162), .B(n_164), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_148), .B(n_510), .Y(n_509) );
BUFx3_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g169 ( .A(n_149), .Y(n_169) );
INVxp67_ASAP7_75t_L g309 ( .A(n_151), .Y(n_309) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
AO21x2_ASAP7_75t_L g152 ( .A1(n_153), .A2(n_154), .B(n_155), .Y(n_152) );
AOI21x1_ASAP7_75t_L g185 ( .A1(n_153), .A2(n_154), .B(n_155), .Y(n_185) );
INVx1_ASAP7_75t_L g311 ( .A(n_156), .Y(n_311) );
AND2x2_ASAP7_75t_L g427 ( .A(n_157), .B(n_294), .Y(n_427) );
OA21x2_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_160), .B(n_177), .Y(n_157) );
INVx1_ASAP7_75t_SL g158 ( .A(n_159), .Y(n_158) );
OAI21x1_ASAP7_75t_L g262 ( .A1(n_160), .A2(n_177), .B(n_263), .Y(n_262) );
OAI21x1_ASAP7_75t_L g160 ( .A1(n_161), .A2(n_166), .B(n_176), .Y(n_160) );
OAI21xp5_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_170), .B(n_173), .Y(n_166) );
INVx1_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
BUFx10_ASAP7_75t_L g213 ( .A(n_169), .Y(n_213) );
INVxp67_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g188 ( .A(n_172), .B(n_189), .Y(n_188) );
INVx1_ASAP7_75t_L g202 ( .A(n_172), .Y(n_202) );
INVx1_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx2_ASAP7_75t_L g235 ( .A(n_175), .Y(n_235) );
OAI21xp5_ASAP7_75t_L g209 ( .A1(n_176), .A2(n_210), .B(n_214), .Y(n_209) );
AND2x2_ASAP7_75t_L g178 ( .A(n_179), .B(n_222), .Y(n_178) );
AND2x2_ASAP7_75t_L g398 ( .A(n_179), .B(n_328), .Y(n_398) );
HB1xp67_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx1_ASAP7_75t_L g451 ( .A(n_180), .Y(n_451) );
AND2x2_ASAP7_75t_L g499 ( .A(n_180), .B(n_338), .Y(n_499) );
AND2x2_ASAP7_75t_L g180 ( .A(n_181), .B(n_205), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_182), .B(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g333 ( .A(n_182), .B(n_334), .Y(n_333) );
AO21x1_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_186), .B(n_203), .Y(n_182) );
AO21x2_ASAP7_75t_L g304 ( .A1(n_183), .A2(n_186), .B(n_203), .Y(n_304) );
HB1xp67_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
NOR2xp33_ASAP7_75t_SL g203 ( .A(n_184), .B(n_204), .Y(n_203) );
INVx2_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_187), .B(n_197), .Y(n_186) );
AOI22xp5_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_190), .B1(n_193), .B2(n_195), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g190 ( .A(n_191), .B(n_192), .Y(n_190) );
NOR3xp33_ASAP7_75t_L g198 ( .A(n_191), .B(n_192), .C(n_199), .Y(n_198) );
INVx2_ASAP7_75t_L g220 ( .A(n_191), .Y(n_220) );
INVx2_ASAP7_75t_L g234 ( .A(n_191), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_192), .B(n_196), .Y(n_195) );
NOR3xp33_ASAP7_75t_L g200 ( .A(n_192), .B(n_196), .C(n_201), .Y(n_200) );
INVx2_ASAP7_75t_L g270 ( .A(n_205), .Y(n_270) );
INVx3_ASAP7_75t_L g312 ( .A(n_205), .Y(n_312) );
INVx1_ASAP7_75t_L g327 ( .A(n_205), .Y(n_327) );
AND2x2_ASAP7_75t_L g332 ( .A(n_205), .B(n_274), .Y(n_332) );
INVx3_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
OAI21x1_ASAP7_75t_L g206 ( .A1(n_207), .A2(n_209), .B(n_221), .Y(n_206) );
OAI21x1_ASAP7_75t_L g225 ( .A1(n_207), .A2(n_226), .B(n_241), .Y(n_225) );
BUFx3_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_212), .B(n_213), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_213), .A2(n_237), .B(n_238), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g254 ( .A1(n_213), .A2(n_255), .B(n_257), .Y(n_254) );
O2A1O1Ixp5_ASAP7_75t_L g214 ( .A1(n_215), .A2(n_216), .B(n_218), .C(n_220), .Y(n_214) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
NOR2x1p5_ASAP7_75t_L g305 ( .A(n_222), .B(n_306), .Y(n_305) );
INVx2_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
OR2x2_ASAP7_75t_L g463 ( .A(n_223), .B(n_433), .Y(n_463) );
INVx1_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
HB1xp67_ASAP7_75t_L g267 ( .A(n_224), .Y(n_267) );
INVx3_ASAP7_75t_L g317 ( .A(n_224), .Y(n_317) );
INVx2_ASAP7_75t_L g334 ( .A(n_224), .Y(n_334) );
AND2x2_ASAP7_75t_L g340 ( .A(n_224), .B(n_303), .Y(n_340) );
AND2x2_ASAP7_75t_L g363 ( .A(n_224), .B(n_274), .Y(n_363) );
AND2x2_ASAP7_75t_L g392 ( .A(n_224), .B(n_304), .Y(n_392) );
INVx1_ASAP7_75t_L g461 ( .A(n_224), .Y(n_461) );
BUFx6f_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
OAI21x1_ASAP7_75t_L g226 ( .A1(n_227), .A2(n_236), .B(n_240), .Y(n_226) );
OAI21xp5_ASAP7_75t_L g227 ( .A1(n_228), .A2(n_230), .B(n_231), .Y(n_227) );
INVxp67_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
INVxp67_ASAP7_75t_L g283 ( .A(n_229), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_232), .B(n_235), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_233), .B(n_234), .Y(n_232) );
OAI21x1_ASAP7_75t_L g248 ( .A1(n_240), .A2(n_249), .B(n_254), .Y(n_248) );
INVx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
OR2x2_ASAP7_75t_L g243 ( .A(n_244), .B(n_259), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
AND2x2_ASAP7_75t_L g293 ( .A(n_245), .B(n_294), .Y(n_293) );
BUFx3_ASAP7_75t_L g354 ( .A(n_245), .Y(n_354) );
AND2x4_ASAP7_75t_L g373 ( .A(n_245), .B(n_298), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_245), .B(n_379), .Y(n_378) );
INVx2_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
HB1xp67_ASAP7_75t_L g495 ( .A(n_246), .Y(n_495) );
OAI21x1_ASAP7_75t_L g246 ( .A1(n_247), .A2(n_248), .B(n_258), .Y(n_246) );
OAI21x1_ASAP7_75t_L g274 ( .A1(n_247), .A2(n_275), .B(n_286), .Y(n_274) );
OAI21x1_ASAP7_75t_L g297 ( .A1(n_247), .A2(n_248), .B(n_258), .Y(n_297) );
INVx2_ASAP7_75t_L g280 ( .A(n_256), .Y(n_280) );
OR2x2_ASAP7_75t_L g414 ( .A(n_259), .B(n_415), .Y(n_414) );
OR2x2_ASAP7_75t_L g468 ( .A(n_259), .B(n_354), .Y(n_468) );
INVx2_ASAP7_75t_SL g486 ( .A(n_259), .Y(n_486) );
AND2x2_ASAP7_75t_L g368 ( .A(n_260), .B(n_297), .Y(n_368) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVxp67_ASAP7_75t_SL g321 ( .A(n_261), .Y(n_321) );
INVx2_ASAP7_75t_L g380 ( .A(n_261), .Y(n_380) );
INVx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
INVx1_ASAP7_75t_SL g264 ( .A(n_265), .Y(n_264) );
OR2x2_ASAP7_75t_L g265 ( .A(n_266), .B(n_268), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
NAND4xp25_ASAP7_75t_L g502 ( .A(n_267), .B(n_344), .C(n_423), .D(n_503), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_269), .B(n_271), .Y(n_268) );
NAND2xp5_ASAP7_75t_SL g497 ( .A(n_269), .B(n_363), .Y(n_497) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_270), .B(n_317), .Y(n_316) );
NOR2xp67_ASAP7_75t_L g375 ( .A(n_270), .B(n_352), .Y(n_375) );
NOR2x1_ASAP7_75t_L g454 ( .A(n_270), .B(n_303), .Y(n_454) );
AND2x2_ASAP7_75t_L g374 ( .A(n_271), .B(n_375), .Y(n_374) );
INVx2_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
OR2x2_ASAP7_75t_L g315 ( .A(n_272), .B(n_316), .Y(n_315) );
NOR5xp2_ASAP7_75t_L g404 ( .A(n_273), .B(n_405), .C(n_406), .D(n_408), .E(n_409), .Y(n_404) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AND2x4_ASAP7_75t_L g386 ( .A(n_274), .B(n_312), .Y(n_386) );
INVx2_ASAP7_75t_L g308 ( .A(n_275), .Y(n_308) );
OAI22x1_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_279), .B1(n_280), .B2(n_281), .Y(n_276) );
INVxp67_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
AO31x2_ASAP7_75t_L g307 ( .A1(n_287), .A2(n_308), .A3(n_309), .B(n_310), .Y(n_307) );
AO31x2_ASAP7_75t_L g339 ( .A1(n_287), .A2(n_308), .A3(n_309), .B(n_310), .Y(n_339) );
AOI22xp5_ASAP7_75t_L g288 ( .A1(n_289), .A2(n_299), .B1(n_313), .B2(n_314), .Y(n_288) );
NAND3xp33_ASAP7_75t_L g289 ( .A(n_290), .B(n_292), .C(n_295), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NAND2x1p5_ASAP7_75t_L g485 ( .A(n_291), .B(n_486), .Y(n_485) );
OR2x2_ASAP7_75t_L g482 ( .A(n_292), .B(n_345), .Y(n_482) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_293), .Y(n_313) );
AND2x2_ASAP7_75t_L g396 ( .A(n_293), .B(n_361), .Y(n_396) );
AND2x2_ASAP7_75t_L g432 ( .A(n_293), .B(n_433), .Y(n_432) );
AND2x4_ASAP7_75t_L g344 ( .A(n_294), .B(n_297), .Y(n_344) );
HB1xp67_ASAP7_75t_L g395 ( .A(n_294), .Y(n_395) );
INVx1_ASAP7_75t_L g407 ( .A(n_294), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_294), .B(n_380), .Y(n_448) );
OAI22xp33_ASAP7_75t_SL g471 ( .A1(n_295), .A2(n_296), .B1(n_315), .B2(n_384), .Y(n_471) );
OAI22xp5_ASAP7_75t_L g487 ( .A1(n_295), .A2(n_330), .B1(n_425), .B2(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g348 ( .A(n_296), .B(n_349), .Y(n_348) );
AND2x4_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
AND2x4_ASAP7_75t_L g435 ( .A(n_297), .B(n_423), .Y(n_435) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_301), .B(n_305), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g326 ( .A(n_302), .B(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_302), .B(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_303), .B(n_312), .Y(n_365) );
BUFx2_ASAP7_75t_L g408 ( .A(n_303), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_303), .B(n_461), .Y(n_460) );
INVx3_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
AOI22xp33_ASAP7_75t_L g371 ( .A1(n_305), .A2(n_372), .B1(n_374), .B2(n_376), .Y(n_371) );
INVx1_ASAP7_75t_L g384 ( .A(n_305), .Y(n_384) );
HB1xp67_ASAP7_75t_L g465 ( .A(n_306), .Y(n_465) );
OR2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_312), .Y(n_306) );
OR2x2_ASAP7_75t_L g329 ( .A(n_307), .B(n_317), .Y(n_329) );
AND2x2_ASAP7_75t_L g507 ( .A(n_310), .B(n_508), .Y(n_507) );
BUFx2_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
AO21x1_ASAP7_75t_L g412 ( .A1(n_316), .A2(n_413), .B(n_416), .Y(n_412) );
INVx2_ASAP7_75t_L g352 ( .A(n_317), .Y(n_352) );
AOI22xp5_ASAP7_75t_L g318 ( .A1(n_319), .A2(n_323), .B1(n_335), .B2(n_341), .Y(n_318) );
BUFx3_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_320), .B(n_354), .Y(n_474) );
AND2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
BUFx2_ASAP7_75t_L g349 ( .A(n_322), .Y(n_349) );
INVx1_ASAP7_75t_L g356 ( .A(n_322), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_324), .B(n_330), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
AOI221xp5_ASAP7_75t_L g490 ( .A1(n_325), .A2(n_491), .B1(n_492), .B2(n_496), .C(n_500), .Y(n_490) );
AND2x4_ASAP7_75t_L g325 ( .A(n_326), .B(n_328), .Y(n_325) );
INVx1_ASAP7_75t_L g504 ( .A(n_327), .Y(n_504) );
INVx2_ASAP7_75t_SL g328 ( .A(n_329), .Y(n_328) );
OR2x2_ASAP7_75t_L g370 ( .A(n_329), .B(n_365), .Y(n_370) );
INVx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g331 ( .A(n_332), .B(n_333), .Y(n_331) );
INVx1_ASAP7_75t_L g357 ( .A(n_332), .Y(n_357) );
AND2x2_ASAP7_75t_L g443 ( .A(n_332), .B(n_392), .Y(n_443) );
AND2x2_ASAP7_75t_L g355 ( .A(n_333), .B(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g420 ( .A(n_333), .B(n_337), .Y(n_420) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_337), .B(n_340), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g391 ( .A(n_338), .B(n_392), .Y(n_391) );
INVx2_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
BUFx3_ASAP7_75t_L g403 ( .A(n_339), .Y(n_403) );
INVxp67_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
OR2x2_ASAP7_75t_L g342 ( .A(n_343), .B(n_345), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
NOR2xp33_ASAP7_75t_L g359 ( .A(n_344), .B(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g388 ( .A(n_344), .B(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g399 ( .A(n_344), .Y(n_399) );
NOR2x1_ASAP7_75t_L g421 ( .A(n_344), .B(n_422), .Y(n_421) );
AND2x2_ASAP7_75t_L g491 ( .A(n_344), .B(n_349), .Y(n_491) );
INVx2_ASAP7_75t_L g429 ( .A(n_345), .Y(n_429) );
OAI211xp5_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_357), .B(n_358), .C(n_371), .Y(n_346) );
AOI21xp5_ASAP7_75t_L g347 ( .A1(n_348), .A2(n_350), .B(n_353), .Y(n_347) );
AND2x2_ASAP7_75t_L g372 ( .A(n_349), .B(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
BUFx2_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
OR2x2_ASAP7_75t_L g450 ( .A(n_352), .B(n_451), .Y(n_450) );
AND2x2_ASAP7_75t_L g353 ( .A(n_354), .B(n_355), .Y(n_353) );
OR2x2_ASAP7_75t_L g413 ( .A(n_354), .B(n_414), .Y(n_413) );
OR2x2_ASAP7_75t_L g377 ( .A(n_356), .B(n_378), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_356), .B(n_417), .Y(n_416) );
HB1xp67_ASAP7_75t_L g472 ( .A(n_356), .Y(n_472) );
AOI22xp33_ASAP7_75t_L g358 ( .A1(n_359), .A2(n_362), .B1(n_366), .B2(n_369), .Y(n_358) );
OR2x2_ASAP7_75t_L g493 ( .A(n_360), .B(n_494), .Y(n_493) );
INVx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
AND2x4_ASAP7_75t_L g362 ( .A(n_363), .B(n_364), .Y(n_362) );
INVx1_ASAP7_75t_L g489 ( .A(n_363), .Y(n_489) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
OR2x2_ASAP7_75t_L g402 ( .A(n_365), .B(n_403), .Y(n_402) );
HB1xp67_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
HB1xp67_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g394 ( .A(n_368), .B(n_395), .Y(n_394) );
AOI221xp5_ASAP7_75t_L g419 ( .A1(n_369), .A2(n_420), .B1(n_421), .B2(n_424), .C(n_430), .Y(n_419) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_373), .B(n_429), .Y(n_428) );
INVx3_ASAP7_75t_R g464 ( .A(n_373), .Y(n_464) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
HB1xp67_ASAP7_75t_L g389 ( .A(n_379), .Y(n_389) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
HB1xp67_ASAP7_75t_L g409 ( .A(n_380), .Y(n_409) );
OAI221xp5_ASAP7_75t_L g381 ( .A1(n_382), .A2(n_387), .B1(n_390), .B2(n_393), .C(n_397), .Y(n_381) );
INVxp67_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_384), .B(n_385), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_386), .B(n_392), .Y(n_436) );
AND2x2_ASAP7_75t_L g440 ( .A(n_386), .B(n_408), .Y(n_440) );
OAI32xp33_ASAP7_75t_L g457 ( .A1(n_386), .A2(n_418), .A3(n_431), .B1(n_453), .B2(n_458), .Y(n_457) );
AND2x2_ASAP7_75t_L g478 ( .A(n_386), .B(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVxp67_ASAP7_75t_SL g400 ( .A(n_389), .Y(n_400) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
AOI221x1_ASAP7_75t_L g480 ( .A1(n_391), .A2(n_481), .B1(n_483), .B2(n_484), .C(n_487), .Y(n_480) );
AND2x2_ASAP7_75t_L g483 ( .A(n_392), .B(n_403), .Y(n_483) );
NOR2xp33_ASAP7_75t_SL g393 ( .A(n_394), .B(n_396), .Y(n_393) );
AOI321xp33_ASAP7_75t_L g397 ( .A1(n_394), .A2(n_398), .A3(n_399), .B1(n_400), .B2(n_401), .C(n_404), .Y(n_397) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
OAI21xp33_ASAP7_75t_L g500 ( .A1(n_402), .A2(n_501), .B(n_502), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_403), .B(n_454), .Y(n_453) );
OR2x2_ASAP7_75t_L g469 ( .A(n_403), .B(n_460), .Y(n_469) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
NOR2x1_ASAP7_75t_L g410 ( .A(n_411), .B(n_455), .Y(n_410) );
NAND3xp33_ASAP7_75t_SL g411 ( .A(n_412), .B(n_419), .C(n_437), .Y(n_411) );
OR2x2_ASAP7_75t_L g501 ( .A(n_415), .B(n_448), .Y(n_501) );
INVx3_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_425), .B(n_428), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
NAND2xp5_ASAP7_75t_SL g466 ( .A(n_427), .B(n_433), .Y(n_466) );
INVx1_ASAP7_75t_L g449 ( .A(n_429), .Y(n_449) );
AOI21xp33_ASAP7_75t_L g430 ( .A1(n_431), .A2(n_434), .B(n_436), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g446 ( .A(n_433), .Y(n_446) );
INVx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
AOI211xp5_ASAP7_75t_L g437 ( .A1(n_438), .A2(n_440), .B(n_441), .C(n_452), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
OAI22xp5_ASAP7_75t_L g441 ( .A1(n_442), .A2(n_444), .B1(n_449), .B2(n_450), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
AND2x4_ASAP7_75t_L g445 ( .A(n_446), .B(n_447), .Y(n_445) );
INVx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
HB1xp67_ASAP7_75t_SL g467 ( .A(n_451), .Y(n_467) );
OR2x2_ASAP7_75t_L g488 ( .A(n_451), .B(n_489), .Y(n_488) );
NAND4xp25_ASAP7_75t_L g455 ( .A(n_456), .B(n_470), .C(n_480), .D(n_490), .Y(n_455) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_457), .B(n_462), .Y(n_456) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVxp67_ASAP7_75t_SL g479 ( .A(n_460), .Y(n_479) );
OAI322xp33_ASAP7_75t_L g462 ( .A1(n_463), .A2(n_464), .A3(n_465), .B1(n_466), .B2(n_467), .C1(n_468), .C2(n_469), .Y(n_462) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_472), .B(n_473), .Y(n_470) );
AOI21xp33_ASAP7_75t_L g473 ( .A1(n_474), .A2(n_475), .B(n_477), .Y(n_473) );
INVx2_ASAP7_75t_SL g475 ( .A(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_497), .B(n_498), .Y(n_496) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
CKINVDCx6p67_ASAP7_75t_R g505 ( .A(n_506), .Y(n_505) );
CKINVDCx20_ASAP7_75t_R g506 ( .A(n_507), .Y(n_506) );
INVxp67_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
AO21x2_ASAP7_75t_L g748 ( .A1(n_509), .A2(n_736), .B(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
OAI221xp5_ASAP7_75t_L g512 ( .A1(n_513), .A2(n_704), .B1(n_727), .B2(n_729), .C(n_738), .Y(n_512) );
AOI22xp5_ASAP7_75t_L g513 ( .A1(n_514), .A2(n_680), .B1(n_681), .B2(n_703), .Y(n_513) );
INVx1_ASAP7_75t_L g703 ( .A(n_514), .Y(n_703) );
XOR2xp5_ASAP7_75t_L g742 ( .A(n_514), .B(n_743), .Y(n_742) );
HB1xp67_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
AOI211xp5_ASAP7_75t_L g515 ( .A1(n_516), .A2(n_522), .B(n_596), .C(n_655), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
CKINVDCx5p33_ASAP7_75t_R g517 ( .A(n_518), .Y(n_517) );
BUFx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
AND2x6_ASAP7_75t_L g638 ( .A(n_520), .B(n_639), .Y(n_638) );
INVx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g602 ( .A(n_521), .Y(n_602) );
OR2x2_ASAP7_75t_L g647 ( .A(n_521), .B(n_648), .Y(n_647) );
NAND5xp2_ASAP7_75t_SL g522 ( .A(n_523), .B(n_540), .C(n_550), .D(n_580), .E(n_586), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_524), .A2(n_525), .B1(n_534), .B2(n_535), .Y(n_523) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
OR2x2_ASAP7_75t_L g526 ( .A(n_527), .B(n_530), .Y(n_526) );
INVx1_ASAP7_75t_L g536 ( .A(n_527), .Y(n_536) );
INVx1_ASAP7_75t_L g584 ( .A(n_527), .Y(n_584) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
AND2x2_ASAP7_75t_L g569 ( .A(n_529), .B(n_570), .Y(n_569) );
OR2x6_ASAP7_75t_L g543 ( .A(n_530), .B(n_544), .Y(n_543) );
BUFx6f_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_532), .B(n_533), .Y(n_531) );
AND2x4_ASAP7_75t_L g538 ( .A(n_532), .B(n_539), .Y(n_538) );
INVx2_ASAP7_75t_L g562 ( .A(n_532), .Y(n_562) );
INVx2_ASAP7_75t_L g539 ( .A(n_533), .Y(n_539) );
INVx2_ASAP7_75t_L g561 ( .A(n_533), .Y(n_561) );
AND2x2_ASAP7_75t_L g535 ( .A(n_536), .B(n_537), .Y(n_535) );
AND2x4_ASAP7_75t_L g547 ( .A(n_536), .B(n_548), .Y(n_547) );
INVx2_ASAP7_75t_L g574 ( .A(n_537), .Y(n_574) );
BUFx6f_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx5_ASAP7_75t_L g557 ( .A(n_538), .Y(n_557) );
INVx1_ASAP7_75t_L g567 ( .A(n_539), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_541), .A2(n_542), .B1(n_546), .B2(n_547), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g643 ( .A1(n_541), .A2(n_593), .B1(n_644), .B2(n_652), .Y(n_643) );
CKINVDCx14_ASAP7_75t_R g542 ( .A(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g595 ( .A(n_544), .Y(n_595) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
AND2x2_ASAP7_75t_L g587 ( .A(n_545), .B(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g590 ( .A(n_545), .B(n_591), .Y(n_590) );
BUFx4f_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
BUFx3_ASAP7_75t_L g554 ( .A(n_549), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_551), .A2(n_558), .B1(n_571), .B2(n_575), .Y(n_550) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx3_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
BUFx3_ASAP7_75t_L g572 ( .A(n_554), .Y(n_572) );
HB1xp67_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx3_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
BUFx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
BUFx2_ASAP7_75t_L g577 ( .A(n_560), .Y(n_577) );
BUFx4f_ASAP7_75t_L g585 ( .A(n_560), .Y(n_585) );
AND2x2_ASAP7_75t_L g594 ( .A(n_560), .B(n_595), .Y(n_594) );
AND2x4_ASAP7_75t_L g560 ( .A(n_561), .B(n_562), .Y(n_560) );
BUFx3_ASAP7_75t_L g588 ( .A(n_561), .Y(n_588) );
INVx1_ASAP7_75t_L g592 ( .A(n_562), .Y(n_592) );
INVx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx5_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
BUFx2_ASAP7_75t_L g576 ( .A(n_565), .Y(n_576) );
AND2x4_ASAP7_75t_L g565 ( .A(n_566), .B(n_567), .Y(n_565) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
BUFx4_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_581), .B(n_582), .Y(n_580) );
OAI22xp33_ASAP7_75t_L g673 ( .A1(n_581), .A2(n_624), .B1(n_674), .B2(n_675), .Y(n_673) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
NAND2x1p5_ASAP7_75t_L g583 ( .A(n_584), .B(n_585), .Y(n_583) );
AOI221xp5_ASAP7_75t_L g586 ( .A1(n_587), .A2(n_589), .B1(n_590), .B2(n_593), .C(n_594), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_589), .A2(n_598), .B1(n_610), .B2(n_611), .Y(n_597) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
NAND3xp33_ASAP7_75t_L g596 ( .A(n_597), .B(n_616), .C(n_643), .Y(n_596) );
INVx2_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_601), .B(n_607), .Y(n_600) );
AND2x4_ASAP7_75t_L g611 ( .A(n_601), .B(n_612), .Y(n_611) );
AND2x4_ASAP7_75t_L g642 ( .A(n_601), .B(n_625), .Y(n_642) );
INVx2_ASAP7_75t_L g679 ( .A(n_601), .Y(n_679) );
AND2x4_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .Y(n_601) );
AND2x6_ASAP7_75t_L g667 ( .A(n_602), .B(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g726 ( .A(n_603), .Y(n_726) );
AND2x2_ASAP7_75t_L g603 ( .A(n_604), .B(n_605), .Y(n_603) );
INVx1_ASAP7_75t_L g641 ( .A(n_604), .Y(n_641) );
OR2x6_ASAP7_75t_L g648 ( .A(n_604), .B(n_606), .Y(n_648) );
AND2x4_ASAP7_75t_L g668 ( .A(n_604), .B(n_640), .Y(n_668) );
OR2x2_ASAP7_75t_L g718 ( .A(n_604), .B(n_605), .Y(n_718) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
BUFx2_ASAP7_75t_L g640 ( .A(n_606), .Y(n_640) );
INVx2_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
HB1xp67_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
AND2x4_ASAP7_75t_L g661 ( .A(n_609), .B(n_615), .Y(n_661) );
INVx1_ASAP7_75t_L g716 ( .A(n_609), .Y(n_716) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
AND2x4_ASAP7_75t_L g637 ( .A(n_615), .B(n_627), .Y(n_637) );
AOI31xp33_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_629), .A3(n_638), .B(n_642), .Y(n_616) );
INVx5_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g620 ( .A(n_621), .B(n_622), .Y(n_620) );
INVx2_ASAP7_75t_L g627 ( .A(n_621), .Y(n_627) );
AND2x2_ASAP7_75t_L g633 ( .A(n_621), .B(n_628), .Y(n_633) );
INVx2_ASAP7_75t_L g628 ( .A(n_622), .Y(n_628) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx2_ASAP7_75t_SL g624 ( .A(n_625), .Y(n_624) );
BUFx6f_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
BUFx6f_ASAP7_75t_L g654 ( .A(n_626), .Y(n_654) );
AND2x4_ASAP7_75t_L g626 ( .A(n_627), .B(n_628), .Y(n_626) );
HB1xp67_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
BUFx12f_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
BUFx6f_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx3_ASAP7_75t_L g665 ( .A(n_633), .Y(n_665) );
INVx2_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx2_ASAP7_75t_SL g635 ( .A(n_636), .Y(n_635) );
BUFx6f_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
BUFx3_ASAP7_75t_L g651 ( .A(n_637), .Y(n_651) );
BUFx12f_ASAP7_75t_L g672 ( .A(n_637), .Y(n_672) );
AND2x2_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .Y(n_639) );
BUFx2_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
AND2x4_ASAP7_75t_L g645 ( .A(n_646), .B(n_649), .Y(n_645) );
AND2x2_ASAP7_75t_L g652 ( .A(n_646), .B(n_653), .Y(n_652) );
AND2x2_ASAP7_75t_L g663 ( .A(n_646), .B(n_664), .Y(n_663) );
INVx2_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
OR2x6_ASAP7_75t_L g659 ( .A(n_647), .B(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
BUFx6f_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_656), .B(n_666), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g656 ( .A1(n_657), .A2(n_658), .B1(n_662), .B2(n_663), .Y(n_656) );
CKINVDCx5p33_ASAP7_75t_R g658 ( .A(n_659), .Y(n_658) );
BUFx3_ASAP7_75t_L g675 ( .A(n_660), .Y(n_675) );
OR2x2_ASAP7_75t_L g678 ( .A(n_660), .B(n_679), .Y(n_678) );
INVx8_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx5_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_669), .B1(n_676), .B2(n_677), .Y(n_666) );
INVxp67_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx2_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
CKINVDCx14_ASAP7_75t_R g680 ( .A(n_681), .Y(n_680) );
AOI22xp5_ASAP7_75t_L g681 ( .A1(n_682), .A2(n_683), .B1(n_693), .B2(n_702), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
XNOR2xp5_ASAP7_75t_L g683 ( .A(n_684), .B(n_689), .Y(n_683) );
AOI22xp5_ASAP7_75t_L g684 ( .A1(n_685), .A2(n_686), .B1(n_687), .B2(n_688), .Y(n_684) );
INVx1_ASAP7_75t_SL g688 ( .A(n_685), .Y(n_688) );
INVx2_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g692 ( .A(n_691), .Y(n_692) );
INVx1_ASAP7_75t_L g702 ( .A(n_693), .Y(n_702) );
OAI22xp5_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_699), .B1(n_700), .B2(n_701), .Y(n_693) );
INVx1_ASAP7_75t_L g700 ( .A(n_694), .Y(n_700) );
OAI22xp5_ASAP7_75t_L g694 ( .A1(n_695), .A2(n_696), .B1(n_697), .B2(n_698), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g701 ( .A(n_699), .Y(n_701) );
BUFx2_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx5_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
AND2x6_ASAP7_75t_L g706 ( .A(n_707), .B(n_719), .Y(n_706) );
NOR2xp33_ASAP7_75t_L g707 ( .A(n_708), .B(n_712), .Y(n_707) );
INVxp67_ASAP7_75t_L g740 ( .A(n_708), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_709), .B(n_710), .Y(n_708) );
INVx1_ASAP7_75t_L g737 ( .A(n_709), .Y(n_737) );
INVx1_ASAP7_75t_L g750 ( .A(n_710), .Y(n_750) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
BUFx2_ASAP7_75t_L g736 ( .A(n_711), .Y(n_736) );
INVxp67_ASAP7_75t_SL g712 ( .A(n_713), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_713), .B(n_723), .Y(n_741) );
NAND3xp33_ASAP7_75t_L g713 ( .A(n_714), .B(n_716), .C(n_717), .Y(n_713) );
INVx2_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
CKINVDCx11_ASAP7_75t_R g721 ( .A(n_715), .Y(n_721) );
AND2x4_ASAP7_75t_L g724 ( .A(n_716), .B(n_725), .Y(n_724) );
BUFx6f_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_720), .B(n_722), .Y(n_719) );
CKINVDCx5p33_ASAP7_75t_R g720 ( .A(n_721), .Y(n_720) );
INVx2_ASAP7_75t_SL g722 ( .A(n_723), .Y(n_722) );
INVx2_ASAP7_75t_SL g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
CKINVDCx20_ASAP7_75t_R g729 ( .A(n_730), .Y(n_729) );
CKINVDCx20_ASAP7_75t_R g730 ( .A(n_731), .Y(n_730) );
INVx3_ASAP7_75t_SL g731 ( .A(n_732), .Y(n_731) );
CKINVDCx20_ASAP7_75t_R g732 ( .A(n_733), .Y(n_732) );
BUFx6f_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_735), .B(n_737), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
AND2x2_ASAP7_75t_L g749 ( .A(n_737), .B(n_750), .Y(n_749) );
AOI22xp5_ASAP7_75t_L g738 ( .A1(n_739), .A2(n_742), .B1(n_745), .B2(n_746), .Y(n_738) );
AND2x2_ASAP7_75t_L g739 ( .A(n_740), .B(n_741), .Y(n_739) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
CKINVDCx20_ASAP7_75t_R g746 ( .A(n_747), .Y(n_746) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_748), .Y(n_747) );
endmodule