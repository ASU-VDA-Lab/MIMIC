module fake_jpeg_29964_n_64 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_64);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_64;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_6),
.B(n_16),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

OA22x2_ASAP7_75t_L g30 ( 
.A1(n_27),
.A2(n_21),
.B1(n_20),
.B2(n_17),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_30),
.A2(n_22),
.B1(n_24),
.B2(n_23),
.Y(n_36)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_22),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_29),
.Y(n_37)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVxp67_ASAP7_75t_SL g42 ( 
.A(n_34),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_25),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_35),
.A2(n_24),
.B1(n_28),
.B2(n_3),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_37),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_SL g48 ( 
.A1(n_38),
.A2(n_30),
.B(n_39),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_31),
.A2(n_13),
.B1(n_12),
.B2(n_10),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_40),
.A2(n_34),
.B1(n_4),
.B2(n_5),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_1),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_2),
.Y(n_49)
);

AO21x1_ASAP7_75t_L g44 ( 
.A1(n_36),
.A2(n_30),
.B(n_33),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_44),
.A2(n_8),
.B1(n_3),
.B2(n_7),
.Y(n_55)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_49),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_30),
.C(n_34),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_9),
.C(n_7),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_48),
.A2(n_8),
.B1(n_47),
.B2(n_46),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_50),
.A2(n_40),
.B1(n_5),
.B2(n_6),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_42),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_51),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g60 ( 
.A(n_52),
.B(n_55),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g59 ( 
.A(n_53),
.B(n_57),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_54),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_58),
.B(n_56),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_61),
.B(n_46),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g63 ( 
.A1(n_62),
.A2(n_53),
.B(n_44),
.Y(n_63)
);

AOI221xp5_ASAP7_75t_L g64 ( 
.A1(n_63),
.A2(n_52),
.B1(n_59),
.B2(n_60),
.C(n_57),
.Y(n_64)
);


endmodule