module fake_aes_6420_n_25 (n_11, n_1, n_2, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_25);
input n_11;
input n_1;
input n_2;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_25;
wire n_20;
wire n_23;
wire n_22;
wire n_16;
wire n_13;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
INVx1_ASAP7_75t_L g13 ( .A(n_0), .Y(n_13) );
CKINVDCx16_ASAP7_75t_R g14 ( .A(n_4), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_3), .Y(n_15) );
BUFx10_ASAP7_75t_L g16 ( .A(n_10), .Y(n_16) );
AOI21x1_ASAP7_75t_SL g17 ( .A1(n_16), .A2(n_0), .B(n_1), .Y(n_17) );
NAND2xp5_ASAP7_75t_L g18 ( .A(n_13), .B(n_1), .Y(n_18) );
NAND3xp33_ASAP7_75t_L g19 ( .A(n_18), .B(n_15), .C(n_14), .Y(n_19) );
AND2x4_ASAP7_75t_L g20 ( .A(n_19), .B(n_2), .Y(n_20) );
AND2x2_ASAP7_75t_L g21 ( .A(n_20), .B(n_16), .Y(n_21) );
O2A1O1Ixp5_ASAP7_75t_L g22 ( .A1(n_21), .A2(n_20), .B(n_17), .C(n_7), .Y(n_22) );
CKINVDCx5p33_ASAP7_75t_R g23 ( .A(n_22), .Y(n_23) );
AO22x2_ASAP7_75t_L g24 ( .A1(n_23), .A2(n_5), .B1(n_6), .B2(n_8), .Y(n_24) );
AOI22xp33_ASAP7_75t_L g25 ( .A1(n_24), .A2(n_9), .B1(n_11), .B2(n_12), .Y(n_25) );
endmodule