module fake_jpeg_1813_n_189 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_189);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_189;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_4),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_14),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_32),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_14),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_7),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_12),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_44),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_63),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_71),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_70),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_47),
.B(n_48),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_0),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_73),
.B(n_57),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_77),
.B(n_57),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_72),
.A2(n_64),
.B1(n_62),
.B2(n_60),
.Y(n_78)
);

AOI32xp33_ASAP7_75t_L g97 ( 
.A1(n_78),
.A2(n_65),
.A3(n_66),
.B1(n_70),
.B2(n_58),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_68),
.A2(n_64),
.B1(n_59),
.B2(n_51),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_80),
.A2(n_68),
.B1(n_72),
.B2(n_51),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_69),
.A2(n_58),
.B1(n_49),
.B2(n_55),
.Y(n_82)
);

AOI21xp33_ASAP7_75t_L g98 ( 
.A1(n_82),
.A2(n_70),
.B(n_52),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_71),
.B(n_56),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_84),
.B(n_85),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_67),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_88),
.Y(n_108)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_83),
.Y(n_89)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_90),
.A2(n_74),
.B1(n_1),
.B2(n_2),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_85),
.B(n_61),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_94),
.Y(n_109)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_93),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_73),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_54),
.Y(n_94)
);

AO22x2_ASAP7_75t_L g96 ( 
.A1(n_78),
.A2(n_69),
.B1(n_66),
.B2(n_65),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_96),
.A2(n_98),
.B1(n_74),
.B2(n_2),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_97),
.B(n_53),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_52),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_100),
.Y(n_120)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_79),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_83),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_102),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_95),
.B(n_79),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_103),
.B(n_111),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_122),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_90),
.A2(n_81),
.B1(n_79),
.B2(n_74),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_106),
.A2(n_114),
.B1(n_10),
.B2(n_11),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_107),
.A2(n_87),
.B1(n_30),
.B2(n_31),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_94),
.B(n_22),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_112),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_91),
.B(n_0),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_100),
.B(n_24),
.Y(n_112)
);

NOR3xp33_ASAP7_75t_L g115 ( 
.A(n_96),
.B(n_1),
.C(n_3),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_117),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_96),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_116),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_89),
.Y(n_117)
);

AOI32xp33_ASAP7_75t_L g119 ( 
.A1(n_96),
.A2(n_5),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_119),
.A2(n_15),
.B(n_16),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_29),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_124),
.A2(n_131),
.B1(n_138),
.B2(n_139),
.Y(n_154)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_121),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_125),
.B(n_126),
.Y(n_145)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_120),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_105),
.A2(n_8),
.B(n_9),
.Y(n_127)
);

OA21x2_ASAP7_75t_L g149 ( 
.A1(n_127),
.A2(n_104),
.B(n_113),
.Y(n_149)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_108),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_128),
.B(n_133),
.Y(n_150)
);

OA21x2_ASAP7_75t_L g129 ( 
.A1(n_106),
.A2(n_33),
.B(n_43),
.Y(n_129)
);

AO21x2_ASAP7_75t_SL g155 ( 
.A1(n_129),
.A2(n_25),
.B(n_28),
.Y(n_155)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_113),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_118),
.Y(n_135)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_135),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_109),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_136)
);

INVxp67_ASAP7_75t_SL g148 ( 
.A(n_136),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_109),
.A2(n_13),
.B1(n_15),
.B2(n_16),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_110),
.A2(n_34),
.B1(n_42),
.B2(n_18),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_140),
.B(n_20),
.Y(n_153)
);

BUFx2_ASAP7_75t_L g141 ( 
.A(n_104),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_141),
.Y(n_143)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_112),
.Y(n_142)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_142),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_134),
.A2(n_127),
.B1(n_130),
.B2(n_129),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_144),
.A2(n_136),
.B1(n_137),
.B2(n_148),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_123),
.B(n_122),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_146),
.Y(n_167)
);

INVx1_ASAP7_75t_SL g168 ( 
.A(n_149),
.Y(n_168)
);

XOR2x2_ASAP7_75t_L g151 ( 
.A(n_134),
.B(n_19),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_151),
.B(n_157),
.C(n_159),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_153),
.Y(n_163)
);

INVx3_ASAP7_75t_SL g162 ( 
.A(n_155),
.Y(n_162)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_141),
.Y(n_156)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_156),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_130),
.B(n_35),
.C(n_36),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_129),
.A2(n_37),
.B1(n_38),
.B2(n_41),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_158),
.A2(n_155),
.B1(n_159),
.B2(n_148),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_132),
.B(n_45),
.C(n_139),
.Y(n_159)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_161),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_150),
.B(n_152),
.Y(n_164)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_164),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_145),
.B(n_149),
.Y(n_165)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_165),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_169),
.B(n_149),
.Y(n_170)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_170),
.Y(n_177)
);

NOR3xp33_ASAP7_75t_SL g171 ( 
.A(n_167),
.B(n_147),
.C(n_151),
.Y(n_171)
);

NAND4xp25_ASAP7_75t_L g179 ( 
.A(n_171),
.B(n_155),
.C(n_169),
.D(n_164),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_163),
.B(n_143),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_173),
.B(n_174),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_160),
.B(n_144),
.C(n_157),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_175),
.B(n_165),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_178),
.B(n_176),
.C(n_161),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_179),
.A2(n_162),
.B1(n_168),
.B2(n_172),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_181),
.A2(n_182),
.B(n_176),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_183),
.A2(n_180),
.B(n_162),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_184),
.B(n_168),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_185),
.B(n_178),
.Y(n_186)
);

AOI21x1_ASAP7_75t_L g187 ( 
.A1(n_186),
.A2(n_177),
.B(n_160),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_187),
.B(n_154),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_188),
.B(n_166),
.Y(n_189)
);


endmodule