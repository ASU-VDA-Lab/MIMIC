module fake_jpeg_29971_n_421 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_421);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_421;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_19;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_16),
.B(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx6_ASAP7_75t_SL g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_16),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_12),
.B(n_1),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx16f_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_43),
.Y(n_121)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_44),
.Y(n_93)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_45),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_48),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_34),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_49),
.B(n_50),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_25),
.B(n_16),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_34),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_51),
.B(n_53),
.Y(n_107)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_52),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g53 ( 
.A(n_34),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_54),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_55),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_29),
.Y(n_56)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_58),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_59),
.Y(n_103)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_60),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_34),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_61),
.B(n_63),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

INVx3_ASAP7_75t_SL g99 ( 
.A(n_62),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_20),
.B(n_15),
.Y(n_63)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_64),
.Y(n_129)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_65),
.Y(n_128)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_66),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_20),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_67),
.B(n_76),
.Y(n_123)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_68),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g119 ( 
.A(n_69),
.Y(n_119)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_70),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_71),
.Y(n_125)
);

BUFx10_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

INVx5_ASAP7_75t_SL g111 ( 
.A(n_72),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_32),
.Y(n_73)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_73),
.Y(n_131)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_30),
.Y(n_74)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_74),
.Y(n_120)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_30),
.Y(n_75)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_75),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_25),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_77),
.Y(n_135)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_31),
.Y(n_78)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_78),
.Y(n_136)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_33),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_80),
.Y(n_132)
);

NAND2x1_ASAP7_75t_SL g81 ( 
.A(n_23),
.B(n_0),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_81),
.B(n_23),
.Y(n_114)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_38),
.Y(n_82)
);

INVx2_ASAP7_75t_SL g112 ( 
.A(n_82),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_32),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g122 ( 
.A(n_83),
.Y(n_122)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_33),
.Y(n_84)
);

INVx4_ASAP7_75t_SL g98 ( 
.A(n_84),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_50),
.B(n_27),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_86),
.B(n_102),
.Y(n_143)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g173 ( 
.A(n_87),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_81),
.B(n_41),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_88),
.B(n_91),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_72),
.B(n_41),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_24),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_94),
.B(n_97),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_74),
.A2(n_35),
.B1(n_27),
.B2(n_18),
.Y(n_95)
);

OA22x2_ASAP7_75t_L g169 ( 
.A1(n_95),
.A2(n_22),
.B1(n_36),
.B2(n_17),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_71),
.A2(n_32),
.B1(n_35),
.B2(n_18),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_57),
.B(n_24),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_80),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_104),
.Y(n_165)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_60),
.Y(n_110)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_110),
.Y(n_147)
);

BUFx5_ASAP7_75t_L g113 ( 
.A(n_46),
.Y(n_113)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_113),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_114),
.A2(n_28),
.B(n_39),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_58),
.B(n_28),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_117),
.B(n_124),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_82),
.B(n_39),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_59),
.B(n_39),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_127),
.B(n_130),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_75),
.B(n_28),
.Y(n_130)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_116),
.Y(n_138)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_138),
.Y(n_176)
);

CKINVDCx9p33_ASAP7_75t_R g139 ( 
.A(n_111),
.Y(n_139)
);

CKINVDCx14_ASAP7_75t_R g192 ( 
.A(n_139),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_140),
.Y(n_187)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_92),
.Y(n_142)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_142),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_111),
.A2(n_36),
.B1(n_22),
.B2(n_70),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_145),
.A2(n_149),
.B1(n_162),
.B2(n_170),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_123),
.B(n_38),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_146),
.B(n_151),
.Y(n_174)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_128),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_101),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_150),
.Y(n_188)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_133),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_121),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_152),
.B(n_153),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_123),
.B(n_38),
.Y(n_153)
);

CKINVDCx12_ASAP7_75t_R g154 ( 
.A(n_107),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_154),
.Y(n_194)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_135),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_155),
.B(n_160),
.Y(n_181)
);

A2O1A1O1Ixp25_ASAP7_75t_L g157 ( 
.A1(n_105),
.A2(n_36),
.B(n_22),
.C(n_17),
.D(n_38),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_157),
.B(n_166),
.Y(n_179)
);

CKINVDCx12_ASAP7_75t_R g158 ( 
.A(n_107),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_158),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_R g159 ( 
.A(n_114),
.B(n_40),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_159),
.B(n_167),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_118),
.Y(n_160)
);

INVx8_ASAP7_75t_L g162 ( 
.A(n_128),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_126),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_163),
.B(n_164),
.Y(n_193)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_106),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_124),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_136),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_115),
.B(n_105),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_168),
.B(n_169),
.Y(n_186)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_125),
.Y(n_170)
);

CKINVDCx12_ASAP7_75t_R g171 ( 
.A(n_87),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_171),
.B(n_172),
.Y(n_190)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_131),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_144),
.A2(n_156),
.B1(n_159),
.B2(n_169),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_180),
.A2(n_183),
.B1(n_98),
.B2(n_73),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_144),
.A2(n_129),
.B1(n_64),
.B2(n_44),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_148),
.B(n_115),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_185),
.B(n_189),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_148),
.B(n_127),
.C(n_120),
.Y(n_189)
);

OAI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_169),
.A2(n_129),
.B1(n_119),
.B2(n_96),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_191),
.A2(n_119),
.B1(n_98),
.B2(n_151),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_169),
.A2(n_17),
.B(n_112),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_195),
.B(n_99),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_174),
.B(n_143),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_196),
.B(n_202),
.Y(n_229)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_193),
.Y(n_197)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_197),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_195),
.A2(n_139),
.B1(n_96),
.B2(n_134),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_198),
.A2(n_203),
.B1(n_192),
.B2(n_177),
.Y(n_217)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_193),
.Y(n_200)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_200),
.Y(n_219)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_181),
.Y(n_201)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_201),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_186),
.B(n_150),
.Y(n_202)
);

INVx5_ASAP7_75t_L g204 ( 
.A(n_176),
.Y(n_204)
);

BUFx2_ASAP7_75t_L g233 ( 
.A(n_204),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_186),
.B(n_141),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_205),
.B(n_206),
.Y(n_230)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_176),
.Y(n_207)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_207),
.Y(n_220)
);

INVx13_ASAP7_75t_L g208 ( 
.A(n_192),
.Y(n_208)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_208),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_209),
.A2(n_182),
.B(n_177),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_185),
.B(n_140),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_210),
.B(n_211),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_180),
.A2(n_195),
.B1(n_186),
.B2(n_183),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_185),
.B(n_157),
.Y(n_212)
);

BUFx24_ASAP7_75t_SL g237 ( 
.A(n_212),
.Y(n_237)
);

AOI21xp33_ASAP7_75t_L g213 ( 
.A1(n_179),
.A2(n_147),
.B(n_173),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_213),
.B(n_182),
.Y(n_234)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_178),
.Y(n_214)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_214),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_179),
.B(n_38),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_215),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_190),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_216),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_217),
.A2(n_224),
.B1(n_191),
.B2(n_175),
.Y(n_254)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_197),
.Y(n_222)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_222),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_198),
.A2(n_180),
.B1(n_183),
.B2(n_186),
.Y(n_224)
);

AND2x4_ASAP7_75t_L g238 ( 
.A(n_225),
.B(n_209),
.Y(n_238)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_200),
.Y(n_226)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_226),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_209),
.A2(n_182),
.B(n_187),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_228),
.B(n_182),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_234),
.A2(n_202),
.B(n_209),
.Y(n_242)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_201),
.Y(n_235)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_235),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_238),
.B(n_248),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_236),
.B(n_199),
.C(n_189),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_239),
.B(n_241),
.C(n_245),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_236),
.B(n_199),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_242),
.B(n_249),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_243),
.B(n_251),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_218),
.B(n_211),
.Y(n_244)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_244),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_229),
.B(n_205),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_233),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_247),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_230),
.A2(n_203),
.B1(n_206),
.B2(n_189),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_229),
.B(n_196),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_234),
.B(n_210),
.C(n_212),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_250),
.B(n_228),
.C(n_219),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_231),
.B(n_174),
.Y(n_251)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_218),
.Y(n_253)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_253),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_254),
.A2(n_257),
.B1(n_227),
.B2(n_221),
.Y(n_260)
);

AND2x6_ASAP7_75t_L g255 ( 
.A(n_237),
.B(n_213),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_255),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_233),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_256),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_224),
.A2(n_215),
.B1(n_175),
.B2(n_188),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_254),
.A2(n_230),
.B1(n_222),
.B2(n_226),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_259),
.A2(n_260),
.B1(n_264),
.B2(n_223),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_244),
.A2(n_219),
.B1(n_235),
.B2(n_221),
.Y(n_264)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_240),
.Y(n_267)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_267),
.Y(n_282)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_240),
.Y(n_268)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_268),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_269),
.B(n_260),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_257),
.A2(n_231),
.B1(n_217),
.B2(n_184),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_270),
.A2(n_274),
.B1(n_223),
.B2(n_190),
.Y(n_291)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_246),
.Y(n_272)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_272),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_246),
.A2(n_252),
.B1(n_253),
.B2(n_239),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_252),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_275),
.Y(n_293)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_248),
.Y(n_277)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_277),
.Y(n_300)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_242),
.Y(n_278)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_278),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_271),
.B(n_245),
.Y(n_279)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_279),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_241),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_280),
.B(n_287),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_262),
.A2(n_238),
.B1(n_255),
.B2(n_250),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_281),
.A2(n_291),
.B1(n_294),
.B2(n_204),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_271),
.B(n_181),
.Y(n_283)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_283),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_265),
.B(n_225),
.C(n_238),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_284),
.B(n_292),
.C(n_258),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_285),
.B(n_266),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_SL g304 ( 
.A(n_286),
.B(n_278),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_276),
.B(n_238),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_263),
.B(n_184),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_288),
.B(n_289),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_269),
.B(n_194),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_259),
.A2(n_238),
.B1(n_247),
.B2(n_256),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_290),
.A2(n_273),
.B1(n_261),
.B2(n_268),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_277),
.B(n_214),
.C(n_207),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_262),
.A2(n_188),
.B1(n_233),
.B2(n_232),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_275),
.B(n_178),
.Y(n_295)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_295),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_258),
.A2(n_232),
.B(n_220),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_296),
.B(n_161),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_264),
.B(n_220),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_298),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_302),
.B(n_304),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_305),
.A2(n_310),
.B1(n_172),
.B2(n_170),
.Y(n_346)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_300),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_306),
.B(n_312),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_281),
.A2(n_273),
.B1(n_261),
.B2(n_267),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_307),
.A2(n_318),
.B1(n_321),
.B2(n_299),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_280),
.B(n_272),
.C(n_266),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_309),
.B(n_311),
.C(n_320),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_286),
.B(n_284),
.C(n_292),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_293),
.B(n_214),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_287),
.B(n_207),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_313),
.B(n_317),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_301),
.A2(n_167),
.B(n_164),
.Y(n_315)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_315),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_SL g317 ( 
.A(n_285),
.B(n_208),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_293),
.A2(n_208),
.B1(n_204),
.B2(n_162),
.Y(n_319)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_319),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_301),
.B(n_149),
.C(n_138),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_300),
.A2(n_89),
.B1(n_103),
.B2(n_99),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g337 ( 
.A(n_322),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_282),
.B(n_14),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g332 ( 
.A(n_324),
.B(n_15),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_311),
.B(n_309),
.C(n_302),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_327),
.B(n_333),
.C(n_335),
.Y(n_349)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_325),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_328),
.B(n_343),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_314),
.A2(n_290),
.B1(n_298),
.B2(n_297),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_329),
.A2(n_137),
.B1(n_85),
.B2(n_165),
.Y(n_348)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_332),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_323),
.B(n_296),
.C(n_299),
.Y(n_333)
);

INVxp67_ASAP7_75t_SL g358 ( 
.A(n_334),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_323),
.B(n_304),
.C(n_307),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_308),
.A2(n_297),
.B(n_282),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_338),
.B(n_345),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_313),
.B(n_155),
.C(n_163),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_340),
.B(n_112),
.C(n_93),
.Y(n_350)
);

OAI321xp33_ASAP7_75t_L g341 ( 
.A1(n_316),
.A2(n_10),
.A3(n_109),
.B1(n_134),
.B2(n_108),
.C(n_161),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_341),
.A2(n_100),
.B1(n_132),
.B2(n_69),
.Y(n_355)
);

NAND2xp33_ASAP7_75t_L g343 ( 
.A(n_303),
.B(n_173),
.Y(n_343)
);

NAND2xp33_ASAP7_75t_SL g344 ( 
.A(n_317),
.B(n_165),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_SL g359 ( 
.A(n_344),
.B(n_104),
.Y(n_359)
);

OAI21x1_ASAP7_75t_L g345 ( 
.A1(n_320),
.A2(n_173),
.B(n_142),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_346),
.B(n_93),
.Y(n_352)
);

BUFx12_ASAP7_75t_L g347 ( 
.A(n_321),
.Y(n_347)
);

HB1xp67_ASAP7_75t_L g357 ( 
.A(n_347),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_348),
.B(n_353),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_350),
.B(n_360),
.Y(n_371)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_352),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_337),
.A2(n_109),
.B1(n_108),
.B2(n_83),
.Y(n_353)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_355),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_330),
.B(n_10),
.Y(n_356)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_356),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_359),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_327),
.B(n_90),
.C(n_54),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_326),
.B(n_56),
.C(n_55),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_361),
.B(n_363),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_336),
.B(n_122),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_SL g364 ( 
.A(n_336),
.B(n_10),
.Y(n_364)
);

NAND3xp33_ASAP7_75t_L g367 ( 
.A(n_364),
.B(n_331),
.C(n_1),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_335),
.B(n_122),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_365),
.B(n_326),
.C(n_333),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_366),
.B(n_0),
.Y(n_391)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_367),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_357),
.B(n_349),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_SL g383 ( 
.A(n_368),
.B(n_378),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_349),
.B(n_339),
.C(n_342),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_375),
.B(n_38),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_357),
.A2(n_347),
.B1(n_346),
.B2(n_344),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_377),
.A2(n_350),
.B1(n_48),
.B2(n_84),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_362),
.B(n_339),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_SL g379 ( 
.A1(n_351),
.A2(n_358),
.B(n_347),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_379),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_SL g380 ( 
.A1(n_375),
.A2(n_358),
.B(n_340),
.Y(n_380)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_380),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_SL g381 ( 
.A1(n_373),
.A2(n_359),
.B(n_354),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_SL g393 ( 
.A1(n_381),
.A2(n_391),
.B(n_384),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_382),
.B(n_385),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_SL g385 ( 
.A1(n_366),
.A2(n_122),
.B(n_1),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_368),
.A2(n_371),
.B(n_370),
.Y(n_386)
);

OR2x2_ASAP7_75t_L g396 ( 
.A(n_386),
.B(n_387),
.Y(n_396)
);

INVx11_ASAP7_75t_L g387 ( 
.A(n_379),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_388),
.B(n_389),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_369),
.A2(n_33),
.B1(n_1),
.B2(n_2),
.Y(n_389)
);

NOR3xp33_ASAP7_75t_SL g392 ( 
.A(n_387),
.B(n_372),
.C(n_376),
.Y(n_392)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_392),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_393),
.B(n_3),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_384),
.A2(n_377),
.B1(n_378),
.B2(n_374),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_394),
.B(n_0),
.C(n_2),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_383),
.B(n_19),
.C(n_26),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_397),
.A2(n_398),
.B(n_399),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_390),
.B(n_19),
.C(n_26),
.Y(n_398)
);

NOR2xp67_ASAP7_75t_L g399 ( 
.A(n_381),
.B(n_0),
.Y(n_399)
);

MAJx2_ASAP7_75t_L g409 ( 
.A(n_403),
.B(n_405),
.C(n_400),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_395),
.B(n_19),
.C(n_26),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_406),
.B(n_26),
.C(n_19),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_SL g407 ( 
.A1(n_396),
.A2(n_3),
.B(n_4),
.Y(n_407)
);

AOI322xp5_ASAP7_75t_L g410 ( 
.A1(n_407),
.A2(n_399),
.A3(n_401),
.B1(n_7),
.B2(n_8),
.C1(n_5),
.C2(n_6),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g408 ( 
.A1(n_401),
.A2(n_3),
.B(n_4),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_SL g411 ( 
.A1(n_408),
.A2(n_5),
.B(n_6),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_409),
.B(n_410),
.C(n_413),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_L g415 ( 
.A1(n_411),
.A2(n_412),
.B(n_6),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_SL g412 ( 
.A(n_402),
.B(n_404),
.Y(n_412)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_415),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_L g416 ( 
.A1(n_412),
.A2(n_19),
.B(n_8),
.Y(n_416)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_416),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_418),
.B(n_414),
.C(n_26),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_419),
.B(n_7),
.Y(n_420)
);

AOI21xp5_ASAP7_75t_L g421 ( 
.A1(n_420),
.A2(n_417),
.B(n_8),
.Y(n_421)
);


endmodule