module real_jpeg_6819_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_14;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_1),
.A2(n_106),
.B1(n_193),
.B2(n_194),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_1),
.Y(n_193)
);

OAI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_1),
.A2(n_193),
.B1(n_231),
.B2(n_233),
.Y(n_230)
);

OAI22xp33_ASAP7_75t_SL g330 ( 
.A1(n_1),
.A2(n_157),
.B1(n_193),
.B2(n_331),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_L g352 ( 
.A1(n_1),
.A2(n_193),
.B1(n_353),
.B2(n_356),
.Y(n_352)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_2),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_3),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.Y(n_28)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_3),
.A2(n_32),
.B1(n_155),
.B2(n_157),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_3),
.A2(n_32),
.B1(n_185),
.B2(n_188),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_3),
.B(n_92),
.Y(n_260)
);

O2A1O1Ixp33_ASAP7_75t_L g318 ( 
.A1(n_3),
.A2(n_319),
.B(n_321),
.C(n_325),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_3),
.B(n_343),
.C(n_345),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_3),
.B(n_121),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_3),
.B(n_377),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_3),
.B(n_57),
.Y(n_382)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_4),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_5),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_5),
.Y(n_370)
);

INVx8_ASAP7_75t_L g378 ( 
.A(n_5),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_6),
.A2(n_68),
.B1(n_69),
.B2(n_71),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_6),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_6),
.A2(n_68),
.B1(n_147),
.B2(n_150),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_6),
.A2(n_68),
.B1(n_175),
.B2(n_177),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_6),
.A2(n_68),
.B1(n_203),
.B2(n_205),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_7),
.Y(n_85)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_7),
.Y(n_89)
);

BUFx5_ASAP7_75t_L g102 ( 
.A(n_7),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g243 ( 
.A(n_7),
.Y(n_243)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_8),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_9),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_9),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_9),
.Y(n_106)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_9),
.Y(n_194)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_9),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_9),
.Y(n_206)
);

BUFx5_ASAP7_75t_L g244 ( 
.A(n_9),
.Y(n_244)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_10),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_11),
.A2(n_37),
.B1(n_43),
.B2(n_44),
.Y(n_36)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_11),
.A2(n_43),
.B1(n_114),
.B2(n_117),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_11),
.A2(n_43),
.B1(n_252),
.B2(n_254),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_217),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_215),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_195),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_15),
.B(n_195),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_110),
.C(n_163),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_16),
.A2(n_110),
.B1(n_111),
.B2(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_16),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_74),
.B2(n_75),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_17),
.A2(n_76),
.B(n_78),
.Y(n_214)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_35),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_19),
.A2(n_76),
.B1(n_77),
.B2(n_78),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_19),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_19),
.A2(n_35),
.B1(n_76),
.B2(n_299),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_19),
.B(n_318),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_19),
.A2(n_76),
.B1(n_318),
.B2(n_394),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_25),
.B(n_28),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_20),
.B(n_174),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_20),
.B(n_28),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_20),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_20),
.B(n_352),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_23),
.Y(n_20)
);

BUFx8_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_22),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_23),
.B(n_174),
.Y(n_263)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_28),
.Y(n_171)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_31),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_32),
.A2(n_106),
.B(n_107),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_32),
.B(n_108),
.Y(n_107)
);

OAI21xp33_ASAP7_75t_L g321 ( 
.A1(n_32),
.A2(n_322),
.B(n_324),
.Y(n_321)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_35),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_46),
.B(n_66),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_36),
.A2(n_159),
.B(n_161),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_39),
.Y(n_324)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_42),
.Y(n_127)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_42),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_46),
.A2(n_153),
.B(n_159),
.Y(n_210)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_47),
.B(n_67),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_47),
.B(n_154),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_47),
.B(n_330),
.Y(n_329)
);

NOR2x1_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_57),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_51),
.B1(n_53),
.B2(n_55),
.Y(n_48)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_50),
.A2(n_123),
.B1(n_126),
.B2(n_128),
.Y(n_122)
);

AO22x1_ASAP7_75t_SL g57 ( 
.A1(n_51),
.A2(n_58),
.B1(n_60),
.B2(n_64),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_52),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_57),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_57),
.B(n_330),
.Y(n_347)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_61),
.Y(n_356)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_63),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_63),
.Y(n_178)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_65),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_65),
.Y(n_375)
);

AND2x2_ASAP7_75t_SL g269 ( 
.A(n_66),
.B(n_270),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_66),
.B(n_329),
.Y(n_358)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_70),
.Y(n_156)
);

INVx6_ASAP7_75t_L g341 ( 
.A(n_70),
.Y(n_341)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_103),
.B(n_104),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_80),
.B(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_80),
.B(n_105),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_80),
.B(n_202),
.Y(n_289)
);

NOR2x1_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_92),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_84),
.B1(n_86),
.B2(n_90),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_85),
.Y(n_249)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_89),
.Y(n_94)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_92),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_92),
.B(n_105),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_92),
.B(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_92),
.B(n_192),
.Y(n_225)
);

AO22x1_ASAP7_75t_SL g92 ( 
.A1(n_93),
.A2(n_95),
.B1(n_98),
.B2(n_101),
.Y(n_92)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_95),
.Y(n_247)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_97),
.Y(n_100)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_97),
.Y(n_116)
);

BUFx5_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_97),
.Y(n_144)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_97),
.Y(n_241)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_100),
.Y(n_232)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_106),
.Y(n_109)
);

INVxp33_ASAP7_75t_L g245 ( 
.A(n_107),
.Y(n_245)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_151),
.B(n_162),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_112),
.B(n_151),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_121),
.B(n_131),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_113),
.A2(n_183),
.B(n_212),
.Y(n_211)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_114),
.Y(n_325)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g138 ( 
.A(n_116),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_116),
.Y(n_187)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g150 ( 
.A(n_120),
.Y(n_150)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_120),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_121),
.B(n_146),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_121),
.B(n_230),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_121),
.A2(n_183),
.B(n_184),
.Y(n_287)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_122),
.B(n_133),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_122),
.B(n_278),
.Y(n_277)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_125),
.Y(n_130)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_125),
.Y(n_136)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_125),
.Y(n_140)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_125),
.Y(n_323)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_127),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_130),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_131),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_145),
.Y(n_131)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_132),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_137),
.B1(n_139),
.B2(n_141),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_144),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_144),
.Y(n_188)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_160),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_152),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_153),
.B(n_159),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVxp67_ASAP7_75t_SL g160 ( 
.A(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_161),
.B(n_347),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_162),
.A2(n_197),
.B1(n_198),
.B2(n_213),
.Y(n_196)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_162),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_163),
.B(n_302),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_180),
.C(n_189),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_164),
.A2(n_165),
.B1(n_296),
.B2(n_297),
.Y(n_295)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_179),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_166),
.B(n_179),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_172),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_167),
.B(n_350),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_171),
.Y(n_167)
);

INVx3_ASAP7_75t_SL g168 ( 
.A(n_169),
.Y(n_168)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_170),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_172),
.B(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_173),
.A2(n_251),
.B(n_255),
.Y(n_250)
);

BUFx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_176),
.Y(n_253)
);

INVx4_ASAP7_75t_L g254 ( 
.A(n_177),
.Y(n_254)
);

INVx8_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_180),
.B(n_189),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_181),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_181),
.B(n_258),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_182),
.B(n_229),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_183),
.B(n_230),
.Y(n_258)
);

INVxp67_ASAP7_75t_SL g278 ( 
.A(n_184),
.Y(n_278)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_191),
.B(n_201),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_214),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_200),
.B1(n_208),
.B2(n_209),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_207),
.Y(n_200)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_207),
.B(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_210),
.A2(n_227),
.B1(n_235),
.B2(n_236),
.Y(n_226)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_210),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_210),
.B(n_224),
.C(n_227),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_403),
.Y(n_218)
);

NAND3xp33_ASAP7_75t_SL g219 ( 
.A(n_220),
.B(n_292),
.C(n_308),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_279),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_264),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_222),
.B(n_264),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_237),
.C(n_256),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_223),
.B(n_311),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_224),
.B(n_226),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_225),
.B(n_289),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_227),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

INVx8_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_237),
.A2(n_238),
.B1(n_256),
.B2(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_250),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_239),
.B(n_250),
.Y(n_272)
);

AOI32xp33_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_242),
.A3(n_244),
.B1(n_245),
.B2(n_246),
.Y(n_239)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

NAND2xp33_ASAP7_75t_SL g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_251),
.A2(n_263),
.B(n_268),
.Y(n_267)
);

BUFx3_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_256),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_259),
.C(n_261),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_257),
.B(n_315),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_258),
.B(n_276),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_259),
.A2(n_260),
.B1(n_261),
.B2(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g316 ( 
.A(n_261),
.Y(n_316)
);

OR2x2_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_262),
.B(n_368),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_SL g381 ( 
.A(n_263),
.B(n_351),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_264),
.B(n_280),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_264),
.B(n_280),
.Y(n_407)
);

FAx1_ASAP7_75t_SL g264 ( 
.A(n_265),
.B(n_266),
.CI(n_271),
.CON(n_264),
.SN(n_264)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_269),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_267),
.B(n_269),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_270),
.B(n_347),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_SL g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_272),
.B(n_274),
.C(n_275),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g405 ( 
.A1(n_279),
.A2(n_406),
.B(n_407),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_281),
.B(n_283),
.C(n_284),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_285),
.B(n_288),
.C(n_290),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_288),
.B1(n_290),
.B2(n_291),
.Y(n_286)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_287),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_288),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_304),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_293),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_301),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_294),
.B(n_301),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_298),
.C(n_300),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_295),
.B(n_298),
.Y(n_306)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_300),
.B(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_304),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_307),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_305),
.B(n_307),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_309),
.A2(n_334),
.B(n_402),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_310),
.B(n_313),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_310),
.B(n_313),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_317),
.C(n_326),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_314),
.B(n_398),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_317),
.A2(n_326),
.B1(n_327),
.B2(n_399),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_317),
.Y(n_399)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_318),
.Y(n_394)
);

BUFx3_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx6_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_329),
.Y(n_327)
);

INVx5_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx3_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_335),
.A2(n_396),
.B(n_401),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_336),
.A2(n_386),
.B(n_395),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_337),
.A2(n_362),
.B(n_385),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_348),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_338),
.B(n_348),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_346),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_339),
.A2(n_340),
.B1(n_346),
.B2(n_365),
.Y(n_364)
);

CKINVDCx16_ASAP7_75t_R g339 ( 
.A(n_340),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_342),
.Y(n_340)
);

INVx4_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_346),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_357),
.Y(n_348)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_349),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_352),
.B(n_369),
.Y(n_368)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx6_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_358),
.A2(n_359),
.B1(n_360),
.B2(n_361),
.Y(n_357)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_358),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_359),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_359),
.B(n_360),
.C(n_388),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_SL g362 ( 
.A1(n_363),
.A2(n_371),
.B(n_384),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_SL g363 ( 
.A(n_364),
.B(n_366),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_364),
.B(n_366),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx3_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_372),
.A2(n_380),
.B(n_383),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_379),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_376),
.Y(n_373)
);

INVx4_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx4_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_381),
.B(n_382),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_381),
.B(n_382),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_389),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_387),
.B(n_389),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_393),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_392),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_391),
.B(n_392),
.C(n_393),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_397),
.B(n_400),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_397),
.B(n_400),
.Y(n_401)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g403 ( 
.A1(n_404),
.A2(n_405),
.B(n_408),
.C(n_409),
.D(n_410),
.Y(n_403)
);


endmodule