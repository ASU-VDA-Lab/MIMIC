module fake_netlist_5_1709_n_104 (n_8, n_10, n_4, n_5, n_7, n_0, n_12, n_9, n_14, n_2, n_16, n_13, n_3, n_11, n_15, n_6, n_1, n_104);

input n_8;
input n_10;
input n_4;
input n_5;
input n_7;
input n_0;
input n_12;
input n_9;
input n_14;
input n_2;
input n_16;
input n_13;
input n_3;
input n_11;
input n_15;
input n_6;
input n_1;

output n_104;

wire n_91;
wire n_82;
wire n_24;
wire n_86;
wire n_83;
wire n_61;
wire n_90;
wire n_75;
wire n_101;
wire n_78;
wire n_65;
wire n_74;
wire n_57;
wire n_96;
wire n_37;
wire n_31;
wire n_66;
wire n_98;
wire n_60;
wire n_43;
wire n_58;
wire n_69;
wire n_18;
wire n_42;
wire n_22;
wire n_45;
wire n_46;
wire n_21;
wire n_94;
wire n_38;
wire n_80;
wire n_35;
wire n_73;
wire n_17;
wire n_92;
wire n_19;
wire n_30;
wire n_33;
wire n_84;
wire n_23;
wire n_29;
wire n_79;
wire n_47;
wire n_25;
wire n_53;
wire n_44;
wire n_40;
wire n_34;
wire n_100;
wire n_62;
wire n_71;
wire n_85;
wire n_95;
wire n_59;
wire n_26;
wire n_55;
wire n_99;
wire n_49;
wire n_20;
wire n_39;
wire n_54;
wire n_67;
wire n_36;
wire n_76;
wire n_87;
wire n_27;
wire n_64;
wire n_77;
wire n_102;
wire n_81;
wire n_28;
wire n_89;
wire n_70;
wire n_68;
wire n_93;
wire n_72;
wire n_32;
wire n_41;
wire n_103;
wire n_56;
wire n_51;
wire n_63;
wire n_97;
wire n_48;
wire n_50;
wire n_52;
wire n_88;

INVxp67_ASAP7_75t_SL g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVxp67_ASAP7_75t_SL g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVxp67_ASAP7_75t_SL g28 ( 
.A(n_4),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_25),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_23),
.Y(n_35)
);

CKINVDCx5p33_ASAP7_75t_R g36 ( 
.A(n_24),
.Y(n_36)
);

CKINVDCx5p33_ASAP7_75t_R g37 ( 
.A(n_20),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_22),
.B(n_2),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_42),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

NAND3xp33_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_30),
.C(n_29),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_28),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_19),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

CKINVDCx5p33_ASAP7_75t_R g54 ( 
.A(n_47),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_52),
.B(n_37),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_54),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_58),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_61),
.A2(n_35),
.B1(n_45),
.B2(n_17),
.Y(n_64)
);

NAND2x1p5_ASAP7_75t_L g65 ( 
.A(n_62),
.B(n_57),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

CKINVDCx5p33_ASAP7_75t_R g67 ( 
.A(n_59),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_61),
.A2(n_45),
.B1(n_51),
.B2(n_56),
.Y(n_68)
);

INVxp67_ASAP7_75t_R g69 ( 
.A(n_64),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_L g70 ( 
.A1(n_67),
.A2(n_60),
.B1(n_31),
.B2(n_34),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_68),
.A2(n_63),
.B1(n_62),
.B2(n_21),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_69),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_71),
.B(n_48),
.Y(n_73)
);

CKINVDCx5p33_ASAP7_75t_R g74 ( 
.A(n_70),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_71),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_72),
.B(n_74),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_72),
.B(n_44),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_75),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_75),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_74),
.B(n_73),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_79),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_79),
.B(n_66),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_76),
.B(n_47),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_78),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_77),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_83),
.A2(n_80),
.B1(n_29),
.B2(n_26),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_85),
.B(n_40),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_81),
.Y(n_88)
);

NOR3xp33_ASAP7_75t_L g89 ( 
.A(n_87),
.B(n_82),
.C(n_84),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_88),
.Y(n_90)
);

NAND2xp33_ASAP7_75t_SL g91 ( 
.A(n_90),
.B(n_86),
.Y(n_91)
);

AOI21xp33_ASAP7_75t_L g92 ( 
.A1(n_89),
.A2(n_82),
.B(n_26),
.Y(n_92)
);

XNOR2x2_ASAP7_75t_L g93 ( 
.A(n_90),
.B(n_33),
.Y(n_93)
);

OAI211xp5_ASAP7_75t_L g94 ( 
.A1(n_91),
.A2(n_41),
.B(n_38),
.C(n_3),
.Y(n_94)
);

NAND2xp33_ASAP7_75t_R g95 ( 
.A(n_93),
.B(n_3),
.Y(n_95)
);

AO22x2_ASAP7_75t_L g96 ( 
.A1(n_94),
.A2(n_95),
.B1(n_92),
.B2(n_57),
.Y(n_96)
);

OAI221xp5_ASAP7_75t_L g97 ( 
.A1(n_95),
.A2(n_52),
.B1(n_65),
.B2(n_43),
.C(n_49),
.Y(n_97)
);

NOR3xp33_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_66),
.C(n_6),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_96),
.A2(n_63),
.B1(n_62),
.B2(n_49),
.Y(n_99)
);

NOR2x1p5_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_49),
.Y(n_100)
);

AND3x1_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_98),
.C(n_7),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_101),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_102),
.Y(n_103)
);

AOI221xp5_ASAP7_75t_L g104 ( 
.A1(n_103),
.A2(n_63),
.B1(n_9),
.B2(n_13),
.C(n_15),
.Y(n_104)
);


endmodule