module fake_jpeg_19750_n_314 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_314);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_314;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx8_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

OR2x2_ASAP7_75t_L g32 ( 
.A(n_5),
.B(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_19),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_37),
.B(n_40),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_20),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_20),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_44),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_16),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_16),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_14),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_41),
.A2(n_32),
.B1(n_24),
.B2(n_29),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_46),
.A2(n_52),
.B1(n_60),
.B2(n_63),
.Y(n_89)
);

NAND2xp33_ASAP7_75t_SL g47 ( 
.A(n_38),
.B(n_43),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_38),
.Y(n_69)
);

A2O1A1Ixp33_ASAP7_75t_L g48 ( 
.A1(n_44),
.A2(n_35),
.B(n_34),
.C(n_28),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_48),
.B(n_65),
.Y(n_93)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_44),
.A2(n_24),
.B1(n_29),
.B2(n_19),
.Y(n_52)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_54),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_37),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_55),
.B(n_67),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_40),
.A2(n_29),
.B1(n_22),
.B2(n_33),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_56),
.A2(n_57),
.B1(n_60),
.B2(n_50),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_40),
.A2(n_22),
.B1(n_26),
.B2(n_27),
.Y(n_57)
);

NAND2x2_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_30),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_42),
.A2(n_27),
.B1(n_26),
.B2(n_33),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_37),
.A2(n_35),
.B1(n_34),
.B2(n_17),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_30),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_23),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_38),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_61),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_68),
.B(n_71),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_69),
.A2(n_85),
.B(n_86),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_58),
.B(n_45),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_55),
.A2(n_43),
.B1(n_39),
.B2(n_31),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_73),
.A2(n_21),
.B1(n_31),
.B2(n_36),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_74),
.B(n_75),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_64),
.B(n_18),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_76),
.A2(n_88),
.B1(n_38),
.B2(n_30),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_65),
.A2(n_43),
.B1(n_39),
.B2(n_17),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_77),
.A2(n_79),
.B1(n_96),
.B2(n_7),
.Y(n_138)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_78),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_58),
.A2(n_39),
.B1(n_21),
.B2(n_23),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_49),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_80),
.B(n_81),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_58),
.B(n_18),
.Y(n_81)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_83),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_SL g84 ( 
.A(n_66),
.B(n_28),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_SL g127 ( 
.A(n_84),
.B(n_36),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_38),
.Y(n_85)
);

NOR4xp25_ASAP7_75t_SL g86 ( 
.A(n_60),
.B(n_14),
.C(n_1),
.D(n_3),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_63),
.B(n_18),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_87),
.B(n_90),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_60),
.A2(n_25),
.B1(n_28),
.B2(n_30),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_46),
.B(n_28),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_51),
.B(n_28),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_91),
.B(n_100),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_92),
.Y(n_125)
);

BUFx12_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

INVx13_ASAP7_75t_L g124 ( 
.A(n_94),
.Y(n_124)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_59),
.Y(n_95)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_95),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_47),
.A2(n_23),
.B1(n_21),
.B2(n_31),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_59),
.Y(n_97)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

INVx2_ASAP7_75t_SL g99 ( 
.A(n_54),
.Y(n_99)
);

INVx11_ASAP7_75t_L g126 ( 
.A(n_99),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_53),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_53),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_102),
.B(n_104),
.Y(n_137)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_59),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_103),
.B(n_25),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_48),
.B(n_13),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_62),
.Y(n_105)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_105),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

INVxp33_ASAP7_75t_L g115 ( 
.A(n_106),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_48),
.B(n_23),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_107),
.B(n_108),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_67),
.B(n_21),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_68),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_109),
.B(n_118),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_110),
.A2(n_131),
.B1(n_82),
.B2(n_103),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_111),
.A2(n_138),
.B1(n_77),
.B2(n_79),
.Y(n_152)
);

AND2x6_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_25),
.Y(n_114)
);

OAI32xp33_ASAP7_75t_L g153 ( 
.A1(n_114),
.A2(n_96),
.A3(n_86),
.B1(n_94),
.B2(n_70),
.Y(n_153)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_116),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_93),
.B(n_36),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_78),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_122),
.B(n_102),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_127),
.B(n_132),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_85),
.B(n_0),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_130),
.B(n_139),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_83),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_82),
.A2(n_4),
.B(n_6),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_69),
.A2(n_7),
.B(n_8),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_134),
.B(n_84),
.C(n_74),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_85),
.B(n_7),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_142),
.A2(n_151),
.B1(n_159),
.B2(n_167),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_117),
.Y(n_144)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_144),
.Y(n_178)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_129),
.Y(n_146)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_146),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_121),
.B(n_80),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_147),
.B(n_150),
.Y(n_191)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_117),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_148),
.B(n_158),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_118),
.B(n_109),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_149),
.B(n_156),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_121),
.B(n_136),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_114),
.A2(n_89),
.B1(n_94),
.B2(n_69),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_152),
.A2(n_120),
.B1(n_131),
.B2(n_116),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_153),
.B(n_157),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_129),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_154),
.B(n_155),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_112),
.B(n_72),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_98),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_114),
.A2(n_89),
.B1(n_72),
.B2(n_100),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_119),
.Y(n_160)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_160),
.Y(n_184)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_119),
.Y(n_161)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_161),
.Y(n_197)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_125),
.Y(n_162)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_162),
.Y(n_201)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_125),
.Y(n_163)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_163),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_112),
.B(n_92),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_164),
.B(n_169),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_113),
.B(n_106),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_165),
.B(n_166),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_113),
.B(n_101),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_137),
.A2(n_135),
.B1(n_123),
.B2(n_110),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_123),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_168),
.Y(n_195)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_122),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_137),
.B(n_95),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_170),
.B(n_126),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_143),
.A2(n_133),
.B(n_135),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_171),
.A2(n_199),
.B(n_186),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_140),
.B(n_133),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_175),
.B(n_181),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_152),
.A2(n_138),
.B1(n_127),
.B2(n_124),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_177),
.A2(n_187),
.B1(n_162),
.B2(n_126),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_141),
.B(n_127),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_179),
.B(n_163),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_140),
.B(n_149),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_156),
.B(n_120),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_183),
.B(n_190),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_143),
.A2(n_139),
.B(n_130),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_186),
.A2(n_8),
.B(n_9),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_159),
.A2(n_151),
.B1(n_153),
.B2(n_168),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_188),
.A2(n_193),
.B1(n_194),
.B2(n_196),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_189),
.B(n_148),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_164),
.B(n_169),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_160),
.A2(n_111),
.B1(n_124),
.B2(n_134),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_161),
.A2(n_124),
.B1(n_132),
.B2(n_105),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_154),
.A2(n_146),
.B1(n_141),
.B2(n_145),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_157),
.A2(n_116),
.B(n_115),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_145),
.B(n_128),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_200),
.B(n_144),
.Y(n_220)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_173),
.Y(n_202)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_202),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_192),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_203),
.B(n_206),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_204),
.B(n_205),
.Y(n_238)
);

MAJx2_ASAP7_75t_L g205 ( 
.A(n_171),
.B(n_101),
.C(n_98),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_207),
.B(n_225),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_185),
.A2(n_128),
.B1(n_126),
.B2(n_99),
.Y(n_209)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_209),
.Y(n_230)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_173),
.Y(n_210)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_210),
.Y(n_231)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_190),
.Y(n_212)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_212),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_213),
.A2(n_215),
.B(n_221),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_214),
.B(n_227),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_188),
.A2(n_99),
.B(n_144),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_201),
.Y(n_216)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_216),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_182),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_218),
.B(n_219),
.Y(n_248)
);

NOR4xp25_ASAP7_75t_L g219 ( 
.A(n_175),
.B(n_10),
.C(n_11),
.D(n_12),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_220),
.B(n_222),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_199),
.A2(n_10),
.B(n_12),
.Y(n_221)
);

OR2x2_ASAP7_75t_L g222 ( 
.A(n_183),
.B(n_97),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_185),
.A2(n_10),
.B(n_13),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_223),
.Y(n_237)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_201),
.Y(n_224)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_224),
.Y(n_243)
);

NAND3xp33_ASAP7_75t_L g225 ( 
.A(n_191),
.B(n_13),
.C(n_15),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_182),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_226),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_172),
.B(n_15),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_184),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_228),
.B(n_174),
.Y(n_247)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_215),
.Y(n_234)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_234),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_217),
.A2(n_177),
.B1(n_176),
.B2(n_181),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_236),
.A2(n_223),
.B1(n_193),
.B2(n_194),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_204),
.B(n_176),
.C(n_179),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_241),
.B(n_242),
.C(n_246),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_214),
.B(n_196),
.C(n_172),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_208),
.B(n_200),
.C(n_197),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_247),
.B(n_222),
.Y(n_251)
);

BUFx2_ASAP7_75t_L g250 ( 
.A(n_235),
.Y(n_250)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_250),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_251),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_237),
.A2(n_217),
.B1(n_212),
.B2(n_202),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_253),
.A2(n_254),
.B1(n_246),
.B2(n_243),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_237),
.A2(n_210),
.B1(n_180),
.B2(n_207),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_241),
.B(n_208),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_255),
.B(n_259),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_247),
.A2(n_240),
.B(n_239),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_256),
.A2(n_239),
.B(n_249),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_248),
.B(n_227),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_257),
.B(n_258),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_242),
.B(n_211),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_238),
.B(n_211),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_238),
.B(n_205),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_260),
.B(n_264),
.Y(n_276)
);

INVxp33_ASAP7_75t_L g261 ( 
.A(n_244),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_261),
.B(n_266),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_240),
.B(n_247),
.Y(n_262)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_262),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_236),
.B(n_221),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_245),
.B(n_213),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_265),
.B(n_245),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_234),
.A2(n_220),
.B1(n_228),
.B2(n_224),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_267),
.A2(n_244),
.B1(n_229),
.B2(n_232),
.Y(n_268)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_268),
.Y(n_289)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_250),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_270),
.B(n_272),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g285 ( 
.A(n_271),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_263),
.A2(n_230),
.B1(n_231),
.B2(n_233),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_267),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_278),
.B(n_279),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_281),
.B(n_252),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_274),
.B(n_264),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_282),
.B(n_283),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_277),
.B(n_252),
.C(n_255),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_286),
.B(n_287),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_277),
.B(n_259),
.C(n_260),
.Y(n_287)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_268),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_290),
.A2(n_278),
.B1(n_273),
.B2(n_272),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_269),
.B(n_195),
.Y(n_291)
);

BUFx24_ASAP7_75t_SL g296 ( 
.A(n_291),
.Y(n_296)
);

BUFx24_ASAP7_75t_SL g292 ( 
.A(n_275),
.Y(n_292)
);

OAI211xp5_ASAP7_75t_SL g300 ( 
.A1(n_292),
.A2(n_288),
.B(n_261),
.C(n_184),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_294),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_285),
.A2(n_280),
.B(n_216),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_295),
.A2(n_198),
.B(n_178),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_289),
.B(n_265),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_297),
.B(n_298),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_283),
.B(n_276),
.C(n_281),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_300),
.B(n_197),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_296),
.B(n_284),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_302),
.B(n_303),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_297),
.A2(n_287),
.B(n_276),
.Y(n_304)
);

MAJx2_ASAP7_75t_L g307 ( 
.A(n_304),
.B(n_305),
.C(n_293),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_307),
.B(n_308),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_306),
.B(n_299),
.C(n_178),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_309),
.A2(n_301),
.B1(n_304),
.B2(n_198),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_311),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_312),
.B(n_310),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_313),
.B(n_16),
.Y(n_314)
);


endmodule