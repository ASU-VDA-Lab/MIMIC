module fake_jpeg_31546_n_279 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_279);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_279;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_12),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_36),
.B(n_37),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_12),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_42),
.Y(n_83)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_47),
.Y(n_50)
);

AO22x1_ASAP7_75t_SL g48 ( 
.A1(n_41),
.A2(n_46),
.B1(n_45),
.B2(n_44),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_48),
.A2(n_70),
.B1(n_76),
.B2(n_15),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_36),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_52),
.B(n_59),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_42),
.A2(n_20),
.B1(n_34),
.B2(n_18),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_54),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_43),
.A2(n_20),
.B1(n_34),
.B2(n_18),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_43),
.A2(n_20),
.B1(n_34),
.B2(n_18),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_39),
.A2(n_34),
.B1(n_18),
.B2(n_22),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_37),
.B(n_16),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_31),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_61),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_16),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_66),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_28),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_63),
.B(n_31),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_16),
.Y(n_66)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_45),
.A2(n_32),
.B1(n_33),
.B2(n_46),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_42),
.A2(n_18),
.B1(n_35),
.B2(n_22),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_72),
.A2(n_77),
.B1(n_26),
.B2(n_1),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_36),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_73),
.B(n_80),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_39),
.A2(n_35),
.B1(n_22),
.B2(n_17),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_42),
.A2(n_18),
.B1(n_35),
.B2(n_32),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_79),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_36),
.B(n_33),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_36),
.B(n_33),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_32),
.Y(n_96)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_63),
.B(n_21),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_86),
.B(n_100),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_61),
.A2(n_21),
.B(n_19),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_89),
.A2(n_49),
.B(n_1),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_52),
.B(n_15),
.C(n_17),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_91),
.B(n_7),
.Y(n_147)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_51),
.Y(n_95)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_95),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_96),
.B(n_99),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_73),
.A2(n_31),
.B1(n_29),
.B2(n_28),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_98),
.A2(n_105),
.B1(n_75),
.B2(n_55),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_74),
.B(n_25),
.Y(n_99)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_76),
.Y(n_101)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_103),
.B(n_118),
.Y(n_139)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_50),
.Y(n_104)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_104),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_51),
.A2(n_29),
.B1(n_28),
.B2(n_15),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_74),
.B(n_29),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_115),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_L g107 ( 
.A1(n_48),
.A2(n_68),
.B1(n_65),
.B2(n_69),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_107),
.A2(n_108),
.B1(n_113),
.B2(n_117),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_61),
.A2(n_21),
.B1(n_19),
.B2(n_17),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_50),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_109),
.Y(n_129)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_55),
.Y(n_110)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_110),
.Y(n_135)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_67),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_111),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_48),
.A2(n_19),
.B1(n_25),
.B2(n_14),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_112),
.A2(n_75),
.B1(n_55),
.B2(n_67),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_79),
.A2(n_26),
.B1(n_27),
.B2(n_12),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_60),
.B(n_27),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_114),
.B(n_49),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_82),
.B(n_26),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_116),
.A2(n_83),
.B1(n_26),
.B2(n_2),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_53),
.A2(n_26),
.B1(n_11),
.B2(n_10),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_83),
.A2(n_65),
.B1(n_71),
.B2(n_78),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_53),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_120),
.B(n_7),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_53),
.B(n_26),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_7),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_122),
.A2(n_133),
.B(n_91),
.Y(n_158)
);

AOI22x1_ASAP7_75t_L g123 ( 
.A1(n_101),
.A2(n_83),
.B1(n_64),
.B2(n_75),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_123),
.A2(n_132),
.B1(n_138),
.B2(n_140),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_119),
.A2(n_64),
.B(n_26),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_125),
.Y(n_171)
);

OR2x2_ASAP7_75t_L g181 ( 
.A(n_127),
.B(n_111),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_130),
.B(n_145),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_100),
.B(n_67),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_134),
.B(n_144),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_136),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_97),
.A2(n_11),
.B1(n_10),
.B2(n_3),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_112),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_119),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_141),
.A2(n_142),
.B1(n_151),
.B2(n_140),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_103),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_108),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g163 ( 
.A(n_143),
.B(n_152),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_86),
.B(n_4),
.Y(n_144)
);

INVxp33_ASAP7_75t_L g145 ( 
.A(n_118),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_146),
.B(n_154),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_147),
.B(n_102),
.Y(n_183)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_148),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_84),
.B(n_8),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_150),
.B(n_9),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_86),
.A2(n_8),
.B1(n_9),
.B2(n_106),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_85),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_89),
.B(n_9),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_107),
.A2(n_9),
.B1(n_113),
.B2(n_84),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_155),
.A2(n_110),
.B1(n_95),
.B2(n_120),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_129),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_157),
.B(n_162),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_158),
.A2(n_144),
.B(n_125),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_137),
.B(n_115),
.C(n_121),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_160),
.B(n_166),
.C(n_170),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_152),
.B(n_93),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_161),
.B(n_150),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_129),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_164),
.A2(n_184),
.B1(n_132),
.B2(n_139),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_137),
.B(n_90),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_131),
.Y(n_167)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_167),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_137),
.B(n_90),
.C(n_104),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_128),
.B(n_92),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_172),
.B(n_179),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_124),
.B(n_94),
.C(n_109),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_174),
.B(n_176),
.C(n_147),
.Y(n_206)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_131),
.Y(n_175)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_175),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_124),
.B(n_94),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_178),
.B(n_127),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_128),
.B(n_92),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_139),
.A2(n_88),
.B1(n_102),
.B2(n_87),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_180),
.A2(n_181),
.B1(n_149),
.B2(n_135),
.Y(n_204)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_126),
.Y(n_182)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_182),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_183),
.B(n_134),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_153),
.A2(n_88),
.B1(n_87),
.B2(n_111),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_126),
.Y(n_185)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_185),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_148),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_186),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_187),
.B(n_206),
.Y(n_215)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_191),
.Y(n_212)
);

OAI32xp33_ASAP7_75t_L g192 ( 
.A1(n_171),
.A2(n_143),
.A3(n_151),
.B1(n_154),
.B2(n_139),
.Y(n_192)
);

AOI221xp5_ASAP7_75t_L g216 ( 
.A1(n_192),
.A2(n_156),
.B1(n_168),
.B2(n_177),
.C(n_184),
.Y(n_216)
);

AO21x1_ASAP7_75t_L g194 ( 
.A1(n_163),
.A2(n_133),
.B(n_123),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_194),
.A2(n_201),
.B(n_205),
.Y(n_217)
);

NAND2xp33_ASAP7_75t_L g196 ( 
.A(n_163),
.B(n_123),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_196),
.B(n_202),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_163),
.Y(n_198)
);

INVx3_ASAP7_75t_SL g199 ( 
.A(n_181),
.Y(n_199)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_199),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_173),
.A2(n_155),
.B1(n_153),
.B2(n_122),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_200),
.A2(n_204),
.B1(n_164),
.B2(n_165),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_158),
.A2(n_142),
.B(n_138),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_159),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_183),
.B(n_146),
.C(n_149),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_208),
.B(n_170),
.C(n_178),
.Y(n_227)
);

OAI322xp33_ASAP7_75t_L g211 ( 
.A1(n_198),
.A2(n_168),
.A3(n_177),
.B1(n_186),
.B2(n_160),
.C1(n_176),
.C2(n_166),
.Y(n_211)
);

OAI211xp5_ASAP7_75t_L g236 ( 
.A1(n_211),
.A2(n_218),
.B(n_223),
.C(n_194),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_216),
.B(n_207),
.Y(n_238)
);

AOI321xp33_ASAP7_75t_L g218 ( 
.A1(n_192),
.A2(n_187),
.A3(n_195),
.B1(n_189),
.B2(n_205),
.C(n_196),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_193),
.Y(n_219)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_219),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_199),
.B(n_180),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_220),
.Y(n_232)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_221),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_203),
.B(n_157),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_222),
.B(n_224),
.Y(n_233)
);

AOI221xp5_ASAP7_75t_L g223 ( 
.A1(n_201),
.A2(n_156),
.B1(n_185),
.B2(n_182),
.C(n_162),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_207),
.B(n_190),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_195),
.B(n_174),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_225),
.B(n_227),
.C(n_206),
.Y(n_231)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_193),
.Y(n_226)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_226),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_200),
.A2(n_165),
.B1(n_173),
.B2(n_175),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_228),
.A2(n_199),
.B1(n_204),
.B2(n_188),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_229),
.A2(n_230),
.B1(n_243),
.B2(n_221),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_212),
.A2(n_188),
.B1(n_191),
.B2(n_194),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_231),
.B(n_234),
.C(n_227),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_215),
.B(n_208),
.C(n_190),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_236),
.A2(n_218),
.B(n_211),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_238),
.B(n_228),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_214),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_217),
.A2(n_202),
.B(n_210),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_240),
.A2(n_220),
.B(n_213),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_220),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_212),
.A2(n_210),
.B1(n_209),
.B2(n_197),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_244),
.B(n_246),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_245),
.B(n_249),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_234),
.B(n_215),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_233),
.Y(n_247)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_247),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_238),
.B(n_169),
.Y(n_248)
);

AOI31xp67_ASAP7_75t_SL g256 ( 
.A1(n_248),
.A2(n_239),
.A3(n_148),
.B(n_232),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_231),
.B(n_225),
.C(n_217),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_250),
.A2(n_232),
.B1(n_237),
.B2(n_243),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_230),
.B(n_213),
.Y(n_253)
);

OR2x2_ASAP7_75t_L g261 ( 
.A(n_253),
.B(n_242),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_229),
.B(n_214),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_253),
.A2(n_240),
.B(n_241),
.Y(n_255)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_256),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_257),
.B(n_254),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_245),
.A2(n_237),
.B1(n_242),
.B2(n_235),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_258),
.B(n_226),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_263),
.B(n_264),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_257),
.B(n_246),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_260),
.B(n_244),
.C(n_250),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_258),
.B(n_251),
.C(n_249),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_267),
.B(n_268),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_265),
.B(n_262),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_271),
.B(n_261),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_266),
.A2(n_252),
.B(n_259),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_272),
.A2(n_255),
.B(n_263),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_273),
.B(n_274),
.Y(n_276)
);

BUFx24_ASAP7_75t_SL g275 ( 
.A(n_273),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_275),
.B(n_270),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_277),
.A2(n_269),
.B(n_276),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_278),
.B(n_269),
.Y(n_279)
);


endmodule