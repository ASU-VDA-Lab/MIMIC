module fake_ibex_1479_n_3878 (n_151, n_85, n_599, n_778, n_822, n_507, n_743, n_540, n_754, n_395, n_84, n_64, n_171, n_756, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_766, n_688, n_130, n_177, n_707, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_845, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_790, n_452, n_86, n_70, n_664, n_255, n_175, n_586, n_773, n_638, n_398, n_59, n_28, n_125, n_304, n_821, n_191, n_873, n_593, n_5, n_62, n_71, n_153, n_862, n_545, n_583, n_678, n_663, n_194, n_249, n_334, n_634, n_733, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_872, n_423, n_608, n_864, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_336, n_258, n_861, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_727, n_58, n_43, n_216, n_33, n_652, n_781, n_421, n_828, n_738, n_475, n_802, n_166, n_163, n_753, n_645, n_500, n_747, n_542, n_114, n_236, n_34, n_376, n_377, n_584, n_531, n_647, n_15, n_761, n_556, n_748, n_24, n_189, n_498, n_698, n_280, n_317, n_340, n_375, n_708, n_105, n_187, n_667, n_1, n_154, n_682, n_850, n_182, n_196, n_326, n_327, n_879, n_89, n_50, n_723, n_144, n_170, n_270, n_346, n_383, n_113, n_840, n_561, n_117, n_417, n_471, n_846, n_739, n_755, n_265, n_853, n_504, n_158, n_859, n_259, n_276, n_339, n_470, n_770, n_210, n_348, n_220, n_875, n_674, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_671, n_228, n_711, n_876, n_147, n_552, n_251, n_384, n_632, n_373, n_854, n_458, n_244, n_73, n_343, n_310, n_714, n_703, n_426, n_323, n_469, n_829, n_598, n_825, n_143, n_740, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_67, n_453, n_591, n_655, n_333, n_110, n_306, n_400, n_47, n_550, n_736, n_169, n_10, n_673, n_21, n_732, n_798, n_832, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_121, n_527, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_690, n_120, n_835, n_168, n_526, n_785, n_155, n_824, n_315, n_441, n_604, n_13, n_637, n_122, n_523, n_116, n_694, n_787, n_614, n_370, n_431, n_719, n_574, n_0, n_289, n_716, n_865, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_669, n_838, n_750, n_746, n_22, n_136, n_261, n_742, n_521, n_665, n_459, n_30, n_518, n_367, n_221, n_852, n_789, n_654, n_656, n_724, n_437, n_731, n_602, n_842, n_355, n_767, n_474, n_878, n_758, n_594, n_636, n_710, n_720, n_407, n_102, n_490, n_568, n_813, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_156, n_570, n_126, n_623, n_585, n_715, n_791, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_769, n_222, n_660, n_186, n_524, n_349, n_765, n_849, n_857, n_454, n_777, n_295, n_730, n_331, n_576, n_230, n_96, n_759, n_185, n_388, n_625, n_619, n_536, n_611, n_352, n_290, n_558, n_666, n_174, n_467, n_427, n_607, n_827, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_851, n_689, n_793, n_167, n_676, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_771, n_205, n_618, n_488, n_139, n_514, n_705, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_635, n_844, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_783, n_347, n_847, n_830, n_473, n_445, n_629, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_359, n_826, n_299, n_87, n_262, n_433, n_75, n_439, n_704, n_643, n_137, n_679, n_841, n_772, n_810, n_768, n_839, n_338, n_173, n_696, n_796, n_797, n_837, n_477, n_640, n_363, n_402, n_725, n_180, n_369, n_596, n_201, n_699, n_14, n_351, n_368, n_456, n_834, n_257, n_77, n_869, n_718, n_801, n_44, n_672, n_722, n_401, n_553, n_554, n_66, n_735, n_305, n_713, n_307, n_192, n_804, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_721, n_4, n_814, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_763, n_745, n_329, n_447, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_868, n_546, n_199, n_788, n_795, n_592, n_495, n_762, n_410, n_308, n_675, n_800, n_463, n_624, n_706, n_411, n_135, n_520, n_784, n_684, n_775, n_658, n_512, n_615, n_685, n_283, n_366, n_397, n_111, n_803, n_692, n_36, n_627, n_18, n_709, n_322, n_53, n_227, n_499, n_115, n_757, n_11, n_248, n_92, n_702, n_451, n_712, n_101, n_190, n_138, n_650, n_776, n_409, n_582, n_818, n_653, n_214, n_238, n_579, n_843, n_332, n_799, n_517, n_211, n_744, n_817, n_218, n_314, n_691, n_563, n_132, n_277, n_555, n_337, n_522, n_700, n_479, n_534, n_225, n_360, n_272, n_511, n_23, n_734, n_468, n_223, n_381, n_525, n_815, n_780, n_535, n_382, n_502, n_681, n_633, n_532, n_726, n_95, n_405, n_863, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_819, n_161, n_237, n_29, n_203, n_268, n_440, n_858, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_729, n_741, n_603, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_616, n_782, n_833, n_217, n_324, n_391, n_831, n_537, n_728, n_78, n_805, n_670, n_820, n_20, n_69, n_390, n_544, n_39, n_178, n_509, n_695, n_786, n_639, n_303, n_362, n_717, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_680, n_501, n_809, n_752, n_856, n_668, n_779, n_871, n_266, n_42, n_294, n_112, n_485, n_870, n_46, n_284, n_811, n_808, n_80, n_172, n_250, n_493, n_460, n_609, n_476, n_792, n_461, n_575, n_313, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_774, n_72, n_319, n_195, n_513, n_212, n_588, n_877, n_693, n_311, n_860, n_661, n_848, n_406, n_606, n_737, n_97, n_197, n_528, n_181, n_131, n_123, n_631, n_683, n_260, n_620, n_794, n_836, n_462, n_302, n_450, n_443, n_686, n_572, n_867, n_644, n_577, n_344, n_393, n_436, n_428, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_697, n_816, n_874, n_83, n_32, n_107, n_149, n_489, n_677, n_399, n_254, n_213, n_424, n_565, n_823, n_701, n_271, n_241, n_68, n_503, n_292, n_807, n_394, n_79, n_81, n_35, n_364, n_687, n_159, n_202, n_231, n_298, n_587, n_760, n_751, n_806, n_160, n_657, n_764, n_184, n_56, n_492, n_649, n_812, n_855, n_232, n_380, n_749, n_281, n_866, n_559, n_425, n_3878);

input n_151;
input n_85;
input n_599;
input n_778;
input n_822;
input n_507;
input n_743;
input n_540;
input n_754;
input n_395;
input n_84;
input n_64;
input n_171;
input n_756;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_766;
input n_688;
input n_130;
input n_177;
input n_707;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_845;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_790;
input n_452;
input n_86;
input n_70;
input n_664;
input n_255;
input n_175;
input n_586;
input n_773;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_821;
input n_191;
input n_873;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_862;
input n_545;
input n_583;
input n_678;
input n_663;
input n_194;
input n_249;
input n_334;
input n_634;
input n_733;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_872;
input n_423;
input n_608;
input n_864;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_336;
input n_258;
input n_861;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_727;
input n_58;
input n_43;
input n_216;
input n_33;
input n_652;
input n_781;
input n_421;
input n_828;
input n_738;
input n_475;
input n_802;
input n_166;
input n_163;
input n_753;
input n_645;
input n_500;
input n_747;
input n_542;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_761;
input n_556;
input n_748;
input n_24;
input n_189;
input n_498;
input n_698;
input n_280;
input n_317;
input n_340;
input n_375;
input n_708;
input n_105;
input n_187;
input n_667;
input n_1;
input n_154;
input n_682;
input n_850;
input n_182;
input n_196;
input n_326;
input n_327;
input n_879;
input n_89;
input n_50;
input n_723;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_840;
input n_561;
input n_117;
input n_417;
input n_471;
input n_846;
input n_739;
input n_755;
input n_265;
input n_853;
input n_504;
input n_158;
input n_859;
input n_259;
input n_276;
input n_339;
input n_470;
input n_770;
input n_210;
input n_348;
input n_220;
input n_875;
input n_674;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_671;
input n_228;
input n_711;
input n_876;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_373;
input n_854;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_714;
input n_703;
input n_426;
input n_323;
input n_469;
input n_829;
input n_598;
input n_825;
input n_143;
input n_740;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_67;
input n_453;
input n_591;
input n_655;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_736;
input n_169;
input n_10;
input n_673;
input n_21;
input n_732;
input n_798;
input n_832;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_690;
input n_120;
input n_835;
input n_168;
input n_526;
input n_785;
input n_155;
input n_824;
input n_315;
input n_441;
input n_604;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_694;
input n_787;
input n_614;
input n_370;
input n_431;
input n_719;
input n_574;
input n_0;
input n_289;
input n_716;
input n_865;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_669;
input n_838;
input n_750;
input n_746;
input n_22;
input n_136;
input n_261;
input n_742;
input n_521;
input n_665;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_852;
input n_789;
input n_654;
input n_656;
input n_724;
input n_437;
input n_731;
input n_602;
input n_842;
input n_355;
input n_767;
input n_474;
input n_878;
input n_758;
input n_594;
input n_636;
input n_710;
input n_720;
input n_407;
input n_102;
input n_490;
input n_568;
input n_813;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_715;
input n_791;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_769;
input n_222;
input n_660;
input n_186;
input n_524;
input n_349;
input n_765;
input n_849;
input n_857;
input n_454;
input n_777;
input n_295;
input n_730;
input n_331;
input n_576;
input n_230;
input n_96;
input n_759;
input n_185;
input n_388;
input n_625;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_666;
input n_174;
input n_467;
input n_427;
input n_607;
input n_827;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_851;
input n_689;
input n_793;
input n_167;
input n_676;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_771;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_705;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_635;
input n_844;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_783;
input n_347;
input n_847;
input n_830;
input n_473;
input n_445;
input n_629;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_359;
input n_826;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_704;
input n_643;
input n_137;
input n_679;
input n_841;
input n_772;
input n_810;
input n_768;
input n_839;
input n_338;
input n_173;
input n_696;
input n_796;
input n_797;
input n_837;
input n_477;
input n_640;
input n_363;
input n_402;
input n_725;
input n_180;
input n_369;
input n_596;
input n_201;
input n_699;
input n_14;
input n_351;
input n_368;
input n_456;
input n_834;
input n_257;
input n_77;
input n_869;
input n_718;
input n_801;
input n_44;
input n_672;
input n_722;
input n_401;
input n_553;
input n_554;
input n_66;
input n_735;
input n_305;
input n_713;
input n_307;
input n_192;
input n_804;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_721;
input n_4;
input n_814;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_763;
input n_745;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_868;
input n_546;
input n_199;
input n_788;
input n_795;
input n_592;
input n_495;
input n_762;
input n_410;
input n_308;
input n_675;
input n_800;
input n_463;
input n_624;
input n_706;
input n_411;
input n_135;
input n_520;
input n_784;
input n_684;
input n_775;
input n_658;
input n_512;
input n_615;
input n_685;
input n_283;
input n_366;
input n_397;
input n_111;
input n_803;
input n_692;
input n_36;
input n_627;
input n_18;
input n_709;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_757;
input n_11;
input n_248;
input n_92;
input n_702;
input n_451;
input n_712;
input n_101;
input n_190;
input n_138;
input n_650;
input n_776;
input n_409;
input n_582;
input n_818;
input n_653;
input n_214;
input n_238;
input n_579;
input n_843;
input n_332;
input n_799;
input n_517;
input n_211;
input n_744;
input n_817;
input n_218;
input n_314;
input n_691;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_700;
input n_479;
input n_534;
input n_225;
input n_360;
input n_272;
input n_511;
input n_23;
input n_734;
input n_468;
input n_223;
input n_381;
input n_525;
input n_815;
input n_780;
input n_535;
input n_382;
input n_502;
input n_681;
input n_633;
input n_532;
input n_726;
input n_95;
input n_405;
input n_863;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_819;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_858;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_729;
input n_741;
input n_603;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_782;
input n_833;
input n_217;
input n_324;
input n_391;
input n_831;
input n_537;
input n_728;
input n_78;
input n_805;
input n_670;
input n_820;
input n_20;
input n_69;
input n_390;
input n_544;
input n_39;
input n_178;
input n_509;
input n_695;
input n_786;
input n_639;
input n_303;
input n_362;
input n_717;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_680;
input n_501;
input n_809;
input n_752;
input n_856;
input n_668;
input n_779;
input n_871;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_870;
input n_46;
input n_284;
input n_811;
input n_808;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_609;
input n_476;
input n_792;
input n_461;
input n_575;
input n_313;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_774;
input n_72;
input n_319;
input n_195;
input n_513;
input n_212;
input n_588;
input n_877;
input n_693;
input n_311;
input n_860;
input n_661;
input n_848;
input n_406;
input n_606;
input n_737;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_631;
input n_683;
input n_260;
input n_620;
input n_794;
input n_836;
input n_462;
input n_302;
input n_450;
input n_443;
input n_686;
input n_572;
input n_867;
input n_644;
input n_577;
input n_344;
input n_393;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_697;
input n_816;
input n_874;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_677;
input n_399;
input n_254;
input n_213;
input n_424;
input n_565;
input n_823;
input n_701;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_807;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_687;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_760;
input n_751;
input n_806;
input n_160;
input n_657;
input n_764;
input n_184;
input n_56;
input n_492;
input n_649;
input n_812;
input n_855;
input n_232;
input n_380;
input n_749;
input n_281;
input n_866;
input n_559;
input n_425;

output n_3878;

wire n_1084;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_1983;
wire n_2804;
wire n_3150;
wire n_992;
wire n_1582;
wire n_2201;
wire n_3853;
wire n_2512;
wire n_3590;
wire n_2960;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_3548;
wire n_2607;
wire n_1382;
wire n_3610;
wire n_3144;
wire n_2569;
wire n_2949;
wire n_1998;
wire n_2840;
wire n_1596;
wire n_926;
wire n_3319;
wire n_1079;
wire n_3077;
wire n_2835;
wire n_1100;
wire n_3559;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_1234;
wire n_3019;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_2498;
wire n_3817;
wire n_3755;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_3812;
wire n_2017;
wire n_1227;
wire n_962;
wire n_1080;
wire n_909;
wire n_2290;
wire n_3750;
wire n_3838;
wire n_957;
wire n_3255;
wire n_3272;
wire n_3674;
wire n_1652;
wire n_969;
wire n_1859;
wire n_1954;
wire n_2183;
wire n_2074;
wire n_2897;
wire n_1883;
wire n_1125;
wire n_2687;
wire n_3456;
wire n_2037;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_3132;
wire n_1765;
wire n_2392;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2640;
wire n_2682;
wire n_3605;
wire n_930;
wire n_1044;
wire n_3280;
wire n_3105;
wire n_3146;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_3569;
wire n_1614;
wire n_2374;
wire n_3334;
wire n_3819;
wire n_2598;
wire n_1722;
wire n_911;
wire n_2023;
wire n_2720;
wire n_3870;
wire n_3340;
wire n_2322;
wire n_1233;
wire n_2335;
wire n_3025;
wire n_3411;
wire n_2955;
wire n_3458;
wire n_3653;
wire n_3519;
wire n_2276;
wire n_1045;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_2230;
wire n_963;
wire n_1782;
wire n_2889;
wire n_3843;
wire n_2139;
wire n_2847;
wire n_3693;
wire n_3033;
wire n_1308;
wire n_1138;
wire n_2943;
wire n_1096;
wire n_2151;
wire n_2391;
wire n_1391;
wire n_3338;
wire n_3168;
wire n_884;
wire n_2396;
wire n_3440;
wire n_3135;
wire n_3175;
wire n_3729;
wire n_3484;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_3570;
wire n_2179;
wire n_1957;
wire n_2188;
wire n_1144;
wire n_2359;
wire n_2360;
wire n_2506;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_3187;
wire n_3830;
wire n_3598;
wire n_2724;
wire n_3086;
wire n_2475;
wire n_3721;
wire n_948;
wire n_2799;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_3726;
wire n_1730;
wire n_1307;
wire n_1327;
wire n_2644;
wire n_3211;
wire n_3479;
wire n_1840;
wire n_2837;
wire n_3751;
wire n_989;
wire n_3262;
wire n_3407;
wire n_3804;
wire n_1908;
wire n_3315;
wire n_3537;
wire n_1668;
wire n_2343;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_2565;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_3251;
wire n_1681;
wire n_2921;
wire n_3724;
wire n_1636;
wire n_939;
wire n_1687;
wire n_3192;
wire n_3533;
wire n_3753;
wire n_2192;
wire n_1766;
wire n_3184;
wire n_3566;
wire n_3469;
wire n_3170;
wire n_1922;
wire n_2032;
wire n_2820;
wire n_3323;
wire n_2311;
wire n_1937;
wire n_3392;
wire n_3347;
wire n_893;
wire n_3395;
wire n_3242;
wire n_3839;
wire n_1654;
wire n_3577;
wire n_2995;
wire n_3330;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_2707;
wire n_3509;
wire n_3472;
wire n_1749;
wire n_1680;
wire n_1981;
wire n_1195;
wire n_2918;
wire n_3353;
wire n_1945;
wire n_2638;
wire n_2860;
wire n_2448;
wire n_3631;
wire n_2015;
wire n_3807;
wire n_2537;
wire n_1130;
wire n_2643;
wire n_1228;
wire n_2998;
wire n_2336;
wire n_3845;
wire n_3641;
wire n_2163;
wire n_1081;
wire n_2354;
wire n_3639;
wire n_3856;
wire n_1155;
wire n_1292;
wire n_2432;
wire n_2873;
wire n_3043;
wire n_1576;
wire n_1664;
wire n_2273;
wire n_3298;
wire n_1427;
wire n_1133;
wire n_3049;
wire n_2421;
wire n_1926;
wire n_3208;
wire n_904;
wire n_2363;
wire n_2814;
wire n_3237;
wire n_3264;
wire n_3204;
wire n_2003;
wire n_1970;
wire n_3671;
wire n_3727;
wire n_2621;
wire n_3620;
wire n_1778;
wire n_2558;
wire n_2953;
wire n_2922;
wire n_2347;
wire n_3507;
wire n_3103;
wire n_2839;
wire n_1030;
wire n_1698;
wire n_3688;
wire n_1094;
wire n_2462;
wire n_3770;
wire n_1496;
wire n_1910;
wire n_2436;
wire n_1663;
wire n_2705;
wire n_1214;
wire n_1274;
wire n_2333;
wire n_2527;
wire n_1606;
wire n_1595;
wire n_2164;
wire n_3711;
wire n_1509;
wire n_1648;
wire n_1618;
wire n_2944;
wire n_1886;
wire n_2269;
wire n_3748;
wire n_1070;
wire n_1841;
wire n_2472;
wire n_2685;
wire n_2846;
wire n_3197;
wire n_3699;
wire n_1955;
wire n_3668;
wire n_917;
wire n_2249;
wire n_2413;
wire n_2362;
wire n_968;
wire n_3148;
wire n_3022;
wire n_2822;
wire n_3766;
wire n_1253;
wire n_3707;
wire n_1306;
wire n_1484;
wire n_2686;
wire n_1493;
wire n_2597;
wire n_1313;
wire n_2774;
wire n_3151;
wire n_2090;
wire n_2260;
wire n_3722;
wire n_3125;
wire n_2812;
wire n_3802;
wire n_3681;
wire n_2753;
wire n_3603;
wire n_1638;
wire n_2215;
wire n_1071;
wire n_1449;
wire n_1723;
wire n_1960;
wire n_2663;
wire n_3129;
wire n_937;
wire n_2595;
wire n_2116;
wire n_3714;
wire n_3592;
wire n_1645;
wire n_3186;
wire n_973;
wire n_1038;
wire n_2280;
wire n_1943;
wire n_3541;
wire n_1863;
wire n_2844;
wire n_1269;
wire n_2393;
wire n_2773;
wire n_3565;
wire n_2906;
wire n_3030;
wire n_3097;
wire n_3809;
wire n_979;
wire n_1309;
wire n_1999;
wire n_3810;
wire n_3718;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_3679;
wire n_3579;
wire n_2777;
wire n_2480;
wire n_3769;
wire n_1445;
wire n_2283;
wire n_2806;
wire n_2813;
wire n_2147;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_3210;
wire n_3221;
wire n_3667;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_1276;
wire n_3822;
wire n_1637;
wire n_3310;
wire n_2900;
wire n_3858;
wire n_1401;
wire n_3764;
wire n_3795;
wire n_1817;
wire n_2951;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_3765;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_2876;
wire n_2242;
wire n_1620;
wire n_1561;
wire n_3301;
wire n_2370;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_3451;
wire n_1219;
wire n_1865;
wire n_3177;
wire n_3518;
wire n_3399;
wire n_1252;
wire n_2022;
wire n_2730;
wire n_1170;
wire n_1927;
wire n_2373;
wire n_1869;
wire n_3842;
wire n_1853;
wire n_2275;
wire n_2980;
wire n_2189;
wire n_2482;
wire n_3799;
wire n_2767;
wire n_3676;
wire n_2899;
wire n_2826;
wire n_2112;
wire n_1753;
wire n_3351;
wire n_1322;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_1248;
wire n_2762;
wire n_2171;
wire n_3307;
wire n_1388;
wire n_2859;
wire n_2564;
wire n_3780;
wire n_3023;
wire n_1653;
wire n_1375;
wire n_3224;
wire n_1356;
wire n_894;
wire n_1118;
wire n_2591;
wire n_1881;
wire n_3762;
wire n_1969;
wire n_3798;
wire n_1296;
wire n_3060;
wire n_1326;
wire n_971;
wire n_1350;
wire n_3627;
wire n_906;
wire n_2957;
wire n_2586;
wire n_1093;
wire n_1764;
wire n_2412;
wire n_2783;
wire n_978;
wire n_3777;
wire n_899;
wire n_1799;
wire n_3293;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_2541;
wire n_2987;
wire n_881;
wire n_3259;
wire n_1702;
wire n_3381;
wire n_3630;
wire n_1558;
wire n_2750;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_2722;
wire n_2509;
wire n_2727;
wire n_3618;
wire n_1794;
wire n_1423;
wire n_3836;
wire n_1239;
wire n_2399;
wire n_1370;
wire n_2719;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_3038;
wire n_3732;
wire n_3779;
wire n_3521;
wire n_3203;
wire n_3295;
wire n_2723;
wire n_1616;
wire n_3199;
wire n_3808;
wire n_3093;
wire n_1569;
wire n_2664;
wire n_1434;
wire n_3716;
wire n_1649;
wire n_2389;
wire n_3450;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_3567;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_3435;
wire n_3530;
wire n_1613;
wire n_1988;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_2401;
wire n_1787;
wire n_2782;
wire n_2511;
wire n_3217;
wire n_1281;
wire n_3094;
wire n_3874;
wire n_1447;
wire n_2166;
wire n_2451;
wire n_2150;
wire n_1549;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_2919;
wire n_1332;
wire n_2660;
wire n_2661;
wire n_2292;
wire n_3573;
wire n_3563;
wire n_3510;
wire n_3560;
wire n_2334;
wire n_1424;
wire n_3467;
wire n_2625;
wire n_2350;
wire n_1742;
wire n_2444;
wire n_3652;
wire n_1818;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_3847;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_2649;
wire n_1040;
wire n_2203;
wire n_2693;
wire n_3194;
wire n_3607;
wire n_3371;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_1154;
wire n_3202;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_3572;
wire n_2646;
wire n_2387;
wire n_3375;
wire n_2397;
wire n_1121;
wire n_2746;
wire n_3241;
wire n_2256;
wire n_3317;
wire n_3800;
wire n_3461;
wire n_2445;
wire n_2729;
wire n_1571;
wire n_1980;
wire n_3355;
wire n_2529;
wire n_3583;
wire n_2019;
wire n_1407;
wire n_3282;
wire n_1235;
wire n_1821;
wire n_3832;
wire n_3508;
wire n_1003;
wire n_889;
wire n_3827;
wire n_2708;
wire n_3156;
wire n_3457;
wire n_2748;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_2697;
wire n_3531;
wire n_3415;
wire n_2470;
wire n_2355;
wire n_2890;
wire n_3698;
wire n_2731;
wire n_1543;
wire n_3466;
wire n_3386;
wire n_2233;
wire n_2499;
wire n_3370;
wire n_1504;
wire n_3814;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_2069;
wire n_2602;
wire n_1441;
wire n_2028;
wire n_3309;
wire n_3678;
wire n_1924;
wire n_2856;
wire n_1921;
wire n_3024;
wire n_1156;
wire n_2857;
wire n_1293;
wire n_1360;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_2070;
wire n_1042;
wire n_1888;
wire n_3471;
wire n_3117;
wire n_3320;
wire n_1786;
wire n_2033;
wire n_3039;
wire n_1319;
wire n_1553;
wire n_3478;
wire n_3701;
wire n_3542;
wire n_1041;
wire n_2766;
wire n_3756;
wire n_2828;
wire n_3754;
wire n_1964;
wire n_1090;
wire n_3720;
wire n_3374;
wire n_1196;
wire n_3704;
wire n_1182;
wire n_1271;
wire n_3811;
wire n_2416;
wire n_3633;
wire n_2786;
wire n_1731;
wire n_1905;
wire n_2962;
wire n_1031;
wire n_3416;
wire n_2879;
wire n_2958;
wire n_3147;
wire n_3694;
wire n_2052;
wire n_3690;
wire n_981;
wire n_3628;
wire n_2425;
wire n_2800;
wire n_3514;
wire n_3091;
wire n_3006;
wire n_3348;
wire n_2118;
wire n_2259;
wire n_3859;
wire n_2162;
wire n_2236;
wire n_3455;
wire n_3660;
wire n_2718;
wire n_2377;
wire n_2577;
wire n_1591;
wire n_3426;
wire n_3165;
wire n_2289;
wire n_2288;
wire n_2841;
wire n_3075;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_3448;
wire n_3634;
wire n_2744;
wire n_2101;
wire n_2795;
wire n_3524;
wire n_3788;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_3520;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_2924;
wire n_3054;
wire n_2456;
wire n_2264;
wire n_2076;
wire n_1036;
wire n_974;
wire n_2599;
wire n_1831;
wire n_3626;
wire n_3733;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_3171;
wire n_1733;
wire n_3365;
wire n_3684;
wire n_1634;
wire n_2853;
wire n_1932;
wire n_3775;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_1508;
wire n_2217;
wire n_3741;
wire n_3854;
wire n_1217;
wire n_3594;
wire n_2866;
wire n_3153;
wire n_3291;
wire n_2655;
wire n_3487;
wire n_2454;
wire n_1715;
wire n_1189;
wire n_3300;
wire n_1713;
wire n_3621;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_2829;
wire n_2968;
wire n_2740;
wire n_3473;
wire n_1700;
wire n_2623;
wire n_2622;
wire n_3232;
wire n_2819;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_3263;
wire n_3815;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_2858;
wire n_3708;
wire n_1056;
wire n_2626;
wire n_1283;
wire n_3007;
wire n_3790;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_1421;
wire n_1203;
wire n_3640;
wire n_3218;
wire n_2821;
wire n_2424;
wire n_1793;
wire n_1237;
wire n_2573;
wire n_2390;
wire n_2880;
wire n_2423;
wire n_3849;
wire n_1109;
wire n_965;
wire n_2741;
wire n_2793;
wire n_3098;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_3299;
wire n_2580;
wire n_3222;
wire n_1711;
wire n_3529;
wire n_3069;
wire n_3107;
wire n_3352;
wire n_3436;
wire n_1051;
wire n_1008;
wire n_3065;
wire n_2964;
wire n_2375;
wire n_1498;
wire n_2312;
wire n_2572;
wire n_2946;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1735;
wire n_1076;
wire n_2063;
wire n_1032;
wire n_936;
wire n_3082;
wire n_1884;
wire n_2176;
wire n_3813;
wire n_1825;
wire n_2805;
wire n_1589;
wire n_2717;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_3757;
wire n_2877;
wire n_1933;
wire n_2522;
wire n_3357;
wire n_3855;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2852;
wire n_2132;
wire n_3110;
wire n_1677;
wire n_1246;
wire n_3364;
wire n_1236;
wire n_2297;
wire n_3429;
wire n_3306;
wire n_3412;
wire n_3037;
wire n_3188;
wire n_2780;
wire n_3787;
wire n_1792;
wire n_1712;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_1877;
wire n_3445;
wire n_1477;
wire n_1184;
wire n_2080;
wire n_2220;
wire n_2585;
wire n_1724;
wire n_2554;
wire n_3155;
wire n_2838;
wire n_1364;
wire n_3183;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_3243;
wire n_2468;
wire n_929;
wire n_3248;
wire n_3214;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_3128;
wire n_1918;
wire n_2606;
wire n_3642;
wire n_2549;
wire n_2461;
wire n_3468;
wire n_2006;
wire n_2440;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_907;
wire n_1179;
wire n_1990;
wire n_3680;
wire n_1153;
wire n_3624;
wire n_1751;
wire n_2787;
wire n_3785;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_3525;
wire n_1737;
wire n_3145;
wire n_2779;
wire n_1117;
wire n_1273;
wire n_3821;
wire n_2547;
wire n_2930;
wire n_2616;
wire n_1748;
wire n_2662;
wire n_1083;
wire n_3205;
wire n_3872;
wire n_1014;
wire n_3801;
wire n_2883;
wire n_938;
wire n_1178;
wire n_2935;
wire n_2441;
wire n_3503;
wire n_2358;
wire n_2490;
wire n_3127;
wire n_3496;
wire n_2361;
wire n_1464;
wire n_1566;
wire n_3568;
wire n_944;
wire n_3312;
wire n_3003;
wire n_1848;
wire n_2062;
wire n_2277;
wire n_3841;
wire n_2650;
wire n_1982;
wire n_2252;
wire n_2888;
wire n_2339;
wire n_3614;
wire n_1334;
wire n_1963;
wire n_3394;
wire n_1695;
wire n_1418;
wire n_3331;
wire n_2402;
wire n_1137;
wire n_2552;
wire n_2910;
wire n_2999;
wire n_2590;
wire n_3119;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_3345;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_2792;
wire n_1602;
wire n_2965;
wire n_1776;
wire n_2372;
wire n_3341;
wire n_2382;
wire n_1852;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_3544;
wire n_3868;
wire n_1279;
wire n_2505;
wire n_931;
wire n_3488;
wire n_3554;
wire n_2481;
wire n_3692;
wire n_1064;
wire n_1408;
wire n_2832;
wire n_1028;
wire n_1264;
wire n_3535;
wire n_3730;
wire n_2808;
wire n_2287;
wire n_3597;
wire n_3396;
wire n_2954;
wire n_3526;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_3367;
wire n_3492;
wire n_1146;
wire n_3558;
wire n_2751;
wire n_2785;
wire n_2142;
wire n_1548;
wire n_3703;
wire n_2977;
wire n_1682;
wire n_1608;
wire n_3776;
wire n_3599;
wire n_1009;
wire n_1260;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2699;
wire n_2234;
wire n_2991;
wire n_1436;
wire n_3239;
wire n_2600;
wire n_1485;
wire n_1069;
wire n_2239;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_3826;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_2715;
wire n_3781;
wire n_1345;
wire n_2434;
wire n_1590;
wire n_2332;
wire n_2971;
wire n_954;
wire n_3578;
wire n_1628;
wire n_1773;
wire n_2133;
wire n_3553;
wire n_3072;
wire n_1545;
wire n_3249;
wire n_3580;
wire n_2369;
wire n_3470;
wire n_3584;
wire n_1471;
wire n_1738;
wire n_3441;
wire n_3797;
wire n_998;
wire n_1395;
wire n_1729;
wire n_1115;
wire n_2551;
wire n_3281;
wire n_2823;
wire n_3274;
wire n_2094;
wire n_2613;
wire n_1479;
wire n_3505;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_3397;
wire n_2934;
wire n_2807;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_2525;
wire n_3829;
wire n_1864;
wire n_943;
wire n_2568;
wire n_3087;
wire n_2629;
wire n_3587;
wire n_1086;
wire n_1523;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2733;
wire n_2241;
wire n_1470;
wire n_2109;
wire n_2098;
wire n_1761;
wire n_3796;
wire n_2648;
wire n_2458;
wire n_1836;
wire n_2398;
wire n_3032;
wire n_3401;
wire n_1593;
wire n_986;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_2833;
wire n_1699;
wire n_3179;
wire n_927;
wire n_1563;
wire n_2905;
wire n_3460;
wire n_2570;
wire n_3123;
wire n_1875;
wire n_3379;
wire n_1615;
wire n_2184;
wire n_2418;
wire n_1087;
wire n_3390;
wire n_3719;
wire n_1599;
wire n_1400;
wire n_1539;
wire n_1806;
wire n_2711;
wire n_3070;
wire n_3477;
wire n_3646;
wire n_2635;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_3074;
wire n_3020;
wire n_3142;
wire n_3164;
wire n_3475;
wire n_1448;
wire n_2077;
wire n_3136;
wire n_2520;
wire n_2193;
wire n_2612;
wire n_3034;
wire n_2095;
wire n_3108;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2908;
wire n_2053;
wire n_2752;
wire n_1580;
wire n_2124;
wire n_1574;
wire n_2200;
wire n_1705;
wire n_3625;
wire n_2304;
wire n_1746;
wire n_2716;
wire n_1439;
wire n_2263;
wire n_2212;
wire n_2352;
wire n_3495;
wire n_2185;
wire n_3169;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2376;
wire n_2979;
wire n_3398;
wire n_1266;
wire n_1300;
wire n_3759;
wire n_2781;
wire n_3419;
wire n_3629;
wire n_2460;
wire n_2170;
wire n_3600;
wire n_1785;
wire n_1870;
wire n_2484;
wire n_2721;
wire n_1405;
wire n_2884;
wire n_3383;
wire n_3167;
wire n_3687;
wire n_997;
wire n_2308;
wire n_3459;
wire n_3498;
wire n_2986;
wire n_3238;
wire n_1428;
wire n_2691;
wire n_2243;
wire n_2400;
wire n_3731;
wire n_3092;
wire n_3555;
wire n_2903;
wire n_891;
wire n_3659;
wire n_3254;
wire n_2507;
wire n_2759;
wire n_3434;
wire n_1528;
wire n_1495;
wire n_3131;
wire n_3682;
wire n_2463;
wire n_2654;
wire n_3840;
wire n_2975;
wire n_1357;
wire n_2503;
wire n_2478;
wire n_3178;
wire n_2794;
wire n_1512;
wire n_3672;
wire n_2496;
wire n_3378;
wire n_3481;
wire n_2974;
wire n_2990;
wire n_2923;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_3449;
wire n_3517;
wire n_3350;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_3877;
wire n_945;
wire n_2925;
wire n_2270;
wire n_3260;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_2776;
wire n_1461;
wire n_3166;
wire n_2695;
wire n_2630;
wire n_903;
wire n_1967;
wire n_2340;
wire n_3385;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_3834;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_3656;
wire n_3257;
wire n_1048;
wire n_2459;
wire n_3137;
wire n_3116;
wire n_1925;
wire n_2439;
wire n_3638;
wire n_2106;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_3816;
wire n_2450;
wire n_1475;
wire n_3337;
wire n_2465;
wire n_1263;
wire n_3316;
wire n_1683;
wire n_1185;
wire n_3575;
wire n_1122;
wire n_2765;
wire n_3387;
wire n_890;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_1514;
wire n_964;
wire n_2728;
wire n_3772;
wire n_2948;
wire n_916;
wire n_3428;
wire n_2298;
wire n_2771;
wire n_3219;
wire n_2936;
wire n_895;
wire n_3867;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_2985;
wire n_1535;
wire n_3158;
wire n_3106;
wire n_2190;
wire n_1127;
wire n_932;
wire n_3657;
wire n_1972;
wire n_3080;
wire n_2772;
wire n_2778;
wire n_947;
wire n_1004;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_1667;
wire n_1845;
wire n_1104;
wire n_2205;
wire n_1011;
wire n_2684;
wire n_2875;
wire n_2524;
wire n_3284;
wire n_1437;
wire n_3835;
wire n_3723;
wire n_2747;
wire n_3389;
wire n_1707;
wire n_1941;
wire n_2422;
wire n_2064;
wire n_3088;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_3564;
wire n_2385;
wire n_3095;
wire n_3864;
wire n_3026;
wire n_2545;
wire n_1578;
wire n_3294;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_2712;
wire n_3695;
wire n_3279;
wire n_2584;
wire n_972;
wire n_1815;
wire n_2500;
wire n_3344;
wire n_1917;
wire n_1444;
wire n_920;
wire n_2442;
wire n_1067;
wire n_3328;
wire n_2763;
wire n_2788;
wire n_994;
wire n_2000;
wire n_2089;
wire n_1857;
wire n_2761;
wire n_1920;
wire n_2696;
wire n_3252;
wire n_887;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_2745;
wire n_1894;
wire n_2110;
wire n_2904;
wire n_2896;
wire n_3064;
wire n_3314;
wire n_3747;
wire n_961;
wire n_991;
wire n_1349;
wire n_1223;
wire n_1331;
wire n_2127;
wire n_3735;
wire n_1323;
wire n_1739;
wire n_3130;
wire n_1777;
wire n_3028;
wire n_3228;
wire n_3710;
wire n_1353;
wire n_3409;
wire n_2386;
wire n_3706;
wire n_3324;
wire n_1429;
wire n_3073;
wire n_2029;
wire n_3209;
wire n_2026;
wire n_1546;
wire n_3588;
wire n_3420;
wire n_1432;
wire n_2103;
wire n_3322;
wire n_1950;
wire n_1320;
wire n_996;
wire n_3632;
wire n_915;
wire n_2238;
wire n_2619;
wire n_3289;
wire n_1174;
wire n_1874;
wire n_1834;
wire n_3372;
wire n_3499;
wire n_3552;
wire n_2862;
wire n_3850;
wire n_3100;
wire n_3405;
wire n_1727;
wire n_3377;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_1601;
wire n_1294;
wire n_900;
wire n_3784;
wire n_3414;
wire n_1351;
wire n_2933;
wire n_2138;
wire n_1380;
wire n_1367;
wire n_3336;
wire n_3240;
wire n_3828;
wire n_1291;
wire n_3763;
wire n_2895;
wire n_1914;
wire n_3833;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_2271;
wire n_2356;
wire n_3339;
wire n_1830;
wire n_2261;
wire n_3016;
wire n_1629;
wire n_3476;
wire n_3673;
wire n_2842;
wire n_2994;
wire n_2011;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2105;
wire n_2187;
wire n_3556;
wire n_1340;
wire n_2694;
wire n_3443;
wire n_2562;
wire n_2642;
wire n_3029;
wire n_3269;
wire n_3609;
wire n_3447;
wire n_3771;
wire n_2647;
wire n_1626;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_2415;
wire n_3876;
wire n_3152;
wire n_3154;
wire n_2344;
wire n_3589;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2683;
wire n_2384;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_3432;
wire n_3523;
wire n_2815;
wire n_1816;
wire n_2446;
wire n_3388;
wire n_1612;
wire n_2318;
wire n_1172;
wire n_2659;
wire n_3616;
wire n_1099;
wire n_2141;
wire n_3113;
wire n_3696;
wire n_2902;
wire n_2909;
wire n_1422;
wire n_1527;
wire n_3174;
wire n_3608;
wire n_3190;
wire n_1524;
wire n_1055;
wire n_2849;
wire n_2947;
wire n_1754;
wire n_3048;
wire n_3686;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2566;
wire n_2679;
wire n_3292;
wire n_2210;
wire n_1517;
wire n_2502;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_982;
wire n_3670;
wire n_1624;
wire n_1952;
wire n_2180;
wire n_3002;
wire n_3376;
wire n_2087;
wire n_2920;
wire n_3290;
wire n_1598;
wire n_2952;
wire n_2617;
wire n_3585;
wire n_977;
wire n_2878;
wire n_1895;
wire n_2250;
wire n_1491;
wire n_1860;
wire n_2831;
wire n_1810;
wire n_1763;
wire n_923;
wire n_3778;
wire n_3818;
wire n_1607;
wire n_2865;
wire n_2075;
wire n_3047;
wire n_1625;
wire n_2959;
wire n_2610;
wire n_2420;
wire n_2380;
wire n_3335;
wire n_3265;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_2120;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_3669;
wire n_3427;
wire n_1289;
wire n_1348;
wire n_2892;
wire n_1021;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_3356;
wire n_1191;
wire n_2004;
wire n_3431;
wire n_3220;
wire n_2024;
wire n_3783;
wire n_2086;
wire n_1503;
wire n_3422;
wire n_1052;
wire n_1942;
wire n_3666;
wire n_3141;
wire n_2309;
wire n_2274;
wire n_2698;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_2330;
wire n_2555;
wire n_2639;
wire n_1259;
wire n_2108;
wire n_3099;
wire n_3712;
wire n_2535;
wire n_1001;
wire n_2945;
wire n_3057;
wire n_2143;
wire n_2410;
wire n_3760;
wire n_1396;
wire n_2916;
wire n_1224;
wire n_1923;
wire n_3206;
wire n_3736;
wire n_2196;
wire n_2739;
wire n_2611;
wire n_1538;
wire n_2528;
wire n_3773;
wire n_2548;
wire n_3216;
wire n_2709;
wire n_3061;
wire n_3717;
wire n_2633;
wire n_1017;
wire n_2244;
wire n_2604;
wire n_3462;
wire n_3424;
wire n_3745;
wire n_2351;
wire n_2437;
wire n_3664;
wire n_2049;
wire n_1456;
wire n_3245;
wire n_1889;
wire n_2113;
wire n_2665;
wire n_1124;
wire n_1690;
wire n_3063;
wire n_2688;
wire n_2881;
wire n_3862;
wire n_3302;
wire n_1673;
wire n_3361;
wire n_2018;
wire n_3134;
wire n_922;
wire n_2817;
wire n_1790;
wire n_993;
wire n_3196;
wire n_2085;
wire n_3304;
wire n_2581;
wire n_1725;
wire n_2809;
wire n_2149;
wire n_2237;
wire n_2268;
wire n_2320;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_1800;
wire n_3277;
wire n_3480;
wire n_2758;
wire n_3746;
wire n_1494;
wire n_1550;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_3474;
wire n_1169;
wire n_1726;
wire n_1946;
wire n_3111;
wire n_1938;
wire n_3452;
wire n_1241;
wire n_3645;
wire n_2589;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_2736;
wire n_1208;
wire n_1604;
wire n_1639;
wire n_2735;
wire n_2845;
wire n_3506;
wire n_1976;
wire n_2154;
wire n_2035;
wire n_1337;
wire n_2732;
wire n_3162;
wire n_2984;
wire n_1906;
wire n_3004;
wire n_1647;
wire n_1901;
wire n_3096;
wire n_3333;
wire n_3705;
wire n_3031;
wire n_1278;
wire n_2059;
wire n_3276;
wire n_1006;
wire n_2956;
wire n_1415;
wire n_1238;
wire n_3743;
wire n_976;
wire n_1710;
wire n_3021;
wire n_1063;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_2891;
wire n_2457;
wire n_3825;
wire n_2144;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_3404;
wire n_2072;
wire n_2737;
wire n_2012;
wire n_2251;
wire n_2963;
wire n_3512;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_3591;
wire n_1880;
wire n_1993;
wire n_3860;
wire n_2137;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_2182;
wire n_2868;
wire n_3044;
wire n_2447;
wire n_3493;
wire n_2818;
wire n_3358;
wire n_3115;
wire n_1057;
wire n_1473;
wire n_3140;
wire n_3486;
wire n_2125;
wire n_2426;
wire n_2894;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_2587;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_2099;
wire n_1202;
wire n_3848;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_3172;
wire n_905;
wire n_2159;
wire n_3410;
wire n_975;
wire n_934;
wire n_3273;
wire n_950;
wire n_2700;
wire n_1222;
wire n_3139;
wire n_1630;
wire n_3408;
wire n_2286;
wire n_3182;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_3734;
wire n_3637;
wire n_1311;
wire n_3393;
wire n_1261;
wire n_2299;
wire n_3538;
wire n_2078;
wire n_3650;
wire n_3327;
wire n_2265;
wire n_1114;
wire n_3513;
wire n_3709;
wire n_3011;
wire n_1167;
wire n_3231;
wire n_2677;
wire n_2531;
wire n_2315;
wire n_3623;
wire n_3647;
wire n_3138;
wire n_2157;
wire n_3212;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_1779;
wire n_3446;
wire n_3619;
wire n_3349;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_3454;
wire n_3058;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_2950;
wire n_919;
wire n_2272;
wire n_1956;
wire n_3574;
wire n_2608;
wire n_3384;
wire n_2983;
wire n_1718;
wire n_2225;
wire n_3229;
wire n_2546;
wire n_3739;
wire n_1411;
wire n_2825;
wire n_1139;
wire n_1018;
wire n_2345;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_2742;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_3540;
wire n_1838;
wire n_3649;
wire n_3604;
wire n_3824;
wire n_2680;
wire n_1343;
wire n_1801;
wire n_3439;
wire n_1371;
wire n_1513;
wire n_3740;
wire n_3001;
wire n_2861;
wire n_2976;
wire n_2161;
wire n_2191;
wire n_3611;
wire n_2329;
wire n_1788;
wire n_2093;
wire n_2576;
wire n_2348;
wire n_2417;
wire n_2675;
wire n_2043;
wire n_3601;
wire n_2366;
wire n_1621;
wire n_2338;
wire n_3571;
wire n_1919;
wire n_1342;
wire n_2756;
wire n_2893;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_3500;
wire n_1416;
wire n_1659;
wire n_2850;
wire n_3465;
wire n_1221;
wire n_3875;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_3846;
wire n_2851;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_2973;
wire n_3651;
wire n_1433;
wire n_1314;
wire n_2567;
wire n_3059;
wire n_3085;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_2810;
wire n_2867;
wire n_3871;
wire n_1085;
wire n_3027;
wire n_2388;
wire n_2981;
wire n_3438;
wire n_2222;
wire n_3112;
wire n_1907;
wire n_3464;
wire n_885;
wire n_1530;
wire n_3215;
wire n_3413;
wire n_2871;
wire n_2135;
wire n_1088;
wire n_896;
wire n_2764;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_3234;
wire n_3648;
wire n_2471;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_2757;
wire n_2714;
wire n_3066;
wire n_2669;
wire n_2869;
wire n_1105;
wire n_1459;
wire n_912;
wire n_2898;
wire n_2232;
wire n_3121;
wire n_2455;
wire n_2121;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_2874;
wire n_995;
wire n_2278;
wire n_1000;
wire n_2284;
wire n_1931;
wire n_2433;
wire n_2803;
wire n_2816;
wire n_3402;
wire n_1256;
wire n_2798;
wire n_3425;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_3308;
wire n_1526;
wire n_1507;
wire n_1809;
wire n_1206;
wire n_2367;
wire n_3236;
wire n_3576;
wire n_3491;
wire n_3109;
wire n_1961;
wire n_3271;
wire n_3013;
wire n_2553;
wire n_1050;
wire n_2218;
wire n_2667;
wire n_3062;
wire n_3806;
wire n_1769;
wire n_2130;
wire n_3256;
wire n_1060;
wire n_3126;
wire n_1372;
wire n_1847;
wire n_1565;
wire n_1257;
wire n_3805;
wire n_2325;
wire n_2406;
wire n_1632;
wire n_2864;
wire n_3346;
wire n_3104;
wire n_3391;
wire n_1547;
wire n_1586;
wire n_1542;
wire n_1362;
wire n_946;
wire n_3497;
wire n_1097;
wire n_3354;
wire n_3288;
wire n_3373;
wire n_3382;
wire n_3122;
wire n_2518;
wire n_2784;
wire n_3012;
wire n_3045;
wire n_1909;
wire n_2543;
wire n_3368;
wire n_2381;
wire n_2313;
wire n_3561;
wire n_3586;
wire n_956;
wire n_2495;
wire n_2992;
wire n_1541;
wire n_2703;
wire n_1812;
wire n_3014;
wire n_1951;
wire n_1330;
wire n_1697;
wire n_2128;
wire n_2574;
wire n_1872;
wire n_1940;
wire n_2690;
wire n_1747;
wire n_3767;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_3400;
wire n_2020;
wire n_3504;
wire n_1978;
wire n_2508;
wire n_3511;
wire n_2540;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_3820;
wire n_3159;
wire n_1768;
wire n_1443;
wire n_3697;
wire n_2068;
wire n_2636;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_3101;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_2593;
wire n_1623;
wire n_2911;
wire n_1828;
wire n_2364;
wire n_1389;
wire n_3303;
wire n_1131;
wire n_2641;
wire n_1798;
wire n_1077;
wire n_3120;
wire n_1554;
wire n_3549;
wire n_1481;
wire n_1584;
wire n_2021;
wire n_1928;
wire n_2713;
wire n_2938;
wire n_3227;
wire n_1438;
wire n_3774;
wire n_3342;
wire n_1973;
wire n_2314;
wire n_2939;
wire n_2156;
wire n_2494;
wire n_2126;
wire n_1147;
wire n_3403;
wire n_1363;
wire n_3863;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_1518;
wire n_1366;
wire n_1361;
wire n_1187;
wire n_2034;
wire n_1693;
wire n_3102;
wire n_2872;
wire n_3173;
wire n_2790;
wire n_2411;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_3539;
wire n_2266;
wire n_2993;
wire n_3433;
wire n_2061;
wire n_3018;
wire n_1373;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_3866;
wire n_3761;
wire n_2526;
wire n_2830;
wire n_1302;
wire n_3803;
wire n_3017;
wire n_3083;
wire n_2083;
wire n_886;
wire n_2119;
wire n_1010;
wire n_3844;
wire n_883;
wire n_2207;
wire n_2044;
wire n_2542;
wire n_2091;
wire n_2843;
wire n_3362;
wire n_3035;
wire n_3191;
wire n_1029;
wire n_3485;
wire n_2394;
wire n_3051;
wire n_1572;
wire n_1635;
wire n_3305;
wire n_3149;
wire n_2827;
wire n_941;
wire n_1245;
wire n_1317;
wire n_3643;
wire n_2615;
wire n_3278;
wire n_2487;
wire n_2701;
wire n_2929;
wire n_3163;
wire n_3343;
wire n_3752;
wire n_3786;
wire n_1329;
wire n_2409;
wire n_2637;
wire n_2337;
wire n_2405;
wire n_2601;
wire n_2513;
wire n_3118;
wire n_1297;
wire n_1912;
wire n_1369;
wire n_3143;
wire n_1734;
wire n_3543;
wire n_3655;
wire n_3742;
wire n_3791;
wire n_1876;
wire n_2666;
wire n_3050;
wire n_2323;
wire n_3532;
wire n_1811;
wire n_898;
wire n_928;
wire n_1285;
wire n_3042;
wire n_2997;
wire n_967;
wire n_2561;
wire n_3725;
wire n_2913;
wire n_2491;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_3522;
wire n_1486;
wire n_1068;
wire n_2914;
wire n_1833;
wire n_3551;
wire n_2371;
wire n_914;
wire n_3444;
wire n_1986;
wire n_3366;
wire n_2882;
wire n_1024;
wire n_3009;
wire n_1141;
wire n_3453;
wire n_3297;
wire n_3176;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2408;
wire n_2429;
wire n_3326;
wire n_1168;
wire n_3581;
wire n_3000;
wire n_2115;
wire n_2013;
wire n_2140;
wire n_2134;
wire n_2483;
wire n_2305;
wire n_1556;
wire n_3547;
wire n_3423;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_3700;
wire n_2514;
wire n_2466;
wire n_3661;
wire n_1759;
wire n_2048;
wire n_2760;
wire n_987;
wire n_1299;
wire n_2942;
wire n_2096;
wire n_3663;
wire n_2129;
wire n_3230;
wire n_3545;
wire n_1101;
wire n_2532;
wire n_3665;
wire n_2079;
wire n_2296;
wire n_3782;
wire n_1720;
wire n_880;
wire n_2671;
wire n_1911;
wire n_2293;
wire n_3296;
wire n_3831;
wire n_1336;
wire n_3068;
wire n_3071;
wire n_3683;
wire n_2734;
wire n_2870;
wire n_1166;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_1358;
wire n_2310;
wire n_3223;
wire n_3318;
wire n_1397;
wire n_1211;
wire n_2674;
wire n_1284;
wire n_2005;
wire n_3794;
wire n_1359;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_3226;
wire n_3702;
wire n_1532;
wire n_2848;
wire n_1419;
wire n_2689;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_3430;
wire n_3200;
wire n_1213;
wire n_2596;
wire n_2801;
wire n_1193;
wire n_980;
wire n_1488;
wire n_2928;
wire n_3067;
wire n_2227;
wire n_2652;
wire n_3225;
wire n_1074;
wire n_3380;
wire n_3557;
wire n_3207;
wire n_3596;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_2627;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_3606;
wire n_3369;
wire n_3823;
wire n_3185;
wire n_2326;
wire n_3869;
wire n_1866;
wire n_3852;
wire n_1220;
wire n_1398;
wire n_2169;
wire n_2111;
wire n_1904;
wire n_1262;
wire n_2966;
wire n_3084;
wire n_3036;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_960;
wire n_1022;
wire n_1760;
wire n_3737;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_3285;
wire n_3160;
wire n_3483;
wire n_1204;
wire n_1151;
wire n_2824;
wire n_1814;
wire n_2982;
wire n_999;
wire n_2634;
wire n_3124;
wire n_3286;
wire n_1092;
wire n_1808;
wire n_2768;
wire n_2668;
wire n_1658;
wire n_1386;
wire n_2588;
wire n_3015;
wire n_2931;
wire n_3321;
wire n_2492;
wire n_3081;
wire n_3636;
wire n_910;
wire n_2291;
wire n_3837;
wire n_3612;
wire n_3046;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_3076;
wire n_1385;
wire n_1142;
wire n_2927;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_3622;
wire n_3857;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_2155;
wire n_2706;
wire n_1868;
wire n_966;
wire n_2148;
wire n_2104;
wire n_949;
wire n_2357;
wire n_2303;
wire n_2618;
wire n_2653;
wire n_2855;
wire n_924;
wire n_2937;
wire n_3728;
wire n_3359;
wire n_3114;
wire n_2331;
wire n_3332;
wire n_1600;
wire n_1661;
wire n_2967;
wire n_1965;
wire n_3005;
wire n_1757;
wire n_2136;
wire n_3617;
wire n_3602;
wire n_2403;
wire n_918;
wire n_3053;
wire n_2056;
wire n_1913;
wire n_2702;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_2407;
wire n_2791;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_2302;
wire n_1450;
wire n_2082;
wire n_2560;
wire n_2453;
wire n_3056;
wire n_3267;
wire n_2092;
wire n_3008;
wire n_1472;
wire n_1365;
wire n_2443;
wire n_2802;
wire n_3189;
wire n_3052;
wire n_2797;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_2066;
wire n_1719;
wire n_1974;
wire n_1158;
wire n_2988;
wire n_1882;
wire n_2770;
wire n_2996;
wire n_2704;
wire n_2961;
wire n_1915;
wire n_2836;
wire n_940;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_3582;
wire n_3689;
wire n_3283;
wire n_1736;
wire n_3421;
wire n_2907;
wire n_3311;
wire n_1160;
wire n_1442;
wire n_2168;
wire n_1948;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1026;
wire n_3247;
wire n_2886;
wire n_1454;
wire n_1033;
wire n_3613;
wire n_990;
wire n_1383;
wire n_3675;
wire n_1968;
wire n_2057;
wire n_2609;
wire n_2378;
wire n_888;
wire n_2749;
wire n_3658;
wire n_1325;
wire n_3133;
wire n_2754;
wire n_3527;
wire n_2014;
wire n_3041;
wire n_1483;
wire n_1703;
wire n_1205;
wire n_1822;
wire n_1953;
wire n_3715;
wire n_1059;
wire n_2969;
wire n_3713;
wire n_2692;
wire n_3261;
wire n_3550;
wire n_1804;
wire n_1581;
wire n_3287;
wire n_3534;
wire n_1837;
wire n_3325;
wire n_1744;
wire n_1975;
wire n_3437;
wire n_3744;
wire n_1414;
wire n_2246;
wire n_2738;
wire n_2324;
wire n_3861;
wire n_3161;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_2940;
wire n_1111;
wire n_1819;
wire n_3313;
wire n_1341;
wire n_1807;
wire n_2670;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_3275;
wire n_1745;
wire n_1714;
wire n_3198;
wire n_3463;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_3516;
wire n_2262;
wire n_3562;
wire n_955;
wire n_1916;
wire n_1333;
wire n_2726;
wire n_2917;
wire n_3873;
wire n_3738;
wire n_2073;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_3157;
wire n_1551;
wire n_3793;
wire n_1533;
wire n_1145;
wire n_2307;
wire n_2515;
wire n_3792;
wire n_3546;
wire n_1511;
wire n_1791;
wire n_1113;
wire n_3089;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3406;
wire n_1468;
wire n_3442;
wire n_2327;
wire n_3758;
wire n_2656;
wire n_913;
wire n_2353;
wire n_1164;
wire n_2258;
wire n_3662;
wire n_3595;
wire n_1732;
wire n_3749;
wire n_2167;
wire n_3079;
wire n_1354;
wire n_3329;
wire n_2039;
wire n_1696;
wire n_1277;
wire n_1016;
wire n_3233;
wire n_1355;
wire n_3691;
wire n_2544;
wire n_3193;
wire n_3501;
wire n_3635;
wire n_2538;
wire n_3270;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_1280;
wire n_2854;
wire n_2932;
wire n_3258;
wire n_1335;
wire n_3266;
wire n_2285;
wire n_3213;
wire n_3789;
wire n_1934;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_3246;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_3418;
wire n_2435;
wire n_1665;
wire n_2583;
wire n_3417;
wire n_1678;
wire n_1091;
wire n_1780;
wire n_2725;
wire n_3865;
wire n_1287;
wire n_2769;
wire n_1482;
wire n_1525;
wire n_3244;
wire n_3195;
wire n_3593;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_2536;
wire n_2474;
wire n_1194;
wire n_1150;
wire n_1399;
wire n_3685;
wire n_3851;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_3768;
wire n_983;
wire n_1417;
wire n_3482;
wire n_2282;
wire n_970;
wire n_3654;
wire n_2430;
wire n_2676;
wire n_921;
wire n_2673;
wire n_3515;
wire n_3489;
wire n_2926;
wire n_1534;
wire n_2912;
wire n_3181;
wire n_908;
wire n_3536;
wire n_1346;
wire n_2834;
wire n_3644;
wire n_3268;
wire n_1123;
wire n_2710;
wire n_1272;
wire n_2497;
wire n_1393;
wire n_2970;
wire n_1655;
wire n_984;
wire n_3040;
wire n_3494;
wire n_2978;
wire n_3615;
wire n_1410;
wire n_988;
wire n_2368;
wire n_3363;
wire n_3528;
wire n_1157;
wire n_3502;
wire n_3677;
wire n_2657;
wire n_1186;
wire n_2065;
wire n_2901;
wire n_3180;
wire n_1743;
wire n_2743;
wire n_1854;
wire n_1506;
wire n_2658;

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_323),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_778),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_261),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_698),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_168),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_375),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_98),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_322),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_642),
.Y(n_888)
);

INVx1_ASAP7_75t_SL g889 ( 
.A(n_725),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_343),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_501),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_791),
.Y(n_892)
);

CKINVDCx20_ASAP7_75t_R g893 ( 
.A(n_704),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_714),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_314),
.Y(n_895)
);

CKINVDCx20_ASAP7_75t_R g896 ( 
.A(n_746),
.Y(n_896)
);

BUFx3_ASAP7_75t_L g897 ( 
.A(n_336),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_76),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_233),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_497),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_818),
.Y(n_901)
);

HB1xp67_ASAP7_75t_L g902 ( 
.A(n_831),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_814),
.Y(n_903)
);

INVx1_ASAP7_75t_SL g904 ( 
.A(n_125),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_276),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_347),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_784),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_862),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_77),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_843),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_57),
.Y(n_911)
);

BUFx5_ASAP7_75t_L g912 ( 
.A(n_84),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_647),
.Y(n_913)
);

CKINVDCx20_ASAP7_75t_R g914 ( 
.A(n_201),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_354),
.Y(n_915)
);

INVx2_ASAP7_75t_SL g916 ( 
.A(n_208),
.Y(n_916)
);

BUFx3_ASAP7_75t_L g917 ( 
.A(n_56),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_101),
.Y(n_918)
);

CKINVDCx16_ASAP7_75t_R g919 ( 
.A(n_688),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_850),
.Y(n_920)
);

INVx3_ASAP7_75t_L g921 ( 
.A(n_10),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_611),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_837),
.Y(n_923)
);

CKINVDCx20_ASAP7_75t_R g924 ( 
.A(n_860),
.Y(n_924)
);

INVx2_ASAP7_75t_SL g925 ( 
.A(n_528),
.Y(n_925)
);

BUFx3_ASAP7_75t_L g926 ( 
.A(n_773),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_155),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_269),
.Y(n_928)
);

INVx1_ASAP7_75t_SL g929 ( 
.A(n_852),
.Y(n_929)
);

INVx2_ASAP7_75t_SL g930 ( 
.A(n_396),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_286),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_647),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_380),
.Y(n_933)
);

BUFx10_ASAP7_75t_L g934 ( 
.A(n_855),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_398),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_115),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_774),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_822),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_811),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_867),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_790),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_291),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_232),
.Y(n_943)
);

CKINVDCx20_ASAP7_75t_R g944 ( 
.A(n_859),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_879),
.Y(n_945)
);

BUFx6f_ASAP7_75t_L g946 ( 
.A(n_675),
.Y(n_946)
);

BUFx10_ASAP7_75t_L g947 ( 
.A(n_37),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_224),
.Y(n_948)
);

BUFx5_ASAP7_75t_L g949 ( 
.A(n_595),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_809),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_111),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_639),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_873),
.Y(n_953)
);

BUFx3_ASAP7_75t_L g954 ( 
.A(n_537),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_820),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_591),
.Y(n_956)
);

INVx1_ASAP7_75t_SL g957 ( 
.A(n_746),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_385),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_694),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_874),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_81),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_564),
.Y(n_962)
);

BUFx2_ASAP7_75t_L g963 ( 
.A(n_378),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_821),
.Y(n_964)
);

BUFx6f_ASAP7_75t_L g965 ( 
.A(n_766),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_695),
.Y(n_966)
);

CKINVDCx16_ASAP7_75t_R g967 ( 
.A(n_854),
.Y(n_967)
);

INVx2_ASAP7_75t_SL g968 ( 
.A(n_290),
.Y(n_968)
);

CKINVDCx20_ASAP7_75t_R g969 ( 
.A(n_30),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_199),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_753),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_619),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_447),
.Y(n_973)
);

INVx1_ASAP7_75t_SL g974 ( 
.A(n_824),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_795),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_302),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_208),
.Y(n_977)
);

CKINVDCx20_ASAP7_75t_R g978 ( 
.A(n_515),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_878),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_646),
.Y(n_980)
);

INVxp67_ASAP7_75t_L g981 ( 
.A(n_423),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_451),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_144),
.Y(n_983)
);

BUFx10_ASAP7_75t_L g984 ( 
.A(n_772),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_275),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_234),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_197),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_414),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_234),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_439),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_121),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_302),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_512),
.Y(n_993)
);

CKINVDCx16_ASAP7_75t_R g994 ( 
.A(n_627),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_166),
.Y(n_995)
);

CKINVDCx20_ASAP7_75t_R g996 ( 
.A(n_308),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_270),
.Y(n_997)
);

HB1xp67_ASAP7_75t_L g998 ( 
.A(n_290),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_202),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_845),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_294),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_720),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_539),
.Y(n_1003)
);

CKINVDCx20_ASAP7_75t_R g1004 ( 
.A(n_693),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_842),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_329),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_82),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_249),
.Y(n_1008)
);

BUFx2_ASAP7_75t_L g1009 ( 
.A(n_354),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_758),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_343),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_789),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_355),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_296),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_817),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_147),
.Y(n_1016)
);

BUFx2_ASAP7_75t_L g1017 ( 
.A(n_787),
.Y(n_1017)
);

HB1xp67_ASAP7_75t_L g1018 ( 
.A(n_695),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_360),
.Y(n_1019)
);

BUFx10_ASAP7_75t_L g1020 ( 
.A(n_296),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_123),
.Y(n_1021)
);

BUFx10_ASAP7_75t_L g1022 ( 
.A(n_221),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_30),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_258),
.Y(n_1024)
);

INVx1_ASAP7_75t_SL g1025 ( 
.A(n_114),
.Y(n_1025)
);

INVxp67_ASAP7_75t_R g1026 ( 
.A(n_189),
.Y(n_1026)
);

BUFx3_ASAP7_75t_L g1027 ( 
.A(n_869),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_675),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_653),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_338),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_853),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_845),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_832),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_170),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_863),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_293),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_867),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_608),
.Y(n_1038)
);

HB1xp67_ASAP7_75t_L g1039 ( 
.A(n_866),
.Y(n_1039)
);

BUFx8_ASAP7_75t_SL g1040 ( 
.A(n_855),
.Y(n_1040)
);

BUFx6f_ASAP7_75t_L g1041 ( 
.A(n_826),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_264),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_524),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_865),
.Y(n_1044)
);

CKINVDCx20_ASAP7_75t_R g1045 ( 
.A(n_801),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_567),
.Y(n_1046)
);

BUFx2_ASAP7_75t_L g1047 ( 
.A(n_541),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_191),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_768),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_767),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_671),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_72),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_23),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_782),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_836),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_802),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_30),
.Y(n_1057)
);

INVx1_ASAP7_75t_SL g1058 ( 
.A(n_558),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_612),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_327),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_281),
.Y(n_1061)
);

INVxp33_ASAP7_75t_R g1062 ( 
.A(n_777),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_796),
.Y(n_1063)
);

INVxp67_ASAP7_75t_L g1064 ( 
.A(n_830),
.Y(n_1064)
);

BUFx10_ASAP7_75t_L g1065 ( 
.A(n_97),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_199),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_553),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_781),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_127),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_562),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_588),
.Y(n_1071)
);

CKINVDCx20_ASAP7_75t_R g1072 ( 
.A(n_751),
.Y(n_1072)
);

BUFx6f_ASAP7_75t_L g1073 ( 
.A(n_571),
.Y(n_1073)
);

CKINVDCx14_ASAP7_75t_R g1074 ( 
.A(n_579),
.Y(n_1074)
);

INVx1_ASAP7_75t_SL g1075 ( 
.A(n_786),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_833),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_265),
.Y(n_1077)
);

BUFx6f_ASAP7_75t_L g1078 ( 
.A(n_140),
.Y(n_1078)
);

CKINVDCx20_ASAP7_75t_R g1079 ( 
.A(n_490),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_466),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_461),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_153),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_64),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_427),
.Y(n_1084)
);

INVx1_ASAP7_75t_SL g1085 ( 
.A(n_28),
.Y(n_1085)
);

CKINVDCx16_ASAP7_75t_R g1086 ( 
.A(n_372),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_858),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_840),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_177),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_436),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_577),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_243),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_625),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_868),
.Y(n_1094)
);

INVx2_ASAP7_75t_SL g1095 ( 
.A(n_390),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_850),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_696),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_597),
.Y(n_1098)
);

BUFx6f_ASAP7_75t_L g1099 ( 
.A(n_632),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_482),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_844),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_257),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_547),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_750),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_715),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_629),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_478),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_88),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_801),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_616),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_718),
.Y(n_1111)
);

HB1xp67_ASAP7_75t_L g1112 ( 
.A(n_582),
.Y(n_1112)
);

CKINVDCx20_ASAP7_75t_R g1113 ( 
.A(n_23),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_385),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_831),
.Y(n_1115)
);

CKINVDCx20_ASAP7_75t_R g1116 ( 
.A(n_825),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_656),
.Y(n_1117)
);

BUFx8_ASAP7_75t_SL g1118 ( 
.A(n_800),
.Y(n_1118)
);

BUFx10_ASAP7_75t_L g1119 ( 
.A(n_545),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_753),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_52),
.Y(n_1121)
);

CKINVDCx20_ASAP7_75t_R g1122 ( 
.A(n_697),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_35),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_626),
.Y(n_1124)
);

BUFx2_ASAP7_75t_L g1125 ( 
.A(n_154),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_22),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_466),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_856),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_583),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_181),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_793),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_648),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_372),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_573),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_875),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_307),
.Y(n_1136)
);

BUFx3_ASAP7_75t_L g1137 ( 
.A(n_634),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_583),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_724),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_125),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_165),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_631),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_478),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_83),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_55),
.Y(n_1145)
);

CKINVDCx20_ASAP7_75t_R g1146 ( 
.A(n_55),
.Y(n_1146)
);

CKINVDCx20_ASAP7_75t_R g1147 ( 
.A(n_584),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_365),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_321),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_643),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_221),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_729),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_851),
.Y(n_1153)
);

BUFx3_ASAP7_75t_L g1154 ( 
.A(n_727),
.Y(n_1154)
);

BUFx6f_ASAP7_75t_L g1155 ( 
.A(n_131),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_829),
.Y(n_1156)
);

INVxp67_ASAP7_75t_L g1157 ( 
.A(n_467),
.Y(n_1157)
);

INVx1_ASAP7_75t_SL g1158 ( 
.A(n_828),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_839),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_815),
.Y(n_1160)
);

CKINVDCx16_ASAP7_75t_R g1161 ( 
.A(n_520),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_791),
.Y(n_1162)
);

BUFx6f_ASAP7_75t_L g1163 ( 
.A(n_803),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_236),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_291),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_701),
.Y(n_1166)
);

BUFx3_ASAP7_75t_L g1167 ( 
.A(n_482),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_85),
.Y(n_1168)
);

BUFx6f_ASAP7_75t_L g1169 ( 
.A(n_208),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_846),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_288),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_841),
.Y(n_1172)
);

BUFx6f_ASAP7_75t_L g1173 ( 
.A(n_598),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_779),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_857),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_667),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_397),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_409),
.Y(n_1178)
);

INVx1_ASAP7_75t_SL g1179 ( 
.A(n_304),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_655),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_428),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_419),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_395),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_239),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_459),
.Y(n_1185)
);

BUFx6f_ASAP7_75t_L g1186 ( 
.A(n_285),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_658),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_7),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_105),
.Y(n_1189)
);

BUFx6f_ASAP7_75t_L g1190 ( 
.A(n_427),
.Y(n_1190)
);

INVxp67_ASAP7_75t_L g1191 ( 
.A(n_770),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_716),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_273),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_28),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_391),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_521),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_654),
.Y(n_1197)
);

CKINVDCx11_ASAP7_75t_R g1198 ( 
.A(n_593),
.Y(n_1198)
);

BUFx6f_ASAP7_75t_L g1199 ( 
.A(n_804),
.Y(n_1199)
);

CKINVDCx20_ASAP7_75t_R g1200 ( 
.A(n_785),
.Y(n_1200)
);

BUFx3_ASAP7_75t_L g1201 ( 
.A(n_439),
.Y(n_1201)
);

INVxp67_ASAP7_75t_L g1202 ( 
.A(n_340),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_26),
.Y(n_1203)
);

BUFx10_ASAP7_75t_L g1204 ( 
.A(n_726),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_805),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_835),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_349),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_31),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_435),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_563),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_639),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_43),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_819),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_477),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_761),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_812),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_699),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_799),
.Y(n_1218)
);

BUFx5_ASAP7_75t_L g1219 ( 
.A(n_769),
.Y(n_1219)
);

CKINVDCx20_ASAP7_75t_R g1220 ( 
.A(n_506),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_430),
.Y(n_1221)
);

CKINVDCx20_ASAP7_75t_R g1222 ( 
.A(n_868),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_398),
.Y(n_1223)
);

INVx1_ASAP7_75t_SL g1224 ( 
.A(n_43),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_487),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_654),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_823),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_116),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_662),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_827),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_700),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_807),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_630),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_15),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_604),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_775),
.Y(n_1236)
);

CKINVDCx20_ASAP7_75t_R g1237 ( 
.A(n_763),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_645),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_714),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_864),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_501),
.Y(n_1241)
);

BUFx10_ASAP7_75t_L g1242 ( 
.A(n_871),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_712),
.Y(n_1243)
);

BUFx3_ASAP7_75t_L g1244 ( 
.A(n_293),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_97),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_161),
.Y(n_1246)
);

CKINVDCx20_ASAP7_75t_R g1247 ( 
.A(n_49),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_16),
.Y(n_1248)
);

INVx1_ASAP7_75t_SL g1249 ( 
.A(n_164),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_691),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_145),
.Y(n_1251)
);

BUFx6f_ASAP7_75t_L g1252 ( 
.A(n_700),
.Y(n_1252)
);

INVx1_ASAP7_75t_SL g1253 ( 
.A(n_783),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_810),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_39),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_639),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_104),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_816),
.Y(n_1258)
);

BUFx6f_ASAP7_75t_L g1259 ( 
.A(n_729),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_638),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_389),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_597),
.Y(n_1262)
);

CKINVDCx20_ASAP7_75t_R g1263 ( 
.A(n_578),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_631),
.Y(n_1264)
);

CKINVDCx5p33_ASAP7_75t_R g1265 ( 
.A(n_828),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_374),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_565),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_764),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_497),
.Y(n_1269)
);

CKINVDCx5p33_ASAP7_75t_R g1270 ( 
.A(n_709),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_135),
.Y(n_1271)
);

INVxp67_ASAP7_75t_L g1272 ( 
.A(n_702),
.Y(n_1272)
);

CKINVDCx5p33_ASAP7_75t_R g1273 ( 
.A(n_21),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_730),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_168),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_739),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_780),
.Y(n_1277)
);

BUFx10_ASAP7_75t_L g1278 ( 
.A(n_530),
.Y(n_1278)
);

CKINVDCx5p33_ASAP7_75t_R g1279 ( 
.A(n_725),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_1),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_865),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_388),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_633),
.Y(n_1283)
);

CKINVDCx16_ASAP7_75t_R g1284 ( 
.A(n_130),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_730),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_95),
.Y(n_1286)
);

CKINVDCx20_ASAP7_75t_R g1287 ( 
.A(n_688),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_848),
.Y(n_1288)
);

CKINVDCx5p33_ASAP7_75t_R g1289 ( 
.A(n_649),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_81),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_350),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_446),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_771),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_672),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_383),
.Y(n_1295)
);

CKINVDCx5p33_ASAP7_75t_R g1296 ( 
.A(n_146),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_564),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_393),
.Y(n_1298)
);

CKINVDCx20_ASAP7_75t_R g1299 ( 
.A(n_870),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_240),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_629),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_759),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_877),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_118),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_482),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_798),
.Y(n_1306)
);

CKINVDCx20_ASAP7_75t_R g1307 ( 
.A(n_61),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_492),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_834),
.Y(n_1309)
);

CKINVDCx16_ASAP7_75t_R g1310 ( 
.A(n_728),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_529),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_847),
.Y(n_1312)
);

CKINVDCx5p33_ASAP7_75t_R g1313 ( 
.A(n_187),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_674),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_92),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_661),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_788),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_567),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_640),
.Y(n_1319)
);

CKINVDCx20_ASAP7_75t_R g1320 ( 
.A(n_351),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_772),
.Y(n_1321)
);

INVx2_ASAP7_75t_L g1322 ( 
.A(n_121),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_274),
.Y(n_1323)
);

CKINVDCx5p33_ASAP7_75t_R g1324 ( 
.A(n_741),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_588),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_433),
.Y(n_1326)
);

INVxp33_ASAP7_75t_L g1327 ( 
.A(n_681),
.Y(n_1327)
);

INVx1_ASAP7_75t_SL g1328 ( 
.A(n_390),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_808),
.Y(n_1329)
);

BUFx3_ASAP7_75t_L g1330 ( 
.A(n_806),
.Y(n_1330)
);

CKINVDCx5p33_ASAP7_75t_R g1331 ( 
.A(n_760),
.Y(n_1331)
);

CKINVDCx20_ASAP7_75t_R g1332 ( 
.A(n_307),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_697),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_359),
.Y(n_1334)
);

CKINVDCx5p33_ASAP7_75t_R g1335 ( 
.A(n_132),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_679),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_44),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_860),
.Y(n_1338)
);

CKINVDCx20_ASAP7_75t_R g1339 ( 
.A(n_750),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_756),
.Y(n_1340)
);

CKINVDCx20_ASAP7_75t_R g1341 ( 
.A(n_642),
.Y(n_1341)
);

CKINVDCx5p33_ASAP7_75t_R g1342 ( 
.A(n_861),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_163),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_872),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_792),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_797),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_132),
.Y(n_1347)
);

INVx1_ASAP7_75t_SL g1348 ( 
.A(n_762),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_407),
.Y(n_1349)
);

BUFx2_ASAP7_75t_L g1350 ( 
.A(n_667),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_189),
.Y(n_1351)
);

BUFx10_ASAP7_75t_L g1352 ( 
.A(n_837),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_506),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_530),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_328),
.Y(n_1355)
);

CKINVDCx5p33_ASAP7_75t_R g1356 ( 
.A(n_357),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_585),
.Y(n_1357)
);

CKINVDCx20_ASAP7_75t_R g1358 ( 
.A(n_338),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_652),
.Y(n_1359)
);

CKINVDCx5p33_ASAP7_75t_R g1360 ( 
.A(n_766),
.Y(n_1360)
);

CKINVDCx5p33_ASAP7_75t_R g1361 ( 
.A(n_636),
.Y(n_1361)
);

BUFx2_ASAP7_75t_L g1362 ( 
.A(n_472),
.Y(n_1362)
);

CKINVDCx5p33_ASAP7_75t_R g1363 ( 
.A(n_315),
.Y(n_1363)
);

CKINVDCx5p33_ASAP7_75t_R g1364 ( 
.A(n_15),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_662),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_239),
.Y(n_1366)
);

CKINVDCx5p33_ASAP7_75t_R g1367 ( 
.A(n_54),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_123),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_518),
.Y(n_1369)
);

BUFx6f_ASAP7_75t_L g1370 ( 
.A(n_765),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_528),
.Y(n_1371)
);

CKINVDCx5p33_ASAP7_75t_R g1372 ( 
.A(n_776),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_876),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_745),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_692),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_32),
.Y(n_1376)
);

BUFx6f_ASAP7_75t_L g1377 ( 
.A(n_838),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_348),
.Y(n_1378)
);

CKINVDCx5p33_ASAP7_75t_R g1379 ( 
.A(n_538),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_427),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_608),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_739),
.Y(n_1382)
);

CKINVDCx5p33_ASAP7_75t_R g1383 ( 
.A(n_849),
.Y(n_1383)
);

BUFx2_ASAP7_75t_L g1384 ( 
.A(n_406),
.Y(n_1384)
);

INVx1_ASAP7_75t_SL g1385 ( 
.A(n_635),
.Y(n_1385)
);

CKINVDCx5p33_ASAP7_75t_R g1386 ( 
.A(n_794),
.Y(n_1386)
);

CKINVDCx5p33_ASAP7_75t_R g1387 ( 
.A(n_857),
.Y(n_1387)
);

CKINVDCx20_ASAP7_75t_R g1388 ( 
.A(n_851),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_741),
.Y(n_1389)
);

CKINVDCx5p33_ASAP7_75t_R g1390 ( 
.A(n_691),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_248),
.Y(n_1391)
);

CKINVDCx5p33_ASAP7_75t_R g1392 ( 
.A(n_217),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_424),
.Y(n_1393)
);

CKINVDCx5p33_ASAP7_75t_R g1394 ( 
.A(n_687),
.Y(n_1394)
);

BUFx10_ASAP7_75t_L g1395 ( 
.A(n_331),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_813),
.Y(n_1396)
);

INVx2_ASAP7_75t_SL g1397 ( 
.A(n_49),
.Y(n_1397)
);

INVx2_ASAP7_75t_SL g1398 ( 
.A(n_752),
.Y(n_1398)
);

CKINVDCx5p33_ASAP7_75t_R g1399 ( 
.A(n_1198),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_916),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_925),
.Y(n_1401)
);

CKINVDCx5p33_ASAP7_75t_R g1402 ( 
.A(n_1198),
.Y(n_1402)
);

BUFx2_ASAP7_75t_L g1403 ( 
.A(n_1074),
.Y(n_1403)
);

INVxp67_ASAP7_75t_L g1404 ( 
.A(n_963),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_930),
.Y(n_1405)
);

NOR2xp33_ASAP7_75t_L g1406 ( 
.A(n_1017),
.B(n_0),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_1074),
.Y(n_1407)
);

INVxp67_ASAP7_75t_SL g1408 ( 
.A(n_921),
.Y(n_1408)
);

CKINVDCx5p33_ASAP7_75t_R g1409 ( 
.A(n_1040),
.Y(n_1409)
);

CKINVDCx20_ASAP7_75t_R g1410 ( 
.A(n_914),
.Y(n_1410)
);

NOR2xp33_ASAP7_75t_L g1411 ( 
.A(n_1350),
.B(n_0),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_968),
.Y(n_1412)
);

CKINVDCx20_ASAP7_75t_R g1413 ( 
.A(n_914),
.Y(n_1413)
);

HB1xp67_ASAP7_75t_L g1414 ( 
.A(n_998),
.Y(n_1414)
);

BUFx3_ASAP7_75t_L g1415 ( 
.A(n_926),
.Y(n_1415)
);

INVxp67_ASAP7_75t_SL g1416 ( 
.A(n_921),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1095),
.Y(n_1417)
);

INVxp67_ASAP7_75t_L g1418 ( 
.A(n_1009),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1397),
.Y(n_1419)
);

CKINVDCx20_ASAP7_75t_R g1420 ( 
.A(n_969),
.Y(n_1420)
);

INVxp67_ASAP7_75t_L g1421 ( 
.A(n_1047),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1125),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1362),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1384),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1112),
.Y(n_1425)
);

HB1xp67_ASAP7_75t_L g1426 ( 
.A(n_902),
.Y(n_1426)
);

CKINVDCx5p33_ASAP7_75t_R g1427 ( 
.A(n_1040),
.Y(n_1427)
);

INVx1_ASAP7_75t_SL g1428 ( 
.A(n_880),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_1118),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_899),
.Y(n_1430)
);

HB1xp67_ASAP7_75t_L g1431 ( 
.A(n_1018),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_900),
.Y(n_1432)
);

CKINVDCx20_ASAP7_75t_R g1433 ( 
.A(n_969),
.Y(n_1433)
);

BUFx2_ASAP7_75t_L g1434 ( 
.A(n_994),
.Y(n_1434)
);

NOR2xp33_ASAP7_75t_L g1435 ( 
.A(n_1327),
.B(n_0),
.Y(n_1435)
);

HB1xp67_ASAP7_75t_L g1436 ( 
.A(n_1039),
.Y(n_1436)
);

CKINVDCx5p33_ASAP7_75t_R g1437 ( 
.A(n_1086),
.Y(n_1437)
);

BUFx6f_ASAP7_75t_L g1438 ( 
.A(n_1073),
.Y(n_1438)
);

CKINVDCx20_ASAP7_75t_R g1439 ( 
.A(n_1146),
.Y(n_1439)
);

CKINVDCx5p33_ASAP7_75t_R g1440 ( 
.A(n_1161),
.Y(n_1440)
);

CKINVDCx5p33_ASAP7_75t_R g1441 ( 
.A(n_1284),
.Y(n_1441)
);

CKINVDCx5p33_ASAP7_75t_R g1442 ( 
.A(n_884),
.Y(n_1442)
);

CKINVDCx5p33_ASAP7_75t_R g1443 ( 
.A(n_885),
.Y(n_1443)
);

CKINVDCx5p33_ASAP7_75t_R g1444 ( 
.A(n_886),
.Y(n_1444)
);

CKINVDCx16_ASAP7_75t_R g1445 ( 
.A(n_919),
.Y(n_1445)
);

HB1xp67_ASAP7_75t_L g1446 ( 
.A(n_981),
.Y(n_1446)
);

NOR2xp33_ASAP7_75t_L g1447 ( 
.A(n_1327),
.B(n_1),
.Y(n_1447)
);

CKINVDCx5p33_ASAP7_75t_R g1448 ( 
.A(n_887),
.Y(n_1448)
);

NOR2xp33_ASAP7_75t_L g1449 ( 
.A(n_1398),
.B(n_1),
.Y(n_1449)
);

CKINVDCx5p33_ASAP7_75t_R g1450 ( 
.A(n_888),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_905),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_927),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_932),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_933),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_943),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_948),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_970),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_972),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1219),
.Y(n_1459)
);

CKINVDCx5p33_ASAP7_75t_R g1460 ( 
.A(n_890),
.Y(n_1460)
);

NOR2xp33_ASAP7_75t_R g1461 ( 
.A(n_891),
.B(n_2),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_977),
.Y(n_1462)
);

BUFx2_ASAP7_75t_L g1463 ( 
.A(n_897),
.Y(n_1463)
);

INVxp67_ASAP7_75t_SL g1464 ( 
.A(n_897),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_985),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_999),
.Y(n_1466)
);

CKINVDCx5p33_ASAP7_75t_R g1467 ( 
.A(n_895),
.Y(n_1467)
);

CKINVDCx20_ASAP7_75t_R g1468 ( 
.A(n_1147),
.Y(n_1468)
);

CKINVDCx5p33_ASAP7_75t_R g1469 ( 
.A(n_898),
.Y(n_1469)
);

INVxp67_ASAP7_75t_SL g1470 ( 
.A(n_917),
.Y(n_1470)
);

INVxp33_ASAP7_75t_SL g1471 ( 
.A(n_1026),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_906),
.B(n_2),
.Y(n_1472)
);

BUFx6f_ASAP7_75t_L g1473 ( 
.A(n_1073),
.Y(n_1473)
);

HB1xp67_ASAP7_75t_L g1474 ( 
.A(n_1157),
.Y(n_1474)
);

CKINVDCx5p33_ASAP7_75t_R g1475 ( 
.A(n_909),
.Y(n_1475)
);

CKINVDCx5p33_ASAP7_75t_R g1476 ( 
.A(n_911),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1014),
.Y(n_1477)
);

CKINVDCx5p33_ASAP7_75t_R g1478 ( 
.A(n_913),
.Y(n_1478)
);

CKINVDCx5p33_ASAP7_75t_R g1479 ( 
.A(n_915),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1019),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1023),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1024),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1029),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1030),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1034),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1042),
.Y(n_1486)
);

CKINVDCx5p33_ASAP7_75t_R g1487 ( 
.A(n_918),
.Y(n_1487)
);

NOR2xp33_ASAP7_75t_L g1488 ( 
.A(n_1064),
.B(n_2),
.Y(n_1488)
);

CKINVDCx5p33_ASAP7_75t_R g1489 ( 
.A(n_928),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_931),
.Y(n_1490)
);

CKINVDCx5p33_ASAP7_75t_R g1491 ( 
.A(n_935),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1046),
.Y(n_1492)
);

INVxp67_ASAP7_75t_L g1493 ( 
.A(n_917),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1048),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1219),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1052),
.Y(n_1496)
);

HB1xp67_ASAP7_75t_L g1497 ( 
.A(n_1202),
.Y(n_1497)
);

NOR2xp33_ASAP7_75t_L g1498 ( 
.A(n_1191),
.B(n_3),
.Y(n_1498)
);

CKINVDCx20_ASAP7_75t_R g1499 ( 
.A(n_1220),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1053),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1057),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1059),
.Y(n_1502)
);

CKINVDCx5p33_ASAP7_75t_R g1503 ( 
.A(n_936),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1067),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1071),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1081),
.Y(n_1506)
);

CKINVDCx5p33_ASAP7_75t_R g1507 ( 
.A(n_942),
.Y(n_1507)
);

INVxp67_ASAP7_75t_SL g1508 ( 
.A(n_954),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_951),
.B(n_3),
.Y(n_1509)
);

CKINVDCx20_ASAP7_75t_R g1510 ( 
.A(n_1220),
.Y(n_1510)
);

INVx4_ASAP7_75t_L g1511 ( 
.A(n_1403),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1463),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1493),
.Y(n_1513)
);

INVxp67_ASAP7_75t_L g1514 ( 
.A(n_1434),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1493),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1415),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1408),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1416),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1464),
.Y(n_1519)
);

HB1xp67_ASAP7_75t_L g1520 ( 
.A(n_1414),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1495),
.Y(n_1521)
);

HB1xp67_ASAP7_75t_L g1522 ( 
.A(n_1428),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1404),
.B(n_952),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1404),
.B(n_956),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1470),
.Y(n_1525)
);

NOR2xp33_ASAP7_75t_L g1526 ( 
.A(n_1400),
.B(n_1272),
.Y(n_1526)
);

BUFx6f_ASAP7_75t_L g1527 ( 
.A(n_1438),
.Y(n_1527)
);

BUFx6f_ASAP7_75t_L g1528 ( 
.A(n_1438),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1508),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1401),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1405),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1412),
.Y(n_1532)
);

INVxp67_ASAP7_75t_L g1533 ( 
.A(n_1446),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1417),
.Y(n_1534)
);

INVx2_ASAP7_75t_SL g1535 ( 
.A(n_1442),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1418),
.B(n_947),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1419),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1418),
.B(n_958),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1430),
.Y(n_1539)
);

INVxp67_ASAP7_75t_L g1540 ( 
.A(n_1474),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1432),
.Y(n_1541)
);

BUFx6f_ASAP7_75t_L g1542 ( 
.A(n_1438),
.Y(n_1542)
);

CKINVDCx20_ASAP7_75t_R g1543 ( 
.A(n_1410),
.Y(n_1543)
);

NAND2xp33_ASAP7_75t_L g1544 ( 
.A(n_1407),
.B(n_912),
.Y(n_1544)
);

OAI22xp5_ASAP7_75t_SL g1545 ( 
.A1(n_1413),
.A2(n_978),
.B1(n_1079),
.B2(n_996),
.Y(n_1545)
);

INVx4_ASAP7_75t_L g1546 ( 
.A(n_1443),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1451),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1452),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1421),
.B(n_1497),
.Y(n_1549)
);

NOR2xp33_ASAP7_75t_L g1550 ( 
.A(n_1471),
.B(n_967),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1421),
.B(n_961),
.Y(n_1551)
);

AND2x4_ASAP7_75t_L g1552 ( 
.A(n_1422),
.B(n_926),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1453),
.Y(n_1553)
);

HB1xp67_ASAP7_75t_L g1554 ( 
.A(n_1444),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1454),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1426),
.B(n_947),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1455),
.Y(n_1557)
);

NAND2x1_ASAP7_75t_L g1558 ( 
.A(n_1456),
.B(n_882),
.Y(n_1558)
);

HB1xp67_ASAP7_75t_L g1559 ( 
.A(n_1448),
.Y(n_1559)
);

BUFx8_ASAP7_75t_L g1560 ( 
.A(n_1425),
.Y(n_1560)
);

AND2x4_ASAP7_75t_L g1561 ( 
.A(n_1423),
.B(n_1027),
.Y(n_1561)
);

OA21x2_ASAP7_75t_L g1562 ( 
.A1(n_1457),
.A2(n_922),
.B(n_882),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1431),
.B(n_1020),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1436),
.B(n_1424),
.Y(n_1564)
);

AND2x4_ASAP7_75t_L g1565 ( 
.A(n_1458),
.B(n_1462),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1465),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1466),
.Y(n_1567)
);

BUFx6f_ASAP7_75t_L g1568 ( 
.A(n_1473),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1445),
.B(n_1020),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1477),
.B(n_962),
.Y(n_1570)
);

BUFx3_ASAP7_75t_L g1571 ( 
.A(n_1450),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_1480),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1481),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1482),
.Y(n_1574)
);

BUFx6f_ASAP7_75t_L g1575 ( 
.A(n_1473),
.Y(n_1575)
);

OA21x2_ASAP7_75t_L g1576 ( 
.A1(n_1483),
.A2(n_973),
.B(n_922),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1484),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1485),
.Y(n_1578)
);

AND2x4_ASAP7_75t_L g1579 ( 
.A(n_1486),
.B(n_1027),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1492),
.Y(n_1580)
);

HB1xp67_ASAP7_75t_L g1581 ( 
.A(n_1460),
.Y(n_1581)
);

INVx3_ASAP7_75t_L g1582 ( 
.A(n_1494),
.Y(n_1582)
);

BUFx3_ASAP7_75t_L g1583 ( 
.A(n_1467),
.Y(n_1583)
);

INVx3_ASAP7_75t_L g1584 ( 
.A(n_1496),
.Y(n_1584)
);

AOI22xp5_ASAP7_75t_L g1585 ( 
.A1(n_1469),
.A2(n_980),
.B1(n_983),
.B2(n_982),
.Y(n_1585)
);

AND2x6_ASAP7_75t_L g1586 ( 
.A(n_1435),
.B(n_954),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1500),
.Y(n_1587)
);

AND2x4_ASAP7_75t_L g1588 ( 
.A(n_1501),
.B(n_1154),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1475),
.B(n_1022),
.Y(n_1589)
);

CKINVDCx8_ASAP7_75t_R g1590 ( 
.A(n_1399),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1502),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1504),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1505),
.Y(n_1593)
);

HB1xp67_ASAP7_75t_L g1594 ( 
.A(n_1476),
.Y(n_1594)
);

NAND2xp33_ASAP7_75t_SL g1595 ( 
.A(n_1402),
.B(n_986),
.Y(n_1595)
);

AOI22xp5_ASAP7_75t_L g1596 ( 
.A1(n_1478),
.A2(n_988),
.B1(n_989),
.B2(n_987),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1506),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1449),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1479),
.B(n_990),
.Y(n_1599)
);

BUFx2_ASAP7_75t_L g1600 ( 
.A(n_1487),
.Y(n_1600)
);

BUFx6f_ASAP7_75t_L g1601 ( 
.A(n_1473),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1447),
.Y(n_1602)
);

BUFx3_ASAP7_75t_L g1603 ( 
.A(n_1489),
.Y(n_1603)
);

AND2x4_ASAP7_75t_L g1604 ( 
.A(n_1472),
.B(n_1154),
.Y(n_1604)
);

INVx3_ASAP7_75t_L g1605 ( 
.A(n_1490),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1509),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1491),
.B(n_1022),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1488),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1498),
.Y(n_1609)
);

AND2x4_ASAP7_75t_L g1610 ( 
.A(n_1406),
.B(n_1330),
.Y(n_1610)
);

AND2x4_ASAP7_75t_L g1611 ( 
.A(n_1411),
.B(n_1330),
.Y(n_1611)
);

BUFx6f_ASAP7_75t_L g1612 ( 
.A(n_1503),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_1507),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1461),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1437),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1440),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1441),
.B(n_991),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1409),
.B(n_992),
.Y(n_1618)
);

BUFx6f_ASAP7_75t_L g1619 ( 
.A(n_1427),
.Y(n_1619)
);

BUFx6f_ASAP7_75t_L g1620 ( 
.A(n_1429),
.Y(n_1620)
);

BUFx6f_ASAP7_75t_L g1621 ( 
.A(n_1420),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1433),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1439),
.B(n_993),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1468),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1499),
.B(n_1065),
.Y(n_1625)
);

INVx1_ASAP7_75t_SL g1626 ( 
.A(n_1510),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1415),
.Y(n_1627)
);

INVx3_ASAP7_75t_L g1628 ( 
.A(n_1415),
.Y(n_1628)
);

BUFx3_ASAP7_75t_L g1629 ( 
.A(n_1463),
.Y(n_1629)
);

HB1xp67_ASAP7_75t_L g1630 ( 
.A(n_1434),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1463),
.Y(n_1631)
);

AOI22xp5_ASAP7_75t_L g1632 ( 
.A1(n_1471),
.A2(n_997),
.B1(n_1003),
.B2(n_995),
.Y(n_1632)
);

AND2x4_ASAP7_75t_L g1633 ( 
.A(n_1403),
.B(n_1137),
.Y(n_1633)
);

AOI22xp5_ASAP7_75t_SL g1634 ( 
.A1(n_1410),
.A2(n_1116),
.B1(n_1122),
.B2(n_944),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1463),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1403),
.B(n_1006),
.Y(n_1636)
);

HB1xp67_ASAP7_75t_L g1637 ( 
.A(n_1434),
.Y(n_1637)
);

OR2x2_ASAP7_75t_L g1638 ( 
.A(n_1414),
.B(n_1310),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1403),
.B(n_1007),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1463),
.Y(n_1640)
);

BUFx6f_ASAP7_75t_L g1641 ( 
.A(n_1438),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1403),
.B(n_1008),
.Y(n_1642)
);

CKINVDCx5p33_ASAP7_75t_R g1643 ( 
.A(n_1399),
.Y(n_1643)
);

NOR2xp33_ASAP7_75t_L g1644 ( 
.A(n_1403),
.B(n_1011),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1463),
.Y(n_1645)
);

BUFx3_ASAP7_75t_L g1646 ( 
.A(n_1463),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1463),
.Y(n_1647)
);

INVx2_ASAP7_75t_SL g1648 ( 
.A(n_1403),
.Y(n_1648)
);

AND2x2_ASAP7_75t_SL g1649 ( 
.A(n_1434),
.B(n_945),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1463),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1463),
.Y(n_1651)
);

BUFx2_ASAP7_75t_L g1652 ( 
.A(n_1403),
.Y(n_1652)
);

AND2x4_ASAP7_75t_L g1653 ( 
.A(n_1403),
.B(n_1137),
.Y(n_1653)
);

BUFx2_ASAP7_75t_L g1654 ( 
.A(n_1403),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1404),
.B(n_1065),
.Y(n_1655)
);

AND2x4_ASAP7_75t_L g1656 ( 
.A(n_1403),
.B(n_1167),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1415),
.Y(n_1657)
);

HB1xp67_ASAP7_75t_L g1658 ( 
.A(n_1434),
.Y(n_1658)
);

BUFx8_ASAP7_75t_L g1659 ( 
.A(n_1434),
.Y(n_1659)
);

BUFx3_ASAP7_75t_L g1660 ( 
.A(n_1463),
.Y(n_1660)
);

HB1xp67_ASAP7_75t_L g1661 ( 
.A(n_1434),
.Y(n_1661)
);

CKINVDCx8_ASAP7_75t_R g1662 ( 
.A(n_1399),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1415),
.Y(n_1663)
);

OAI21x1_ASAP7_75t_L g1664 ( 
.A1(n_1459),
.A2(n_1001),
.B(n_976),
.Y(n_1664)
);

BUFx8_ASAP7_75t_L g1665 ( 
.A(n_1434),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1403),
.B(n_1013),
.Y(n_1666)
);

INVx3_ASAP7_75t_L g1667 ( 
.A(n_1415),
.Y(n_1667)
);

BUFx6f_ASAP7_75t_L g1668 ( 
.A(n_1438),
.Y(n_1668)
);

CKINVDCx6p67_ASAP7_75t_R g1669 ( 
.A(n_1445),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1463),
.Y(n_1670)
);

CKINVDCx6p67_ASAP7_75t_R g1671 ( 
.A(n_1445),
.Y(n_1671)
);

BUFx2_ASAP7_75t_L g1672 ( 
.A(n_1403),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1415),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1403),
.B(n_1016),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1415),
.Y(n_1675)
);

BUFx6f_ASAP7_75t_L g1676 ( 
.A(n_1438),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1463),
.Y(n_1677)
);

HB1xp67_ASAP7_75t_L g1678 ( 
.A(n_1434),
.Y(n_1678)
);

INVx3_ASAP7_75t_L g1679 ( 
.A(n_1415),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1463),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1463),
.Y(n_1681)
);

AND2x6_ASAP7_75t_L g1682 ( 
.A(n_1425),
.B(n_1201),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_SL g1683 ( 
.A(n_1403),
.B(n_912),
.Y(n_1683)
);

BUFx6f_ASAP7_75t_L g1684 ( 
.A(n_1438),
.Y(n_1684)
);

INVx6_ASAP7_75t_L g1685 ( 
.A(n_1415),
.Y(n_1685)
);

OA21x2_ASAP7_75t_L g1686 ( 
.A1(n_1459),
.A2(n_1077),
.B(n_1001),
.Y(n_1686)
);

BUFx8_ASAP7_75t_L g1687 ( 
.A(n_1434),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1415),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1463),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1404),
.B(n_1119),
.Y(n_1690)
);

INVx4_ASAP7_75t_L g1691 ( 
.A(n_1403),
.Y(n_1691)
);

INVxp67_ASAP7_75t_L g1692 ( 
.A(n_1522),
.Y(n_1692)
);

AND2x4_ASAP7_75t_L g1693 ( 
.A(n_1633),
.B(n_883),
.Y(n_1693)
);

OAI22xp33_ASAP7_75t_L g1694 ( 
.A1(n_1533),
.A2(n_1113),
.B1(n_1263),
.B2(n_1247),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_SL g1695 ( 
.A(n_1565),
.B(n_1077),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1531),
.Y(n_1696)
);

OR2x6_ASAP7_75t_L g1697 ( 
.A(n_1600),
.B(n_1062),
.Y(n_1697)
);

BUFx4f_ASAP7_75t_L g1698 ( 
.A(n_1669),
.Y(n_1698)
);

BUFx3_ASAP7_75t_L g1699 ( 
.A(n_1600),
.Y(n_1699)
);

INVx4_ASAP7_75t_L g1700 ( 
.A(n_1682),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1537),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1664),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1562),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1562),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_SL g1705 ( 
.A(n_1565),
.B(n_1110),
.Y(n_1705)
);

CKINVDCx5p33_ASAP7_75t_R g1706 ( 
.A(n_1659),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_SL g1707 ( 
.A(n_1536),
.B(n_1110),
.Y(n_1707)
);

BUFx4f_ASAP7_75t_L g1708 ( 
.A(n_1671),
.Y(n_1708)
);

CKINVDCx5p33_ASAP7_75t_R g1709 ( 
.A(n_1659),
.Y(n_1709)
);

INVx3_ASAP7_75t_L g1710 ( 
.A(n_1685),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1576),
.Y(n_1711)
);

NOR3xp33_ASAP7_75t_L g1712 ( 
.A(n_1545),
.B(n_1025),
.C(n_904),
.Y(n_1712)
);

OR2x2_ASAP7_75t_L g1713 ( 
.A(n_1520),
.B(n_1058),
.Y(n_1713)
);

AND3x1_ASAP7_75t_L g1714 ( 
.A(n_1625),
.B(n_901),
.C(n_892),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1576),
.Y(n_1715)
);

INVx2_ASAP7_75t_SL g1716 ( 
.A(n_1629),
.Y(n_1716)
);

INVx2_ASAP7_75t_SL g1717 ( 
.A(n_1646),
.Y(n_1717)
);

INVx4_ASAP7_75t_L g1718 ( 
.A(n_1682),
.Y(n_1718)
);

OR2x2_ASAP7_75t_L g1719 ( 
.A(n_1540),
.B(n_1085),
.Y(n_1719)
);

AND2x6_ASAP7_75t_L g1720 ( 
.A(n_1602),
.B(n_1244),
.Y(n_1720)
);

NOR2xp33_ASAP7_75t_L g1721 ( 
.A(n_1598),
.B(n_1021),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1686),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1686),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1582),
.Y(n_1724)
);

CKINVDCx20_ASAP7_75t_R g1725 ( 
.A(n_1687),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_SL g1726 ( 
.A(n_1655),
.B(n_1140),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1584),
.Y(n_1727)
);

INVx1_ASAP7_75t_SL g1728 ( 
.A(n_1652),
.Y(n_1728)
);

INVx4_ASAP7_75t_L g1729 ( 
.A(n_1682),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_SL g1730 ( 
.A(n_1690),
.B(n_1140),
.Y(n_1730)
);

INVx2_ASAP7_75t_SL g1731 ( 
.A(n_1660),
.Y(n_1731)
);

AOI22xp33_ASAP7_75t_L g1732 ( 
.A1(n_1608),
.A2(n_1092),
.B1(n_1098),
.B2(n_1084),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1516),
.Y(n_1733)
);

INVx3_ASAP7_75t_L g1734 ( 
.A(n_1685),
.Y(n_1734)
);

INVx2_ASAP7_75t_SL g1735 ( 
.A(n_1511),
.Y(n_1735)
);

AOI22xp33_ASAP7_75t_L g1736 ( 
.A1(n_1519),
.A2(n_1102),
.B1(n_1121),
.B2(n_1100),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1627),
.Y(n_1737)
);

OAI22x1_ASAP7_75t_L g1738 ( 
.A1(n_1626),
.A2(n_1036),
.B1(n_1043),
.B2(n_1038),
.Y(n_1738)
);

INVx4_ASAP7_75t_L g1739 ( 
.A(n_1546),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1513),
.B(n_1515),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1530),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1532),
.Y(n_1742)
);

OR2x2_ASAP7_75t_L g1743 ( 
.A(n_1549),
.B(n_1179),
.Y(n_1743)
);

INVx2_ASAP7_75t_L g1744 ( 
.A(n_1657),
.Y(n_1744)
);

CKINVDCx5p33_ASAP7_75t_R g1745 ( 
.A(n_1687),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1604),
.B(n_912),
.Y(n_1746)
);

INVx5_ASAP7_75t_L g1747 ( 
.A(n_1628),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1534),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1558),
.Y(n_1749)
);

INVx1_ASAP7_75t_SL g1750 ( 
.A(n_1652),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1579),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1663),
.Y(n_1752)
);

INVx4_ASAP7_75t_SL g1753 ( 
.A(n_1586),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1579),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1588),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1588),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1525),
.Y(n_1757)
);

BUFx6f_ASAP7_75t_L g1758 ( 
.A(n_1571),
.Y(n_1758)
);

NOR2xp33_ASAP7_75t_L g1759 ( 
.A(n_1691),
.B(n_1060),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1556),
.B(n_1278),
.Y(n_1760)
);

BUFx6f_ASAP7_75t_L g1761 ( 
.A(n_1583),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1673),
.Y(n_1762)
);

OR2x6_ASAP7_75t_L g1763 ( 
.A(n_1569),
.B(n_1603),
.Y(n_1763)
);

OR2x6_ASAP7_75t_L g1764 ( 
.A(n_1612),
.B(n_1307),
.Y(n_1764)
);

HB1xp67_ASAP7_75t_L g1765 ( 
.A(n_1630),
.Y(n_1765)
);

AOI22xp33_ASAP7_75t_L g1766 ( 
.A1(n_1529),
.A2(n_1123),
.B1(n_1127),
.B2(n_1124),
.Y(n_1766)
);

NOR3xp33_ASAP7_75t_L g1767 ( 
.A(n_1623),
.B(n_1249),
.C(n_1224),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1675),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1517),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_1563),
.B(n_1278),
.Y(n_1770)
);

INVx2_ASAP7_75t_SL g1771 ( 
.A(n_1654),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1518),
.Y(n_1772)
);

INVx3_ASAP7_75t_L g1773 ( 
.A(n_1667),
.Y(n_1773)
);

OR2x2_ASAP7_75t_L g1774 ( 
.A(n_1638),
.B(n_1328),
.Y(n_1774)
);

OAI22xp5_ASAP7_75t_L g1775 ( 
.A1(n_1523),
.A2(n_1066),
.B1(n_1069),
.B2(n_1061),
.Y(n_1775)
);

NOR2xp33_ASAP7_75t_L g1776 ( 
.A(n_1636),
.B(n_1070),
.Y(n_1776)
);

BUFx2_ASAP7_75t_L g1777 ( 
.A(n_1637),
.Y(n_1777)
);

OAI22xp33_ASAP7_75t_L g1778 ( 
.A1(n_1654),
.A2(n_1332),
.B1(n_1341),
.B2(n_1320),
.Y(n_1778)
);

NOR2xp33_ASAP7_75t_L g1779 ( 
.A(n_1639),
.B(n_1080),
.Y(n_1779)
);

INVx3_ASAP7_75t_L g1780 ( 
.A(n_1679),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1570),
.B(n_949),
.Y(n_1781)
);

NOR2xp33_ASAP7_75t_L g1782 ( 
.A(n_1642),
.B(n_1082),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1541),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1609),
.B(n_949),
.Y(n_1784)
);

CKINVDCx5p33_ASAP7_75t_R g1785 ( 
.A(n_1665),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1547),
.Y(n_1786)
);

NOR2xp33_ASAP7_75t_SL g1787 ( 
.A(n_1554),
.B(n_944),
.Y(n_1787)
);

INVx2_ASAP7_75t_L g1788 ( 
.A(n_1688),
.Y(n_1788)
);

OR2x2_ASAP7_75t_L g1789 ( 
.A(n_1658),
.B(n_1661),
.Y(n_1789)
);

BUFx2_ASAP7_75t_L g1790 ( 
.A(n_1678),
.Y(n_1790)
);

OR2x6_ASAP7_75t_L g1791 ( 
.A(n_1612),
.B(n_1358),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1548),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1572),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1524),
.B(n_949),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1538),
.B(n_949),
.Y(n_1795)
);

INVx2_ASAP7_75t_L g1796 ( 
.A(n_1592),
.Y(n_1796)
);

NOR2xp33_ASAP7_75t_L g1797 ( 
.A(n_1666),
.B(n_1083),
.Y(n_1797)
);

INVx3_ASAP7_75t_L g1798 ( 
.A(n_1552),
.Y(n_1798)
);

INVx3_ASAP7_75t_L g1799 ( 
.A(n_1552),
.Y(n_1799)
);

INVx3_ASAP7_75t_L g1800 ( 
.A(n_1561),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_SL g1801 ( 
.A(n_1599),
.B(n_1633),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1593),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1672),
.B(n_1395),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_SL g1804 ( 
.A(n_1653),
.B(n_1656),
.Y(n_1804)
);

AND3x2_ASAP7_75t_L g1805 ( 
.A(n_1514),
.B(n_1122),
.C(n_1116),
.Y(n_1805)
);

BUFx4f_ASAP7_75t_L g1806 ( 
.A(n_1619),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1539),
.Y(n_1807)
);

NAND2xp33_ASAP7_75t_L g1808 ( 
.A(n_1586),
.B(n_949),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_SL g1809 ( 
.A(n_1653),
.B(n_1151),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1553),
.Y(n_1810)
);

INVx2_ASAP7_75t_L g1811 ( 
.A(n_1555),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1551),
.B(n_1089),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1672),
.B(n_1395),
.Y(n_1813)
);

OAI22xp33_ASAP7_75t_L g1814 ( 
.A1(n_1632),
.A2(n_1222),
.B1(n_1237),
.B2(n_1200),
.Y(n_1814)
);

BUFx4f_ASAP7_75t_L g1815 ( 
.A(n_1619),
.Y(n_1815)
);

INVx2_ASAP7_75t_SL g1816 ( 
.A(n_1656),
.Y(n_1816)
);

INVx2_ASAP7_75t_L g1817 ( 
.A(n_1557),
.Y(n_1817)
);

BUFx2_ASAP7_75t_L g1818 ( 
.A(n_1559),
.Y(n_1818)
);

BUFx2_ASAP7_75t_L g1819 ( 
.A(n_1581),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1566),
.B(n_1090),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_L g1821 ( 
.A(n_1567),
.B(n_1091),
.Y(n_1821)
);

HB1xp67_ASAP7_75t_L g1822 ( 
.A(n_1594),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1573),
.Y(n_1823)
);

INVx2_ASAP7_75t_L g1824 ( 
.A(n_1574),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1577),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1578),
.Y(n_1826)
);

OR2x2_ASAP7_75t_L g1827 ( 
.A(n_1564),
.B(n_1385),
.Y(n_1827)
);

AND2x6_ASAP7_75t_L g1828 ( 
.A(n_1589),
.B(n_1151),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1580),
.Y(n_1829)
);

INVx3_ASAP7_75t_L g1830 ( 
.A(n_1561),
.Y(n_1830)
);

INVx2_ASAP7_75t_L g1831 ( 
.A(n_1587),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1591),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1597),
.Y(n_1833)
);

AOI22xp5_ASAP7_75t_L g1834 ( 
.A1(n_1649),
.A2(n_1103),
.B1(n_1106),
.B2(n_1093),
.Y(n_1834)
);

NOR2xp33_ASAP7_75t_L g1835 ( 
.A(n_1674),
.B(n_1107),
.Y(n_1835)
);

HB1xp67_ASAP7_75t_L g1836 ( 
.A(n_1560),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1607),
.B(n_934),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1610),
.B(n_1108),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1610),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1611),
.Y(n_1840)
);

INVx4_ASAP7_75t_L g1841 ( 
.A(n_1605),
.Y(n_1841)
);

NOR2xp33_ASAP7_75t_L g1842 ( 
.A(n_1644),
.B(n_1114),
.Y(n_1842)
);

NOR2xp33_ASAP7_75t_L g1843 ( 
.A(n_1648),
.B(n_1117),
.Y(n_1843)
);

NAND3xp33_ASAP7_75t_L g1844 ( 
.A(n_1596),
.B(n_1130),
.C(n_1126),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1611),
.B(n_1132),
.Y(n_1845)
);

INVx2_ASAP7_75t_L g1846 ( 
.A(n_1521),
.Y(n_1846)
);

INVx2_ASAP7_75t_SL g1847 ( 
.A(n_1614),
.Y(n_1847)
);

BUFx3_ASAP7_75t_L g1848 ( 
.A(n_1620),
.Y(n_1848)
);

BUFx10_ASAP7_75t_L g1849 ( 
.A(n_1550),
.Y(n_1849)
);

NOR2xp33_ASAP7_75t_L g1850 ( 
.A(n_1512),
.B(n_1133),
.Y(n_1850)
);

INVx2_ASAP7_75t_L g1851 ( 
.A(n_1527),
.Y(n_1851)
);

BUFx2_ASAP7_75t_L g1852 ( 
.A(n_1595),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1526),
.Y(n_1853)
);

AND3x2_ASAP7_75t_L g1854 ( 
.A(n_1622),
.B(n_1222),
.C(n_1200),
.Y(n_1854)
);

BUFx3_ASAP7_75t_L g1855 ( 
.A(n_1620),
.Y(n_1855)
);

INVx2_ASAP7_75t_L g1856 ( 
.A(n_1527),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_SL g1857 ( 
.A(n_1613),
.B(n_1322),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_SL g1858 ( 
.A(n_1617),
.B(n_1618),
.Y(n_1858)
);

AOI22xp33_ASAP7_75t_L g1859 ( 
.A1(n_1631),
.A2(n_1134),
.B1(n_1136),
.B2(n_1129),
.Y(n_1859)
);

INVx2_ASAP7_75t_SL g1860 ( 
.A(n_1635),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1683),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1640),
.Y(n_1862)
);

INVxp67_ASAP7_75t_SL g1863 ( 
.A(n_1645),
.Y(n_1863)
);

AND2x4_ASAP7_75t_L g1864 ( 
.A(n_1535),
.B(n_908),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1647),
.B(n_1650),
.Y(n_1865)
);

NOR2x1p5_ASAP7_75t_L g1866 ( 
.A(n_1643),
.B(n_1141),
.Y(n_1866)
);

OR2x6_ASAP7_75t_L g1867 ( 
.A(n_1621),
.B(n_1237),
.Y(n_1867)
);

INVx2_ASAP7_75t_SL g1868 ( 
.A(n_1651),
.Y(n_1868)
);

INVx4_ASAP7_75t_SL g1869 ( 
.A(n_1615),
.Y(n_1869)
);

BUFx6f_ASAP7_75t_L g1870 ( 
.A(n_1590),
.Y(n_1870)
);

INVxp67_ASAP7_75t_L g1871 ( 
.A(n_1621),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1670),
.Y(n_1872)
);

INVx2_ASAP7_75t_L g1873 ( 
.A(n_1528),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1677),
.Y(n_1874)
);

INVx2_ASAP7_75t_L g1875 ( 
.A(n_1528),
.Y(n_1875)
);

NOR2xp33_ASAP7_75t_L g1876 ( 
.A(n_1680),
.B(n_1142),
.Y(n_1876)
);

NOR2xp33_ASAP7_75t_L g1877 ( 
.A(n_1681),
.B(n_1145),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1689),
.Y(n_1878)
);

AND2x2_ASAP7_75t_L g1879 ( 
.A(n_1616),
.B(n_934),
.Y(n_1879)
);

NOR2xp33_ASAP7_75t_SL g1880 ( 
.A(n_1662),
.B(n_1388),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_SL g1881 ( 
.A(n_1544),
.B(n_1322),
.Y(n_1881)
);

INVx2_ASAP7_75t_L g1882 ( 
.A(n_1542),
.Y(n_1882)
);

INVx8_ASAP7_75t_L g1883 ( 
.A(n_1543),
.Y(n_1883)
);

AND2x6_ASAP7_75t_L g1884 ( 
.A(n_1624),
.B(n_1393),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_SL g1885 ( 
.A(n_1542),
.B(n_1326),
.Y(n_1885)
);

OR2x6_ASAP7_75t_L g1886 ( 
.A(n_1634),
.B(n_945),
.Y(n_1886)
);

INVx3_ASAP7_75t_L g1887 ( 
.A(n_1568),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1568),
.Y(n_1888)
);

AND2x6_ASAP7_75t_L g1889 ( 
.A(n_1684),
.B(n_1393),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1575),
.Y(n_1890)
);

INVx2_ASAP7_75t_L g1891 ( 
.A(n_1575),
.Y(n_1891)
);

BUFx4f_ASAP7_75t_L g1892 ( 
.A(n_1601),
.Y(n_1892)
);

NAND2xp33_ASAP7_75t_L g1893 ( 
.A(n_1601),
.B(n_1219),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1641),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1668),
.B(n_1392),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_L g1896 ( 
.A(n_1676),
.B(n_1148),
.Y(n_1896)
);

AOI22xp33_ASAP7_75t_L g1897 ( 
.A1(n_1676),
.A2(n_1143),
.B1(n_1144),
.B2(n_1138),
.Y(n_1897)
);

INVx4_ASAP7_75t_L g1898 ( 
.A(n_1684),
.Y(n_1898)
);

NOR2xp33_ASAP7_75t_L g1899 ( 
.A(n_1598),
.B(n_1150),
.Y(n_1899)
);

INVx2_ASAP7_75t_SL g1900 ( 
.A(n_1522),
.Y(n_1900)
);

BUFx6f_ASAP7_75t_L g1901 ( 
.A(n_1562),
.Y(n_1901)
);

NOR2xp33_ASAP7_75t_L g1902 ( 
.A(n_1598),
.B(n_1164),
.Y(n_1902)
);

INVx4_ASAP7_75t_L g1903 ( 
.A(n_1682),
.Y(n_1903)
);

NOR2xp33_ASAP7_75t_L g1904 ( 
.A(n_1598),
.B(n_1165),
.Y(n_1904)
);

NAND2xp33_ASAP7_75t_L g1905 ( 
.A(n_1682),
.B(n_1219),
.Y(n_1905)
);

BUFx6f_ASAP7_75t_L g1906 ( 
.A(n_1562),
.Y(n_1906)
);

INVx2_ASAP7_75t_SL g1907 ( 
.A(n_1522),
.Y(n_1907)
);

BUFx6f_ASAP7_75t_L g1908 ( 
.A(n_1562),
.Y(n_1908)
);

INVx2_ASAP7_75t_L g1909 ( 
.A(n_1664),
.Y(n_1909)
);

INVx2_ASAP7_75t_L g1910 ( 
.A(n_1664),
.Y(n_1910)
);

INVx3_ASAP7_75t_L g1911 ( 
.A(n_1685),
.Y(n_1911)
);

BUFx6f_ASAP7_75t_L g1912 ( 
.A(n_1562),
.Y(n_1912)
);

INVx4_ASAP7_75t_L g1913 ( 
.A(n_1682),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1531),
.Y(n_1914)
);

OR2x2_ASAP7_75t_L g1915 ( 
.A(n_1520),
.B(n_1171),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_SL g1916 ( 
.A(n_1565),
.B(n_1326),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_SL g1917 ( 
.A(n_1565),
.B(n_1349),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1531),
.Y(n_1918)
);

OR2x6_ASAP7_75t_L g1919 ( 
.A(n_1600),
.B(n_1010),
.Y(n_1919)
);

INVx2_ASAP7_75t_L g1920 ( 
.A(n_1664),
.Y(n_1920)
);

INVx2_ASAP7_75t_L g1921 ( 
.A(n_1664),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1606),
.B(n_1177),
.Y(n_1922)
);

OR2x6_ASAP7_75t_L g1923 ( 
.A(n_1600),
.B(n_1010),
.Y(n_1923)
);

AOI22xp33_ASAP7_75t_L g1924 ( 
.A1(n_1606),
.A2(n_1168),
.B1(n_1178),
.B2(n_1149),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_SL g1925 ( 
.A(n_1565),
.B(n_1349),
.Y(n_1925)
);

INVx3_ASAP7_75t_L g1926 ( 
.A(n_1685),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1531),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1531),
.Y(n_1928)
);

BUFx6f_ASAP7_75t_L g1929 ( 
.A(n_1562),
.Y(n_1929)
);

AND2x2_ASAP7_75t_L g1930 ( 
.A(n_1533),
.B(n_984),
.Y(n_1930)
);

AND2x2_ASAP7_75t_L g1931 ( 
.A(n_1533),
.B(n_984),
.Y(n_1931)
);

NOR2xp33_ASAP7_75t_L g1932 ( 
.A(n_1598),
.B(n_1183),
.Y(n_1932)
);

AOI22xp33_ASAP7_75t_L g1933 ( 
.A1(n_1606),
.A2(n_1181),
.B1(n_1182),
.B2(n_1180),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1531),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_SL g1935 ( 
.A(n_1565),
.B(n_1378),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1531),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1531),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1606),
.B(n_1379),
.Y(n_1938)
);

NAND3xp33_ASAP7_75t_L g1939 ( 
.A(n_1585),
.B(n_1188),
.C(n_1185),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_SL g1940 ( 
.A(n_1900),
.B(n_1197),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_L g1941 ( 
.A(n_1743),
.B(n_1189),
.Y(n_1941)
);

HB1xp67_ASAP7_75t_L g1942 ( 
.A(n_1907),
.Y(n_1942)
);

INVxp33_ASAP7_75t_L g1943 ( 
.A(n_1765),
.Y(n_1943)
);

NOR2xp33_ASAP7_75t_L g1944 ( 
.A(n_1692),
.B(n_1196),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_SL g1945 ( 
.A(n_1718),
.B(n_1729),
.Y(n_1945)
);

OR2x6_ASAP7_75t_L g1946 ( 
.A(n_1697),
.B(n_1028),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1769),
.Y(n_1947)
);

NOR2xp33_ASAP7_75t_L g1948 ( 
.A(n_1837),
.B(n_1203),
.Y(n_1948)
);

BUFx12f_ASAP7_75t_L g1949 ( 
.A(n_1785),
.Y(n_1949)
);

NAND2xp5_ASAP7_75t_L g1950 ( 
.A(n_1922),
.B(n_1207),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_L g1951 ( 
.A(n_1938),
.B(n_1209),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1772),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1757),
.Y(n_1953)
);

NAND2xp33_ASAP7_75t_L g1954 ( 
.A(n_1720),
.B(n_1238),
.Y(n_1954)
);

INVx2_ASAP7_75t_SL g1955 ( 
.A(n_1699),
.Y(n_1955)
);

BUFx8_ASAP7_75t_L g1956 ( 
.A(n_1870),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1751),
.Y(n_1957)
);

INVxp33_ASAP7_75t_L g1958 ( 
.A(n_1713),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_SL g1959 ( 
.A(n_1718),
.B(n_1286),
.Y(n_1959)
);

INVx2_ASAP7_75t_L g1960 ( 
.A(n_1703),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1754),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1755),
.Y(n_1962)
);

INVx2_ASAP7_75t_L g1963 ( 
.A(n_1704),
.Y(n_1963)
);

NAND3xp33_ASAP7_75t_L g1964 ( 
.A(n_1843),
.B(n_1212),
.C(n_1210),
.Y(n_1964)
);

AOI22xp33_ASAP7_75t_L g1965 ( 
.A1(n_1853),
.A2(n_1228),
.B1(n_1241),
.B2(n_1226),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1721),
.B(n_1245),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1756),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1899),
.B(n_1246),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1902),
.B(n_1248),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_SL g1970 ( 
.A(n_1729),
.B(n_1295),
.Y(n_1970)
);

AOI22xp33_ASAP7_75t_L g1971 ( 
.A1(n_1904),
.A2(n_1257),
.B1(n_1260),
.B2(n_1256),
.Y(n_1971)
);

AND2x2_ASAP7_75t_L g1972 ( 
.A(n_1728),
.B(n_893),
.Y(n_1972)
);

AND2x4_ASAP7_75t_L g1973 ( 
.A(n_1739),
.B(n_923),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_SL g1974 ( 
.A(n_1903),
.B(n_1700),
.Y(n_1974)
);

INVx2_ASAP7_75t_SL g1975 ( 
.A(n_1777),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1807),
.Y(n_1976)
);

NAND2xp5_ASAP7_75t_L g1977 ( 
.A(n_1932),
.B(n_1261),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_L g1978 ( 
.A(n_1776),
.B(n_1262),
.Y(n_1978)
);

OR2x6_ASAP7_75t_L g1979 ( 
.A(n_1697),
.B(n_1883),
.Y(n_1979)
);

NOR2xp33_ASAP7_75t_L g1980 ( 
.A(n_1774),
.B(n_1264),
.Y(n_1980)
);

BUFx2_ASAP7_75t_L g1981 ( 
.A(n_1777),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1779),
.B(n_1269),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_L g1983 ( 
.A(n_1782),
.B(n_1273),
.Y(n_1983)
);

INVx2_ASAP7_75t_L g1984 ( 
.A(n_1711),
.Y(n_1984)
);

INVx2_ASAP7_75t_L g1985 ( 
.A(n_1715),
.Y(n_1985)
);

NOR2xp33_ASAP7_75t_L g1986 ( 
.A(n_1760),
.B(n_1275),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_SL g1987 ( 
.A(n_1903),
.B(n_1280),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1810),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_L g1989 ( 
.A(n_1797),
.B(n_1282),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_L g1990 ( 
.A(n_1835),
.B(n_1283),
.Y(n_1990)
);

NOR2xp33_ASAP7_75t_SL g1991 ( 
.A(n_1698),
.B(n_896),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_L g1992 ( 
.A(n_1924),
.B(n_1289),
.Y(n_1992)
);

BUFx12f_ASAP7_75t_SL g1993 ( 
.A(n_1764),
.Y(n_1993)
);

INVx2_ASAP7_75t_L g1994 ( 
.A(n_1901),
.Y(n_1994)
);

NOR2xp33_ASAP7_75t_L g1995 ( 
.A(n_1770),
.B(n_1291),
.Y(n_1995)
);

NOR2xp33_ASAP7_75t_L g1996 ( 
.A(n_1804),
.B(n_1915),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1823),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1825),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_SL g1999 ( 
.A(n_1913),
.B(n_1771),
.Y(n_1999)
);

AOI22xp5_ASAP7_75t_L g2000 ( 
.A1(n_1864),
.A2(n_1296),
.B1(n_1297),
.B2(n_1292),
.Y(n_2000)
);

INVx2_ASAP7_75t_L g2001 ( 
.A(n_1906),
.Y(n_2001)
);

AND2x2_ASAP7_75t_L g2002 ( 
.A(n_1750),
.B(n_924),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_L g2003 ( 
.A(n_1933),
.B(n_1298),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1826),
.Y(n_2004)
);

INVx3_ASAP7_75t_L g2005 ( 
.A(n_1739),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1832),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_L g2007 ( 
.A(n_1842),
.B(n_1300),
.Y(n_2007)
);

BUFx6f_ASAP7_75t_L g2008 ( 
.A(n_1906),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1833),
.Y(n_2009)
);

OAI221xp5_ASAP7_75t_L g2010 ( 
.A1(n_1827),
.A2(n_1315),
.B1(n_1318),
.B2(n_1313),
.C(n_1304),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1741),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_L g2012 ( 
.A(n_1812),
.B(n_1319),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_SL g2013 ( 
.A(n_1841),
.B(n_1356),
.Y(n_2013)
);

O2A1O1Ixp33_ASAP7_75t_L g2014 ( 
.A1(n_1707),
.A2(n_1193),
.B(n_1194),
.C(n_1184),
.Y(n_2014)
);

NOR2xp33_ASAP7_75t_L g2015 ( 
.A(n_1930),
.B(n_1323),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_L g2016 ( 
.A(n_1742),
.B(n_1334),
.Y(n_2016)
);

OR2x2_ASAP7_75t_L g2017 ( 
.A(n_1789),
.B(n_1335),
.Y(n_2017)
);

NOR2xp33_ASAP7_75t_L g2018 ( 
.A(n_1931),
.B(n_1347),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1748),
.Y(n_2019)
);

AOI22xp33_ASAP7_75t_L g2020 ( 
.A1(n_1767),
.A2(n_1357),
.B1(n_1361),
.B2(n_1353),
.Y(n_2020)
);

AOI22xp5_ASAP7_75t_L g2021 ( 
.A1(n_1864),
.A2(n_1364),
.B1(n_1366),
.B2(n_1363),
.Y(n_2021)
);

NOR2xp33_ASAP7_75t_L g2022 ( 
.A(n_1803),
.B(n_1367),
.Y(n_2022)
);

OR2x6_ASAP7_75t_L g2023 ( 
.A(n_1883),
.B(n_1028),
.Y(n_2023)
);

INVx2_ASAP7_75t_L g2024 ( 
.A(n_1908),
.Y(n_2024)
);

NAND2xp5_ASAP7_75t_SL g2025 ( 
.A(n_1790),
.B(n_1368),
.Y(n_2025)
);

INVx3_ASAP7_75t_L g2026 ( 
.A(n_1908),
.Y(n_2026)
);

INVx2_ASAP7_75t_SL g2027 ( 
.A(n_1790),
.Y(n_2027)
);

NOR2xp33_ASAP7_75t_L g2028 ( 
.A(n_1813),
.B(n_1371),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_L g2029 ( 
.A(n_1775),
.B(n_1391),
.Y(n_2029)
);

AOI22xp33_ASAP7_75t_L g2030 ( 
.A1(n_1839),
.A2(n_1208),
.B1(n_1211),
.B2(n_1195),
.Y(n_2030)
);

OR2x2_ASAP7_75t_L g2031 ( 
.A(n_1719),
.B(n_889),
.Y(n_2031)
);

AND2x4_ASAP7_75t_L g2032 ( 
.A(n_1869),
.B(n_950),
.Y(n_2032)
);

INVx2_ASAP7_75t_SL g2033 ( 
.A(n_1818),
.Y(n_2033)
);

NAND2xp33_ASAP7_75t_L g2034 ( 
.A(n_1720),
.B(n_1219),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_L g2035 ( 
.A(n_1820),
.B(n_1380),
.Y(n_2035)
);

NAND2xp33_ASAP7_75t_L g2036 ( 
.A(n_1720),
.B(n_1219),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_L g2037 ( 
.A(n_1821),
.B(n_1381),
.Y(n_2037)
);

NOR2xp33_ASAP7_75t_L g2038 ( 
.A(n_1801),
.B(n_1004),
.Y(n_2038)
);

NAND2xp5_ASAP7_75t_SL g2039 ( 
.A(n_1818),
.B(n_881),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_L g2040 ( 
.A(n_1811),
.B(n_1214),
.Y(n_2040)
);

NAND2xp5_ASAP7_75t_L g2041 ( 
.A(n_1817),
.B(n_1221),
.Y(n_2041)
);

NOR2xp33_ASAP7_75t_L g2042 ( 
.A(n_1860),
.B(n_1045),
.Y(n_2042)
);

NAND2xp5_ASAP7_75t_L g2043 ( 
.A(n_1824),
.B(n_1223),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_SL g2044 ( 
.A(n_1819),
.B(n_894),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_L g2045 ( 
.A(n_1829),
.B(n_1225),
.Y(n_2045)
);

AND2x2_ASAP7_75t_L g2046 ( 
.A(n_1819),
.B(n_1072),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_L g2047 ( 
.A(n_1831),
.B(n_1233),
.Y(n_2047)
);

INVx2_ASAP7_75t_L g2048 ( 
.A(n_1912),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1696),
.Y(n_2049)
);

INVx2_ASAP7_75t_SL g2050 ( 
.A(n_1758),
.Y(n_2050)
);

AOI22xp33_ASAP7_75t_L g2051 ( 
.A1(n_1840),
.A2(n_1235),
.B1(n_1251),
.B2(n_1234),
.Y(n_2051)
);

CKINVDCx5p33_ASAP7_75t_R g2052 ( 
.A(n_1706),
.Y(n_2052)
);

NOR2xp33_ASAP7_75t_L g2053 ( 
.A(n_1868),
.B(n_1287),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_1701),
.Y(n_2054)
);

AOI22xp5_ASAP7_75t_L g2055 ( 
.A1(n_1863),
.A2(n_907),
.B1(n_910),
.B2(n_903),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1914),
.Y(n_2056)
);

NAND2xp5_ASAP7_75t_SL g2057 ( 
.A(n_1847),
.B(n_1759),
.Y(n_2057)
);

BUFx6f_ASAP7_75t_SL g2058 ( 
.A(n_1870),
.Y(n_2058)
);

AND2x2_ASAP7_75t_L g2059 ( 
.A(n_1822),
.B(n_1299),
.Y(n_2059)
);

NAND2xp5_ASAP7_75t_L g2060 ( 
.A(n_1732),
.B(n_1918),
.Y(n_2060)
);

INVx2_ASAP7_75t_L g2061 ( 
.A(n_1929),
.Y(n_2061)
);

AOI21xp5_ASAP7_75t_L g2062 ( 
.A1(n_1702),
.A2(n_1378),
.B(n_1266),
.Y(n_2062)
);

INVxp67_ASAP7_75t_L g2063 ( 
.A(n_1787),
.Y(n_2063)
);

INVx2_ASAP7_75t_L g2064 ( 
.A(n_1929),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_1927),
.Y(n_2065)
);

AOI22xp33_ASAP7_75t_L g2066 ( 
.A1(n_1862),
.A2(n_1267),
.B1(n_1271),
.B2(n_1255),
.Y(n_2066)
);

CKINVDCx5p33_ASAP7_75t_R g2067 ( 
.A(n_1709),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_1928),
.B(n_1934),
.Y(n_2068)
);

NOR2xp33_ASAP7_75t_L g2069 ( 
.A(n_1816),
.B(n_1339),
.Y(n_2069)
);

INVx2_ASAP7_75t_SL g2070 ( 
.A(n_1758),
.Y(n_2070)
);

NAND2xp5_ASAP7_75t_L g2071 ( 
.A(n_1936),
.B(n_1290),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_1937),
.Y(n_2072)
);

AOI22xp5_ASAP7_75t_L g2073 ( 
.A1(n_1714),
.A2(n_1850),
.B1(n_1877),
.B2(n_1876),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1746),
.Y(n_2074)
);

NAND2xp5_ASAP7_75t_SL g2075 ( 
.A(n_1753),
.B(n_920),
.Y(n_2075)
);

INVx2_ASAP7_75t_L g2076 ( 
.A(n_1722),
.Y(n_2076)
);

INVx3_ASAP7_75t_L g2077 ( 
.A(n_1792),
.Y(n_2077)
);

NOR2xp33_ASAP7_75t_L g2078 ( 
.A(n_1858),
.B(n_1726),
.Y(n_2078)
);

NAND2xp33_ASAP7_75t_L g2079 ( 
.A(n_1723),
.B(n_937),
.Y(n_2079)
);

INVx2_ASAP7_75t_L g2080 ( 
.A(n_1796),
.Y(n_2080)
);

OR2x2_ASAP7_75t_L g2081 ( 
.A(n_1778),
.B(n_929),
.Y(n_2081)
);

NAND2xp5_ASAP7_75t_L g2082 ( 
.A(n_1740),
.B(n_1301),
.Y(n_2082)
);

O2A1O1Ixp33_ASAP7_75t_L g2083 ( 
.A1(n_1730),
.A2(n_1308),
.B(n_1311),
.C(n_1305),
.Y(n_2083)
);

NAND2xp5_ASAP7_75t_L g2084 ( 
.A(n_1838),
.B(n_1845),
.Y(n_2084)
);

OAI22xp5_ASAP7_75t_L g2085 ( 
.A1(n_1872),
.A2(n_1874),
.B1(n_1878),
.B2(n_1859),
.Y(n_2085)
);

NAND2xp5_ASAP7_75t_SL g2086 ( 
.A(n_1761),
.B(n_938),
.Y(n_2086)
);

NAND2xp5_ASAP7_75t_L g2087 ( 
.A(n_1783),
.B(n_1325),
.Y(n_2087)
);

OR2x6_ASAP7_75t_L g2088 ( 
.A(n_1764),
.B(n_1033),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_SL g2089 ( 
.A(n_1716),
.B(n_939),
.Y(n_2089)
);

NAND2xp5_ASAP7_75t_L g2090 ( 
.A(n_1786),
.B(n_1376),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_1793),
.Y(n_2091)
);

NAND2xp5_ASAP7_75t_L g2092 ( 
.A(n_1802),
.B(n_1337),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_1695),
.Y(n_2093)
);

NAND2xp5_ASAP7_75t_L g2094 ( 
.A(n_1736),
.B(n_1343),
.Y(n_2094)
);

NAND2xp5_ASAP7_75t_L g2095 ( 
.A(n_1766),
.B(n_1351),
.Y(n_2095)
);

NAND2xp5_ASAP7_75t_L g2096 ( 
.A(n_1834),
.B(n_1354),
.Y(n_2096)
);

NAND2xp5_ASAP7_75t_SL g2097 ( 
.A(n_1717),
.B(n_940),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_SL g2098 ( 
.A(n_1731),
.B(n_941),
.Y(n_2098)
);

INVx2_ASAP7_75t_SL g2099 ( 
.A(n_1919),
.Y(n_2099)
);

A2O1A1Ixp33_ASAP7_75t_L g2100 ( 
.A1(n_1784),
.A2(n_1781),
.B(n_1795),
.C(n_1794),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_1705),
.Y(n_2101)
);

NOR2xp33_ASAP7_75t_L g2102 ( 
.A(n_1879),
.B(n_960),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_1916),
.Y(n_2103)
);

BUFx3_ASAP7_75t_L g2104 ( 
.A(n_1725),
.Y(n_2104)
);

INVx8_ASAP7_75t_L g2105 ( 
.A(n_1919),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_L g2106 ( 
.A(n_1693),
.B(n_1355),
.Y(n_2106)
);

NOR2x1p5_ASAP7_75t_L g2107 ( 
.A(n_1745),
.B(n_1387),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_1917),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_L g2109 ( 
.A(n_1693),
.B(n_1359),
.Y(n_2109)
);

INVx3_ASAP7_75t_L g2110 ( 
.A(n_1733),
.Y(n_2110)
);

INVx2_ASAP7_75t_SL g2111 ( 
.A(n_1923),
.Y(n_2111)
);

INVx2_ASAP7_75t_SL g2112 ( 
.A(n_1923),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_L g2113 ( 
.A(n_1865),
.B(n_1369),
.Y(n_2113)
);

INVx2_ASAP7_75t_L g2114 ( 
.A(n_1737),
.Y(n_2114)
);

NAND2xp5_ASAP7_75t_SL g2115 ( 
.A(n_1735),
.B(n_955),
.Y(n_2115)
);

INVx2_ASAP7_75t_L g2116 ( 
.A(n_1744),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_1925),
.Y(n_2117)
);

INVx2_ASAP7_75t_SL g2118 ( 
.A(n_1806),
.Y(n_2118)
);

NOR2xp67_ASAP7_75t_L g2119 ( 
.A(n_1836),
.B(n_3),
.Y(n_2119)
);

AND2x2_ASAP7_75t_L g2120 ( 
.A(n_1763),
.B(n_1204),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_1935),
.Y(n_2121)
);

BUFx6f_ASAP7_75t_L g2122 ( 
.A(n_1892),
.Y(n_2122)
);

AO221x1_ASAP7_75t_L g2123 ( 
.A1(n_1694),
.A2(n_1099),
.B1(n_1155),
.B2(n_1078),
.C(n_1073),
.Y(n_2123)
);

OAI221xp5_ASAP7_75t_L g2124 ( 
.A1(n_1844),
.A2(n_957),
.B1(n_1158),
.B2(n_1075),
.C(n_974),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_1798),
.Y(n_2125)
);

INVx2_ASAP7_75t_L g2126 ( 
.A(n_1752),
.Y(n_2126)
);

INVxp33_ASAP7_75t_L g2127 ( 
.A(n_1880),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_L g2128 ( 
.A(n_1724),
.B(n_966),
.Y(n_2128)
);

INVx2_ASAP7_75t_L g2129 ( 
.A(n_1762),
.Y(n_2129)
);

INVx2_ASAP7_75t_L g2130 ( 
.A(n_1768),
.Y(n_2130)
);

NAND2xp5_ASAP7_75t_L g2131 ( 
.A(n_1727),
.B(n_971),
.Y(n_2131)
);

NAND2xp5_ASAP7_75t_L g2132 ( 
.A(n_1828),
.B(n_979),
.Y(n_2132)
);

INVx2_ASAP7_75t_SL g2133 ( 
.A(n_1815),
.Y(n_2133)
);

A2O1A1Ixp33_ASAP7_75t_L g2134 ( 
.A1(n_1749),
.A2(n_953),
.B(n_964),
.C(n_959),
.Y(n_2134)
);

NOR3xp33_ASAP7_75t_L g2135 ( 
.A(n_1814),
.B(n_1712),
.C(n_1939),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_L g2136 ( 
.A(n_1809),
.B(n_1012),
.Y(n_2136)
);

NAND2xp5_ASAP7_75t_L g2137 ( 
.A(n_1799),
.B(n_1015),
.Y(n_2137)
);

AND2x4_ASAP7_75t_L g2138 ( 
.A(n_1869),
.B(n_975),
.Y(n_2138)
);

AOI22xp5_ASAP7_75t_L g2139 ( 
.A1(n_1884),
.A2(n_1032),
.B1(n_1035),
.B2(n_1031),
.Y(n_2139)
);

NAND2xp5_ASAP7_75t_L g2140 ( 
.A(n_1800),
.B(n_1037),
.Y(n_2140)
);

AND2x2_ASAP7_75t_L g2141 ( 
.A(n_1763),
.B(n_1204),
.Y(n_2141)
);

NAND2xp33_ASAP7_75t_L g2142 ( 
.A(n_1889),
.B(n_1044),
.Y(n_2142)
);

NAND2xp5_ASAP7_75t_L g2143 ( 
.A(n_1830),
.B(n_1049),
.Y(n_2143)
);

NOR3xp33_ASAP7_75t_L g2144 ( 
.A(n_1871),
.B(n_1348),
.C(n_1253),
.Y(n_2144)
);

NAND2xp5_ASAP7_75t_SL g2145 ( 
.A(n_1852),
.B(n_1050),
.Y(n_2145)
);

INVx2_ASAP7_75t_L g2146 ( 
.A(n_1788),
.Y(n_2146)
);

NAND2xp5_ASAP7_75t_L g2147 ( 
.A(n_1857),
.B(n_1055),
.Y(n_2147)
);

OAI22xp5_ASAP7_75t_L g2148 ( 
.A1(n_1861),
.A2(n_1002),
.B1(n_1005),
.B2(n_1000),
.Y(n_2148)
);

INVx4_ASAP7_75t_L g2149 ( 
.A(n_1708),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_1895),
.Y(n_2150)
);

NAND2x1_ASAP7_75t_L g2151 ( 
.A(n_1889),
.B(n_1073),
.Y(n_2151)
);

O2A1O1Ixp33_ASAP7_75t_L g2152 ( 
.A1(n_1905),
.A2(n_1051),
.B(n_1056),
.C(n_1054),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_1896),
.Y(n_2153)
);

NAND2xp5_ASAP7_75t_L g2154 ( 
.A(n_1884),
.B(n_1094),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_L g2155 ( 
.A(n_1846),
.B(n_1101),
.Y(n_2155)
);

INVx2_ASAP7_75t_L g2156 ( 
.A(n_1909),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_1773),
.Y(n_2157)
);

NAND2xp5_ASAP7_75t_SL g2158 ( 
.A(n_1849),
.B(n_1104),
.Y(n_2158)
);

OAI22xp5_ASAP7_75t_L g2159 ( 
.A1(n_1897),
.A2(n_1087),
.B1(n_1088),
.B2(n_1076),
.Y(n_2159)
);

NOR2xp67_ASAP7_75t_L g2160 ( 
.A(n_1738),
.B(n_4),
.Y(n_2160)
);

BUFx6f_ASAP7_75t_L g2161 ( 
.A(n_1889),
.Y(n_2161)
);

NOR2xp33_ASAP7_75t_L g2162 ( 
.A(n_1780),
.B(n_1105),
.Y(n_2162)
);

NAND2xp5_ASAP7_75t_SL g2163 ( 
.A(n_1747),
.B(n_1111),
.Y(n_2163)
);

NOR2xp33_ASAP7_75t_L g2164 ( 
.A(n_1747),
.B(n_1128),
.Y(n_2164)
);

NAND2xp33_ASAP7_75t_SL g2165 ( 
.A(n_1866),
.B(n_1881),
.Y(n_2165)
);

NAND2xp5_ASAP7_75t_SL g2166 ( 
.A(n_1747),
.B(n_1848),
.Y(n_2166)
);

OAI22xp33_ASAP7_75t_L g2167 ( 
.A1(n_1886),
.A2(n_1390),
.B1(n_1394),
.B2(n_1386),
.Y(n_2167)
);

INVxp33_ASAP7_75t_L g2168 ( 
.A(n_1855),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_1910),
.Y(n_2169)
);

INVx2_ASAP7_75t_L g2170 ( 
.A(n_1920),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_1921),
.Y(n_2171)
);

NAND2xp5_ASAP7_75t_L g2172 ( 
.A(n_1808),
.B(n_1135),
.Y(n_2172)
);

NAND2xp5_ASAP7_75t_L g2173 ( 
.A(n_1710),
.B(n_1139),
.Y(n_2173)
);

NOR2xp67_ASAP7_75t_L g2174 ( 
.A(n_1734),
.B(n_4),
.Y(n_2174)
);

NAND2xp5_ASAP7_75t_L g2175 ( 
.A(n_1911),
.B(n_1152),
.Y(n_2175)
);

INVx2_ASAP7_75t_SL g2176 ( 
.A(n_1926),
.Y(n_2176)
);

BUFx3_ASAP7_75t_L g2177 ( 
.A(n_1791),
.Y(n_2177)
);

NAND2xp5_ASAP7_75t_L g2178 ( 
.A(n_1898),
.B(n_1156),
.Y(n_2178)
);

NAND2xp5_ASAP7_75t_SL g2179 ( 
.A(n_1898),
.B(n_1159),
.Y(n_2179)
);

NAND2xp5_ASAP7_75t_SL g2180 ( 
.A(n_1885),
.B(n_1162),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_1886),
.Y(n_2181)
);

INVx4_ASAP7_75t_L g2182 ( 
.A(n_1791),
.Y(n_2182)
);

INVx2_ASAP7_75t_L g2183 ( 
.A(n_1887),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_1893),
.Y(n_2184)
);

NAND2xp5_ASAP7_75t_L g2185 ( 
.A(n_1805),
.B(n_1166),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_L g2186 ( 
.A(n_1854),
.B(n_1170),
.Y(n_2186)
);

NAND2xp5_ASAP7_75t_L g2187 ( 
.A(n_1867),
.B(n_1172),
.Y(n_2187)
);

NOR2xp67_ASAP7_75t_L g2188 ( 
.A(n_1890),
.B(n_5),
.Y(n_2188)
);

NAND2xp33_ASAP7_75t_L g2189 ( 
.A(n_1894),
.B(n_1174),
.Y(n_2189)
);

OAI22xp5_ASAP7_75t_L g2190 ( 
.A1(n_1851),
.A2(n_1096),
.B1(n_1109),
.B2(n_1097),
.Y(n_2190)
);

NAND2xp5_ASAP7_75t_L g2191 ( 
.A(n_1856),
.B(n_1175),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_1873),
.Y(n_2192)
);

BUFx3_ASAP7_75t_L g2193 ( 
.A(n_1875),
.Y(n_2193)
);

BUFx3_ASAP7_75t_L g2194 ( 
.A(n_1882),
.Y(n_2194)
);

A2O1A1Ixp33_ASAP7_75t_L g2195 ( 
.A1(n_1888),
.A2(n_1131),
.B(n_1160),
.C(n_1120),
.Y(n_2195)
);

AND2x4_ASAP7_75t_L g2196 ( 
.A(n_1891),
.B(n_1216),
.Y(n_2196)
);

BUFx6f_ASAP7_75t_L g2197 ( 
.A(n_1901),
.Y(n_2197)
);

O2A1O1Ixp5_ASAP7_75t_L g2198 ( 
.A1(n_1881),
.A2(n_1063),
.B(n_1068),
.C(n_1033),
.Y(n_2198)
);

INVx2_ASAP7_75t_L g2199 ( 
.A(n_1703),
.Y(n_2199)
);

NAND2xp5_ASAP7_75t_L g2200 ( 
.A(n_1743),
.B(n_1176),
.Y(n_2200)
);

AND2x2_ASAP7_75t_L g2201 ( 
.A(n_1900),
.B(n_1242),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_1769),
.Y(n_2202)
);

INVx2_ASAP7_75t_L g2203 ( 
.A(n_1703),
.Y(n_2203)
);

INVxp67_ASAP7_75t_L g2204 ( 
.A(n_1900),
.Y(n_2204)
);

INVx2_ASAP7_75t_SL g2205 ( 
.A(n_1699),
.Y(n_2205)
);

NAND2xp5_ASAP7_75t_SL g2206 ( 
.A(n_1900),
.B(n_1187),
.Y(n_2206)
);

NAND2xp5_ASAP7_75t_SL g2207 ( 
.A(n_1900),
.B(n_1192),
.Y(n_2207)
);

BUFx3_ASAP7_75t_L g2208 ( 
.A(n_1725),
.Y(n_2208)
);

NAND2xp33_ASAP7_75t_R g2209 ( 
.A(n_1706),
.B(n_1205),
.Y(n_2209)
);

NAND2xp33_ASAP7_75t_L g2210 ( 
.A(n_1720),
.B(n_1206),
.Y(n_2210)
);

NAND2xp5_ASAP7_75t_SL g2211 ( 
.A(n_1900),
.B(n_1213),
.Y(n_2211)
);

NOR2xp33_ASAP7_75t_L g2212 ( 
.A(n_1692),
.B(n_1215),
.Y(n_2212)
);

AND2x2_ASAP7_75t_L g2213 ( 
.A(n_1900),
.B(n_1352),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_1769),
.Y(n_2214)
);

AND2x2_ASAP7_75t_L g2215 ( 
.A(n_1900),
.B(n_1352),
.Y(n_2215)
);

NAND2xp5_ASAP7_75t_L g2216 ( 
.A(n_1743),
.B(n_1217),
.Y(n_2216)
);

NAND2xp5_ASAP7_75t_L g2217 ( 
.A(n_1743),
.B(n_1227),
.Y(n_2217)
);

NAND3xp33_ASAP7_75t_L g2218 ( 
.A(n_1843),
.B(n_1230),
.C(n_1229),
.Y(n_2218)
);

INVx3_ASAP7_75t_L g2219 ( 
.A(n_1718),
.Y(n_2219)
);

NAND2xp5_ASAP7_75t_L g2220 ( 
.A(n_1743),
.B(n_1231),
.Y(n_2220)
);

BUFx8_ASAP7_75t_L g2221 ( 
.A(n_1870),
.Y(n_2221)
);

OAI21xp33_ASAP7_75t_L g2222 ( 
.A1(n_1743),
.A2(n_1372),
.B(n_1360),
.Y(n_2222)
);

NOR2xp33_ASAP7_75t_L g2223 ( 
.A(n_1692),
.B(n_1232),
.Y(n_2223)
);

NAND2xp5_ASAP7_75t_SL g2224 ( 
.A(n_1900),
.B(n_1236),
.Y(n_2224)
);

NAND2xp33_ASAP7_75t_L g2225 ( 
.A(n_1720),
.B(n_1240),
.Y(n_2225)
);

NAND2xp5_ASAP7_75t_SL g2226 ( 
.A(n_1900),
.B(n_1250),
.Y(n_2226)
);

NAND2xp33_ASAP7_75t_L g2227 ( 
.A(n_1720),
.B(n_1265),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_1769),
.Y(n_2228)
);

OAI22xp5_ASAP7_75t_L g2229 ( 
.A1(n_1692),
.A2(n_1243),
.B1(n_1254),
.B2(n_1218),
.Y(n_2229)
);

NAND2xp5_ASAP7_75t_SL g2230 ( 
.A(n_1900),
.B(n_1270),
.Y(n_2230)
);

INVx3_ASAP7_75t_L g2231 ( 
.A(n_1718),
.Y(n_2231)
);

NOR2xp33_ASAP7_75t_L g2232 ( 
.A(n_1692),
.B(n_1277),
.Y(n_2232)
);

NAND2xp5_ASAP7_75t_SL g2233 ( 
.A(n_1900),
.B(n_1279),
.Y(n_2233)
);

NAND2xp5_ASAP7_75t_L g2234 ( 
.A(n_1743),
.B(n_1281),
.Y(n_2234)
);

NAND2xp5_ASAP7_75t_SL g2235 ( 
.A(n_1900),
.B(n_1288),
.Y(n_2235)
);

NAND2xp5_ASAP7_75t_L g2236 ( 
.A(n_1743),
.B(n_1294),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_1769),
.Y(n_2237)
);

AOI21xp5_ASAP7_75t_L g2238 ( 
.A1(n_1702),
.A2(n_1268),
.B(n_1258),
.Y(n_2238)
);

INVx5_ASAP7_75t_L g2239 ( 
.A(n_1889),
.Y(n_2239)
);

NAND2xp5_ASAP7_75t_L g2240 ( 
.A(n_1743),
.B(n_1302),
.Y(n_2240)
);

INVx2_ASAP7_75t_L g2241 ( 
.A(n_1703),
.Y(n_2241)
);

AOI22xp33_ASAP7_75t_L g2242 ( 
.A1(n_1853),
.A2(n_1099),
.B1(n_1155),
.B2(n_1078),
.Y(n_2242)
);

BUFx12f_ASAP7_75t_SL g2243 ( 
.A(n_1697),
.Y(n_2243)
);

AND2x2_ASAP7_75t_L g2244 ( 
.A(n_1900),
.B(n_1303),
.Y(n_2244)
);

NAND2xp33_ASAP7_75t_L g2245 ( 
.A(n_1720),
.B(n_1306),
.Y(n_2245)
);

NAND2xp5_ASAP7_75t_L g2246 ( 
.A(n_1743),
.B(n_1312),
.Y(n_2246)
);

NAND2xp5_ASAP7_75t_L g2247 ( 
.A(n_1743),
.B(n_1324),
.Y(n_2247)
);

NAND2xp5_ASAP7_75t_L g2248 ( 
.A(n_1743),
.B(n_1329),
.Y(n_2248)
);

NAND2xp5_ASAP7_75t_SL g2249 ( 
.A(n_1975),
.B(n_1383),
.Y(n_2249)
);

OAI21xp5_ASAP7_75t_L g2250 ( 
.A1(n_2062),
.A2(n_1276),
.B(n_1274),
.Y(n_2250)
);

NAND2xp5_ASAP7_75t_L g2251 ( 
.A(n_2085),
.B(n_1331),
.Y(n_2251)
);

NAND2xp5_ASAP7_75t_SL g2252 ( 
.A(n_2027),
.B(n_1338),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_1952),
.Y(n_2253)
);

NOR2xp33_ASAP7_75t_L g2254 ( 
.A(n_1958),
.B(n_1943),
.Y(n_2254)
);

INVx2_ASAP7_75t_L g2255 ( 
.A(n_2169),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_1953),
.Y(n_2256)
);

AOI22xp5_ASAP7_75t_L g2257 ( 
.A1(n_2135),
.A2(n_1344),
.B1(n_1345),
.B2(n_1342),
.Y(n_2257)
);

CKINVDCx5p33_ASAP7_75t_R g2258 ( 
.A(n_1949),
.Y(n_2258)
);

INVx4_ASAP7_75t_L g2259 ( 
.A(n_2105),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_2202),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_2214),
.Y(n_2261)
);

A2O1A1Ixp33_ASAP7_75t_L g2262 ( 
.A1(n_2152),
.A2(n_1293),
.B(n_1314),
.C(n_1285),
.Y(n_2262)
);

AOI21xp5_ASAP7_75t_L g2263 ( 
.A1(n_2100),
.A2(n_2171),
.B(n_2170),
.Y(n_2263)
);

INVx3_ASAP7_75t_L g2264 ( 
.A(n_2161),
.Y(n_2264)
);

OAI21xp5_ASAP7_75t_L g2265 ( 
.A1(n_2238),
.A2(n_1317),
.B(n_1316),
.Y(n_2265)
);

INVx4_ASAP7_75t_L g2266 ( 
.A(n_2105),
.Y(n_2266)
);

BUFx6f_ASAP7_75t_L g2267 ( 
.A(n_2008),
.Y(n_2267)
);

NAND2xp5_ASAP7_75t_L g2268 ( 
.A(n_2033),
.B(n_1382),
.Y(n_2268)
);

NOR2xp33_ASAP7_75t_SL g2269 ( 
.A(n_2161),
.B(n_2239),
.Y(n_2269)
);

AOI21x1_ASAP7_75t_L g2270 ( 
.A1(n_2156),
.A2(n_1068),
.B(n_1063),
.Y(n_2270)
);

INVx3_ASAP7_75t_L g2271 ( 
.A(n_2161),
.Y(n_2271)
);

O2A1O1Ixp5_ASAP7_75t_L g2272 ( 
.A1(n_2198),
.A2(n_1153),
.B(n_1239),
.C(n_1115),
.Y(n_2272)
);

OAI21xp33_ASAP7_75t_L g2273 ( 
.A1(n_1980),
.A2(n_1333),
.B(n_1321),
.Y(n_2273)
);

OAI21xp5_ASAP7_75t_L g2274 ( 
.A1(n_2074),
.A2(n_1340),
.B(n_1336),
.Y(n_2274)
);

AOI21xp5_ASAP7_75t_L g2275 ( 
.A1(n_2076),
.A2(n_1365),
.B(n_1346),
.Y(n_2275)
);

INVx2_ASAP7_75t_L g2276 ( 
.A(n_1960),
.Y(n_2276)
);

NOR2xp33_ASAP7_75t_L g2277 ( 
.A(n_2042),
.B(n_1396),
.Y(n_2277)
);

O2A1O1Ixp33_ASAP7_75t_L g2278 ( 
.A1(n_2134),
.A2(n_1374),
.B(n_1375),
.C(n_1373),
.Y(n_2278)
);

AOI22xp33_ASAP7_75t_L g2279 ( 
.A1(n_1981),
.A2(n_1099),
.B1(n_1155),
.B2(n_1078),
.Y(n_2279)
);

OAI321xp33_ASAP7_75t_L g2280 ( 
.A1(n_2073),
.A2(n_1389),
.A3(n_1078),
.B1(n_1155),
.B2(n_1173),
.C(n_1169),
.Y(n_2280)
);

O2A1O1Ixp33_ASAP7_75t_L g2281 ( 
.A1(n_2010),
.A2(n_1153),
.B(n_1239),
.C(n_1115),
.Y(n_2281)
);

INVx2_ASAP7_75t_L g2282 ( 
.A(n_1963),
.Y(n_2282)
);

NAND2xp5_ASAP7_75t_L g2283 ( 
.A(n_2228),
.B(n_1309),
.Y(n_2283)
);

NAND2xp5_ASAP7_75t_L g2284 ( 
.A(n_2237),
.B(n_1309),
.Y(n_2284)
);

AO21x1_ASAP7_75t_L g2285 ( 
.A1(n_2079),
.A2(n_658),
.B(n_657),
.Y(n_2285)
);

OAI21xp33_ASAP7_75t_L g2286 ( 
.A1(n_1941),
.A2(n_1169),
.B(n_1099),
.Y(n_2286)
);

NAND2xp5_ASAP7_75t_L g2287 ( 
.A(n_1976),
.B(n_6),
.Y(n_2287)
);

AOI22xp33_ASAP7_75t_L g2288 ( 
.A1(n_1996),
.A2(n_1173),
.B1(n_1186),
.B2(n_1169),
.Y(n_2288)
);

AOI21x1_ASAP7_75t_L g2289 ( 
.A1(n_2188),
.A2(n_1186),
.B(n_1173),
.Y(n_2289)
);

AOI221xp5_ASAP7_75t_L g2290 ( 
.A1(n_2229),
.A2(n_1190),
.B1(n_1186),
.B2(n_1041),
.C(n_1163),
.Y(n_2290)
);

INVx2_ASAP7_75t_L g2291 ( 
.A(n_1984),
.Y(n_2291)
);

AND2x4_ASAP7_75t_L g2292 ( 
.A(n_1942),
.B(n_6),
.Y(n_2292)
);

AOI21xp5_ASAP7_75t_L g2293 ( 
.A1(n_1985),
.A2(n_2203),
.B(n_2199),
.Y(n_2293)
);

NOR2xp33_ASAP7_75t_L g2294 ( 
.A(n_2053),
.B(n_6),
.Y(n_2294)
);

BUFx4f_ASAP7_75t_L g2295 ( 
.A(n_1979),
.Y(n_2295)
);

AOI21x1_ASAP7_75t_L g2296 ( 
.A1(n_1994),
.A2(n_1190),
.B(n_965),
.Y(n_2296)
);

NOR2xp33_ASAP7_75t_L g2297 ( 
.A(n_2038),
.B(n_7),
.Y(n_2297)
);

INVx11_ASAP7_75t_L g2298 ( 
.A(n_1956),
.Y(n_2298)
);

CKINVDCx5p33_ASAP7_75t_R g2299 ( 
.A(n_2243),
.Y(n_2299)
);

OAI21xp5_ASAP7_75t_L g2300 ( 
.A1(n_2241),
.A2(n_965),
.B(n_946),
.Y(n_2300)
);

BUFx4f_ASAP7_75t_L g2301 ( 
.A(n_1979),
.Y(n_2301)
);

NAND2x1p5_ASAP7_75t_L g2302 ( 
.A(n_2239),
.B(n_1041),
.Y(n_2302)
);

AOI21xp33_ASAP7_75t_L g2303 ( 
.A1(n_1944),
.A2(n_1163),
.B(n_1041),
.Y(n_2303)
);

NOR2x2_ASAP7_75t_L g2304 ( 
.A(n_1946),
.B(n_8),
.Y(n_2304)
);

BUFx3_ASAP7_75t_L g2305 ( 
.A(n_1956),
.Y(n_2305)
);

NAND2xp5_ASAP7_75t_L g2306 ( 
.A(n_1988),
.B(n_8),
.Y(n_2306)
);

HB1xp67_ASAP7_75t_L g2307 ( 
.A(n_1972),
.Y(n_2307)
);

INVx6_ASAP7_75t_L g2308 ( 
.A(n_2221),
.Y(n_2308)
);

AOI21x1_ASAP7_75t_L g2309 ( 
.A1(n_2001),
.A2(n_1252),
.B(n_1199),
.Y(n_2309)
);

NAND2xp5_ASAP7_75t_L g2310 ( 
.A(n_1997),
.B(n_9),
.Y(n_2310)
);

NAND2xp5_ASAP7_75t_L g2311 ( 
.A(n_1998),
.B(n_9),
.Y(n_2311)
);

NOR2xp33_ASAP7_75t_SL g2312 ( 
.A(n_1993),
.B(n_1252),
.Y(n_2312)
);

NAND2xp5_ASAP7_75t_L g2313 ( 
.A(n_2004),
.B(n_2006),
.Y(n_2313)
);

NAND2xp5_ASAP7_75t_L g2314 ( 
.A(n_2009),
.B(n_9),
.Y(n_2314)
);

AOI21xp5_ASAP7_75t_L g2315 ( 
.A1(n_1950),
.A2(n_1951),
.B(n_2024),
.Y(n_2315)
);

AOI21xp5_ASAP7_75t_L g2316 ( 
.A1(n_2048),
.A2(n_1370),
.B(n_1259),
.Y(n_2316)
);

NAND2xp5_ASAP7_75t_L g2317 ( 
.A(n_2011),
.B(n_10),
.Y(n_2317)
);

NOR2xp67_ASAP7_75t_L g2318 ( 
.A(n_2149),
.B(n_10),
.Y(n_2318)
);

INVx2_ASAP7_75t_L g2319 ( 
.A(n_2019),
.Y(n_2319)
);

AOI21xp5_ASAP7_75t_L g2320 ( 
.A1(n_2061),
.A2(n_1370),
.B(n_1259),
.Y(n_2320)
);

AOI21xp5_ASAP7_75t_L g2321 ( 
.A1(n_2064),
.A2(n_1377),
.B(n_1370),
.Y(n_2321)
);

AND2x6_ASAP7_75t_L g2322 ( 
.A(n_2219),
.B(n_1377),
.Y(n_2322)
);

NOR2xp33_ASAP7_75t_L g2323 ( 
.A(n_2046),
.B(n_11),
.Y(n_2323)
);

AOI21xp5_ASAP7_75t_L g2324 ( 
.A1(n_2035),
.A2(n_1377),
.B(n_11),
.Y(n_2324)
);

NAND2xp5_ASAP7_75t_L g2325 ( 
.A(n_2000),
.B(n_2021),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_SL g2326 ( 
.A(n_2204),
.B(n_1377),
.Y(n_2326)
);

AOI21xp5_ASAP7_75t_L g2327 ( 
.A1(n_2037),
.A2(n_2068),
.B(n_2012),
.Y(n_2327)
);

AOI21xp5_ASAP7_75t_L g2328 ( 
.A1(n_2057),
.A2(n_11),
.B(n_12),
.Y(n_2328)
);

INVx3_ASAP7_75t_L g2329 ( 
.A(n_2239),
.Y(n_2329)
);

AOI21xp5_ASAP7_75t_L g2330 ( 
.A1(n_2016),
.A2(n_2060),
.B(n_2082),
.Y(n_2330)
);

AOI22xp33_ASAP7_75t_L g2331 ( 
.A1(n_2181),
.A2(n_14),
.B1(n_12),
.B2(n_13),
.Y(n_2331)
);

OAI21x1_ASAP7_75t_L g2332 ( 
.A1(n_2026),
.A2(n_659),
.B(n_657),
.Y(n_2332)
);

INVx3_ASAP7_75t_L g2333 ( 
.A(n_2219),
.Y(n_2333)
);

AND2x2_ASAP7_75t_L g2334 ( 
.A(n_2002),
.B(n_12),
.Y(n_2334)
);

INVxp67_ASAP7_75t_L g2335 ( 
.A(n_1991),
.Y(n_2335)
);

AOI22xp5_ASAP7_75t_L g2336 ( 
.A1(n_2078),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.Y(n_2336)
);

O2A1O1Ixp33_ASAP7_75t_L g2337 ( 
.A1(n_2195),
.A2(n_16),
.B(n_13),
.C(n_14),
.Y(n_2337)
);

NAND2xp5_ASAP7_75t_L g2338 ( 
.A(n_2066),
.B(n_16),
.Y(n_2338)
);

INVx4_ASAP7_75t_L g2339 ( 
.A(n_2058),
.Y(n_2339)
);

NAND2xp5_ASAP7_75t_L g2340 ( 
.A(n_2030),
.B(n_17),
.Y(n_2340)
);

NAND2xp5_ASAP7_75t_SL g2341 ( 
.A(n_1955),
.B(n_18),
.Y(n_2341)
);

BUFx2_ASAP7_75t_L g2342 ( 
.A(n_2088),
.Y(n_2342)
);

BUFx4f_ASAP7_75t_L g2343 ( 
.A(n_1946),
.Y(n_2343)
);

NAND2xp5_ASAP7_75t_L g2344 ( 
.A(n_2051),
.B(n_17),
.Y(n_2344)
);

O2A1O1Ixp33_ASAP7_75t_L g2345 ( 
.A1(n_2124),
.A2(n_19),
.B(n_17),
.C(n_18),
.Y(n_2345)
);

NAND2xp5_ASAP7_75t_SL g2346 ( 
.A(n_2205),
.B(n_19),
.Y(n_2346)
);

AOI21xp33_ASAP7_75t_L g2347 ( 
.A1(n_2022),
.A2(n_18),
.B(n_19),
.Y(n_2347)
);

CKINVDCx5p33_ASAP7_75t_R g2348 ( 
.A(n_2052),
.Y(n_2348)
);

AND2x4_ASAP7_75t_L g2349 ( 
.A(n_2149),
.B(n_20),
.Y(n_2349)
);

NOR2x1_ASAP7_75t_R g2350 ( 
.A(n_2182),
.B(n_20),
.Y(n_2350)
);

O2A1O1Ixp33_ASAP7_75t_L g2351 ( 
.A1(n_1966),
.A2(n_22),
.B(n_20),
.C(n_21),
.Y(n_2351)
);

NOR2xp33_ASAP7_75t_SL g2352 ( 
.A(n_2182),
.B(n_21),
.Y(n_2352)
);

CKINVDCx11_ASAP7_75t_R g2353 ( 
.A(n_2104),
.Y(n_2353)
);

NAND2xp5_ASAP7_75t_L g2354 ( 
.A(n_2096),
.B(n_22),
.Y(n_2354)
);

A2O1A1Ixp33_ASAP7_75t_L g2355 ( 
.A1(n_2014),
.A2(n_25),
.B(n_23),
.C(n_24),
.Y(n_2355)
);

NOR2x1_ASAP7_75t_L g2356 ( 
.A(n_2177),
.B(n_24),
.Y(n_2356)
);

NAND2xp5_ASAP7_75t_L g2357 ( 
.A(n_2017),
.B(n_27),
.Y(n_2357)
);

AND2x2_ASAP7_75t_L g2358 ( 
.A(n_2059),
.B(n_27),
.Y(n_2358)
);

NOR2xp33_ASAP7_75t_L g2359 ( 
.A(n_2099),
.B(n_27),
.Y(n_2359)
);

OAI21xp5_ASAP7_75t_L g2360 ( 
.A1(n_2080),
.A2(n_28),
.B(n_29),
.Y(n_2360)
);

BUFx6f_ASAP7_75t_L g2361 ( 
.A(n_2008),
.Y(n_2361)
);

NOR2xp33_ASAP7_75t_L g2362 ( 
.A(n_2111),
.B(n_29),
.Y(n_2362)
);

NAND2xp5_ASAP7_75t_L g2363 ( 
.A(n_2028),
.B(n_29),
.Y(n_2363)
);

NAND2xp5_ASAP7_75t_L g2364 ( 
.A(n_2029),
.B(n_31),
.Y(n_2364)
);

INVx1_ASAP7_75t_L g2365 ( 
.A(n_2049),
.Y(n_2365)
);

NOR2xp33_ASAP7_75t_L g2366 ( 
.A(n_2112),
.B(n_31),
.Y(n_2366)
);

AND2x2_ASAP7_75t_L g2367 ( 
.A(n_2031),
.B(n_32),
.Y(n_2367)
);

NAND2x1p5_ASAP7_75t_L g2368 ( 
.A(n_2122),
.B(n_32),
.Y(n_2368)
);

AOI22xp33_ASAP7_75t_L g2369 ( 
.A1(n_1986),
.A2(n_35),
.B1(n_33),
.B2(n_34),
.Y(n_2369)
);

A2O1A1Ixp33_ASAP7_75t_L g2370 ( 
.A1(n_2083),
.A2(n_2150),
.B(n_2153),
.C(n_2007),
.Y(n_2370)
);

AOI22xp5_ASAP7_75t_L g2371 ( 
.A1(n_2113),
.A2(n_35),
.B1(n_33),
.B2(n_34),
.Y(n_2371)
);

OR2x6_ASAP7_75t_L g2372 ( 
.A(n_2088),
.B(n_36),
.Y(n_2372)
);

INVx2_ASAP7_75t_L g2373 ( 
.A(n_2054),
.Y(n_2373)
);

AOI211xp5_ASAP7_75t_L g2374 ( 
.A1(n_2160),
.A2(n_40),
.B(n_38),
.C(n_39),
.Y(n_2374)
);

NAND2xp5_ASAP7_75t_L g2375 ( 
.A(n_2094),
.B(n_2095),
.Y(n_2375)
);

INVx2_ASAP7_75t_SL g2376 ( 
.A(n_2221),
.Y(n_2376)
);

AOI21xp5_ASAP7_75t_L g2377 ( 
.A1(n_1978),
.A2(n_40),
.B(n_41),
.Y(n_2377)
);

NAND2xp5_ASAP7_75t_SL g2378 ( 
.A(n_2063),
.B(n_42),
.Y(n_2378)
);

A2O1A1Ixp33_ASAP7_75t_L g2379 ( 
.A1(n_1982),
.A2(n_43),
.B(n_41),
.C(n_42),
.Y(n_2379)
);

O2A1O1Ixp33_ASAP7_75t_L g2380 ( 
.A1(n_1968),
.A2(n_44),
.B(n_41),
.C(n_42),
.Y(n_2380)
);

AND2x2_ASAP7_75t_L g2381 ( 
.A(n_2244),
.B(n_44),
.Y(n_2381)
);

AOI21xp5_ASAP7_75t_L g2382 ( 
.A1(n_1983),
.A2(n_45),
.B(n_46),
.Y(n_2382)
);

BUFx6f_ASAP7_75t_L g2383 ( 
.A(n_2008),
.Y(n_2383)
);

AND2x2_ASAP7_75t_L g2384 ( 
.A(n_1995),
.B(n_45),
.Y(n_2384)
);

NOR2x1_ASAP7_75t_L g2385 ( 
.A(n_2107),
.B(n_45),
.Y(n_2385)
);

NAND2xp5_ASAP7_75t_L g2386 ( 
.A(n_2200),
.B(n_46),
.Y(n_2386)
);

NAND2xp5_ASAP7_75t_SL g2387 ( 
.A(n_2139),
.B(n_47),
.Y(n_2387)
);

BUFx3_ASAP7_75t_L g2388 ( 
.A(n_2208),
.Y(n_2388)
);

AND2x2_ASAP7_75t_L g2389 ( 
.A(n_2216),
.B(n_47),
.Y(n_2389)
);

NOR2xp33_ASAP7_75t_L g2390 ( 
.A(n_2069),
.B(n_47),
.Y(n_2390)
);

NAND2xp5_ASAP7_75t_L g2391 ( 
.A(n_2217),
.B(n_48),
.Y(n_2391)
);

NAND2xp5_ASAP7_75t_L g2392 ( 
.A(n_2220),
.B(n_2234),
.Y(n_2392)
);

INVx2_ASAP7_75t_L g2393 ( 
.A(n_2056),
.Y(n_2393)
);

AOI21x1_ASAP7_75t_L g2394 ( 
.A1(n_2174),
.A2(n_2184),
.B(n_2041),
.Y(n_2394)
);

AOI22xp5_ASAP7_75t_L g2395 ( 
.A1(n_2106),
.A2(n_50),
.B1(n_48),
.B2(n_49),
.Y(n_2395)
);

INVx1_ASAP7_75t_L g2396 ( 
.A(n_2065),
.Y(n_2396)
);

AOI21xp5_ASAP7_75t_L g2397 ( 
.A1(n_1989),
.A2(n_48),
.B(n_50),
.Y(n_2397)
);

AOI21xp5_ASAP7_75t_L g2398 ( 
.A1(n_1990),
.A2(n_50),
.B(n_51),
.Y(n_2398)
);

NOR2xp33_ASAP7_75t_L g2399 ( 
.A(n_2025),
.B(n_51),
.Y(n_2399)
);

NAND2xp5_ASAP7_75t_L g2400 ( 
.A(n_2236),
.B(n_51),
.Y(n_2400)
);

AO21x1_ASAP7_75t_L g2401 ( 
.A1(n_2034),
.A2(n_660),
.B(n_659),
.Y(n_2401)
);

NAND2xp5_ASAP7_75t_SL g2402 ( 
.A(n_2122),
.B(n_53),
.Y(n_2402)
);

HB1xp67_ASAP7_75t_L g2403 ( 
.A(n_2023),
.Y(n_2403)
);

AOI21xp5_ASAP7_75t_L g2404 ( 
.A1(n_1969),
.A2(n_52),
.B(n_53),
.Y(n_2404)
);

AOI21xp5_ASAP7_75t_L g2405 ( 
.A1(n_1977),
.A2(n_52),
.B(n_53),
.Y(n_2405)
);

INVx4_ASAP7_75t_L g2406 ( 
.A(n_2058),
.Y(n_2406)
);

NAND2xp5_ASAP7_75t_L g2407 ( 
.A(n_2240),
.B(n_54),
.Y(n_2407)
);

AOI22xp5_ASAP7_75t_L g2408 ( 
.A1(n_2109),
.A2(n_56),
.B1(n_54),
.B2(n_55),
.Y(n_2408)
);

INVx2_ASAP7_75t_SL g2409 ( 
.A(n_2122),
.Y(n_2409)
);

OAI321xp33_ASAP7_75t_L g2410 ( 
.A1(n_2167),
.A2(n_59),
.A3(n_61),
.B1(n_57),
.B2(n_58),
.C(n_60),
.Y(n_2410)
);

AOI22xp5_ASAP7_75t_L g2411 ( 
.A1(n_2222),
.A2(n_60),
.B1(n_58),
.B2(n_59),
.Y(n_2411)
);

AOI21xp5_ASAP7_75t_L g2412 ( 
.A1(n_2172),
.A2(n_58),
.B(n_59),
.Y(n_2412)
);

NAND2xp5_ASAP7_75t_L g2413 ( 
.A(n_2246),
.B(n_60),
.Y(n_2413)
);

NAND2xp5_ASAP7_75t_SL g2414 ( 
.A(n_2055),
.B(n_62),
.Y(n_2414)
);

INVx1_ASAP7_75t_L g2415 ( 
.A(n_2072),
.Y(n_2415)
);

BUFx6f_ASAP7_75t_L g2416 ( 
.A(n_2197),
.Y(n_2416)
);

NAND2xp5_ASAP7_75t_L g2417 ( 
.A(n_2247),
.B(n_62),
.Y(n_2417)
);

OAI22xp5_ASAP7_75t_L g2418 ( 
.A1(n_2091),
.A2(n_65),
.B1(n_63),
.B2(n_64),
.Y(n_2418)
);

INVxp67_ASAP7_75t_L g2419 ( 
.A(n_2209),
.Y(n_2419)
);

OAI21xp5_ASAP7_75t_L g2420 ( 
.A1(n_1964),
.A2(n_63),
.B(n_64),
.Y(n_2420)
);

NAND2xp5_ASAP7_75t_L g2421 ( 
.A(n_2248),
.B(n_63),
.Y(n_2421)
);

INVx2_ASAP7_75t_SL g2422 ( 
.A(n_2067),
.Y(n_2422)
);

NAND2xp5_ASAP7_75t_L g2423 ( 
.A(n_1957),
.B(n_65),
.Y(n_2423)
);

INVx2_ASAP7_75t_L g2424 ( 
.A(n_2114),
.Y(n_2424)
);

NAND2xp5_ASAP7_75t_L g2425 ( 
.A(n_1961),
.B(n_65),
.Y(n_2425)
);

AOI21xp5_ASAP7_75t_L g2426 ( 
.A1(n_2128),
.A2(n_66),
.B(n_67),
.Y(n_2426)
);

O2A1O1Ixp33_ASAP7_75t_SL g2427 ( 
.A1(n_2151),
.A2(n_68),
.B(n_66),
.C(n_67),
.Y(n_2427)
);

INVx11_ASAP7_75t_L g2428 ( 
.A(n_2168),
.Y(n_2428)
);

AND2x4_ASAP7_75t_L g2429 ( 
.A(n_2005),
.B(n_66),
.Y(n_2429)
);

NAND2xp5_ASAP7_75t_L g2430 ( 
.A(n_1962),
.B(n_67),
.Y(n_2430)
);

INVx1_ASAP7_75t_L g2431 ( 
.A(n_1967),
.Y(n_2431)
);

OR2x2_ASAP7_75t_L g2432 ( 
.A(n_2081),
.B(n_68),
.Y(n_2432)
);

NAND2xp5_ASAP7_75t_L g2433 ( 
.A(n_1992),
.B(n_68),
.Y(n_2433)
);

OAI21xp5_ASAP7_75t_L g2434 ( 
.A1(n_2040),
.A2(n_69),
.B(n_70),
.Y(n_2434)
);

NOR2xp33_ASAP7_75t_L g2435 ( 
.A(n_1948),
.B(n_69),
.Y(n_2435)
);

AOI21x1_ASAP7_75t_L g2436 ( 
.A1(n_2043),
.A2(n_69),
.B(n_70),
.Y(n_2436)
);

O2A1O1Ixp5_ASAP7_75t_L g2437 ( 
.A1(n_2165),
.A2(n_72),
.B(n_70),
.C(n_71),
.Y(n_2437)
);

OAI21xp5_ASAP7_75t_L g2438 ( 
.A1(n_2045),
.A2(n_71),
.B(n_72),
.Y(n_2438)
);

INVx4_ASAP7_75t_L g2439 ( 
.A(n_2023),
.Y(n_2439)
);

NAND2xp5_ASAP7_75t_L g2440 ( 
.A(n_2003),
.B(n_71),
.Y(n_2440)
);

NAND2xp5_ASAP7_75t_SL g2441 ( 
.A(n_2005),
.B(n_74),
.Y(n_2441)
);

INVx2_ASAP7_75t_L g2442 ( 
.A(n_2116),
.Y(n_2442)
);

OAI21xp5_ASAP7_75t_L g2443 ( 
.A1(n_2047),
.A2(n_73),
.B(n_74),
.Y(n_2443)
);

AOI21xp5_ASAP7_75t_L g2444 ( 
.A1(n_2131),
.A2(n_73),
.B(n_74),
.Y(n_2444)
);

BUFx6f_ASAP7_75t_L g2445 ( 
.A(n_2197),
.Y(n_2445)
);

INVx3_ASAP7_75t_L g2446 ( 
.A(n_2231),
.Y(n_2446)
);

OAI21xp5_ASAP7_75t_L g2447 ( 
.A1(n_2126),
.A2(n_75),
.B(n_76),
.Y(n_2447)
);

AOI21xp5_ASAP7_75t_L g2448 ( 
.A1(n_2155),
.A2(n_75),
.B(n_76),
.Y(n_2448)
);

BUFx12f_ASAP7_75t_L g2449 ( 
.A(n_2118),
.Y(n_2449)
);

NAND2xp5_ASAP7_75t_L g2450 ( 
.A(n_2015),
.B(n_77),
.Y(n_2450)
);

OAI21xp5_ASAP7_75t_L g2451 ( 
.A1(n_2129),
.A2(n_78),
.B(n_79),
.Y(n_2451)
);

NOR2xp33_ASAP7_75t_SL g2452 ( 
.A(n_2127),
.B(n_78),
.Y(n_2452)
);

NAND3xp33_ASAP7_75t_L g2453 ( 
.A(n_2036),
.B(n_79),
.C(n_80),
.Y(n_2453)
);

NAND2xp5_ASAP7_75t_L g2454 ( 
.A(n_2018),
.B(n_80),
.Y(n_2454)
);

OAI21xp5_ASAP7_75t_L g2455 ( 
.A1(n_2130),
.A2(n_80),
.B(n_81),
.Y(n_2455)
);

AOI21xp5_ASAP7_75t_L g2456 ( 
.A1(n_2013),
.A2(n_1970),
.B(n_1959),
.Y(n_2456)
);

INVx1_ASAP7_75t_L g2457 ( 
.A(n_2071),
.Y(n_2457)
);

NAND2xp5_ASAP7_75t_SL g2458 ( 
.A(n_2201),
.B(n_83),
.Y(n_2458)
);

OAI21xp5_ASAP7_75t_L g2459 ( 
.A1(n_2146),
.A2(n_82),
.B(n_83),
.Y(n_2459)
);

NAND2xp5_ASAP7_75t_SL g2460 ( 
.A(n_2213),
.B(n_84),
.Y(n_2460)
);

AOI21xp5_ASAP7_75t_L g2461 ( 
.A1(n_1987),
.A2(n_82),
.B(n_84),
.Y(n_2461)
);

AOI21xp5_ASAP7_75t_L g2462 ( 
.A1(n_1945),
.A2(n_2090),
.B(n_2087),
.Y(n_2462)
);

NAND2xp5_ASAP7_75t_L g2463 ( 
.A(n_1971),
.B(n_85),
.Y(n_2463)
);

INVx2_ASAP7_75t_L g2464 ( 
.A(n_2077),
.Y(n_2464)
);

INVx1_ASAP7_75t_L g2465 ( 
.A(n_2092),
.Y(n_2465)
);

AND2x4_ASAP7_75t_L g2466 ( 
.A(n_2050),
.B(n_86),
.Y(n_2466)
);

BUFx6f_ASAP7_75t_L g2467 ( 
.A(n_2231),
.Y(n_2467)
);

A2O1A1Ixp33_ASAP7_75t_L g2468 ( 
.A1(n_2102),
.A2(n_89),
.B(n_87),
.C(n_88),
.Y(n_2468)
);

INVx2_ASAP7_75t_L g2469 ( 
.A(n_2077),
.Y(n_2469)
);

NAND2xp5_ASAP7_75t_L g2470 ( 
.A(n_1965),
.B(n_87),
.Y(n_2470)
);

AOI22xp5_ASAP7_75t_L g2471 ( 
.A1(n_1954),
.A2(n_2148),
.B1(n_2159),
.B2(n_2020),
.Y(n_2471)
);

NAND2xp5_ASAP7_75t_L g2472 ( 
.A(n_2093),
.B(n_88),
.Y(n_2472)
);

OAI22xp5_ASAP7_75t_L g2473 ( 
.A1(n_2101),
.A2(n_91),
.B1(n_89),
.B2(n_90),
.Y(n_2473)
);

NAND2xp5_ASAP7_75t_L g2474 ( 
.A(n_2103),
.B(n_89),
.Y(n_2474)
);

AND2x2_ASAP7_75t_L g2475 ( 
.A(n_2215),
.B(n_90),
.Y(n_2475)
);

NAND2xp5_ASAP7_75t_L g2476 ( 
.A(n_2108),
.B(n_90),
.Y(n_2476)
);

NAND2xp5_ASAP7_75t_L g2477 ( 
.A(n_2117),
.B(n_91),
.Y(n_2477)
);

INVx1_ASAP7_75t_L g2478 ( 
.A(n_2196),
.Y(n_2478)
);

NAND2xp5_ASAP7_75t_L g2479 ( 
.A(n_2121),
.B(n_91),
.Y(n_2479)
);

INVx2_ASAP7_75t_L g2480 ( 
.A(n_2110),
.Y(n_2480)
);

NOR2xp33_ASAP7_75t_SL g2481 ( 
.A(n_2119),
.B(n_92),
.Y(n_2481)
);

NOR2xp33_ASAP7_75t_L g2482 ( 
.A(n_2039),
.B(n_2044),
.Y(n_2482)
);

CKINVDCx6p67_ASAP7_75t_R g2483 ( 
.A(n_2086),
.Y(n_2483)
);

AND2x4_ASAP7_75t_L g2484 ( 
.A(n_2070),
.B(n_93),
.Y(n_2484)
);

INVx1_ASAP7_75t_L g2485 ( 
.A(n_2125),
.Y(n_2485)
);

NOR2x1_ASAP7_75t_L g2486 ( 
.A(n_2158),
.B(n_94),
.Y(n_2486)
);

NAND2xp5_ASAP7_75t_SL g2487 ( 
.A(n_1973),
.B(n_95),
.Y(n_2487)
);

NAND2xp5_ASAP7_75t_L g2488 ( 
.A(n_1973),
.B(n_94),
.Y(n_2488)
);

NAND2xp5_ASAP7_75t_L g2489 ( 
.A(n_2212),
.B(n_95),
.Y(n_2489)
);

AOI21xp5_ASAP7_75t_L g2490 ( 
.A1(n_1974),
.A2(n_96),
.B(n_97),
.Y(n_2490)
);

AOI21xp5_ASAP7_75t_L g2491 ( 
.A1(n_2192),
.A2(n_96),
.B(n_98),
.Y(n_2491)
);

OAI21xp5_ASAP7_75t_L g2492 ( 
.A1(n_2218),
.A2(n_96),
.B(n_98),
.Y(n_2492)
);

INVx1_ASAP7_75t_L g2493 ( 
.A(n_2190),
.Y(n_2493)
);

NOR2xp33_ASAP7_75t_L g2494 ( 
.A(n_1940),
.B(n_99),
.Y(n_2494)
);

NAND2xp5_ASAP7_75t_L g2495 ( 
.A(n_2223),
.B(n_99),
.Y(n_2495)
);

NAND2xp5_ASAP7_75t_L g2496 ( 
.A(n_2232),
.B(n_99),
.Y(n_2496)
);

INVx2_ASAP7_75t_L g2497 ( 
.A(n_2193),
.Y(n_2497)
);

AO21x1_ASAP7_75t_L g2498 ( 
.A1(n_2210),
.A2(n_661),
.B(n_660),
.Y(n_2498)
);

NAND2xp5_ASAP7_75t_SL g2499 ( 
.A(n_2154),
.B(n_101),
.Y(n_2499)
);

AOI21xp5_ASAP7_75t_L g2500 ( 
.A1(n_2191),
.A2(n_100),
.B(n_101),
.Y(n_2500)
);

AND2x2_ASAP7_75t_L g2501 ( 
.A(n_2144),
.B(n_100),
.Y(n_2501)
);

NAND2xp5_ASAP7_75t_SL g2502 ( 
.A(n_2132),
.B(n_103),
.Y(n_2502)
);

AOI21xp5_ASAP7_75t_L g2503 ( 
.A1(n_1999),
.A2(n_102),
.B(n_104),
.Y(n_2503)
);

AOI21xp5_ASAP7_75t_L g2504 ( 
.A1(n_2178),
.A2(n_102),
.B(n_105),
.Y(n_2504)
);

AO21x1_ASAP7_75t_L g2505 ( 
.A1(n_2225),
.A2(n_664),
.B(n_663),
.Y(n_2505)
);

OAI21xp5_ASAP7_75t_L g2506 ( 
.A1(n_2242),
.A2(n_102),
.B(n_106),
.Y(n_2506)
);

NAND2xp5_ASAP7_75t_L g2507 ( 
.A(n_2145),
.B(n_106),
.Y(n_2507)
);

AOI21xp5_ASAP7_75t_L g2508 ( 
.A1(n_2137),
.A2(n_107),
.B(n_108),
.Y(n_2508)
);

NOR2xp33_ASAP7_75t_L g2509 ( 
.A(n_2206),
.B(n_108),
.Y(n_2509)
);

AND2x4_ASAP7_75t_L g2510 ( 
.A(n_2163),
.B(n_108),
.Y(n_2510)
);

NOR2xp33_ASAP7_75t_L g2511 ( 
.A(n_2207),
.B(n_2211),
.Y(n_2511)
);

INVx2_ASAP7_75t_L g2512 ( 
.A(n_2194),
.Y(n_2512)
);

AND2x4_ASAP7_75t_L g2513 ( 
.A(n_2075),
.B(n_2157),
.Y(n_2513)
);

NAND2xp5_ASAP7_75t_SL g2514 ( 
.A(n_2162),
.B(n_2032),
.Y(n_2514)
);

NAND2xp5_ASAP7_75t_L g2515 ( 
.A(n_2224),
.B(n_109),
.Y(n_2515)
);

OAI21xp5_ASAP7_75t_L g2516 ( 
.A1(n_2136),
.A2(n_2143),
.B(n_2140),
.Y(n_2516)
);

O2A1O1Ixp33_ASAP7_75t_L g2517 ( 
.A1(n_2185),
.A2(n_111),
.B(n_109),
.C(n_110),
.Y(n_2517)
);

INVx2_ASAP7_75t_L g2518 ( 
.A(n_2183),
.Y(n_2518)
);

OAI21xp5_ASAP7_75t_L g2519 ( 
.A1(n_2147),
.A2(n_110),
.B(n_112),
.Y(n_2519)
);

NOR2xp33_ASAP7_75t_L g2520 ( 
.A(n_2226),
.B(n_112),
.Y(n_2520)
);

BUFx8_ASAP7_75t_L g2521 ( 
.A(n_2133),
.Y(n_2521)
);

INVx4_ASAP7_75t_L g2522 ( 
.A(n_2138),
.Y(n_2522)
);

AOI21xp5_ASAP7_75t_L g2523 ( 
.A1(n_2230),
.A2(n_112),
.B(n_113),
.Y(n_2523)
);

OAI21xp5_ASAP7_75t_L g2524 ( 
.A1(n_2180),
.A2(n_113),
.B(n_114),
.Y(n_2524)
);

AOI21xp5_ASAP7_75t_L g2525 ( 
.A1(n_2233),
.A2(n_2235),
.B(n_2115),
.Y(n_2525)
);

NAND2xp5_ASAP7_75t_SL g2526 ( 
.A(n_2164),
.B(n_114),
.Y(n_2526)
);

OR2x6_ASAP7_75t_L g2527 ( 
.A(n_2120),
.B(n_113),
.Y(n_2527)
);

A2O1A1Ixp33_ASAP7_75t_L g2528 ( 
.A1(n_2227),
.A2(n_117),
.B(n_115),
.C(n_116),
.Y(n_2528)
);

BUFx2_ASAP7_75t_L g2529 ( 
.A(n_2141),
.Y(n_2529)
);

INVx3_ASAP7_75t_L g2530 ( 
.A(n_2176),
.Y(n_2530)
);

NAND2xp5_ASAP7_75t_L g2531 ( 
.A(n_2245),
.B(n_118),
.Y(n_2531)
);

BUFx6f_ASAP7_75t_L g2532 ( 
.A(n_2166),
.Y(n_2532)
);

INVx2_ASAP7_75t_L g2533 ( 
.A(n_2123),
.Y(n_2533)
);

NAND2xp5_ASAP7_75t_L g2534 ( 
.A(n_2089),
.B(n_2097),
.Y(n_2534)
);

NAND2xp5_ASAP7_75t_L g2535 ( 
.A(n_2098),
.B(n_119),
.Y(n_2535)
);

NAND2xp5_ASAP7_75t_L g2536 ( 
.A(n_2187),
.B(n_119),
.Y(n_2536)
);

INVx2_ASAP7_75t_L g2537 ( 
.A(n_2179),
.Y(n_2537)
);

AOI21xp5_ASAP7_75t_L g2538 ( 
.A1(n_2189),
.A2(n_120),
.B(n_122),
.Y(n_2538)
);

INVx1_ASAP7_75t_L g2539 ( 
.A(n_2173),
.Y(n_2539)
);

INVx4_ASAP7_75t_L g2540 ( 
.A(n_2142),
.Y(n_2540)
);

NOR2xp33_ASAP7_75t_L g2541 ( 
.A(n_2175),
.B(n_120),
.Y(n_2541)
);

INVx2_ASAP7_75t_L g2542 ( 
.A(n_2186),
.Y(n_2542)
);

AOI21xp5_ASAP7_75t_L g2543 ( 
.A1(n_2100),
.A2(n_122),
.B(n_123),
.Y(n_2543)
);

NOR2xp33_ASAP7_75t_L g2544 ( 
.A(n_1958),
.B(n_122),
.Y(n_2544)
);

INVx3_ASAP7_75t_L g2545 ( 
.A(n_2161),
.Y(n_2545)
);

AOI21xp5_ASAP7_75t_L g2546 ( 
.A1(n_2100),
.A2(n_124),
.B(n_125),
.Y(n_2546)
);

BUFx12f_ASAP7_75t_L g2547 ( 
.A(n_1956),
.Y(n_2547)
);

AOI21xp5_ASAP7_75t_L g2548 ( 
.A1(n_2100),
.A2(n_124),
.B(n_126),
.Y(n_2548)
);

A2O1A1Ixp33_ASAP7_75t_L g2549 ( 
.A1(n_2152),
.A2(n_128),
.B(n_126),
.C(n_127),
.Y(n_2549)
);

INVx2_ASAP7_75t_L g2550 ( 
.A(n_2169),
.Y(n_2550)
);

NAND2xp5_ASAP7_75t_L g2551 ( 
.A(n_2085),
.B(n_127),
.Y(n_2551)
);

NOR2xp33_ASAP7_75t_L g2552 ( 
.A(n_1958),
.B(n_128),
.Y(n_2552)
);

AOI21xp5_ASAP7_75t_L g2553 ( 
.A1(n_2100),
.A2(n_129),
.B(n_130),
.Y(n_2553)
);

AOI21xp5_ASAP7_75t_L g2554 ( 
.A1(n_2100),
.A2(n_131),
.B(n_132),
.Y(n_2554)
);

NAND2xp5_ASAP7_75t_L g2555 ( 
.A(n_2085),
.B(n_133),
.Y(n_2555)
);

BUFx2_ASAP7_75t_L g2556 ( 
.A(n_1981),
.Y(n_2556)
);

AO21x1_ASAP7_75t_L g2557 ( 
.A1(n_2079),
.A2(n_665),
.B(n_664),
.Y(n_2557)
);

NOR2xp67_ASAP7_75t_L g2558 ( 
.A(n_2149),
.B(n_133),
.Y(n_2558)
);

INVx2_ASAP7_75t_SL g2559 ( 
.A(n_2105),
.Y(n_2559)
);

NAND2xp5_ASAP7_75t_SL g2560 ( 
.A(n_1975),
.B(n_135),
.Y(n_2560)
);

NAND2xp5_ASAP7_75t_L g2561 ( 
.A(n_2085),
.B(n_134),
.Y(n_2561)
);

OAI21xp5_ASAP7_75t_L g2562 ( 
.A1(n_2062),
.A2(n_136),
.B(n_137),
.Y(n_2562)
);

O2A1O1Ixp33_ASAP7_75t_L g2563 ( 
.A1(n_2084),
.A2(n_138),
.B(n_136),
.C(n_137),
.Y(n_2563)
);

AOI21x1_ASAP7_75t_L g2564 ( 
.A1(n_2169),
.A2(n_136),
.B(n_137),
.Y(n_2564)
);

NOR2xp33_ASAP7_75t_SL g2565 ( 
.A(n_2243),
.B(n_139),
.Y(n_2565)
);

NAND2xp5_ASAP7_75t_L g2566 ( 
.A(n_2085),
.B(n_140),
.Y(n_2566)
);

NAND2xp5_ASAP7_75t_L g2567 ( 
.A(n_2085),
.B(n_141),
.Y(n_2567)
);

AO21x1_ASAP7_75t_L g2568 ( 
.A1(n_2079),
.A2(n_668),
.B(n_666),
.Y(n_2568)
);

AOI22xp5_ASAP7_75t_L g2569 ( 
.A1(n_2135),
.A2(n_143),
.B1(n_141),
.B2(n_142),
.Y(n_2569)
);

NAND2xp5_ASAP7_75t_L g2570 ( 
.A(n_2085),
.B(n_142),
.Y(n_2570)
);

CKINVDCx5p33_ASAP7_75t_R g2571 ( 
.A(n_1949),
.Y(n_2571)
);

BUFx4f_ASAP7_75t_L g2572 ( 
.A(n_1949),
.Y(n_2572)
);

O2A1O1Ixp33_ASAP7_75t_L g2573 ( 
.A1(n_2084),
.A2(n_145),
.B(n_143),
.C(n_144),
.Y(n_2573)
);

OAI21xp5_ASAP7_75t_L g2574 ( 
.A1(n_2062),
.A2(n_144),
.B(n_145),
.Y(n_2574)
);

NAND2xp5_ASAP7_75t_L g2575 ( 
.A(n_2085),
.B(n_146),
.Y(n_2575)
);

CKINVDCx10_ASAP7_75t_R g2576 ( 
.A(n_2058),
.Y(n_2576)
);

NAND2xp5_ASAP7_75t_SL g2577 ( 
.A(n_1975),
.B(n_147),
.Y(n_2577)
);

AOI21xp5_ASAP7_75t_L g2578 ( 
.A1(n_2100),
.A2(n_146),
.B(n_147),
.Y(n_2578)
);

BUFx4f_ASAP7_75t_L g2579 ( 
.A(n_1949),
.Y(n_2579)
);

INVx2_ASAP7_75t_L g2580 ( 
.A(n_2169),
.Y(n_2580)
);

AOI21xp5_ASAP7_75t_L g2581 ( 
.A1(n_2100),
.A2(n_148),
.B(n_149),
.Y(n_2581)
);

NOR2xp33_ASAP7_75t_L g2582 ( 
.A(n_1958),
.B(n_148),
.Y(n_2582)
);

NAND2xp5_ASAP7_75t_L g2583 ( 
.A(n_2085),
.B(n_149),
.Y(n_2583)
);

NAND2xp5_ASAP7_75t_L g2584 ( 
.A(n_2085),
.B(n_150),
.Y(n_2584)
);

NAND2xp5_ASAP7_75t_L g2585 ( 
.A(n_2085),
.B(n_150),
.Y(n_2585)
);

NAND2xp5_ASAP7_75t_L g2586 ( 
.A(n_2085),
.B(n_150),
.Y(n_2586)
);

CKINVDCx6p67_ASAP7_75t_R g2587 ( 
.A(n_1949),
.Y(n_2587)
);

O2A1O1Ixp33_ASAP7_75t_L g2588 ( 
.A1(n_2084),
.A2(n_153),
.B(n_151),
.C(n_152),
.Y(n_2588)
);

A2O1A1Ixp33_ASAP7_75t_L g2589 ( 
.A1(n_2152),
.A2(n_156),
.B(n_154),
.C(n_155),
.Y(n_2589)
);

BUFx2_ASAP7_75t_L g2590 ( 
.A(n_1981),
.Y(n_2590)
);

AOI21x1_ASAP7_75t_L g2591 ( 
.A1(n_2169),
.A2(n_154),
.B(n_156),
.Y(n_2591)
);

AOI21xp5_ASAP7_75t_L g2592 ( 
.A1(n_2100),
.A2(n_156),
.B(n_157),
.Y(n_2592)
);

NAND2xp5_ASAP7_75t_L g2593 ( 
.A(n_2085),
.B(n_157),
.Y(n_2593)
);

NAND2xp5_ASAP7_75t_SL g2594 ( 
.A(n_1975),
.B(n_158),
.Y(n_2594)
);

INVxp33_ASAP7_75t_L g2595 ( 
.A(n_1972),
.Y(n_2595)
);

A2O1A1Ixp33_ASAP7_75t_L g2596 ( 
.A1(n_2152),
.A2(n_160),
.B(n_158),
.C(n_159),
.Y(n_2596)
);

NOR2x2_ASAP7_75t_L g2597 ( 
.A(n_1979),
.B(n_158),
.Y(n_2597)
);

AOI21xp5_ASAP7_75t_L g2598 ( 
.A1(n_2100),
.A2(n_159),
.B(n_160),
.Y(n_2598)
);

OAI21xp5_ASAP7_75t_L g2599 ( 
.A1(n_2062),
.A2(n_160),
.B(n_161),
.Y(n_2599)
);

AOI21xp5_ASAP7_75t_L g2600 ( 
.A1(n_2100),
.A2(n_161),
.B(n_162),
.Y(n_2600)
);

NAND2xp5_ASAP7_75t_L g2601 ( 
.A(n_2085),
.B(n_162),
.Y(n_2601)
);

AOI21xp5_ASAP7_75t_L g2602 ( 
.A1(n_2100),
.A2(n_163),
.B(n_164),
.Y(n_2602)
);

AOI21xp5_ASAP7_75t_L g2603 ( 
.A1(n_2100),
.A2(n_163),
.B(n_164),
.Y(n_2603)
);

INVx1_ASAP7_75t_L g2604 ( 
.A(n_1947),
.Y(n_2604)
);

OAI21xp5_ASAP7_75t_L g2605 ( 
.A1(n_2062),
.A2(n_166),
.B(n_167),
.Y(n_2605)
);

OAI22x1_ASAP7_75t_L g2606 ( 
.A1(n_2182),
.A2(n_169),
.B1(n_167),
.B2(n_168),
.Y(n_2606)
);

NAND2xp5_ASAP7_75t_L g2607 ( 
.A(n_2085),
.B(n_169),
.Y(n_2607)
);

NAND2xp5_ASAP7_75t_L g2608 ( 
.A(n_2085),
.B(n_170),
.Y(n_2608)
);

AOI21xp5_ASAP7_75t_L g2609 ( 
.A1(n_2100),
.A2(n_171),
.B(n_172),
.Y(n_2609)
);

AO21x1_ASAP7_75t_L g2610 ( 
.A1(n_2079),
.A2(n_669),
.B(n_668),
.Y(n_2610)
);

INVx5_ASAP7_75t_L g2611 ( 
.A(n_2161),
.Y(n_2611)
);

AOI21x1_ASAP7_75t_L g2612 ( 
.A1(n_2169),
.A2(n_171),
.B(n_172),
.Y(n_2612)
);

NAND2xp5_ASAP7_75t_L g2613 ( 
.A(n_2085),
.B(n_171),
.Y(n_2613)
);

BUFx3_ASAP7_75t_L g2614 ( 
.A(n_1956),
.Y(n_2614)
);

NOR2xp33_ASAP7_75t_L g2615 ( 
.A(n_1958),
.B(n_172),
.Y(n_2615)
);

NOR2xp33_ASAP7_75t_SL g2616 ( 
.A(n_2243),
.B(n_173),
.Y(n_2616)
);

BUFx12f_ASAP7_75t_L g2617 ( 
.A(n_1956),
.Y(n_2617)
);

NOR2xp33_ASAP7_75t_L g2618 ( 
.A(n_1958),
.B(n_173),
.Y(n_2618)
);

NAND2xp5_ASAP7_75t_L g2619 ( 
.A(n_2085),
.B(n_174),
.Y(n_2619)
);

AOI22xp33_ASAP7_75t_L g2620 ( 
.A1(n_2135),
.A2(n_177),
.B1(n_175),
.B2(n_176),
.Y(n_2620)
);

INVx1_ASAP7_75t_L g2621 ( 
.A(n_1947),
.Y(n_2621)
);

OAI21xp5_ASAP7_75t_L g2622 ( 
.A1(n_2062),
.A2(n_175),
.B(n_176),
.Y(n_2622)
);

NAND2xp5_ASAP7_75t_L g2623 ( 
.A(n_2085),
.B(n_175),
.Y(n_2623)
);

OAI22xp5_ASAP7_75t_L g2624 ( 
.A1(n_2068),
.A2(n_178),
.B1(n_176),
.B2(n_177),
.Y(n_2624)
);

INVx3_ASAP7_75t_L g2625 ( 
.A(n_2161),
.Y(n_2625)
);

OAI21xp5_ASAP7_75t_L g2626 ( 
.A1(n_2062),
.A2(n_178),
.B(n_179),
.Y(n_2626)
);

NAND2xp5_ASAP7_75t_L g2627 ( 
.A(n_2085),
.B(n_178),
.Y(n_2627)
);

A2O1A1Ixp33_ASAP7_75t_L g2628 ( 
.A1(n_2152),
.A2(n_181),
.B(n_179),
.C(n_180),
.Y(n_2628)
);

OAI21xp5_ASAP7_75t_L g2629 ( 
.A1(n_2062),
.A2(n_179),
.B(n_180),
.Y(n_2629)
);

NOR2xp33_ASAP7_75t_L g2630 ( 
.A(n_1958),
.B(n_180),
.Y(n_2630)
);

AOI21xp5_ASAP7_75t_L g2631 ( 
.A1(n_2100),
.A2(n_182),
.B(n_183),
.Y(n_2631)
);

NOR2xp33_ASAP7_75t_SL g2632 ( 
.A(n_2161),
.B(n_184),
.Y(n_2632)
);

OAI22xp5_ASAP7_75t_L g2633 ( 
.A1(n_2068),
.A2(n_186),
.B1(n_184),
.B2(n_185),
.Y(n_2633)
);

NOR2xp33_ASAP7_75t_L g2634 ( 
.A(n_1958),
.B(n_185),
.Y(n_2634)
);

NAND2xp5_ASAP7_75t_SL g2635 ( 
.A(n_1975),
.B(n_186),
.Y(n_2635)
);

AND2x2_ASAP7_75t_L g2636 ( 
.A(n_2033),
.B(n_185),
.Y(n_2636)
);

NAND2xp5_ASAP7_75t_L g2637 ( 
.A(n_2085),
.B(n_188),
.Y(n_2637)
);

NAND2xp5_ASAP7_75t_L g2638 ( 
.A(n_2085),
.B(n_190),
.Y(n_2638)
);

NAND2xp5_ASAP7_75t_SL g2639 ( 
.A(n_1975),
.B(n_193),
.Y(n_2639)
);

NAND2xp5_ASAP7_75t_L g2640 ( 
.A(n_2085),
.B(n_192),
.Y(n_2640)
);

NAND2xp5_ASAP7_75t_SL g2641 ( 
.A(n_1975),
.B(n_193),
.Y(n_2641)
);

AOI21xp5_ASAP7_75t_L g2642 ( 
.A1(n_2100),
.A2(n_192),
.B(n_193),
.Y(n_2642)
);

NAND2xp5_ASAP7_75t_SL g2643 ( 
.A(n_1975),
.B(n_195),
.Y(n_2643)
);

INVx3_ASAP7_75t_L g2644 ( 
.A(n_2161),
.Y(n_2644)
);

NAND2xp5_ASAP7_75t_L g2645 ( 
.A(n_2085),
.B(n_194),
.Y(n_2645)
);

AOI21xp5_ASAP7_75t_L g2646 ( 
.A1(n_2100),
.A2(n_195),
.B(n_196),
.Y(n_2646)
);

O2A1O1Ixp33_ASAP7_75t_L g2647 ( 
.A1(n_2084),
.A2(n_197),
.B(n_195),
.C(n_196),
.Y(n_2647)
);

NOR2xp33_ASAP7_75t_L g2648 ( 
.A(n_1958),
.B(n_196),
.Y(n_2648)
);

BUFx6f_ASAP7_75t_L g2649 ( 
.A(n_2008),
.Y(n_2649)
);

AOI33xp33_ASAP7_75t_L g2650 ( 
.A1(n_2020),
.A2(n_199),
.A3(n_201),
.B1(n_197),
.B2(n_198),
.B3(n_200),
.Y(n_2650)
);

NAND2xp5_ASAP7_75t_L g2651 ( 
.A(n_2085),
.B(n_198),
.Y(n_2651)
);

OAI21xp5_ASAP7_75t_L g2652 ( 
.A1(n_2062),
.A2(n_198),
.B(n_200),
.Y(n_2652)
);

NOR2xp67_ASAP7_75t_L g2653 ( 
.A(n_2149),
.B(n_200),
.Y(n_2653)
);

NAND2xp5_ASAP7_75t_L g2654 ( 
.A(n_2085),
.B(n_201),
.Y(n_2654)
);

AOI21xp5_ASAP7_75t_L g2655 ( 
.A1(n_2100),
.A2(n_202),
.B(n_203),
.Y(n_2655)
);

NAND2xp5_ASAP7_75t_SL g2656 ( 
.A(n_1975),
.B(n_203),
.Y(n_2656)
);

NOR2xp33_ASAP7_75t_L g2657 ( 
.A(n_1958),
.B(n_204),
.Y(n_2657)
);

INVx6_ASAP7_75t_L g2658 ( 
.A(n_1956),
.Y(n_2658)
);

AOI22xp33_ASAP7_75t_L g2659 ( 
.A1(n_2135),
.A2(n_207),
.B1(n_205),
.B2(n_206),
.Y(n_2659)
);

NAND2xp5_ASAP7_75t_L g2660 ( 
.A(n_2085),
.B(n_206),
.Y(n_2660)
);

AND2x4_ASAP7_75t_L g2661 ( 
.A(n_1975),
.B(n_207),
.Y(n_2661)
);

CKINVDCx5p33_ASAP7_75t_R g2662 ( 
.A(n_1949),
.Y(n_2662)
);

NOR2xp33_ASAP7_75t_SL g2663 ( 
.A(n_2161),
.B(n_207),
.Y(n_2663)
);

INVx3_ASAP7_75t_L g2664 ( 
.A(n_2161),
.Y(n_2664)
);

AOI21xp5_ASAP7_75t_L g2665 ( 
.A1(n_2100),
.A2(n_209),
.B(n_210),
.Y(n_2665)
);

INVx1_ASAP7_75t_SL g2666 ( 
.A(n_1981),
.Y(n_2666)
);

NOR2xp33_ASAP7_75t_L g2667 ( 
.A(n_1958),
.B(n_209),
.Y(n_2667)
);

BUFx3_ASAP7_75t_L g2668 ( 
.A(n_1956),
.Y(n_2668)
);

NOR2xp33_ASAP7_75t_L g2669 ( 
.A(n_1958),
.B(n_210),
.Y(n_2669)
);

O2A1O1Ixp33_ASAP7_75t_L g2670 ( 
.A1(n_2084),
.A2(n_213),
.B(n_211),
.C(n_212),
.Y(n_2670)
);

INVx2_ASAP7_75t_SL g2671 ( 
.A(n_2105),
.Y(n_2671)
);

NAND2xp5_ASAP7_75t_L g2672 ( 
.A(n_2085),
.B(n_211),
.Y(n_2672)
);

NAND2xp5_ASAP7_75t_L g2673 ( 
.A(n_2085),
.B(n_212),
.Y(n_2673)
);

INVx1_ASAP7_75t_L g2674 ( 
.A(n_1947),
.Y(n_2674)
);

NAND2xp5_ASAP7_75t_L g2675 ( 
.A(n_2085),
.B(n_213),
.Y(n_2675)
);

NOR2xp33_ASAP7_75t_L g2676 ( 
.A(n_1958),
.B(n_214),
.Y(n_2676)
);

OAI21xp5_ASAP7_75t_L g2677 ( 
.A1(n_2062),
.A2(n_214),
.B(n_215),
.Y(n_2677)
);

O2A1O1Ixp33_ASAP7_75t_L g2678 ( 
.A1(n_2084),
.A2(n_217),
.B(n_215),
.C(n_216),
.Y(n_2678)
);

NAND2xp5_ASAP7_75t_L g2679 ( 
.A(n_2085),
.B(n_216),
.Y(n_2679)
);

BUFx4f_ASAP7_75t_L g2680 ( 
.A(n_1949),
.Y(n_2680)
);

NAND2xp5_ASAP7_75t_L g2681 ( 
.A(n_2085),
.B(n_218),
.Y(n_2681)
);

O2A1O1Ixp33_ASAP7_75t_L g2682 ( 
.A1(n_2084),
.A2(n_220),
.B(n_218),
.C(n_219),
.Y(n_2682)
);

BUFx12f_ASAP7_75t_L g2683 ( 
.A(n_1956),
.Y(n_2683)
);

AOI21xp5_ASAP7_75t_L g2684 ( 
.A1(n_2100),
.A2(n_220),
.B(n_221),
.Y(n_2684)
);

INVx1_ASAP7_75t_L g2685 ( 
.A(n_1947),
.Y(n_2685)
);

A2O1A1Ixp33_ASAP7_75t_L g2686 ( 
.A1(n_2152),
.A2(n_224),
.B(n_222),
.C(n_223),
.Y(n_2686)
);

NOR2xp33_ASAP7_75t_L g2687 ( 
.A(n_1958),
.B(n_222),
.Y(n_2687)
);

NAND2xp5_ASAP7_75t_L g2688 ( 
.A(n_2085),
.B(n_222),
.Y(n_2688)
);

NAND2xp5_ASAP7_75t_SL g2689 ( 
.A(n_1975),
.B(n_224),
.Y(n_2689)
);

AOI21xp5_ASAP7_75t_L g2690 ( 
.A1(n_2100),
.A2(n_223),
.B(n_225),
.Y(n_2690)
);

INVx1_ASAP7_75t_L g2691 ( 
.A(n_1947),
.Y(n_2691)
);

BUFx2_ASAP7_75t_L g2692 ( 
.A(n_1981),
.Y(n_2692)
);

NAND2xp5_ASAP7_75t_L g2693 ( 
.A(n_2085),
.B(n_225),
.Y(n_2693)
);

AOI21x1_ASAP7_75t_L g2694 ( 
.A1(n_2169),
.A2(n_226),
.B(n_227),
.Y(n_2694)
);

INVx5_ASAP7_75t_L g2695 ( 
.A(n_2161),
.Y(n_2695)
);

OAI321xp33_ASAP7_75t_L g2696 ( 
.A1(n_2073),
.A2(n_228),
.A3(n_230),
.B1(n_226),
.B2(n_227),
.C(n_229),
.Y(n_2696)
);

OAI21xp5_ASAP7_75t_L g2697 ( 
.A1(n_2062),
.A2(n_226),
.B(n_227),
.Y(n_2697)
);

INVx2_ASAP7_75t_L g2698 ( 
.A(n_2169),
.Y(n_2698)
);

NAND2xp5_ASAP7_75t_SL g2699 ( 
.A(n_1975),
.B(n_229),
.Y(n_2699)
);

AOI21xp5_ASAP7_75t_L g2700 ( 
.A1(n_2100),
.A2(n_228),
.B(n_230),
.Y(n_2700)
);

HB1xp67_ASAP7_75t_L g2701 ( 
.A(n_1981),
.Y(n_2701)
);

AOI21xp5_ASAP7_75t_L g2702 ( 
.A1(n_2100),
.A2(n_231),
.B(n_232),
.Y(n_2702)
);

AND2x4_ASAP7_75t_L g2703 ( 
.A(n_1975),
.B(n_231),
.Y(n_2703)
);

NOR2xp33_ASAP7_75t_L g2704 ( 
.A(n_1958),
.B(n_233),
.Y(n_2704)
);

CKINVDCx5p33_ASAP7_75t_R g2705 ( 
.A(n_1949),
.Y(n_2705)
);

INVx1_ASAP7_75t_SL g2706 ( 
.A(n_1981),
.Y(n_2706)
);

NAND2xp5_ASAP7_75t_L g2707 ( 
.A(n_2085),
.B(n_233),
.Y(n_2707)
);

O2A1O1Ixp5_ASAP7_75t_L g2708 ( 
.A1(n_2100),
.A2(n_236),
.B(n_234),
.C(n_235),
.Y(n_2708)
);

NOR2xp33_ASAP7_75t_L g2709 ( 
.A(n_1958),
.B(n_235),
.Y(n_2709)
);

OAI21xp5_ASAP7_75t_L g2710 ( 
.A1(n_2062),
.A2(n_235),
.B(n_236),
.Y(n_2710)
);

INVxp67_ASAP7_75t_L g2711 ( 
.A(n_1981),
.Y(n_2711)
);

INVx4_ASAP7_75t_L g2712 ( 
.A(n_2105),
.Y(n_2712)
);

NAND2xp5_ASAP7_75t_L g2713 ( 
.A(n_2085),
.B(n_237),
.Y(n_2713)
);

NAND2xp5_ASAP7_75t_L g2714 ( 
.A(n_2085),
.B(n_237),
.Y(n_2714)
);

O2A1O1Ixp33_ASAP7_75t_L g2715 ( 
.A1(n_2084),
.A2(n_241),
.B(n_238),
.C(n_240),
.Y(n_2715)
);

NAND2xp5_ASAP7_75t_L g2716 ( 
.A(n_2085),
.B(n_238),
.Y(n_2716)
);

AOI22xp5_ASAP7_75t_L g2717 ( 
.A1(n_2135),
.A2(n_244),
.B1(n_242),
.B2(n_243),
.Y(n_2717)
);

AOI21xp5_ASAP7_75t_L g2718 ( 
.A1(n_2100),
.A2(n_244),
.B(n_245),
.Y(n_2718)
);

NOR2xp67_ASAP7_75t_L g2719 ( 
.A(n_2149),
.B(n_244),
.Y(n_2719)
);

NAND2xp5_ASAP7_75t_L g2720 ( 
.A(n_2085),
.B(n_245),
.Y(n_2720)
);

AND2x2_ASAP7_75t_L g2721 ( 
.A(n_2033),
.B(n_245),
.Y(n_2721)
);

NOR2xp33_ASAP7_75t_SL g2722 ( 
.A(n_2243),
.B(n_246),
.Y(n_2722)
);

HB1xp67_ASAP7_75t_L g2723 ( 
.A(n_1981),
.Y(n_2723)
);

BUFx6f_ASAP7_75t_L g2724 ( 
.A(n_2008),
.Y(n_2724)
);

A2O1A1Ixp33_ASAP7_75t_L g2725 ( 
.A1(n_2152),
.A2(n_248),
.B(n_246),
.C(n_247),
.Y(n_2725)
);

INVx1_ASAP7_75t_L g2726 ( 
.A(n_1947),
.Y(n_2726)
);

INVxp67_ASAP7_75t_L g2727 ( 
.A(n_1981),
.Y(n_2727)
);

NAND2x1p5_ASAP7_75t_L g2728 ( 
.A(n_2239),
.B(n_249),
.Y(n_2728)
);

CKINVDCx20_ASAP7_75t_R g2729 ( 
.A(n_1956),
.Y(n_2729)
);

INVx1_ASAP7_75t_L g2730 ( 
.A(n_1947),
.Y(n_2730)
);

INVx1_ASAP7_75t_L g2731 ( 
.A(n_1947),
.Y(n_2731)
);

NAND2xp5_ASAP7_75t_L g2732 ( 
.A(n_2085),
.B(n_250),
.Y(n_2732)
);

CKINVDCx5p33_ASAP7_75t_R g2733 ( 
.A(n_1949),
.Y(n_2733)
);

INVx3_ASAP7_75t_L g2734 ( 
.A(n_2161),
.Y(n_2734)
);

A2O1A1Ixp33_ASAP7_75t_L g2735 ( 
.A1(n_2152),
.A2(n_252),
.B(n_250),
.C(n_251),
.Y(n_2735)
);

AOI21xp5_ASAP7_75t_L g2736 ( 
.A1(n_2100),
.A2(n_250),
.B(n_251),
.Y(n_2736)
);

NAND2xp5_ASAP7_75t_L g2737 ( 
.A(n_2085),
.B(n_252),
.Y(n_2737)
);

NOR2xp33_ASAP7_75t_R g2738 ( 
.A(n_2729),
.B(n_253),
.Y(n_2738)
);

AOI22xp33_ASAP7_75t_L g2739 ( 
.A1(n_2372),
.A2(n_255),
.B1(n_253),
.B2(n_254),
.Y(n_2739)
);

NAND2xp5_ASAP7_75t_L g2740 ( 
.A(n_2457),
.B(n_254),
.Y(n_2740)
);

NAND2xp5_ASAP7_75t_L g2741 ( 
.A(n_2465),
.B(n_255),
.Y(n_2741)
);

NAND2xp5_ASAP7_75t_L g2742 ( 
.A(n_2325),
.B(n_255),
.Y(n_2742)
);

BUFx6f_ASAP7_75t_L g2743 ( 
.A(n_2267),
.Y(n_2743)
);

AOI22xp33_ASAP7_75t_L g2744 ( 
.A1(n_2372),
.A2(n_258),
.B1(n_256),
.B2(n_257),
.Y(n_2744)
);

INVx2_ASAP7_75t_L g2745 ( 
.A(n_2276),
.Y(n_2745)
);

INVxp33_ASAP7_75t_SL g2746 ( 
.A(n_2350),
.Y(n_2746)
);

NOR2xp33_ASAP7_75t_L g2747 ( 
.A(n_2595),
.B(n_256),
.Y(n_2747)
);

INVx2_ASAP7_75t_L g2748 ( 
.A(n_2282),
.Y(n_2748)
);

AOI21xp5_ASAP7_75t_L g2749 ( 
.A1(n_2330),
.A2(n_256),
.B(n_257),
.Y(n_2749)
);

INVx2_ASAP7_75t_L g2750 ( 
.A(n_2291),
.Y(n_2750)
);

NAND3xp33_ASAP7_75t_SL g2751 ( 
.A(n_2565),
.B(n_2722),
.C(n_2616),
.Y(n_2751)
);

OR2x6_ASAP7_75t_L g2752 ( 
.A(n_2547),
.B(n_258),
.Y(n_2752)
);

AOI21xp5_ASAP7_75t_L g2753 ( 
.A1(n_2327),
.A2(n_259),
.B(n_260),
.Y(n_2753)
);

AOI21xp5_ASAP7_75t_L g2754 ( 
.A1(n_2263),
.A2(n_259),
.B(n_260),
.Y(n_2754)
);

AOI21xp5_ASAP7_75t_L g2755 ( 
.A1(n_2315),
.A2(n_259),
.B(n_260),
.Y(n_2755)
);

AOI21xp5_ASAP7_75t_L g2756 ( 
.A1(n_2462),
.A2(n_261),
.B(n_262),
.Y(n_2756)
);

OAI22x1_ASAP7_75t_L g2757 ( 
.A1(n_2569),
.A2(n_2717),
.B1(n_2336),
.B2(n_2439),
.Y(n_2757)
);

OAI21xp33_ASAP7_75t_L g2758 ( 
.A1(n_2273),
.A2(n_262),
.B(n_263),
.Y(n_2758)
);

INVx1_ASAP7_75t_L g2759 ( 
.A(n_2319),
.Y(n_2759)
);

AOI21xp5_ASAP7_75t_L g2760 ( 
.A1(n_2293),
.A2(n_263),
.B(n_264),
.Y(n_2760)
);

NAND2xp5_ASAP7_75t_L g2761 ( 
.A(n_2392),
.B(n_264),
.Y(n_2761)
);

NAND2xp5_ASAP7_75t_L g2762 ( 
.A(n_2253),
.B(n_265),
.Y(n_2762)
);

INVx1_ASAP7_75t_L g2763 ( 
.A(n_2256),
.Y(n_2763)
);

NAND3xp33_ASAP7_75t_SL g2764 ( 
.A(n_2374),
.B(n_265),
.C(n_266),
.Y(n_2764)
);

AOI22xp5_ASAP7_75t_L g2765 ( 
.A1(n_2471),
.A2(n_268),
.B1(n_266),
.B2(n_267),
.Y(n_2765)
);

INVx2_ASAP7_75t_SL g2766 ( 
.A(n_2298),
.Y(n_2766)
);

BUFx3_ASAP7_75t_L g2767 ( 
.A(n_2617),
.Y(n_2767)
);

CKINVDCx14_ASAP7_75t_R g2768 ( 
.A(n_2587),
.Y(n_2768)
);

AOI21xp5_ASAP7_75t_L g2769 ( 
.A1(n_2370),
.A2(n_268),
.B(n_269),
.Y(n_2769)
);

NAND2xp5_ASAP7_75t_L g2770 ( 
.A(n_2260),
.B(n_2261),
.Y(n_2770)
);

A2O1A1Ixp33_ASAP7_75t_L g2771 ( 
.A1(n_2435),
.A2(n_273),
.B(n_271),
.C(n_272),
.Y(n_2771)
);

INVx3_ASAP7_75t_L g2772 ( 
.A(n_2611),
.Y(n_2772)
);

INVx2_ASAP7_75t_L g2773 ( 
.A(n_2373),
.Y(n_2773)
);

O2A1O1Ixp5_ASAP7_75t_L g2774 ( 
.A1(n_2533),
.A2(n_273),
.B(n_271),
.C(n_272),
.Y(n_2774)
);

BUFx2_ASAP7_75t_L g2775 ( 
.A(n_2556),
.Y(n_2775)
);

AOI22xp33_ASAP7_75t_L g2776 ( 
.A1(n_2323),
.A2(n_276),
.B1(n_274),
.B2(n_275),
.Y(n_2776)
);

AOI21x1_ASAP7_75t_L g2777 ( 
.A1(n_2394),
.A2(n_274),
.B(n_275),
.Y(n_2777)
);

HB1xp67_ASAP7_75t_L g2778 ( 
.A(n_2666),
.Y(n_2778)
);

BUFx12f_ASAP7_75t_L g2779 ( 
.A(n_2683),
.Y(n_2779)
);

NAND2xp5_ASAP7_75t_SL g2780 ( 
.A(n_2343),
.B(n_669),
.Y(n_2780)
);

OR2x6_ASAP7_75t_L g2781 ( 
.A(n_2308),
.B(n_276),
.Y(n_2781)
);

O2A1O1Ixp33_ASAP7_75t_L g2782 ( 
.A1(n_2262),
.A2(n_279),
.B(n_277),
.C(n_278),
.Y(n_2782)
);

NOR2xp67_ASAP7_75t_SL g2783 ( 
.A(n_2305),
.B(n_277),
.Y(n_2783)
);

NOR2xp33_ASAP7_75t_SL g2784 ( 
.A(n_2572),
.B(n_278),
.Y(n_2784)
);

AO32x1_ASAP7_75t_L g2785 ( 
.A1(n_2473),
.A2(n_280),
.A3(n_278),
.B1(n_279),
.B2(n_281),
.Y(n_2785)
);

BUFx6f_ASAP7_75t_L g2786 ( 
.A(n_2267),
.Y(n_2786)
);

NAND2xp5_ASAP7_75t_L g2787 ( 
.A(n_2604),
.B(n_280),
.Y(n_2787)
);

NOR2xp33_ASAP7_75t_L g2788 ( 
.A(n_2706),
.B(n_281),
.Y(n_2788)
);

NOR2xp33_ASAP7_75t_L g2789 ( 
.A(n_2307),
.B(n_282),
.Y(n_2789)
);

BUFx6f_ASAP7_75t_L g2790 ( 
.A(n_2267),
.Y(n_2790)
);

NAND2xp5_ASAP7_75t_SL g2791 ( 
.A(n_2343),
.B(n_670),
.Y(n_2791)
);

CKINVDCx8_ASAP7_75t_R g2792 ( 
.A(n_2576),
.Y(n_2792)
);

NAND2xp5_ASAP7_75t_SL g2793 ( 
.A(n_2312),
.B(n_670),
.Y(n_2793)
);

INVx2_ASAP7_75t_L g2794 ( 
.A(n_2393),
.Y(n_2794)
);

NAND2xp5_ASAP7_75t_L g2795 ( 
.A(n_2621),
.B(n_282),
.Y(n_2795)
);

NOR2xp33_ASAP7_75t_L g2796 ( 
.A(n_2439),
.B(n_282),
.Y(n_2796)
);

NAND2xp5_ASAP7_75t_SL g2797 ( 
.A(n_2295),
.B(n_671),
.Y(n_2797)
);

NAND3xp33_ASAP7_75t_SL g2798 ( 
.A(n_2374),
.B(n_283),
.C(n_284),
.Y(n_2798)
);

AOI221xp5_ASAP7_75t_L g2799 ( 
.A1(n_2273),
.A2(n_285),
.B1(n_283),
.B2(n_284),
.C(n_286),
.Y(n_2799)
);

NAND2xp5_ASAP7_75t_L g2800 ( 
.A(n_2674),
.B(n_283),
.Y(n_2800)
);

AND2x4_ASAP7_75t_L g2801 ( 
.A(n_2522),
.B(n_284),
.Y(n_2801)
);

NAND2xp5_ASAP7_75t_L g2802 ( 
.A(n_2685),
.B(n_285),
.Y(n_2802)
);

NOR2xp33_ASAP7_75t_R g2803 ( 
.A(n_2299),
.B(n_286),
.Y(n_2803)
);

AND2x4_ASAP7_75t_L g2804 ( 
.A(n_2522),
.B(n_287),
.Y(n_2804)
);

AOI22xp5_ASAP7_75t_L g2805 ( 
.A1(n_2471),
.A2(n_2297),
.B1(n_2254),
.B2(n_2277),
.Y(n_2805)
);

NAND2xp5_ASAP7_75t_SL g2806 ( 
.A(n_2295),
.B(n_672),
.Y(n_2806)
);

INVx3_ASAP7_75t_L g2807 ( 
.A(n_2611),
.Y(n_2807)
);

AOI21xp5_ASAP7_75t_L g2808 ( 
.A1(n_2286),
.A2(n_287),
.B(n_288),
.Y(n_2808)
);

NAND2xp5_ASAP7_75t_SL g2809 ( 
.A(n_2301),
.B(n_673),
.Y(n_2809)
);

NAND2xp5_ASAP7_75t_L g2810 ( 
.A(n_2691),
.B(n_289),
.Y(n_2810)
);

NOR2xp33_ASAP7_75t_SL g2811 ( 
.A(n_2572),
.B(n_2579),
.Y(n_2811)
);

AO21x2_ASAP7_75t_L g2812 ( 
.A1(n_2300),
.A2(n_289),
.B(n_290),
.Y(n_2812)
);

BUFx6f_ASAP7_75t_L g2813 ( 
.A(n_2361),
.Y(n_2813)
);

NOR2xp33_ASAP7_75t_L g2814 ( 
.A(n_2711),
.B(n_289),
.Y(n_2814)
);

NAND2x1_ASAP7_75t_L g2815 ( 
.A(n_2322),
.B(n_291),
.Y(n_2815)
);

NOR2xp67_ASAP7_75t_L g2816 ( 
.A(n_2259),
.B(n_292),
.Y(n_2816)
);

NOR2xp33_ASAP7_75t_R g2817 ( 
.A(n_2258),
.B(n_293),
.Y(n_2817)
);

A2O1A1Ixp33_ASAP7_75t_L g2818 ( 
.A1(n_2736),
.A2(n_296),
.B(n_294),
.C(n_295),
.Y(n_2818)
);

INVx2_ASAP7_75t_L g2819 ( 
.A(n_2255),
.Y(n_2819)
);

O2A1O1Ixp33_ASAP7_75t_L g2820 ( 
.A1(n_2468),
.A2(n_297),
.B(n_294),
.C(n_295),
.Y(n_2820)
);

INVx3_ASAP7_75t_L g2821 ( 
.A(n_2611),
.Y(n_2821)
);

AOI22xp5_ASAP7_75t_L g2822 ( 
.A1(n_2292),
.A2(n_298),
.B1(n_295),
.B2(n_297),
.Y(n_2822)
);

BUFx6f_ASAP7_75t_L g2823 ( 
.A(n_2361),
.Y(n_2823)
);

NOR2xp33_ASAP7_75t_L g2824 ( 
.A(n_2727),
.B(n_297),
.Y(n_2824)
);

INVx2_ASAP7_75t_L g2825 ( 
.A(n_2550),
.Y(n_2825)
);

NAND2xp5_ASAP7_75t_L g2826 ( 
.A(n_2726),
.B(n_298),
.Y(n_2826)
);

O2A1O1Ixp33_ASAP7_75t_L g2827 ( 
.A1(n_2363),
.A2(n_301),
.B(n_299),
.C(n_300),
.Y(n_2827)
);

O2A1O1Ixp33_ASAP7_75t_L g2828 ( 
.A1(n_2345),
.A2(n_302),
.B(n_300),
.C(n_301),
.Y(n_2828)
);

A2O1A1Ixp33_ASAP7_75t_L g2829 ( 
.A1(n_2543),
.A2(n_305),
.B(n_303),
.C(n_304),
.Y(n_2829)
);

NOR2xp33_ASAP7_75t_L g2830 ( 
.A(n_2529),
.B(n_303),
.Y(n_2830)
);

NOR2xp33_ASAP7_75t_L g2831 ( 
.A(n_2342),
.B(n_303),
.Y(n_2831)
);

NAND2xp5_ASAP7_75t_L g2832 ( 
.A(n_2730),
.B(n_304),
.Y(n_2832)
);

NAND2xp5_ASAP7_75t_SL g2833 ( 
.A(n_2301),
.B(n_673),
.Y(n_2833)
);

O2A1O1Ixp33_ASAP7_75t_L g2834 ( 
.A1(n_2347),
.A2(n_2454),
.B(n_2450),
.C(n_2489),
.Y(n_2834)
);

OAI22xp5_ASAP7_75t_SL g2835 ( 
.A1(n_2527),
.A2(n_307),
.B1(n_305),
.B2(n_306),
.Y(n_2835)
);

AOI21xp5_ASAP7_75t_L g2836 ( 
.A1(n_2280),
.A2(n_308),
.B(n_309),
.Y(n_2836)
);

OAI22xp5_ASAP7_75t_L g2837 ( 
.A1(n_2527),
.A2(n_2336),
.B1(n_2371),
.B2(n_2357),
.Y(n_2837)
);

NAND2xp5_ASAP7_75t_L g2838 ( 
.A(n_2731),
.B(n_309),
.Y(n_2838)
);

BUFx2_ASAP7_75t_L g2839 ( 
.A(n_2590),
.Y(n_2839)
);

NOR3xp33_ASAP7_75t_SL g2840 ( 
.A(n_2571),
.B(n_310),
.C(n_311),
.Y(n_2840)
);

AO21x1_ASAP7_75t_L g2841 ( 
.A1(n_2481),
.A2(n_676),
.B(n_674),
.Y(n_2841)
);

BUFx6f_ASAP7_75t_L g2842 ( 
.A(n_2361),
.Y(n_2842)
);

BUFx3_ASAP7_75t_L g2843 ( 
.A(n_2614),
.Y(n_2843)
);

A2O1A1Ixp33_ASAP7_75t_L g2844 ( 
.A1(n_2546),
.A2(n_312),
.B(n_310),
.C(n_311),
.Y(n_2844)
);

AND2x4_ASAP7_75t_L g2845 ( 
.A(n_2259),
.B(n_312),
.Y(n_2845)
);

NAND2xp5_ASAP7_75t_L g2846 ( 
.A(n_2313),
.B(n_312),
.Y(n_2846)
);

NOR2xp67_ASAP7_75t_L g2847 ( 
.A(n_2266),
.B(n_313),
.Y(n_2847)
);

O2A1O1Ixp33_ASAP7_75t_L g2848 ( 
.A1(n_2495),
.A2(n_315),
.B(n_313),
.C(n_314),
.Y(n_2848)
);

BUFx6f_ASAP7_75t_L g2849 ( 
.A(n_2383),
.Y(n_2849)
);

OAI22xp5_ASAP7_75t_L g2850 ( 
.A1(n_2371),
.A2(n_2408),
.B1(n_2395),
.B2(n_2429),
.Y(n_2850)
);

AND2x2_ASAP7_75t_L g2851 ( 
.A(n_2358),
.B(n_315),
.Y(n_2851)
);

AO32x1_ASAP7_75t_L g2852 ( 
.A1(n_2624),
.A2(n_318),
.A3(n_316),
.B1(n_317),
.B2(n_319),
.Y(n_2852)
);

INVx3_ASAP7_75t_L g2853 ( 
.A(n_2695),
.Y(n_2853)
);

INVx6_ASAP7_75t_L g2854 ( 
.A(n_2521),
.Y(n_2854)
);

NOR2xp33_ASAP7_75t_L g2855 ( 
.A(n_2403),
.B(n_316),
.Y(n_2855)
);

INVx2_ASAP7_75t_L g2856 ( 
.A(n_2580),
.Y(n_2856)
);

NOR2xp33_ASAP7_75t_L g2857 ( 
.A(n_2692),
.B(n_316),
.Y(n_2857)
);

AOI21xp5_ASAP7_75t_L g2858 ( 
.A1(n_2375),
.A2(n_317),
.B(n_318),
.Y(n_2858)
);

NAND2xp5_ASAP7_75t_SL g2859 ( 
.A(n_2352),
.B(n_676),
.Y(n_2859)
);

NAND2xp5_ASAP7_75t_L g2860 ( 
.A(n_2367),
.B(n_317),
.Y(n_2860)
);

OAI22xp5_ASAP7_75t_L g2861 ( 
.A1(n_2395),
.A2(n_320),
.B1(n_318),
.B2(n_319),
.Y(n_2861)
);

NOR3xp33_ASAP7_75t_L g2862 ( 
.A(n_2294),
.B(n_320),
.C(n_321),
.Y(n_2862)
);

O2A1O1Ixp33_ASAP7_75t_L g2863 ( 
.A1(n_2496),
.A2(n_322),
.B(n_320),
.C(n_321),
.Y(n_2863)
);

BUFx6f_ASAP7_75t_L g2864 ( 
.A(n_2383),
.Y(n_2864)
);

A2O1A1Ixp33_ASAP7_75t_L g2865 ( 
.A1(n_2548),
.A2(n_324),
.B(n_322),
.C(n_323),
.Y(n_2865)
);

NAND2xp5_ASAP7_75t_L g2866 ( 
.A(n_2493),
.B(n_323),
.Y(n_2866)
);

AOI22xp33_ASAP7_75t_L g2867 ( 
.A1(n_2544),
.A2(n_326),
.B1(n_324),
.B2(n_325),
.Y(n_2867)
);

AOI22xp33_ASAP7_75t_L g2868 ( 
.A1(n_2552),
.A2(n_327),
.B1(n_325),
.B2(n_326),
.Y(n_2868)
);

OAI21xp5_ASAP7_75t_L g2869 ( 
.A1(n_2272),
.A2(n_326),
.B(n_327),
.Y(n_2869)
);

AOI22xp5_ASAP7_75t_L g2870 ( 
.A1(n_2292),
.A2(n_330),
.B1(n_328),
.B2(n_329),
.Y(n_2870)
);

HAxp5_ASAP7_75t_L g2871 ( 
.A(n_2597),
.B(n_330),
.CON(n_2871),
.SN(n_2871)
);

INVx1_ASAP7_75t_L g2872 ( 
.A(n_2365),
.Y(n_2872)
);

INVx1_ASAP7_75t_SL g2873 ( 
.A(n_2701),
.Y(n_2873)
);

NOR2xp67_ASAP7_75t_SL g2874 ( 
.A(n_2668),
.B(n_331),
.Y(n_2874)
);

INVxp67_ASAP7_75t_L g2875 ( 
.A(n_2723),
.Y(n_2875)
);

CKINVDCx5p33_ASAP7_75t_R g2876 ( 
.A(n_2579),
.Y(n_2876)
);

NAND2xp5_ASAP7_75t_L g2877 ( 
.A(n_2384),
.B(n_332),
.Y(n_2877)
);

NAND2xp5_ASAP7_75t_SL g2878 ( 
.A(n_2632),
.B(n_677),
.Y(n_2878)
);

AOI21x1_ASAP7_75t_L g2879 ( 
.A1(n_2289),
.A2(n_333),
.B(n_334),
.Y(n_2879)
);

O2A1O1Ixp33_ASAP7_75t_SL g2880 ( 
.A1(n_2528),
.A2(n_335),
.B(n_333),
.C(n_334),
.Y(n_2880)
);

NOR2xp33_ASAP7_75t_L g2881 ( 
.A(n_2257),
.B(n_334),
.Y(n_2881)
);

NAND2xp5_ASAP7_75t_L g2882 ( 
.A(n_2396),
.B(n_335),
.Y(n_2882)
);

INVxp67_ASAP7_75t_SL g2883 ( 
.A(n_2632),
.Y(n_2883)
);

CKINVDCx20_ASAP7_75t_R g2884 ( 
.A(n_2353),
.Y(n_2884)
);

NAND2xp5_ASAP7_75t_SL g2885 ( 
.A(n_2663),
.B(n_677),
.Y(n_2885)
);

INVx1_ASAP7_75t_L g2886 ( 
.A(n_2415),
.Y(n_2886)
);

OAI21xp5_ASAP7_75t_L g2887 ( 
.A1(n_2274),
.A2(n_336),
.B(n_337),
.Y(n_2887)
);

O2A1O1Ixp33_ASAP7_75t_L g2888 ( 
.A1(n_2281),
.A2(n_339),
.B(n_337),
.C(n_338),
.Y(n_2888)
);

BUFx3_ASAP7_75t_L g2889 ( 
.A(n_2308),
.Y(n_2889)
);

NAND2xp5_ASAP7_75t_L g2890 ( 
.A(n_2431),
.B(n_337),
.Y(n_2890)
);

AOI21xp5_ASAP7_75t_L g2891 ( 
.A1(n_2516),
.A2(n_339),
.B(n_340),
.Y(n_2891)
);

AOI21xp5_ASAP7_75t_L g2892 ( 
.A1(n_2553),
.A2(n_339),
.B(n_340),
.Y(n_2892)
);

AND2x2_ASAP7_75t_L g2893 ( 
.A(n_2334),
.B(n_341),
.Y(n_2893)
);

AND2x4_ASAP7_75t_L g2894 ( 
.A(n_2266),
.B(n_2712),
.Y(n_2894)
);

BUFx6f_ASAP7_75t_L g2895 ( 
.A(n_2383),
.Y(n_2895)
);

OR2x6_ASAP7_75t_L g2896 ( 
.A(n_2658),
.B(n_341),
.Y(n_2896)
);

AND2x2_ASAP7_75t_L g2897 ( 
.A(n_2381),
.B(n_341),
.Y(n_2897)
);

INVx6_ASAP7_75t_L g2898 ( 
.A(n_2658),
.Y(n_2898)
);

OAI22x1_ASAP7_75t_L g2899 ( 
.A1(n_2569),
.A2(n_344),
.B1(n_342),
.B2(n_343),
.Y(n_2899)
);

NOR2xp33_ASAP7_75t_R g2900 ( 
.A(n_2662),
.B(n_342),
.Y(n_2900)
);

NAND2xp5_ASAP7_75t_SL g2901 ( 
.A(n_2663),
.B(n_678),
.Y(n_2901)
);

INVx2_ASAP7_75t_SL g2902 ( 
.A(n_2680),
.Y(n_2902)
);

NAND2xp33_ASAP7_75t_R g2903 ( 
.A(n_2348),
.B(n_342),
.Y(n_2903)
);

NOR3xp33_ASAP7_75t_SL g2904 ( 
.A(n_2705),
.B(n_344),
.C(n_345),
.Y(n_2904)
);

O2A1O1Ixp5_ASAP7_75t_L g2905 ( 
.A1(n_2303),
.A2(n_346),
.B(n_344),
.C(n_345),
.Y(n_2905)
);

INVx2_ASAP7_75t_L g2906 ( 
.A(n_2698),
.Y(n_2906)
);

AND2x2_ASAP7_75t_L g2907 ( 
.A(n_2501),
.B(n_346),
.Y(n_2907)
);

INVx3_ASAP7_75t_L g2908 ( 
.A(n_2695),
.Y(n_2908)
);

NAND2xp5_ASAP7_75t_SL g2909 ( 
.A(n_2481),
.B(n_2661),
.Y(n_2909)
);

HB1xp67_ASAP7_75t_L g2910 ( 
.A(n_2661),
.Y(n_2910)
);

AOI21xp5_ASAP7_75t_L g2911 ( 
.A1(n_2554),
.A2(n_347),
.B(n_348),
.Y(n_2911)
);

NAND2xp5_ASAP7_75t_L g2912 ( 
.A(n_2389),
.B(n_349),
.Y(n_2912)
);

AND2x4_ASAP7_75t_L g2913 ( 
.A(n_2712),
.B(n_349),
.Y(n_2913)
);

NAND2xp5_ASAP7_75t_SL g2914 ( 
.A(n_2703),
.B(n_678),
.Y(n_2914)
);

NAND2xp5_ASAP7_75t_L g2915 ( 
.A(n_2539),
.B(n_350),
.Y(n_2915)
);

AOI22xp5_ASAP7_75t_L g2916 ( 
.A1(n_2390),
.A2(n_353),
.B1(n_351),
.B2(n_352),
.Y(n_2916)
);

INVx2_ASAP7_75t_L g2917 ( 
.A(n_2424),
.Y(n_2917)
);

OAI22xp5_ASAP7_75t_L g2918 ( 
.A1(n_2429),
.A2(n_356),
.B1(n_353),
.B2(n_355),
.Y(n_2918)
);

INVx1_ASAP7_75t_L g2919 ( 
.A(n_2703),
.Y(n_2919)
);

NAND2xp5_ASAP7_75t_SL g2920 ( 
.A(n_2452),
.B(n_679),
.Y(n_2920)
);

OAI22xp5_ASAP7_75t_L g2921 ( 
.A1(n_2717),
.A2(n_358),
.B1(n_356),
.B2(n_357),
.Y(n_2921)
);

NAND2xp5_ASAP7_75t_SL g2922 ( 
.A(n_2335),
.B(n_680),
.Y(n_2922)
);

INVx1_ASAP7_75t_L g2923 ( 
.A(n_2287),
.Y(n_2923)
);

OAI21x1_ASAP7_75t_L g2924 ( 
.A1(n_2296),
.A2(n_356),
.B(n_357),
.Y(n_2924)
);

O2A1O1Ixp5_ASAP7_75t_L g2925 ( 
.A1(n_2526),
.A2(n_360),
.B(n_358),
.C(n_359),
.Y(n_2925)
);

NOR2xp33_ASAP7_75t_L g2926 ( 
.A(n_2458),
.B(n_361),
.Y(n_2926)
);

INVx2_ASAP7_75t_L g2927 ( 
.A(n_2442),
.Y(n_2927)
);

O2A1O1Ixp5_ASAP7_75t_L g2928 ( 
.A1(n_2285),
.A2(n_364),
.B(n_362),
.C(n_363),
.Y(n_2928)
);

AND2x6_ASAP7_75t_SL g2929 ( 
.A(n_2680),
.B(n_363),
.Y(n_2929)
);

OR2x6_ASAP7_75t_L g2930 ( 
.A(n_2376),
.B(n_363),
.Y(n_2930)
);

NOR2xp33_ASAP7_75t_L g2931 ( 
.A(n_2460),
.B(n_364),
.Y(n_2931)
);

OAI21xp33_ASAP7_75t_SL g2932 ( 
.A1(n_2650),
.A2(n_364),
.B(n_365),
.Y(n_2932)
);

NAND2xp5_ASAP7_75t_L g2933 ( 
.A(n_2432),
.B(n_365),
.Y(n_2933)
);

NOR2xp33_ASAP7_75t_L g2934 ( 
.A(n_2482),
.B(n_2514),
.Y(n_2934)
);

NAND2xp5_ASAP7_75t_L g2935 ( 
.A(n_2475),
.B(n_366),
.Y(n_2935)
);

O2A1O1Ixp33_ASAP7_75t_L g2936 ( 
.A1(n_2379),
.A2(n_368),
.B(n_366),
.C(n_367),
.Y(n_2936)
);

AO32x2_ASAP7_75t_L g2937 ( 
.A1(n_2418),
.A2(n_369),
.A3(n_367),
.B1(n_368),
.B2(n_370),
.Y(n_2937)
);

NOR2xp33_ASAP7_75t_SL g2938 ( 
.A(n_2733),
.B(n_369),
.Y(n_2938)
);

NOR2xp33_ASAP7_75t_L g2939 ( 
.A(n_2542),
.B(n_370),
.Y(n_2939)
);

O2A1O1Ixp33_ASAP7_75t_L g2940 ( 
.A1(n_2414),
.A2(n_373),
.B(n_371),
.C(n_372),
.Y(n_2940)
);

BUFx2_ASAP7_75t_L g2941 ( 
.A(n_2388),
.Y(n_2941)
);

OR2x2_ASAP7_75t_L g2942 ( 
.A(n_2268),
.B(n_371),
.Y(n_2942)
);

A2O1A1Ixp33_ASAP7_75t_L g2943 ( 
.A1(n_2578),
.A2(n_375),
.B(n_373),
.C(n_374),
.Y(n_2943)
);

NAND2xp5_ASAP7_75t_SL g2944 ( 
.A(n_2540),
.B(n_680),
.Y(n_2944)
);

NOR2xp33_ASAP7_75t_R g2945 ( 
.A(n_2559),
.B(n_2671),
.Y(n_2945)
);

AOI21xp5_ASAP7_75t_L g2946 ( 
.A1(n_2581),
.A2(n_376),
.B(n_377),
.Y(n_2946)
);

O2A1O1Ixp33_ASAP7_75t_L g2947 ( 
.A1(n_2549),
.A2(n_379),
.B(n_377),
.C(n_378),
.Y(n_2947)
);

A2O1A1Ixp33_ASAP7_75t_L g2948 ( 
.A1(n_2592),
.A2(n_380),
.B(n_377),
.C(n_379),
.Y(n_2948)
);

NAND2xp5_ASAP7_75t_L g2949 ( 
.A(n_2478),
.B(n_379),
.Y(n_2949)
);

INVx1_ASAP7_75t_L g2950 ( 
.A(n_2306),
.Y(n_2950)
);

NOR2xp33_ASAP7_75t_L g2951 ( 
.A(n_2511),
.B(n_380),
.Y(n_2951)
);

NOR2xp67_ASAP7_75t_SL g2952 ( 
.A(n_2449),
.B(n_2339),
.Y(n_2952)
);

AOI21xp5_ASAP7_75t_L g2953 ( 
.A1(n_2598),
.A2(n_381),
.B(n_382),
.Y(n_2953)
);

NOR2x1_ASAP7_75t_L g2954 ( 
.A(n_2339),
.B(n_381),
.Y(n_2954)
);

NOR2xp33_ASAP7_75t_L g2955 ( 
.A(n_2249),
.B(n_381),
.Y(n_2955)
);

NAND2xp5_ASAP7_75t_SL g2956 ( 
.A(n_2467),
.B(n_682),
.Y(n_2956)
);

INVx2_ASAP7_75t_SL g2957 ( 
.A(n_2428),
.Y(n_2957)
);

INVx3_ASAP7_75t_L g2958 ( 
.A(n_2695),
.Y(n_2958)
);

AOI21xp5_ASAP7_75t_L g2959 ( 
.A1(n_2600),
.A2(n_382),
.B(n_383),
.Y(n_2959)
);

NOR2xp33_ASAP7_75t_L g2960 ( 
.A(n_2252),
.B(n_382),
.Y(n_2960)
);

O2A1O1Ixp33_ASAP7_75t_L g2961 ( 
.A1(n_2589),
.A2(n_387),
.B(n_384),
.C(n_386),
.Y(n_2961)
);

AOI21xp5_ASAP7_75t_L g2962 ( 
.A1(n_2602),
.A2(n_384),
.B(n_386),
.Y(n_2962)
);

AOI21xp5_ASAP7_75t_L g2963 ( 
.A1(n_2603),
.A2(n_384),
.B(n_386),
.Y(n_2963)
);

NOR2xp33_ASAP7_75t_L g2964 ( 
.A(n_2534),
.B(n_387),
.Y(n_2964)
);

NAND2xp5_ASAP7_75t_L g2965 ( 
.A(n_2636),
.B(n_387),
.Y(n_2965)
);

INVx2_ASAP7_75t_L g2966 ( 
.A(n_2332),
.Y(n_2966)
);

OR2x2_ASAP7_75t_L g2967 ( 
.A(n_2488),
.B(n_388),
.Y(n_2967)
);

INVx5_ASAP7_75t_L g2968 ( 
.A(n_2322),
.Y(n_2968)
);

INVx1_ASAP7_75t_L g2969 ( 
.A(n_2310),
.Y(n_2969)
);

INVxp67_ASAP7_75t_L g2970 ( 
.A(n_2582),
.Y(n_2970)
);

AOI21xp5_ASAP7_75t_L g2971 ( 
.A1(n_2609),
.A2(n_389),
.B(n_390),
.Y(n_2971)
);

INVx1_ASAP7_75t_L g2972 ( 
.A(n_2311),
.Y(n_2972)
);

INVx1_ASAP7_75t_L g2973 ( 
.A(n_2314),
.Y(n_2973)
);

CKINVDCx8_ASAP7_75t_R g2974 ( 
.A(n_2349),
.Y(n_2974)
);

INVx3_ASAP7_75t_SL g2975 ( 
.A(n_2304),
.Y(n_2975)
);

O2A1O1Ixp33_ASAP7_75t_L g2976 ( 
.A1(n_2596),
.A2(n_394),
.B(n_392),
.C(n_393),
.Y(n_2976)
);

HB1xp67_ASAP7_75t_L g2977 ( 
.A(n_2466),
.Y(n_2977)
);

INVxp67_ASAP7_75t_L g2978 ( 
.A(n_2615),
.Y(n_2978)
);

NOR3xp33_ASAP7_75t_L g2979 ( 
.A(n_2385),
.B(n_392),
.C(n_394),
.Y(n_2979)
);

A2O1A1Ixp33_ASAP7_75t_L g2980 ( 
.A1(n_2631),
.A2(n_396),
.B(n_394),
.C(n_395),
.Y(n_2980)
);

INVx4_ASAP7_75t_L g2981 ( 
.A(n_2406),
.Y(n_2981)
);

INVx2_ASAP7_75t_L g2982 ( 
.A(n_2436),
.Y(n_2982)
);

OR2x6_ASAP7_75t_L g2983 ( 
.A(n_2406),
.B(n_395),
.Y(n_2983)
);

AOI22xp33_ASAP7_75t_L g2984 ( 
.A1(n_2618),
.A2(n_399),
.B1(n_397),
.B2(n_398),
.Y(n_2984)
);

BUFx3_ASAP7_75t_L g2985 ( 
.A(n_2422),
.Y(n_2985)
);

AOI21xp33_ASAP7_75t_L g2986 ( 
.A1(n_2386),
.A2(n_399),
.B(n_400),
.Y(n_2986)
);

O2A1O1Ixp33_ASAP7_75t_L g2987 ( 
.A1(n_2628),
.A2(n_401),
.B(n_399),
.C(n_400),
.Y(n_2987)
);

O2A1O1Ixp33_ASAP7_75t_L g2988 ( 
.A1(n_2686),
.A2(n_402),
.B(n_400),
.C(n_401),
.Y(n_2988)
);

INVxp67_ASAP7_75t_L g2989 ( 
.A(n_2630),
.Y(n_2989)
);

NAND2xp5_ASAP7_75t_L g2990 ( 
.A(n_2721),
.B(n_401),
.Y(n_2990)
);

OAI22xp5_ASAP7_75t_L g2991 ( 
.A1(n_2551),
.A2(n_404),
.B1(n_402),
.B2(n_403),
.Y(n_2991)
);

NAND2xp5_ASAP7_75t_L g2992 ( 
.A(n_2364),
.B(n_402),
.Y(n_2992)
);

OAI22xp5_ASAP7_75t_L g2993 ( 
.A1(n_2555),
.A2(n_405),
.B1(n_403),
.B2(n_404),
.Y(n_2993)
);

OR2x6_ASAP7_75t_L g2994 ( 
.A(n_2728),
.B(n_405),
.Y(n_2994)
);

AND2x2_ASAP7_75t_SL g2995 ( 
.A(n_2484),
.B(n_405),
.Y(n_2995)
);

NAND3xp33_ASAP7_75t_L g2996 ( 
.A(n_2708),
.B(n_406),
.C(n_407),
.Y(n_2996)
);

A2O1A1Ixp33_ASAP7_75t_L g2997 ( 
.A1(n_2642),
.A2(n_408),
.B(n_406),
.C(n_407),
.Y(n_2997)
);

NOR3xp33_ASAP7_75t_SL g2998 ( 
.A(n_2696),
.B(n_408),
.C(n_409),
.Y(n_2998)
);

A2O1A1Ixp33_ASAP7_75t_L g2999 ( 
.A1(n_2646),
.A2(n_410),
.B(n_408),
.C(n_409),
.Y(n_2999)
);

NAND2xp5_ASAP7_75t_L g3000 ( 
.A(n_2391),
.B(n_410),
.Y(n_3000)
);

INVx2_ASAP7_75t_L g3001 ( 
.A(n_2564),
.Y(n_3001)
);

OR2x4_ASAP7_75t_L g3002 ( 
.A(n_2399),
.B(n_410),
.Y(n_3002)
);

A2O1A1Ixp33_ASAP7_75t_L g3003 ( 
.A1(n_2655),
.A2(n_413),
.B(n_411),
.C(n_412),
.Y(n_3003)
);

INVx2_ASAP7_75t_L g3004 ( 
.A(n_2591),
.Y(n_3004)
);

OR2x6_ASAP7_75t_L g3005 ( 
.A(n_2728),
.B(n_411),
.Y(n_3005)
);

O2A1O1Ixp33_ASAP7_75t_L g3006 ( 
.A1(n_2725),
.A2(n_415),
.B(n_413),
.C(n_414),
.Y(n_3006)
);

A2O1A1Ixp33_ASAP7_75t_L g3007 ( 
.A1(n_2665),
.A2(n_416),
.B(n_414),
.C(n_415),
.Y(n_3007)
);

OAI22xp5_ASAP7_75t_L g3008 ( 
.A1(n_2561),
.A2(n_418),
.B1(n_416),
.B2(n_417),
.Y(n_3008)
);

O2A1O1Ixp33_ASAP7_75t_SL g3009 ( 
.A1(n_2735),
.A2(n_418),
.B(n_416),
.C(n_417),
.Y(n_3009)
);

INVx2_ASAP7_75t_L g3010 ( 
.A(n_2612),
.Y(n_3010)
);

O2A1O1Ixp5_ASAP7_75t_L g3011 ( 
.A1(n_2557),
.A2(n_419),
.B(n_417),
.C(n_418),
.Y(n_3011)
);

O2A1O1Ixp33_ASAP7_75t_SL g3012 ( 
.A1(n_2355),
.A2(n_421),
.B(n_419),
.C(n_420),
.Y(n_3012)
);

AND2x4_ASAP7_75t_L g3013 ( 
.A(n_2513),
.B(n_420),
.Y(n_3013)
);

NAND2xp5_ASAP7_75t_L g3014 ( 
.A(n_2400),
.B(n_420),
.Y(n_3014)
);

INVx2_ASAP7_75t_L g3015 ( 
.A(n_2694),
.Y(n_3015)
);

HB1xp67_ASAP7_75t_L g3016 ( 
.A(n_2510),
.Y(n_3016)
);

INVx2_ASAP7_75t_SL g3017 ( 
.A(n_2409),
.Y(n_3017)
);

NAND2xp5_ASAP7_75t_L g3018 ( 
.A(n_2407),
.B(n_421),
.Y(n_3018)
);

O2A1O1Ixp33_ASAP7_75t_L g3019 ( 
.A1(n_2487),
.A2(n_423),
.B(n_421),
.C(n_422),
.Y(n_3019)
);

NOR2xp33_ASAP7_75t_L g3020 ( 
.A(n_2537),
.B(n_422),
.Y(n_3020)
);

INVx2_ASAP7_75t_L g3021 ( 
.A(n_2270),
.Y(n_3021)
);

AND2x2_ASAP7_75t_L g3022 ( 
.A(n_2634),
.B(n_423),
.Y(n_3022)
);

NOR2xp67_ASAP7_75t_SL g3023 ( 
.A(n_2410),
.B(n_424),
.Y(n_3023)
);

BUFx2_ASAP7_75t_L g3024 ( 
.A(n_2322),
.Y(n_3024)
);

OAI21xp5_ASAP7_75t_L g3025 ( 
.A1(n_2413),
.A2(n_424),
.B(n_425),
.Y(n_3025)
);

INVx4_ASAP7_75t_L g3026 ( 
.A(n_2322),
.Y(n_3026)
);

OAI21xp33_ASAP7_75t_L g3027 ( 
.A1(n_2541),
.A2(n_425),
.B(n_426),
.Y(n_3027)
);

BUFx12f_ASAP7_75t_L g3028 ( 
.A(n_2368),
.Y(n_3028)
);

NAND2xp5_ASAP7_75t_SL g3029 ( 
.A(n_2318),
.B(n_683),
.Y(n_3029)
);

O2A1O1Ixp5_ASAP7_75t_L g3030 ( 
.A1(n_2568),
.A2(n_428),
.B(n_425),
.C(n_426),
.Y(n_3030)
);

NOR2xp33_ASAP7_75t_L g3031 ( 
.A(n_2419),
.B(n_426),
.Y(n_3031)
);

NOR2xp33_ASAP7_75t_L g3032 ( 
.A(n_2648),
.B(n_428),
.Y(n_3032)
);

CKINVDCx14_ASAP7_75t_R g3033 ( 
.A(n_2483),
.Y(n_3033)
);

NAND2xp5_ASAP7_75t_L g3034 ( 
.A(n_2417),
.B(n_429),
.Y(n_3034)
);

NOR2xp33_ASAP7_75t_L g3035 ( 
.A(n_2657),
.B(n_429),
.Y(n_3035)
);

O2A1O1Ixp33_ASAP7_75t_L g3036 ( 
.A1(n_2378),
.A2(n_431),
.B(n_429),
.C(n_430),
.Y(n_3036)
);

INVx3_ASAP7_75t_L g3037 ( 
.A(n_2329),
.Y(n_3037)
);

INVx1_ASAP7_75t_L g3038 ( 
.A(n_2317),
.Y(n_3038)
);

AOI22xp33_ASAP7_75t_SL g3039 ( 
.A1(n_2368),
.A2(n_434),
.B1(n_432),
.B2(n_433),
.Y(n_3039)
);

OAI22xp5_ASAP7_75t_L g3040 ( 
.A1(n_2566),
.A2(n_434),
.B1(n_432),
.B2(n_433),
.Y(n_3040)
);

NAND2xp5_ASAP7_75t_L g3041 ( 
.A(n_2421),
.B(n_434),
.Y(n_3041)
);

OAI22xp5_ASAP7_75t_L g3042 ( 
.A1(n_2567),
.A2(n_437),
.B1(n_435),
.B2(n_436),
.Y(n_3042)
);

INVx2_ASAP7_75t_L g3043 ( 
.A(n_2485),
.Y(n_3043)
);

AOI21xp5_ASAP7_75t_L g3044 ( 
.A1(n_2684),
.A2(n_437),
.B(n_438),
.Y(n_3044)
);

HB1xp67_ASAP7_75t_L g3045 ( 
.A(n_2560),
.Y(n_3045)
);

INVx2_ASAP7_75t_SL g3046 ( 
.A(n_2530),
.Y(n_3046)
);

O2A1O1Ixp33_ASAP7_75t_L g3047 ( 
.A1(n_2470),
.A2(n_439),
.B(n_437),
.C(n_438),
.Y(n_3047)
);

AOI21x1_ASAP7_75t_L g3048 ( 
.A1(n_2309),
.A2(n_438),
.B(n_440),
.Y(n_3048)
);

AOI21x1_ASAP7_75t_L g3049 ( 
.A1(n_2570),
.A2(n_440),
.B(n_441),
.Y(n_3049)
);

NAND2xp5_ASAP7_75t_SL g3050 ( 
.A(n_2558),
.B(n_683),
.Y(n_3050)
);

AOI21xp5_ASAP7_75t_L g3051 ( 
.A1(n_2690),
.A2(n_440),
.B(n_441),
.Y(n_3051)
);

NAND2xp5_ASAP7_75t_SL g3052 ( 
.A(n_2653),
.B(n_684),
.Y(n_3052)
);

NAND2xp5_ASAP7_75t_SL g3053 ( 
.A(n_2719),
.B(n_684),
.Y(n_3053)
);

OAI22x1_ASAP7_75t_L g3054 ( 
.A1(n_2356),
.A2(n_443),
.B1(n_441),
.B2(n_442),
.Y(n_3054)
);

NAND2xp5_ASAP7_75t_SL g3055 ( 
.A(n_2269),
.B(n_685),
.Y(n_3055)
);

INVx1_ASAP7_75t_L g3056 ( 
.A(n_2423),
.Y(n_3056)
);

NOR3xp33_ASAP7_75t_SL g3057 ( 
.A(n_2494),
.B(n_442),
.C(n_443),
.Y(n_3057)
);

A2O1A1Ixp33_ASAP7_75t_L g3058 ( 
.A1(n_2700),
.A2(n_444),
.B(n_442),
.C(n_443),
.Y(n_3058)
);

INVx1_ASAP7_75t_L g3059 ( 
.A(n_2425),
.Y(n_3059)
);

NOR2xp33_ASAP7_75t_L g3060 ( 
.A(n_2667),
.B(n_444),
.Y(n_3060)
);

AOI22xp5_ASAP7_75t_L g3061 ( 
.A1(n_2669),
.A2(n_447),
.B1(n_445),
.B2(n_446),
.Y(n_3061)
);

NAND2xp5_ASAP7_75t_L g3062 ( 
.A(n_2278),
.B(n_445),
.Y(n_3062)
);

AOI21xp5_ASAP7_75t_L g3063 ( 
.A1(n_2702),
.A2(n_447),
.B(n_448),
.Y(n_3063)
);

INVx1_ASAP7_75t_L g3064 ( 
.A(n_2430),
.Y(n_3064)
);

HB1xp67_ASAP7_75t_L g3065 ( 
.A(n_2577),
.Y(n_3065)
);

O2A1O1Ixp33_ASAP7_75t_L g3066 ( 
.A1(n_2463),
.A2(n_450),
.B(n_448),
.C(n_449),
.Y(n_3066)
);

NAND2xp5_ASAP7_75t_L g3067 ( 
.A(n_2340),
.B(n_449),
.Y(n_3067)
);

INVx1_ASAP7_75t_L g3068 ( 
.A(n_2472),
.Y(n_3068)
);

BUFx6f_ASAP7_75t_L g3069 ( 
.A(n_2416),
.Y(n_3069)
);

INVx1_ASAP7_75t_L g3070 ( 
.A(n_2474),
.Y(n_3070)
);

A2O1A1Ixp33_ASAP7_75t_L g3071 ( 
.A1(n_2718),
.A2(n_452),
.B(n_450),
.C(n_451),
.Y(n_3071)
);

AOI22xp33_ASAP7_75t_L g3072 ( 
.A1(n_2676),
.A2(n_454),
.B1(n_452),
.B2(n_453),
.Y(n_3072)
);

AOI21x1_ASAP7_75t_L g3073 ( 
.A1(n_2575),
.A2(n_452),
.B(n_453),
.Y(n_3073)
);

INVx1_ASAP7_75t_L g3074 ( 
.A(n_2476),
.Y(n_3074)
);

BUFx2_ASAP7_75t_SL g3075 ( 
.A(n_2329),
.Y(n_3075)
);

OAI22xp5_ASAP7_75t_L g3076 ( 
.A1(n_2583),
.A2(n_455),
.B1(n_453),
.B2(n_454),
.Y(n_3076)
);

INVx1_ASAP7_75t_L g3077 ( 
.A(n_2477),
.Y(n_3077)
);

OAI22xp5_ASAP7_75t_L g3078 ( 
.A1(n_2584),
.A2(n_456),
.B1(n_454),
.B2(n_455),
.Y(n_3078)
);

NAND3xp33_ASAP7_75t_L g3079 ( 
.A(n_2288),
.B(n_455),
.C(n_456),
.Y(n_3079)
);

AOI21xp5_ASAP7_75t_L g3080 ( 
.A1(n_2316),
.A2(n_456),
.B(n_457),
.Y(n_3080)
);

INVx1_ASAP7_75t_L g3081 ( 
.A(n_2479),
.Y(n_3081)
);

AOI21xp5_ASAP7_75t_L g3082 ( 
.A1(n_2320),
.A2(n_458),
.B(n_459),
.Y(n_3082)
);

AOI22xp5_ASAP7_75t_L g3083 ( 
.A1(n_2687),
.A2(n_460),
.B1(n_458),
.B2(n_459),
.Y(n_3083)
);

O2A1O1Ixp5_ASAP7_75t_L g3084 ( 
.A1(n_2610),
.A2(n_462),
.B(n_460),
.C(n_461),
.Y(n_3084)
);

INVx1_ASAP7_75t_SL g3085 ( 
.A(n_2497),
.Y(n_3085)
);

OAI22xp5_ASAP7_75t_L g3086 ( 
.A1(n_2585),
.A2(n_462),
.B1(n_460),
.B2(n_461),
.Y(n_3086)
);

NOR2xp67_ASAP7_75t_L g3087 ( 
.A(n_2704),
.B(n_462),
.Y(n_3087)
);

NAND2xp5_ASAP7_75t_L g3088 ( 
.A(n_2344),
.B(n_463),
.Y(n_3088)
);

AOI21xp5_ASAP7_75t_L g3089 ( 
.A1(n_2321),
.A2(n_463),
.B(n_464),
.Y(n_3089)
);

INVx1_ASAP7_75t_L g3090 ( 
.A(n_2283),
.Y(n_3090)
);

NOR3xp33_ASAP7_75t_SL g3091 ( 
.A(n_2509),
.B(n_463),
.C(n_464),
.Y(n_3091)
);

NOR2xp33_ASAP7_75t_L g3092 ( 
.A(n_2709),
.B(n_464),
.Y(n_3092)
);

NAND2xp5_ASAP7_75t_L g3093 ( 
.A(n_2354),
.B(n_465),
.Y(n_3093)
);

HB1xp67_ASAP7_75t_L g3094 ( 
.A(n_2594),
.Y(n_3094)
);

BUFx2_ASAP7_75t_L g3095 ( 
.A(n_2486),
.Y(n_3095)
);

NOR2xp33_ASAP7_75t_L g3096 ( 
.A(n_2536),
.B(n_465),
.Y(n_3096)
);

INVx4_ASAP7_75t_L g3097 ( 
.A(n_2416),
.Y(n_3097)
);

NAND2xp5_ASAP7_75t_L g3098 ( 
.A(n_2338),
.B(n_465),
.Y(n_3098)
);

INVx2_ASAP7_75t_L g3099 ( 
.A(n_2518),
.Y(n_3099)
);

AND2x4_ASAP7_75t_L g3100 ( 
.A(n_2512),
.B(n_466),
.Y(n_3100)
);

AOI22xp33_ASAP7_75t_L g3101 ( 
.A1(n_2387),
.A2(n_469),
.B1(n_467),
.B2(n_468),
.Y(n_3101)
);

INVx3_ASAP7_75t_L g3102 ( 
.A(n_2445),
.Y(n_3102)
);

NOR3xp33_ASAP7_75t_SL g3103 ( 
.A(n_2520),
.B(n_467),
.C(n_468),
.Y(n_3103)
);

INVx1_ASAP7_75t_L g3104 ( 
.A(n_2284),
.Y(n_3104)
);

BUFx12f_ASAP7_75t_L g3105 ( 
.A(n_2532),
.Y(n_3105)
);

CKINVDCx20_ASAP7_75t_R g3106 ( 
.A(n_2411),
.Y(n_3106)
);

NAND2xp5_ASAP7_75t_SL g3107 ( 
.A(n_2269),
.B(n_685),
.Y(n_3107)
);

A2O1A1Ixp33_ASAP7_75t_L g3108 ( 
.A1(n_2377),
.A2(n_470),
.B(n_468),
.C(n_469),
.Y(n_3108)
);

NOR2xp33_ASAP7_75t_L g3109 ( 
.A(n_2525),
.B(n_470),
.Y(n_3109)
);

AO32x2_ASAP7_75t_L g3110 ( 
.A1(n_2633),
.A2(n_472),
.A3(n_470),
.B1(n_471),
.B2(n_473),
.Y(n_3110)
);

AND2x4_ASAP7_75t_L g3111 ( 
.A(n_2264),
.B(n_471),
.Y(n_3111)
);

OAI22xp5_ASAP7_75t_L g3112 ( 
.A1(n_2586),
.A2(n_473),
.B1(n_471),
.B2(n_472),
.Y(n_3112)
);

BUFx6f_ASAP7_75t_L g3113 ( 
.A(n_2445),
.Y(n_3113)
);

A2O1A1Ixp33_ASAP7_75t_L g3114 ( 
.A1(n_2382),
.A2(n_475),
.B(n_473),
.C(n_474),
.Y(n_3114)
);

AND2x2_ASAP7_75t_L g3115 ( 
.A(n_2359),
.B(n_474),
.Y(n_3115)
);

A2O1A1Ixp33_ASAP7_75t_L g3116 ( 
.A1(n_2397),
.A2(n_476),
.B(n_474),
.C(n_475),
.Y(n_3116)
);

NOR2x1p5_ASAP7_75t_L g3117 ( 
.A(n_2531),
.B(n_475),
.Y(n_3117)
);

BUFx2_ASAP7_75t_L g3118 ( 
.A(n_2264),
.Y(n_3118)
);

BUFx2_ASAP7_75t_L g3119 ( 
.A(n_2271),
.Y(n_3119)
);

NAND2xp5_ASAP7_75t_L g3120 ( 
.A(n_2593),
.B(n_476),
.Y(n_3120)
);

OR2x6_ASAP7_75t_L g3121 ( 
.A(n_2606),
.B(n_477),
.Y(n_3121)
);

INVx2_ASAP7_75t_L g3122 ( 
.A(n_2464),
.Y(n_3122)
);

HB1xp67_ASAP7_75t_L g3123 ( 
.A(n_2635),
.Y(n_3123)
);

INVx3_ASAP7_75t_L g3124 ( 
.A(n_2445),
.Y(n_3124)
);

O2A1O1Ixp33_ASAP7_75t_L g3125 ( 
.A1(n_2639),
.A2(n_481),
.B(n_479),
.C(n_480),
.Y(n_3125)
);

NAND2xp5_ASAP7_75t_SL g3126 ( 
.A(n_2649),
.B(n_686),
.Y(n_3126)
);

BUFx12f_ASAP7_75t_L g3127 ( 
.A(n_2532),
.Y(n_3127)
);

OAI22xp5_ASAP7_75t_L g3128 ( 
.A1(n_2601),
.A2(n_481),
.B1(n_479),
.B2(n_480),
.Y(n_3128)
);

AOI22xp5_ASAP7_75t_L g3129 ( 
.A1(n_2362),
.A2(n_481),
.B1(n_479),
.B2(n_480),
.Y(n_3129)
);

NAND2xp5_ASAP7_75t_SL g3130 ( 
.A(n_2649),
.B(n_686),
.Y(n_3130)
);

OAI22xp5_ASAP7_75t_L g3131 ( 
.A1(n_2607),
.A2(n_485),
.B1(n_483),
.B2(n_484),
.Y(n_3131)
);

CKINVDCx5p33_ASAP7_75t_R g3132 ( 
.A(n_2366),
.Y(n_3132)
);

INVx6_ASAP7_75t_L g3133 ( 
.A(n_2532),
.Y(n_3133)
);

AOI22xp5_ASAP7_75t_L g3134 ( 
.A1(n_2641),
.A2(n_485),
.B1(n_483),
.B2(n_484),
.Y(n_3134)
);

INVx2_ASAP7_75t_L g3135 ( 
.A(n_2469),
.Y(n_3135)
);

INVx2_ASAP7_75t_L g3136 ( 
.A(n_2480),
.Y(n_3136)
);

BUFx2_ASAP7_75t_L g3137 ( 
.A(n_2271),
.Y(n_3137)
);

OR2x6_ASAP7_75t_L g3138 ( 
.A(n_2302),
.B(n_486),
.Y(n_3138)
);

OAI21xp33_ASAP7_75t_L g3139 ( 
.A1(n_2251),
.A2(n_486),
.B(n_487),
.Y(n_3139)
);

A2O1A1Ixp33_ASAP7_75t_L g3140 ( 
.A1(n_2398),
.A2(n_2573),
.B(n_2588),
.C(n_2563),
.Y(n_3140)
);

NAND2xp5_ASAP7_75t_L g3141 ( 
.A(n_2737),
.B(n_486),
.Y(n_3141)
);

AO22x1_ASAP7_75t_L g3142 ( 
.A1(n_2434),
.A2(n_489),
.B1(n_487),
.B2(n_488),
.Y(n_3142)
);

O2A1O1Ixp5_ASAP7_75t_L g3143 ( 
.A1(n_2608),
.A2(n_2714),
.B(n_2716),
.C(n_2713),
.Y(n_3143)
);

NAND2xp5_ASAP7_75t_L g3144 ( 
.A(n_2613),
.B(n_2619),
.Y(n_3144)
);

AOI21xp5_ASAP7_75t_L g3145 ( 
.A1(n_2433),
.A2(n_488),
.B(n_489),
.Y(n_3145)
);

NOR2xp33_ASAP7_75t_SL g3146 ( 
.A(n_2302),
.B(n_488),
.Y(n_3146)
);

A2O1A1Ixp33_ASAP7_75t_L g3147 ( 
.A1(n_2647),
.A2(n_491),
.B(n_489),
.C(n_490),
.Y(n_3147)
);

NAND2xp5_ASAP7_75t_L g3148 ( 
.A(n_2623),
.B(n_490),
.Y(n_3148)
);

O2A1O1Ixp5_ASAP7_75t_L g3149 ( 
.A1(n_2627),
.A2(n_493),
.B(n_491),
.C(n_492),
.Y(n_3149)
);

OAI21xp5_ASAP7_75t_L g3150 ( 
.A1(n_2440),
.A2(n_2275),
.B(n_2637),
.Y(n_3150)
);

NOR2xp33_ASAP7_75t_L g3151 ( 
.A(n_2515),
.B(n_492),
.Y(n_3151)
);

BUFx10_ASAP7_75t_L g3152 ( 
.A(n_2854),
.Y(n_3152)
);

AO31x2_ASAP7_75t_L g3153 ( 
.A1(n_2966),
.A2(n_2401),
.A3(n_2505),
.B(n_2498),
.Y(n_3153)
);

BUFx12f_ASAP7_75t_L g3154 ( 
.A(n_2779),
.Y(n_3154)
);

OAI22xp5_ASAP7_75t_L g3155 ( 
.A1(n_2850),
.A2(n_2453),
.B1(n_2369),
.B2(n_2620),
.Y(n_3155)
);

OA21x2_ASAP7_75t_L g3156 ( 
.A1(n_3001),
.A2(n_3010),
.B(n_3004),
.Y(n_3156)
);

OR2x2_ASAP7_75t_L g3157 ( 
.A(n_2873),
.B(n_2638),
.Y(n_3157)
);

AO31x2_ASAP7_75t_L g3158 ( 
.A1(n_3015),
.A2(n_2645),
.A3(n_2651),
.B(n_2640),
.Y(n_3158)
);

NAND2xp5_ASAP7_75t_L g3159 ( 
.A(n_2805),
.B(n_2679),
.Y(n_3159)
);

OAI21x1_ASAP7_75t_SL g3160 ( 
.A1(n_3026),
.A2(n_2447),
.B(n_2360),
.Y(n_3160)
);

OAI21xp5_ASAP7_75t_L g3161 ( 
.A1(n_3143),
.A2(n_2453),
.B(n_2538),
.Y(n_3161)
);

INVx1_ASAP7_75t_L g3162 ( 
.A(n_2763),
.Y(n_3162)
);

BUFx2_ASAP7_75t_L g3163 ( 
.A(n_2945),
.Y(n_3163)
);

INVx2_ASAP7_75t_L g3164 ( 
.A(n_2773),
.Y(n_3164)
);

BUFx3_ASAP7_75t_L g3165 ( 
.A(n_2854),
.Y(n_3165)
);

O2A1O1Ixp33_ASAP7_75t_L g3166 ( 
.A1(n_2837),
.A2(n_2346),
.B(n_2341),
.C(n_2643),
.Y(n_3166)
);

AOI22xp5_ASAP7_75t_L g3167 ( 
.A1(n_2995),
.A2(n_2656),
.B1(n_2699),
.B2(n_2689),
.Y(n_3167)
);

INVx2_ASAP7_75t_L g3168 ( 
.A(n_2794),
.Y(n_3168)
);

AOI21xp5_ASAP7_75t_L g3169 ( 
.A1(n_2883),
.A2(n_2724),
.B(n_2660),
.Y(n_3169)
);

OR2x6_ASAP7_75t_L g3170 ( 
.A(n_2781),
.B(n_2523),
.Y(n_3170)
);

AOI21x1_ASAP7_75t_L g3171 ( 
.A1(n_2909),
.A2(n_2672),
.B(n_2654),
.Y(n_3171)
);

AO31x2_ASAP7_75t_L g3172 ( 
.A1(n_2982),
.A2(n_2675),
.A3(n_2681),
.B(n_2673),
.Y(n_3172)
);

NOR2xp33_ASAP7_75t_L g3173 ( 
.A(n_2974),
.B(n_2535),
.Y(n_3173)
);

NAND3xp33_ASAP7_75t_SL g3174 ( 
.A(n_2784),
.B(n_2738),
.C(n_2817),
.Y(n_3174)
);

OAI21x1_ASAP7_75t_L g3175 ( 
.A1(n_3021),
.A2(n_2924),
.B(n_3048),
.Y(n_3175)
);

CKINVDCx20_ASAP7_75t_R g3176 ( 
.A(n_2768),
.Y(n_3176)
);

INVx2_ASAP7_75t_L g3177 ( 
.A(n_2819),
.Y(n_3177)
);

OAI21xp5_ASAP7_75t_L g3178 ( 
.A1(n_3140),
.A2(n_2420),
.B(n_2492),
.Y(n_3178)
);

HB1xp67_ASAP7_75t_L g3179 ( 
.A(n_2778),
.Y(n_3179)
);

OAI21xp5_ASAP7_75t_L g3180 ( 
.A1(n_2769),
.A2(n_2324),
.B(n_2404),
.Y(n_3180)
);

BUFx6f_ASAP7_75t_L g3181 ( 
.A(n_2843),
.Y(n_3181)
);

AOI21xp5_ASAP7_75t_L g3182 ( 
.A1(n_2834),
.A2(n_2693),
.B(n_2688),
.Y(n_3182)
);

AOI221xp5_ASAP7_75t_L g3183 ( 
.A1(n_2921),
.A2(n_2351),
.B1(n_2380),
.B2(n_2678),
.C(n_2670),
.Y(n_3183)
);

BUFx2_ASAP7_75t_L g3184 ( 
.A(n_3028),
.Y(n_3184)
);

AO31x2_ASAP7_75t_L g3185 ( 
.A1(n_2757),
.A2(n_2707),
.A3(n_2732),
.B(n_2720),
.Y(n_3185)
);

AND2x2_ASAP7_75t_L g3186 ( 
.A(n_2871),
.B(n_2331),
.Y(n_3186)
);

INVx1_ASAP7_75t_L g3187 ( 
.A(n_2872),
.Y(n_3187)
);

AOI221x1_ASAP7_75t_L g3188 ( 
.A1(n_2899),
.A2(n_2758),
.B1(n_3027),
.B2(n_3139),
.C(n_3054),
.Y(n_3188)
);

BUFx10_ASAP7_75t_L g3189 ( 
.A(n_2876),
.Y(n_3189)
);

AOI21xp5_ASAP7_75t_L g3190 ( 
.A1(n_3150),
.A2(n_2455),
.B(n_2451),
.Y(n_3190)
);

AOI21xp5_ASAP7_75t_L g3191 ( 
.A1(n_3144),
.A2(n_2459),
.B(n_2250),
.Y(n_3191)
);

OAI21x1_ASAP7_75t_L g3192 ( 
.A1(n_2777),
.A2(n_2625),
.B(n_2545),
.Y(n_3192)
);

AOI22xp5_ASAP7_75t_L g3193 ( 
.A1(n_2751),
.A2(n_2502),
.B1(n_2499),
.B2(n_2402),
.Y(n_3193)
);

OAI22xp5_ASAP7_75t_L g3194 ( 
.A1(n_2994),
.A2(n_2659),
.B1(n_2443),
.B2(n_2438),
.Y(n_3194)
);

AND2x4_ASAP7_75t_L g3195 ( 
.A(n_2894),
.B(n_2456),
.Y(n_3195)
);

INVx1_ASAP7_75t_L g3196 ( 
.A(n_2886),
.Y(n_3196)
);

NOR2xp33_ASAP7_75t_L g3197 ( 
.A(n_2746),
.B(n_2507),
.Y(n_3197)
);

NOR2xp33_ASAP7_75t_L g3198 ( 
.A(n_2975),
.B(n_3132),
.Y(n_3198)
);

INVx2_ASAP7_75t_L g3199 ( 
.A(n_2825),
.Y(n_3199)
);

AO31x2_ASAP7_75t_L g3200 ( 
.A1(n_2841),
.A2(n_2448),
.A3(n_2405),
.B(n_2491),
.Y(n_3200)
);

INVx3_ASAP7_75t_SL g3201 ( 
.A(n_2766),
.Y(n_3201)
);

AND2x2_ASAP7_75t_L g3202 ( 
.A(n_2851),
.B(n_2893),
.Y(n_3202)
);

AOI221x1_ASAP7_75t_L g3203 ( 
.A1(n_2808),
.A2(n_2519),
.B1(n_2574),
.B2(n_2599),
.C(n_2562),
.Y(n_3203)
);

AOI21xp5_ASAP7_75t_L g3204 ( 
.A1(n_2878),
.A2(n_2629),
.B(n_2626),
.Y(n_3204)
);

O2A1O1Ixp33_ASAP7_75t_SL g3205 ( 
.A1(n_2815),
.A2(n_2622),
.B(n_2652),
.C(n_2605),
.Y(n_3205)
);

AOI221x1_ASAP7_75t_L g3206 ( 
.A1(n_2764),
.A2(n_2710),
.B1(n_2697),
.B2(n_2677),
.C(n_2504),
.Y(n_3206)
);

OAI21x1_ASAP7_75t_L g3207 ( 
.A1(n_3102),
.A2(n_2625),
.B(n_2545),
.Y(n_3207)
);

A2O1A1Ixp33_ASAP7_75t_L g3208 ( 
.A1(n_2828),
.A2(n_2682),
.B(n_2715),
.C(n_2337),
.Y(n_3208)
);

AO21x1_ASAP7_75t_L g3209 ( 
.A1(n_3146),
.A2(n_2517),
.B(n_2441),
.Y(n_3209)
);

OAI221xp5_ASAP7_75t_L g3210 ( 
.A1(n_2970),
.A2(n_2978),
.B1(n_2989),
.B2(n_2979),
.C(n_3057),
.Y(n_3210)
);

OAI21xp5_ASAP7_75t_L g3211 ( 
.A1(n_2996),
.A2(n_2461),
.B(n_2437),
.Y(n_3211)
);

AO21x2_ASAP7_75t_L g3212 ( 
.A1(n_2869),
.A2(n_2506),
.B(n_2524),
.Y(n_3212)
);

BUFx4_ASAP7_75t_R g3213 ( 
.A(n_2767),
.Y(n_3213)
);

BUFx6f_ASAP7_75t_L g3214 ( 
.A(n_2894),
.Y(n_3214)
);

OAI21x1_ASAP7_75t_L g3215 ( 
.A1(n_3102),
.A2(n_2664),
.B(n_2644),
.Y(n_3215)
);

OAI21x1_ASAP7_75t_L g3216 ( 
.A1(n_3124),
.A2(n_2664),
.B(n_2644),
.Y(n_3216)
);

BUFx4f_ASAP7_75t_SL g3217 ( 
.A(n_2884),
.Y(n_3217)
);

OAI21xp5_ASAP7_75t_L g3218 ( 
.A1(n_2932),
.A2(n_2444),
.B(n_2426),
.Y(n_3218)
);

INVx2_ASAP7_75t_L g3219 ( 
.A(n_2856),
.Y(n_3219)
);

INVxp67_ASAP7_75t_SL g3220 ( 
.A(n_2910),
.Y(n_3220)
);

AOI22xp5_ASAP7_75t_L g3221 ( 
.A1(n_2835),
.A2(n_2290),
.B1(n_2508),
.B2(n_2328),
.Y(n_3221)
);

OAI22xp5_ASAP7_75t_L g3222 ( 
.A1(n_2994),
.A2(n_2279),
.B1(n_2500),
.B2(n_2503),
.Y(n_3222)
);

AOI21xp5_ASAP7_75t_L g3223 ( 
.A1(n_2885),
.A2(n_2326),
.B(n_2265),
.Y(n_3223)
);

OAI21xp5_ASAP7_75t_L g3224 ( 
.A1(n_2925),
.A2(n_2490),
.B(n_2412),
.Y(n_3224)
);

INVx3_ASAP7_75t_L g3225 ( 
.A(n_2981),
.Y(n_3225)
);

OA21x2_ASAP7_75t_L g3226 ( 
.A1(n_2755),
.A2(n_2427),
.B(n_2333),
.Y(n_3226)
);

NAND2xp5_ASAP7_75t_L g3227 ( 
.A(n_2770),
.B(n_2333),
.Y(n_3227)
);

AOI21xp5_ASAP7_75t_L g3228 ( 
.A1(n_2901),
.A2(n_2446),
.B(n_2734),
.Y(n_3228)
);

AOI221xp5_ASAP7_75t_L g3229 ( 
.A1(n_2789),
.A2(n_2446),
.B1(n_2734),
.B2(n_496),
.C(n_494),
.Y(n_3229)
);

BUFx6f_ASAP7_75t_L g3230 ( 
.A(n_2889),
.Y(n_3230)
);

INVx2_ASAP7_75t_SL g3231 ( 
.A(n_2898),
.Y(n_3231)
);

A2O1A1Ixp33_ASAP7_75t_L g3232 ( 
.A1(n_2887),
.A2(n_498),
.B(n_495),
.C(n_496),
.Y(n_3232)
);

A2O1A1Ixp33_ASAP7_75t_L g3233 ( 
.A1(n_2820),
.A2(n_499),
.B(n_495),
.C(n_498),
.Y(n_3233)
);

AOI221x1_ASAP7_75t_L g3234 ( 
.A1(n_2798),
.A2(n_500),
.B1(n_495),
.B2(n_499),
.C(n_501),
.Y(n_3234)
);

AOI21xp5_ASAP7_75t_L g3235 ( 
.A1(n_2742),
.A2(n_499),
.B(n_500),
.Y(n_3235)
);

OAI21x1_ASAP7_75t_L g3236 ( 
.A1(n_2879),
.A2(n_503),
.B(n_502),
.Y(n_3236)
);

BUFx10_ASAP7_75t_L g3237 ( 
.A(n_2752),
.Y(n_3237)
);

AO31x2_ASAP7_75t_L g3238 ( 
.A1(n_2749),
.A2(n_503),
.A3(n_500),
.B(n_502),
.Y(n_3238)
);

AOI21xp5_ASAP7_75t_L g3239 ( 
.A1(n_3068),
.A2(n_502),
.B(n_504),
.Y(n_3239)
);

AND2x2_ASAP7_75t_L g3240 ( 
.A(n_2897),
.B(n_504),
.Y(n_3240)
);

O2A1O1Ixp33_ASAP7_75t_L g3241 ( 
.A1(n_3147),
.A2(n_506),
.B(n_504),
.C(n_505),
.Y(n_3241)
);

A2O1A1Ixp33_ASAP7_75t_L g3242 ( 
.A1(n_2947),
.A2(n_508),
.B(n_505),
.C(n_507),
.Y(n_3242)
);

AO31x2_ASAP7_75t_L g3243 ( 
.A1(n_2754),
.A2(n_508),
.A3(n_505),
.B(n_507),
.Y(n_3243)
);

NOR2xp33_ASAP7_75t_L g3244 ( 
.A(n_3002),
.B(n_507),
.Y(n_3244)
);

INVx5_ASAP7_75t_L g3245 ( 
.A(n_2781),
.Y(n_3245)
);

NOR2xp33_ASAP7_75t_L g3246 ( 
.A(n_2934),
.B(n_508),
.Y(n_3246)
);

AOI221xp5_ASAP7_75t_L g3247 ( 
.A1(n_2861),
.A2(n_511),
.B1(n_509),
.B2(n_510),
.C(n_512),
.Y(n_3247)
);

AND2x4_ASAP7_75t_L g3248 ( 
.A(n_2902),
.B(n_509),
.Y(n_3248)
);

NOR2xp67_ASAP7_75t_SL g3249 ( 
.A(n_2968),
.B(n_509),
.Y(n_3249)
);

NAND3xp33_ASAP7_75t_SL g3250 ( 
.A(n_2900),
.B(n_510),
.C(n_511),
.Y(n_3250)
);

AO31x2_ASAP7_75t_L g3251 ( 
.A1(n_2753),
.A2(n_2756),
.A3(n_2829),
.B(n_2818),
.Y(n_3251)
);

AND2x2_ASAP7_75t_L g3252 ( 
.A(n_2907),
.B(n_510),
.Y(n_3252)
);

HB1xp67_ASAP7_75t_L g3253 ( 
.A(n_2775),
.Y(n_3253)
);

OAI21x1_ASAP7_75t_L g3254 ( 
.A1(n_3049),
.A2(n_514),
.B(n_513),
.Y(n_3254)
);

OAI21x1_ASAP7_75t_L g3255 ( 
.A1(n_3073),
.A2(n_514),
.B(n_513),
.Y(n_3255)
);

NAND2xp5_ASAP7_75t_L g3256 ( 
.A(n_2923),
.B(n_512),
.Y(n_3256)
);

A2O1A1Ixp33_ASAP7_75t_L g3257 ( 
.A1(n_2961),
.A2(n_515),
.B(n_513),
.C(n_514),
.Y(n_3257)
);

CKINVDCx20_ASAP7_75t_R g3258 ( 
.A(n_2792),
.Y(n_3258)
);

A2O1A1Ixp33_ASAP7_75t_L g3259 ( 
.A1(n_2976),
.A2(n_517),
.B(n_515),
.C(n_516),
.Y(n_3259)
);

AOI21x1_ASAP7_75t_SL g3260 ( 
.A1(n_3062),
.A2(n_516),
.B(n_517),
.Y(n_3260)
);

OAI21x1_ASAP7_75t_L g3261 ( 
.A1(n_3037),
.A2(n_520),
.B(n_519),
.Y(n_3261)
);

AO31x2_ASAP7_75t_L g3262 ( 
.A1(n_2844),
.A2(n_520),
.A3(n_518),
.B(n_519),
.Y(n_3262)
);

AO31x2_ASAP7_75t_L g3263 ( 
.A1(n_2865),
.A2(n_522),
.A3(n_519),
.B(n_521),
.Y(n_3263)
);

A2O1A1Ixp33_ASAP7_75t_L g3264 ( 
.A1(n_2987),
.A2(n_524),
.B(n_522),
.C(n_523),
.Y(n_3264)
);

INVx6_ASAP7_75t_SL g3265 ( 
.A(n_2752),
.Y(n_3265)
);

CKINVDCx5p33_ASAP7_75t_R g3266 ( 
.A(n_3033),
.Y(n_3266)
);

INVx1_ASAP7_75t_L g3267 ( 
.A(n_2759),
.Y(n_3267)
);

BUFx2_ASAP7_75t_L g3268 ( 
.A(n_2896),
.Y(n_3268)
);

NAND2xp5_ASAP7_75t_SL g3269 ( 
.A(n_2968),
.B(n_523),
.Y(n_3269)
);

O2A1O1Ixp33_ASAP7_75t_L g3270 ( 
.A1(n_2797),
.A2(n_525),
.B(n_523),
.C(n_524),
.Y(n_3270)
);

AOI21xp5_ASAP7_75t_L g3271 ( 
.A1(n_3070),
.A2(n_3077),
.B(n_3074),
.Y(n_3271)
);

AOI21xp5_ASAP7_75t_L g3272 ( 
.A1(n_3081),
.A2(n_525),
.B(n_526),
.Y(n_3272)
);

OAI21x1_ASAP7_75t_L g3273 ( 
.A1(n_3037),
.A2(n_527),
.B(n_526),
.Y(n_3273)
);

CKINVDCx16_ASAP7_75t_R g3274 ( 
.A(n_2811),
.Y(n_3274)
);

AOI221x1_ASAP7_75t_L g3275 ( 
.A1(n_2836),
.A2(n_527),
.B1(n_525),
.B2(n_526),
.C(n_528),
.Y(n_3275)
);

OAI21xp5_ASAP7_75t_SL g3276 ( 
.A1(n_2739),
.A2(n_536),
.B(n_529),
.Y(n_3276)
);

INVx1_ASAP7_75t_SL g3277 ( 
.A(n_2941),
.Y(n_3277)
);

OAI22xp5_ASAP7_75t_L g3278 ( 
.A1(n_3005),
.A2(n_533),
.B1(n_531),
.B2(n_532),
.Y(n_3278)
);

NAND2xp5_ASAP7_75t_L g3279 ( 
.A(n_2950),
.B(n_531),
.Y(n_3279)
);

INVx1_ASAP7_75t_L g3280 ( 
.A(n_3043),
.Y(n_3280)
);

NAND3xp33_ASAP7_75t_L g3281 ( 
.A(n_2840),
.B(n_531),
.C(n_532),
.Y(n_3281)
);

NAND3xp33_ASAP7_75t_L g3282 ( 
.A(n_2904),
.B(n_532),
.C(n_533),
.Y(n_3282)
);

INVx1_ASAP7_75t_L g3283 ( 
.A(n_2906),
.Y(n_3283)
);

HB1xp67_ASAP7_75t_L g3284 ( 
.A(n_2839),
.Y(n_3284)
);

NAND2xp33_ASAP7_75t_L g3285 ( 
.A(n_2968),
.B(n_533),
.Y(n_3285)
);

BUFx10_ASAP7_75t_L g3286 ( 
.A(n_2896),
.Y(n_3286)
);

OAI21xp5_ASAP7_75t_L g3287 ( 
.A1(n_3079),
.A2(n_534),
.B(n_535),
.Y(n_3287)
);

A2O1A1Ixp33_ASAP7_75t_L g3288 ( 
.A1(n_2988),
.A2(n_536),
.B(n_534),
.C(n_535),
.Y(n_3288)
);

A2O1A1Ixp33_ASAP7_75t_L g3289 ( 
.A1(n_3006),
.A2(n_539),
.B(n_537),
.C(n_538),
.Y(n_3289)
);

INVx3_ASAP7_75t_L g3290 ( 
.A(n_2981),
.Y(n_3290)
);

BUFx3_ASAP7_75t_L g3291 ( 
.A(n_2985),
.Y(n_3291)
);

AOI21xp5_ASAP7_75t_L g3292 ( 
.A1(n_3138),
.A2(n_540),
.B(n_541),
.Y(n_3292)
);

OAI22xp5_ASAP7_75t_L g3293 ( 
.A1(n_3005),
.A2(n_543),
.B1(n_540),
.B2(n_542),
.Y(n_3293)
);

AOI21xp5_ASAP7_75t_L g3294 ( 
.A1(n_3138),
.A2(n_2972),
.B(n_2969),
.Y(n_3294)
);

AOI31xp67_ASAP7_75t_L g3295 ( 
.A1(n_3126),
.A2(n_544),
.A3(n_542),
.B(n_543),
.Y(n_3295)
);

AOI22x1_ASAP7_75t_L g3296 ( 
.A1(n_3026),
.A2(n_545),
.B1(n_543),
.B2(n_544),
.Y(n_3296)
);

AOI31xp67_ASAP7_75t_L g3297 ( 
.A1(n_3130),
.A2(n_546),
.A3(n_544),
.B(n_545),
.Y(n_3297)
);

NAND2xp5_ASAP7_75t_SL g3298 ( 
.A(n_3024),
.B(n_546),
.Y(n_3298)
);

NAND2x1p5_ASAP7_75t_L g3299 ( 
.A(n_2952),
.B(n_547),
.Y(n_3299)
);

INVx1_ASAP7_75t_L g3300 ( 
.A(n_3099),
.Y(n_3300)
);

OAI22x1_ASAP7_75t_L g3301 ( 
.A1(n_2845),
.A2(n_549),
.B1(n_547),
.B2(n_548),
.Y(n_3301)
);

AOI221x1_ASAP7_75t_L g3302 ( 
.A1(n_2862),
.A2(n_550),
.B1(n_548),
.B2(n_549),
.C(n_551),
.Y(n_3302)
);

NAND2xp5_ASAP7_75t_L g3303 ( 
.A(n_2973),
.B(n_550),
.Y(n_3303)
);

BUFx10_ASAP7_75t_L g3304 ( 
.A(n_2930),
.Y(n_3304)
);

INVx1_ASAP7_75t_L g3305 ( 
.A(n_2762),
.Y(n_3305)
);

OAI22xp5_ASAP7_75t_L g3306 ( 
.A1(n_3106),
.A2(n_553),
.B1(n_551),
.B2(n_552),
.Y(n_3306)
);

A2O1A1Ixp33_ASAP7_75t_L g3307 ( 
.A1(n_2936),
.A2(n_554),
.B(n_552),
.C(n_553),
.Y(n_3307)
);

OAI22xp5_ASAP7_75t_L g3308 ( 
.A1(n_2765),
.A2(n_555),
.B1(n_552),
.B2(n_554),
.Y(n_3308)
);

NOR2xp67_ASAP7_75t_L g3309 ( 
.A(n_2957),
.B(n_554),
.Y(n_3309)
);

OAI21xp5_ASAP7_75t_L g3310 ( 
.A1(n_2905),
.A2(n_555),
.B(n_556),
.Y(n_3310)
);

O2A1O1Ixp33_ASAP7_75t_L g3311 ( 
.A1(n_2806),
.A2(n_557),
.B(n_555),
.C(n_556),
.Y(n_3311)
);

AOI21xp5_ASAP7_75t_L g3312 ( 
.A1(n_3038),
.A2(n_556),
.B(n_557),
.Y(n_3312)
);

A2O1A1Ixp33_ASAP7_75t_L g3313 ( 
.A1(n_2888),
.A2(n_559),
.B(n_557),
.C(n_558),
.Y(n_3313)
);

NAND2xp5_ASAP7_75t_L g3314 ( 
.A(n_3056),
.B(n_558),
.Y(n_3314)
);

O2A1O1Ixp33_ASAP7_75t_L g3315 ( 
.A1(n_2809),
.A2(n_561),
.B(n_559),
.C(n_560),
.Y(n_3315)
);

INVx2_ASAP7_75t_L g3316 ( 
.A(n_2745),
.Y(n_3316)
);

NAND2xp5_ASAP7_75t_L g3317 ( 
.A(n_3059),
.B(n_559),
.Y(n_3317)
);

AOI21xp5_ASAP7_75t_L g3318 ( 
.A1(n_3064),
.A2(n_560),
.B(n_561),
.Y(n_3318)
);

AO32x2_ASAP7_75t_L g3319 ( 
.A1(n_2918),
.A2(n_564),
.A3(n_562),
.B1(n_563),
.B2(n_565),
.Y(n_3319)
);

NAND2xp5_ASAP7_75t_L g3320 ( 
.A(n_2761),
.B(n_563),
.Y(n_3320)
);

OAI21xp5_ASAP7_75t_L g3321 ( 
.A1(n_3096),
.A2(n_565),
.B(n_566),
.Y(n_3321)
);

OAI21x1_ASAP7_75t_L g3322 ( 
.A1(n_2928),
.A2(n_568),
.B(n_569),
.Y(n_3322)
);

NOR4xp25_ASAP7_75t_L g3323 ( 
.A(n_2744),
.B(n_570),
.C(n_568),
.D(n_569),
.Y(n_3323)
);

BUFx3_ASAP7_75t_L g3324 ( 
.A(n_3105),
.Y(n_3324)
);

AOI22xp5_ASAP7_75t_L g3325 ( 
.A1(n_2881),
.A2(n_2951),
.B1(n_3035),
.B2(n_3032),
.Y(n_3325)
);

OAI21x1_ASAP7_75t_L g3326 ( 
.A1(n_3011),
.A2(n_569),
.B(n_570),
.Y(n_3326)
);

OAI21x1_ASAP7_75t_L g3327 ( 
.A1(n_3030),
.A2(n_570),
.B(n_571),
.Y(n_3327)
);

INVx2_ASAP7_75t_L g3328 ( 
.A(n_2748),
.Y(n_3328)
);

INVx2_ASAP7_75t_SL g3329 ( 
.A(n_3127),
.Y(n_3329)
);

NAND3xp33_ASAP7_75t_SL g3330 ( 
.A(n_2938),
.B(n_571),
.C(n_572),
.Y(n_3330)
);

NAND3xp33_ASAP7_75t_SL g3331 ( 
.A(n_2803),
.B(n_2870),
.C(n_2822),
.Y(n_3331)
);

INVxp67_ASAP7_75t_L g3332 ( 
.A(n_2930),
.Y(n_3332)
);

INVx1_ASAP7_75t_L g3333 ( 
.A(n_2787),
.Y(n_3333)
);

AOI21xp5_ASAP7_75t_L g3334 ( 
.A1(n_3093),
.A2(n_572),
.B(n_573),
.Y(n_3334)
);

AOI22xp33_ASAP7_75t_L g3335 ( 
.A1(n_3060),
.A2(n_3092),
.B1(n_3016),
.B2(n_3117),
.Y(n_3335)
);

OAI21x1_ASAP7_75t_L g3336 ( 
.A1(n_3084),
.A2(n_572),
.B(n_574),
.Y(n_3336)
);

OR2x2_ASAP7_75t_L g3337 ( 
.A(n_2875),
.B(n_574),
.Y(n_3337)
);

AND2x2_ASAP7_75t_L g3338 ( 
.A(n_2845),
.B(n_574),
.Y(n_3338)
);

BUFx6f_ASAP7_75t_L g3339 ( 
.A(n_2743),
.Y(n_3339)
);

INVx2_ASAP7_75t_L g3340 ( 
.A(n_2750),
.Y(n_3340)
);

AOI221x1_ASAP7_75t_L g3341 ( 
.A1(n_2891),
.A2(n_577),
.B1(n_575),
.B2(n_576),
.C(n_578),
.Y(n_3341)
);

AO32x2_ASAP7_75t_L g3342 ( 
.A1(n_2991),
.A2(n_577),
.A3(n_575),
.B1(n_576),
.B2(n_578),
.Y(n_3342)
);

BUFx2_ASAP7_75t_L g3343 ( 
.A(n_2772),
.Y(n_3343)
);

INVx5_ASAP7_75t_L g3344 ( 
.A(n_2983),
.Y(n_3344)
);

INVx1_ASAP7_75t_L g3345 ( 
.A(n_2795),
.Y(n_3345)
);

OAI21x1_ASAP7_75t_L g3346 ( 
.A1(n_2866),
.A2(n_575),
.B(n_576),
.Y(n_3346)
);

AOI21xp5_ASAP7_75t_L g3347 ( 
.A1(n_3012),
.A2(n_579),
.B(n_580),
.Y(n_3347)
);

AOI21xp5_ASAP7_75t_L g3348 ( 
.A1(n_2992),
.A2(n_579),
.B(n_580),
.Y(n_3348)
);

A2O1A1Ixp33_ASAP7_75t_L g3349 ( 
.A1(n_2782),
.A2(n_582),
.B(n_580),
.C(n_581),
.Y(n_3349)
);

A2O1A1Ixp33_ASAP7_75t_L g3350 ( 
.A1(n_2940),
.A2(n_583),
.B(n_581),
.C(n_582),
.Y(n_3350)
);

AND2x2_ASAP7_75t_L g3351 ( 
.A(n_2913),
.B(n_581),
.Y(n_3351)
);

AOI21xp5_ASAP7_75t_L g3352 ( 
.A1(n_3009),
.A2(n_584),
.B(n_585),
.Y(n_3352)
);

INVx1_ASAP7_75t_L g3353 ( 
.A(n_2800),
.Y(n_3353)
);

AOI21xp5_ASAP7_75t_L g3354 ( 
.A1(n_3000),
.A2(n_584),
.B(n_585),
.Y(n_3354)
);

NAND3xp33_ASAP7_75t_L g3355 ( 
.A(n_3091),
.B(n_586),
.C(n_587),
.Y(n_3355)
);

INVx1_ASAP7_75t_L g3356 ( 
.A(n_2802),
.Y(n_3356)
);

A2O1A1Ixp33_ASAP7_75t_L g3357 ( 
.A1(n_2827),
.A2(n_588),
.B(n_586),
.C(n_587),
.Y(n_3357)
);

OAI21xp5_ASAP7_75t_SL g3358 ( 
.A1(n_3039),
.A2(n_586),
.B(n_589),
.Y(n_3358)
);

NOR2xp33_ASAP7_75t_L g3359 ( 
.A(n_2830),
.B(n_589),
.Y(n_3359)
);

OR2x6_ASAP7_75t_L g3360 ( 
.A(n_2983),
.B(n_589),
.Y(n_3360)
);

BUFx10_ASAP7_75t_L g3361 ( 
.A(n_2929),
.Y(n_3361)
);

AOI21x1_ASAP7_75t_L g3362 ( 
.A1(n_3142),
.A2(n_689),
.B(n_687),
.Y(n_3362)
);

AOI21x1_ASAP7_75t_L g3363 ( 
.A1(n_2944),
.A2(n_690),
.B(n_689),
.Y(n_3363)
);

BUFx2_ASAP7_75t_L g3364 ( 
.A(n_2772),
.Y(n_3364)
);

AOI21xp5_ASAP7_75t_L g3365 ( 
.A1(n_3014),
.A2(n_590),
.B(n_591),
.Y(n_3365)
);

AOI21xp5_ASAP7_75t_L g3366 ( 
.A1(n_3018),
.A2(n_591),
.B(n_592),
.Y(n_3366)
);

OAI21xp5_ASAP7_75t_SL g3367 ( 
.A1(n_2954),
.A2(n_592),
.B(n_593),
.Y(n_3367)
);

INVx1_ASAP7_75t_L g3368 ( 
.A(n_2810),
.Y(n_3368)
);

AOI21xp5_ASAP7_75t_L g3369 ( 
.A1(n_3034),
.A2(n_3041),
.B(n_2880),
.Y(n_3369)
);

BUFx2_ASAP7_75t_L g3370 ( 
.A(n_2807),
.Y(n_3370)
);

OAI21x1_ASAP7_75t_L g3371 ( 
.A1(n_2821),
.A2(n_594),
.B(n_595),
.Y(n_3371)
);

OAI21x1_ASAP7_75t_L g3372 ( 
.A1(n_2853),
.A2(n_596),
.B(n_597),
.Y(n_3372)
);

AOI21xp5_ASAP7_75t_SL g3373 ( 
.A1(n_2859),
.A2(n_596),
.B(n_598),
.Y(n_3373)
);

O2A1O1Ixp33_ASAP7_75t_L g3374 ( 
.A1(n_2833),
.A2(n_599),
.B(n_596),
.C(n_598),
.Y(n_3374)
);

AOI21xp5_ASAP7_75t_L g3375 ( 
.A1(n_3120),
.A2(n_599),
.B(n_600),
.Y(n_3375)
);

BUFx6f_ASAP7_75t_L g3376 ( 
.A(n_2743),
.Y(n_3376)
);

A2O1A1Ixp33_ASAP7_75t_L g3377 ( 
.A1(n_2848),
.A2(n_601),
.B(n_599),
.C(n_600),
.Y(n_3377)
);

BUFx2_ASAP7_75t_R g3378 ( 
.A(n_2780),
.Y(n_3378)
);

CKINVDCx11_ASAP7_75t_R g3379 ( 
.A(n_3121),
.Y(n_3379)
);

AOI22xp5_ASAP7_75t_L g3380 ( 
.A1(n_3013),
.A2(n_602),
.B1(n_600),
.B2(n_601),
.Y(n_3380)
);

HB1xp67_ASAP7_75t_L g3381 ( 
.A(n_2977),
.Y(n_3381)
);

AOI21xp5_ASAP7_75t_L g3382 ( 
.A1(n_3141),
.A2(n_601),
.B(n_602),
.Y(n_3382)
);

AOI21xp5_ASAP7_75t_L g3383 ( 
.A1(n_3148),
.A2(n_603),
.B(n_604),
.Y(n_3383)
);

A2O1A1Ixp33_ASAP7_75t_L g3384 ( 
.A1(n_2863),
.A2(n_605),
.B(n_603),
.C(n_604),
.Y(n_3384)
);

A2O1A1Ixp33_ASAP7_75t_L g3385 ( 
.A1(n_3066),
.A2(n_606),
.B(n_603),
.C(n_605),
.Y(n_3385)
);

OAI21x1_ASAP7_75t_L g3386 ( 
.A1(n_2908),
.A2(n_606),
.B(n_607),
.Y(n_3386)
);

AND2x4_ASAP7_75t_L g3387 ( 
.A(n_2801),
.B(n_606),
.Y(n_3387)
);

NOR2xp33_ASAP7_75t_L g3388 ( 
.A(n_2857),
.B(n_607),
.Y(n_3388)
);

NOR2xp33_ASAP7_75t_SL g3389 ( 
.A(n_2783),
.B(n_607),
.Y(n_3389)
);

HB1xp67_ASAP7_75t_L g3390 ( 
.A(n_2801),
.Y(n_3390)
);

AOI22xp33_ASAP7_75t_L g3391 ( 
.A1(n_3121),
.A2(n_610),
.B1(n_608),
.B2(n_609),
.Y(n_3391)
);

OAI21xp33_ASAP7_75t_L g3392 ( 
.A1(n_2998),
.A2(n_3103),
.B(n_3109),
.Y(n_3392)
);

INVx1_ASAP7_75t_SL g3393 ( 
.A(n_3075),
.Y(n_3393)
);

AOI21xp5_ASAP7_75t_L g3394 ( 
.A1(n_3090),
.A2(n_609),
.B(n_610),
.Y(n_3394)
);

AOI21x1_ASAP7_75t_L g3395 ( 
.A1(n_3023),
.A2(n_692),
.B(n_690),
.Y(n_3395)
);

AOI21xp5_ASAP7_75t_L g3396 ( 
.A1(n_3104),
.A2(n_611),
.B(n_612),
.Y(n_3396)
);

AOI21xp5_ASAP7_75t_L g3397 ( 
.A1(n_2812),
.A2(n_3088),
.B(n_3067),
.Y(n_3397)
);

BUFx2_ASAP7_75t_L g3398 ( 
.A(n_2958),
.Y(n_3398)
);

NOR2xp67_ASAP7_75t_SL g3399 ( 
.A(n_2958),
.B(n_613),
.Y(n_3399)
);

A2O1A1Ixp33_ASAP7_75t_L g3400 ( 
.A1(n_3047),
.A2(n_615),
.B(n_613),
.C(n_614),
.Y(n_3400)
);

BUFx4f_ASAP7_75t_L g3401 ( 
.A(n_3154),
.Y(n_3401)
);

INVx4_ASAP7_75t_L g3402 ( 
.A(n_3213),
.Y(n_3402)
);

INVx2_ASAP7_75t_SL g3403 ( 
.A(n_3184),
.Y(n_3403)
);

NAND2x1p5_ASAP7_75t_L g3404 ( 
.A(n_3163),
.B(n_2874),
.Y(n_3404)
);

AOI22xp33_ASAP7_75t_L g3405 ( 
.A1(n_3331),
.A2(n_2804),
.B1(n_3087),
.B2(n_3022),
.Y(n_3405)
);

BUFx3_ASAP7_75t_L g3406 ( 
.A(n_3324),
.Y(n_3406)
);

OAI22xp33_ASAP7_75t_L g3407 ( 
.A1(n_3360),
.A2(n_2903),
.B1(n_2847),
.B2(n_2816),
.Y(n_3407)
);

OAI22xp5_ASAP7_75t_L g3408 ( 
.A1(n_3360),
.A2(n_2916),
.B1(n_3100),
.B2(n_2776),
.Y(n_3408)
);

CKINVDCx11_ASAP7_75t_R g3409 ( 
.A(n_3258),
.Y(n_3409)
);

BUFx6f_ASAP7_75t_L g3410 ( 
.A(n_3214),
.Y(n_3410)
);

OAI22x1_ASAP7_75t_L g3411 ( 
.A1(n_3344),
.A2(n_2796),
.B1(n_2804),
.B2(n_3100),
.Y(n_3411)
);

BUFx12f_ASAP7_75t_L g3412 ( 
.A(n_3237),
.Y(n_3412)
);

AOI22xp33_ASAP7_75t_SL g3413 ( 
.A1(n_3344),
.A2(n_3095),
.B1(n_3045),
.B2(n_3094),
.Y(n_3413)
);

BUFx8_ASAP7_75t_L g3414 ( 
.A(n_3181),
.Y(n_3414)
);

INVx6_ASAP7_75t_L g3415 ( 
.A(n_3152),
.Y(n_3415)
);

BUFx12f_ASAP7_75t_L g3416 ( 
.A(n_3189),
.Y(n_3416)
);

OR2x2_ASAP7_75t_L g3417 ( 
.A(n_3202),
.B(n_3085),
.Y(n_3417)
);

BUFx3_ASAP7_75t_L g3418 ( 
.A(n_3181),
.Y(n_3418)
);

AOI22xp33_ASAP7_75t_SL g3419 ( 
.A1(n_3245),
.A2(n_3065),
.B1(n_3123),
.B2(n_3111),
.Y(n_3419)
);

INVx1_ASAP7_75t_SL g3420 ( 
.A(n_3201),
.Y(n_3420)
);

INVx4_ASAP7_75t_L g3421 ( 
.A(n_3214),
.Y(n_3421)
);

OAI22xp5_ASAP7_75t_SL g3422 ( 
.A1(n_3176),
.A2(n_2831),
.B1(n_2788),
.B2(n_2855),
.Y(n_3422)
);

BUFx6f_ASAP7_75t_L g3423 ( 
.A(n_3230),
.Y(n_3423)
);

AOI22xp33_ASAP7_75t_SL g3424 ( 
.A1(n_3245),
.A2(n_3111),
.B1(n_3025),
.B2(n_2919),
.Y(n_3424)
);

AOI22xp33_ASAP7_75t_L g3425 ( 
.A1(n_3392),
.A2(n_3151),
.B1(n_2926),
.B2(n_2931),
.Y(n_3425)
);

INVx1_ASAP7_75t_L g3426 ( 
.A(n_3162),
.Y(n_3426)
);

BUFx12f_ASAP7_75t_L g3427 ( 
.A(n_3266),
.Y(n_3427)
);

INVx1_ASAP7_75t_L g3428 ( 
.A(n_3187),
.Y(n_3428)
);

INVx4_ASAP7_75t_L g3429 ( 
.A(n_3225),
.Y(n_3429)
);

BUFx12f_ASAP7_75t_L g3430 ( 
.A(n_3379),
.Y(n_3430)
);

AND2x2_ASAP7_75t_L g3431 ( 
.A(n_3240),
.B(n_3115),
.Y(n_3431)
);

HB1xp67_ASAP7_75t_L g3432 ( 
.A(n_3179),
.Y(n_3432)
);

INVx1_ASAP7_75t_L g3433 ( 
.A(n_3196),
.Y(n_3433)
);

INVx6_ASAP7_75t_L g3434 ( 
.A(n_3230),
.Y(n_3434)
);

BUFx12f_ASAP7_75t_L g3435 ( 
.A(n_3361),
.Y(n_3435)
);

OAI22xp5_ASAP7_75t_L g3436 ( 
.A1(n_3325),
.A2(n_2771),
.B1(n_3083),
.B2(n_3061),
.Y(n_3436)
);

CKINVDCx5p33_ASAP7_75t_R g3437 ( 
.A(n_3217),
.Y(n_3437)
);

AOI22xp33_ASAP7_75t_L g3438 ( 
.A1(n_3194),
.A2(n_3186),
.B1(n_3155),
.B2(n_3159),
.Y(n_3438)
);

OAI22xp5_ASAP7_75t_SL g3439 ( 
.A1(n_3274),
.A2(n_2814),
.B1(n_2824),
.B2(n_2747),
.Y(n_3439)
);

CKINVDCx6p67_ASAP7_75t_R g3440 ( 
.A(n_3165),
.Y(n_3440)
);

AOI22xp33_ASAP7_75t_SL g3441 ( 
.A1(n_3268),
.A2(n_3008),
.B1(n_3040),
.B2(n_2993),
.Y(n_3441)
);

INVx3_ASAP7_75t_L g3442 ( 
.A(n_3290),
.Y(n_3442)
);

AOI22xp33_ASAP7_75t_L g3443 ( 
.A1(n_3170),
.A2(n_3031),
.B1(n_2939),
.B2(n_2799),
.Y(n_3443)
);

CKINVDCx11_ASAP7_75t_R g3444 ( 
.A(n_3286),
.Y(n_3444)
);

CKINVDCx20_ASAP7_75t_R g3445 ( 
.A(n_3291),
.Y(n_3445)
);

BUFx3_ASAP7_75t_L g3446 ( 
.A(n_3329),
.Y(n_3446)
);

INVx2_ASAP7_75t_L g3447 ( 
.A(n_3164),
.Y(n_3447)
);

AOI22xp33_ASAP7_75t_L g3448 ( 
.A1(n_3170),
.A2(n_2964),
.B1(n_2914),
.B2(n_2920),
.Y(n_3448)
);

AOI22xp33_ASAP7_75t_L g3449 ( 
.A1(n_3250),
.A2(n_2986),
.B1(n_3076),
.B2(n_3042),
.Y(n_3449)
);

INVx2_ASAP7_75t_L g3450 ( 
.A(n_3168),
.Y(n_3450)
);

INVx6_ASAP7_75t_L g3451 ( 
.A(n_3304),
.Y(n_3451)
);

OAI22xp33_ASAP7_75t_L g3452 ( 
.A1(n_3276),
.A2(n_3129),
.B1(n_3134),
.B2(n_2846),
.Y(n_3452)
);

AOI22xp33_ASAP7_75t_SL g3453 ( 
.A1(n_3390),
.A2(n_3086),
.B1(n_3112),
.B2(n_3078),
.Y(n_3453)
);

BUFx4f_ASAP7_75t_SL g3454 ( 
.A(n_3265),
.Y(n_3454)
);

OAI21xp5_ASAP7_75t_SL g3455 ( 
.A1(n_3174),
.A2(n_3019),
.B(n_3125),
.Y(n_3455)
);

AND2x2_ASAP7_75t_L g3456 ( 
.A(n_3252),
.B(n_3338),
.Y(n_3456)
);

AND2x2_ASAP7_75t_L g3457 ( 
.A(n_3351),
.B(n_2917),
.Y(n_3457)
);

AOI22xp33_ASAP7_75t_SL g3458 ( 
.A1(n_3389),
.A2(n_3285),
.B1(n_3387),
.B2(n_3296),
.Y(n_3458)
);

AOI22xp33_ASAP7_75t_L g3459 ( 
.A1(n_3330),
.A2(n_3131),
.B1(n_3128),
.B2(n_2955),
.Y(n_3459)
);

AOI22xp33_ASAP7_75t_L g3460 ( 
.A1(n_3210),
.A2(n_3335),
.B1(n_3246),
.B2(n_3247),
.Y(n_3460)
);

AOI22xp33_ASAP7_75t_L g3461 ( 
.A1(n_3359),
.A2(n_2960),
.B1(n_2922),
.B2(n_3029),
.Y(n_3461)
);

BUFx6f_ASAP7_75t_L g3462 ( 
.A(n_3339),
.Y(n_3462)
);

AOI22xp33_ASAP7_75t_L g3463 ( 
.A1(n_3183),
.A2(n_3052),
.B1(n_3053),
.B2(n_3050),
.Y(n_3463)
);

AOI22xp33_ASAP7_75t_L g3464 ( 
.A1(n_3388),
.A2(n_2791),
.B1(n_2868),
.B2(n_2867),
.Y(n_3464)
);

AOI22xp33_ASAP7_75t_SL g3465 ( 
.A1(n_3278),
.A2(n_3119),
.B1(n_3137),
.B2(n_3118),
.Y(n_3465)
);

CKINVDCx11_ASAP7_75t_R g3466 ( 
.A(n_3277),
.Y(n_3466)
);

AOI22xp33_ASAP7_75t_SL g3467 ( 
.A1(n_3293),
.A2(n_2877),
.B1(n_2933),
.B2(n_2935),
.Y(n_3467)
);

INVx6_ASAP7_75t_L g3468 ( 
.A(n_3195),
.Y(n_3468)
);

BUFx4_ASAP7_75t_SL g3469 ( 
.A(n_3343),
.Y(n_3469)
);

BUFx2_ASAP7_75t_SL g3470 ( 
.A(n_3309),
.Y(n_3470)
);

BUFx3_ASAP7_75t_L g3471 ( 
.A(n_3231),
.Y(n_3471)
);

BUFx12f_ASAP7_75t_L g3472 ( 
.A(n_3299),
.Y(n_3472)
);

CKINVDCx20_ASAP7_75t_R g3473 ( 
.A(n_3393),
.Y(n_3473)
);

OAI22xp5_ASAP7_75t_L g3474 ( 
.A1(n_3358),
.A2(n_3072),
.B1(n_2984),
.B2(n_3101),
.Y(n_3474)
);

INVx2_ASAP7_75t_L g3475 ( 
.A(n_3177),
.Y(n_3475)
);

OAI22xp33_ASAP7_75t_L g3476 ( 
.A1(n_3367),
.A2(n_2741),
.B1(n_2740),
.B2(n_2793),
.Y(n_3476)
);

AOI22xp33_ASAP7_75t_L g3477 ( 
.A1(n_3308),
.A2(n_3020),
.B1(n_2858),
.B2(n_3145),
.Y(n_3477)
);

BUFx10_ASAP7_75t_L g3478 ( 
.A(n_3198),
.Y(n_3478)
);

INVx4_ASAP7_75t_SL g3479 ( 
.A(n_3248),
.Y(n_3479)
);

INVx2_ASAP7_75t_L g3480 ( 
.A(n_3199),
.Y(n_3480)
);

INVx2_ASAP7_75t_L g3481 ( 
.A(n_3219),
.Y(n_3481)
);

OAI22xp5_ASAP7_75t_L g3482 ( 
.A1(n_3167),
.A2(n_3108),
.B1(n_3116),
.B2(n_3114),
.Y(n_3482)
);

INVx8_ASAP7_75t_L g3483 ( 
.A(n_3339),
.Y(n_3483)
);

BUFx6f_ASAP7_75t_L g3484 ( 
.A(n_3376),
.Y(n_3484)
);

BUFx2_ASAP7_75t_SL g3485 ( 
.A(n_3253),
.Y(n_3485)
);

INVx4_ASAP7_75t_L g3486 ( 
.A(n_3364),
.Y(n_3486)
);

CKINVDCx6p67_ASAP7_75t_R g3487 ( 
.A(n_3301),
.Y(n_3487)
);

BUFx12f_ASAP7_75t_L g3488 ( 
.A(n_3337),
.Y(n_3488)
);

OAI22xp33_ASAP7_75t_L g3489 ( 
.A1(n_3380),
.A2(n_2967),
.B1(n_2915),
.B2(n_3098),
.Y(n_3489)
);

INVx1_ASAP7_75t_L g3490 ( 
.A(n_3267),
.Y(n_3490)
);

BUFx3_ASAP7_75t_L g3491 ( 
.A(n_3370),
.Y(n_3491)
);

OAI22xp5_ASAP7_75t_SL g3492 ( 
.A1(n_3332),
.A2(n_3046),
.B1(n_2942),
.B2(n_2860),
.Y(n_3492)
);

AOI22xp33_ASAP7_75t_L g3493 ( 
.A1(n_3321),
.A2(n_2912),
.B1(n_2892),
.B2(n_2911),
.Y(n_3493)
);

NAND2x1p5_ASAP7_75t_L g3494 ( 
.A(n_3399),
.B(n_3249),
.Y(n_3494)
);

NAND2x1p5_ASAP7_75t_L g3495 ( 
.A(n_3398),
.B(n_3097),
.Y(n_3495)
);

INVx1_ASAP7_75t_L g3496 ( 
.A(n_3280),
.Y(n_3496)
);

BUFx3_ASAP7_75t_L g3497 ( 
.A(n_3284),
.Y(n_3497)
);

INVx6_ASAP7_75t_L g3498 ( 
.A(n_3376),
.Y(n_3498)
);

INVxp67_ASAP7_75t_SL g3499 ( 
.A(n_3294),
.Y(n_3499)
);

HB1xp67_ASAP7_75t_L g3500 ( 
.A(n_3381),
.Y(n_3500)
);

INVx1_ASAP7_75t_L g3501 ( 
.A(n_3283),
.Y(n_3501)
);

AOI22xp33_ASAP7_75t_L g3502 ( 
.A1(n_3244),
.A2(n_2946),
.B1(n_2959),
.B2(n_2953),
.Y(n_3502)
);

INVx1_ASAP7_75t_SL g3503 ( 
.A(n_3378),
.Y(n_3503)
);

NAND2xp33_ASAP7_75t_SL g3504 ( 
.A(n_3306),
.B(n_3097),
.Y(n_3504)
);

AOI22xp33_ASAP7_75t_L g3505 ( 
.A1(n_3229),
.A2(n_2962),
.B1(n_2971),
.B2(n_2963),
.Y(n_3505)
);

INVx2_ASAP7_75t_L g3506 ( 
.A(n_3316),
.Y(n_3506)
);

BUFx3_ASAP7_75t_L g3507 ( 
.A(n_3328),
.Y(n_3507)
);

AOI22xp33_ASAP7_75t_SL g3508 ( 
.A1(n_3160),
.A2(n_3133),
.B1(n_2990),
.B2(n_2965),
.Y(n_3508)
);

INVx2_ASAP7_75t_L g3509 ( 
.A(n_3340),
.Y(n_3509)
);

AOI22xp33_ASAP7_75t_SL g3510 ( 
.A1(n_3220),
.A2(n_3133),
.B1(n_3017),
.B2(n_3113),
.Y(n_3510)
);

AND2x4_ASAP7_75t_L g3511 ( 
.A(n_3185),
.B(n_2743),
.Y(n_3511)
);

INVx2_ASAP7_75t_L g3512 ( 
.A(n_3300),
.Y(n_3512)
);

INVx1_ASAP7_75t_L g3513 ( 
.A(n_3227),
.Y(n_3513)
);

INVx4_ASAP7_75t_L g3514 ( 
.A(n_3157),
.Y(n_3514)
);

AOI22xp33_ASAP7_75t_L g3515 ( 
.A1(n_3355),
.A2(n_3044),
.B1(n_3063),
.B2(n_3051),
.Y(n_3515)
);

INVx2_ASAP7_75t_L g3516 ( 
.A(n_3261),
.Y(n_3516)
);

NAND2xp5_ASAP7_75t_L g3517 ( 
.A(n_3271),
.B(n_3305),
.Y(n_3517)
);

BUFx12f_ASAP7_75t_L g3518 ( 
.A(n_3197),
.Y(n_3518)
);

CKINVDCx6p67_ASAP7_75t_R g3519 ( 
.A(n_3269),
.Y(n_3519)
);

INVx2_ASAP7_75t_L g3520 ( 
.A(n_3273),
.Y(n_3520)
);

OAI22x1_ASAP7_75t_L g3521 ( 
.A1(n_3281),
.A2(n_3107),
.B1(n_3055),
.B2(n_2956),
.Y(n_3521)
);

INVx1_ASAP7_75t_L g3522 ( 
.A(n_3371),
.Y(n_3522)
);

AOI22xp33_ASAP7_75t_L g3523 ( 
.A1(n_3209),
.A2(n_3292),
.B1(n_3222),
.B2(n_3282),
.Y(n_3523)
);

BUFx12f_ASAP7_75t_L g3524 ( 
.A(n_3391),
.Y(n_3524)
);

INVx5_ASAP7_75t_L g3525 ( 
.A(n_3373),
.Y(n_3525)
);

INVx4_ASAP7_75t_SL g3526 ( 
.A(n_3262),
.Y(n_3526)
);

AOI22xp33_ASAP7_75t_L g3527 ( 
.A1(n_3333),
.A2(n_3345),
.B1(n_3356),
.B2(n_3353),
.Y(n_3527)
);

CKINVDCx20_ASAP7_75t_R g3528 ( 
.A(n_3173),
.Y(n_3528)
);

INVxp67_ASAP7_75t_SL g3529 ( 
.A(n_3175),
.Y(n_3529)
);

NAND2xp5_ASAP7_75t_L g3530 ( 
.A(n_3368),
.B(n_2826),
.Y(n_3530)
);

AOI22xp33_ASAP7_75t_SL g3531 ( 
.A1(n_3287),
.A2(n_2786),
.B1(n_2813),
.B2(n_2790),
.Y(n_3531)
);

INVxp67_ASAP7_75t_SL g3532 ( 
.A(n_3156),
.Y(n_3532)
);

INVx1_ASAP7_75t_L g3533 ( 
.A(n_3372),
.Y(n_3533)
);

INVx4_ASAP7_75t_L g3534 ( 
.A(n_3226),
.Y(n_3534)
);

INVx4_ASAP7_75t_L g3535 ( 
.A(n_3212),
.Y(n_3535)
);

BUFx2_ASAP7_75t_L g3536 ( 
.A(n_3185),
.Y(n_3536)
);

BUFx2_ASAP7_75t_L g3537 ( 
.A(n_3192),
.Y(n_3537)
);

CKINVDCx11_ASAP7_75t_R g3538 ( 
.A(n_3260),
.Y(n_3538)
);

AOI22xp5_ASAP7_75t_L g3539 ( 
.A1(n_3193),
.A2(n_2832),
.B1(n_2882),
.B2(n_2838),
.Y(n_3539)
);

AOI22xp33_ASAP7_75t_SL g3540 ( 
.A1(n_3178),
.A2(n_2786),
.B1(n_2813),
.B2(n_2790),
.Y(n_3540)
);

AOI22xp5_ASAP7_75t_SL g3541 ( 
.A1(n_3256),
.A2(n_2890),
.B1(n_2760),
.B2(n_2949),
.Y(n_3541)
);

INVx1_ASAP7_75t_L g3542 ( 
.A(n_3386),
.Y(n_3542)
);

BUFx10_ASAP7_75t_L g3543 ( 
.A(n_3319),
.Y(n_3543)
);

OAI22xp5_ASAP7_75t_L g3544 ( 
.A1(n_3232),
.A2(n_2948),
.B1(n_2980),
.B2(n_2943),
.Y(n_3544)
);

BUFx6f_ASAP7_75t_L g3545 ( 
.A(n_3207),
.Y(n_3545)
);

BUFx6f_ASAP7_75t_L g3546 ( 
.A(n_3215),
.Y(n_3546)
);

BUFx3_ASAP7_75t_L g3547 ( 
.A(n_3216),
.Y(n_3547)
);

INVxp67_ASAP7_75t_SL g3548 ( 
.A(n_3166),
.Y(n_3548)
);

INVx2_ASAP7_75t_SL g3549 ( 
.A(n_3279),
.Y(n_3549)
);

INVx1_ASAP7_75t_L g3550 ( 
.A(n_3303),
.Y(n_3550)
);

INVx1_ASAP7_75t_L g3551 ( 
.A(n_3314),
.Y(n_3551)
);

NAND2xp5_ASAP7_75t_L g3552 ( 
.A(n_3317),
.B(n_2927),
.Y(n_3552)
);

BUFx4f_ASAP7_75t_SL g3553 ( 
.A(n_3298),
.Y(n_3553)
);

OA21x2_ASAP7_75t_L g3554 ( 
.A1(n_3529),
.A2(n_3397),
.B(n_3188),
.Y(n_3554)
);

INVx2_ASAP7_75t_SL g3555 ( 
.A(n_3469),
.Y(n_3555)
);

HB1xp67_ASAP7_75t_L g3556 ( 
.A(n_3507),
.Y(n_3556)
);

INVx1_ASAP7_75t_L g3557 ( 
.A(n_3426),
.Y(n_3557)
);

INVx2_ASAP7_75t_L g3558 ( 
.A(n_3447),
.Y(n_3558)
);

AOI21x1_ASAP7_75t_L g3559 ( 
.A1(n_3411),
.A2(n_3362),
.B(n_3171),
.Y(n_3559)
);

INVx1_ASAP7_75t_L g3560 ( 
.A(n_3428),
.Y(n_3560)
);

INVx2_ASAP7_75t_L g3561 ( 
.A(n_3450),
.Y(n_3561)
);

INVx3_ASAP7_75t_L g3562 ( 
.A(n_3486),
.Y(n_3562)
);

HB1xp67_ASAP7_75t_L g3563 ( 
.A(n_3500),
.Y(n_3563)
);

CKINVDCx20_ASAP7_75t_R g3564 ( 
.A(n_3409),
.Y(n_3564)
);

INVx1_ASAP7_75t_L g3565 ( 
.A(n_3433),
.Y(n_3565)
);

INVx2_ASAP7_75t_L g3566 ( 
.A(n_3475),
.Y(n_3566)
);

AO21x2_ASAP7_75t_L g3567 ( 
.A1(n_3532),
.A2(n_3395),
.B(n_3161),
.Y(n_3567)
);

INVx2_ASAP7_75t_L g3568 ( 
.A(n_3480),
.Y(n_3568)
);

INVx2_ASAP7_75t_L g3569 ( 
.A(n_3481),
.Y(n_3569)
);

INVx3_ASAP7_75t_L g3570 ( 
.A(n_3429),
.Y(n_3570)
);

AND2x2_ASAP7_75t_L g3571 ( 
.A(n_3456),
.B(n_3431),
.Y(n_3571)
);

HB1xp67_ASAP7_75t_L g3572 ( 
.A(n_3432),
.Y(n_3572)
);

INVx1_ASAP7_75t_L g3573 ( 
.A(n_3490),
.Y(n_3573)
);

AO21x2_ASAP7_75t_L g3574 ( 
.A1(n_3407),
.A2(n_3169),
.B(n_3369),
.Y(n_3574)
);

INVx1_ASAP7_75t_L g3575 ( 
.A(n_3496),
.Y(n_3575)
);

INVx2_ASAP7_75t_L g3576 ( 
.A(n_3506),
.Y(n_3576)
);

INVx2_ASAP7_75t_L g3577 ( 
.A(n_3509),
.Y(n_3577)
);

NAND2x1_ASAP7_75t_L g3578 ( 
.A(n_3402),
.B(n_2786),
.Y(n_3578)
);

BUFx10_ASAP7_75t_L g3579 ( 
.A(n_3415),
.Y(n_3579)
);

AOI21xp5_ASAP7_75t_L g3580 ( 
.A1(n_3499),
.A2(n_3190),
.B(n_3205),
.Y(n_3580)
);

INVx1_ASAP7_75t_SL g3581 ( 
.A(n_3420),
.Y(n_3581)
);

AND2x2_ASAP7_75t_L g3582 ( 
.A(n_3417),
.B(n_3158),
.Y(n_3582)
);

INVx1_ASAP7_75t_L g3583 ( 
.A(n_3501),
.Y(n_3583)
);

OR2x2_ASAP7_75t_L g3584 ( 
.A(n_3514),
.B(n_3172),
.Y(n_3584)
);

INVx2_ASAP7_75t_L g3585 ( 
.A(n_3512),
.Y(n_3585)
);

AOI22xp33_ASAP7_75t_L g3586 ( 
.A1(n_3524),
.A2(n_3218),
.B1(n_3191),
.B2(n_3180),
.Y(n_3586)
);

NAND2xp5_ASAP7_75t_L g3587 ( 
.A(n_3513),
.B(n_3323),
.Y(n_3587)
);

AO21x1_ASAP7_75t_L g3588 ( 
.A1(n_3504),
.A2(n_3352),
.B(n_3347),
.Y(n_3588)
);

INVx1_ASAP7_75t_L g3589 ( 
.A(n_3497),
.Y(n_3589)
);

INVx1_ASAP7_75t_L g3590 ( 
.A(n_3522),
.Y(n_3590)
);

AOI21x1_ASAP7_75t_L g3591 ( 
.A1(n_3537),
.A2(n_3363),
.B(n_3182),
.Y(n_3591)
);

INVx1_ASAP7_75t_L g3592 ( 
.A(n_3533),
.Y(n_3592)
);

INVx1_ASAP7_75t_L g3593 ( 
.A(n_3542),
.Y(n_3593)
);

AO21x1_ASAP7_75t_SL g3594 ( 
.A1(n_3523),
.A2(n_3310),
.B(n_3211),
.Y(n_3594)
);

INVx1_ASAP7_75t_L g3595 ( 
.A(n_3517),
.Y(n_3595)
);

AOI22xp33_ASAP7_75t_L g3596 ( 
.A1(n_3438),
.A2(n_3221),
.B1(n_3224),
.B2(n_3235),
.Y(n_3596)
);

INVx3_ASAP7_75t_L g3597 ( 
.A(n_3491),
.Y(n_3597)
);

INVx1_ASAP7_75t_L g3598 ( 
.A(n_3516),
.Y(n_3598)
);

INVx1_ASAP7_75t_L g3599 ( 
.A(n_3485),
.Y(n_3599)
);

INVx3_ASAP7_75t_L g3600 ( 
.A(n_3495),
.Y(n_3600)
);

OAI22xp33_ASAP7_75t_L g3601 ( 
.A1(n_3487),
.A2(n_3302),
.B1(n_3234),
.B2(n_3341),
.Y(n_3601)
);

INVx1_ASAP7_75t_L g3602 ( 
.A(n_3520),
.Y(n_3602)
);

INVx1_ASAP7_75t_L g3603 ( 
.A(n_3526),
.Y(n_3603)
);

INVx1_ASAP7_75t_L g3604 ( 
.A(n_3526),
.Y(n_3604)
);

O2A1O1Ixp33_ASAP7_75t_SL g3605 ( 
.A1(n_3503),
.A2(n_3403),
.B(n_3476),
.C(n_3445),
.Y(n_3605)
);

OAI22xp5_ASAP7_75t_L g3606 ( 
.A1(n_3458),
.A2(n_3377),
.B1(n_3384),
.B2(n_3357),
.Y(n_3606)
);

AOI21xp5_ASAP7_75t_L g3607 ( 
.A1(n_3548),
.A2(n_3204),
.B(n_3223),
.Y(n_3607)
);

INVx2_ASAP7_75t_L g3608 ( 
.A(n_3462),
.Y(n_3608)
);

INVx1_ASAP7_75t_L g3609 ( 
.A(n_3543),
.Y(n_3609)
);

INVx2_ASAP7_75t_L g3610 ( 
.A(n_3484),
.Y(n_3610)
);

BUFx2_ASAP7_75t_L g3611 ( 
.A(n_3442),
.Y(n_3611)
);

AND2x4_ASAP7_75t_L g3612 ( 
.A(n_3479),
.B(n_3158),
.Y(n_3612)
);

INVx2_ASAP7_75t_L g3613 ( 
.A(n_3484),
.Y(n_3613)
);

INVx1_ASAP7_75t_L g3614 ( 
.A(n_3527),
.Y(n_3614)
);

AOI21x1_ASAP7_75t_L g3615 ( 
.A1(n_3537),
.A2(n_3275),
.B(n_3236),
.Y(n_3615)
);

CKINVDCx16_ASAP7_75t_R g3616 ( 
.A(n_3430),
.Y(n_3616)
);

INVx1_ASAP7_75t_L g3617 ( 
.A(n_3550),
.Y(n_3617)
);

CKINVDCx5p33_ASAP7_75t_R g3618 ( 
.A(n_3401),
.Y(n_3618)
);

INVx1_ASAP7_75t_L g3619 ( 
.A(n_3551),
.Y(n_3619)
);

BUFx3_ASAP7_75t_L g3620 ( 
.A(n_3406),
.Y(n_3620)
);

INVx1_ASAP7_75t_SL g3621 ( 
.A(n_3466),
.Y(n_3621)
);

AOI21xp5_ASAP7_75t_L g3622 ( 
.A1(n_3540),
.A2(n_3203),
.B(n_3208),
.Y(n_3622)
);

AND2x2_ASAP7_75t_L g3623 ( 
.A(n_3457),
.B(n_3342),
.Y(n_3623)
);

INVx1_ASAP7_75t_L g3624 ( 
.A(n_3530),
.Y(n_3624)
);

INVx1_ASAP7_75t_L g3625 ( 
.A(n_3552),
.Y(n_3625)
);

INVx2_ASAP7_75t_L g3626 ( 
.A(n_3511),
.Y(n_3626)
);

INVx2_ASAP7_75t_SL g3627 ( 
.A(n_3414),
.Y(n_3627)
);

OAI21x1_ASAP7_75t_L g3628 ( 
.A1(n_3494),
.A2(n_3255),
.B(n_3254),
.Y(n_3628)
);

INVx1_ASAP7_75t_L g3629 ( 
.A(n_3549),
.Y(n_3629)
);

INVx2_ASAP7_75t_L g3630 ( 
.A(n_3511),
.Y(n_3630)
);

INVx2_ASAP7_75t_L g3631 ( 
.A(n_3410),
.Y(n_3631)
);

INVx2_ASAP7_75t_SL g3632 ( 
.A(n_3434),
.Y(n_3632)
);

INVx11_ASAP7_75t_L g3633 ( 
.A(n_3416),
.Y(n_3633)
);

INVx2_ASAP7_75t_SL g3634 ( 
.A(n_3434),
.Y(n_3634)
);

INVx2_ASAP7_75t_L g3635 ( 
.A(n_3410),
.Y(n_3635)
);

OAI21xp5_ASAP7_75t_L g3636 ( 
.A1(n_3455),
.A2(n_2774),
.B(n_3375),
.Y(n_3636)
);

AO21x2_ASAP7_75t_L g3637 ( 
.A1(n_3539),
.A2(n_3320),
.B(n_3382),
.Y(n_3637)
);

INVx2_ASAP7_75t_L g3638 ( 
.A(n_3498),
.Y(n_3638)
);

HB1xp67_ASAP7_75t_L g3639 ( 
.A(n_3479),
.Y(n_3639)
);

AO31x2_ASAP7_75t_L g3640 ( 
.A1(n_3535),
.A2(n_3206),
.A3(n_3400),
.B(n_3385),
.Y(n_3640)
);

A2O1A1Ixp33_ASAP7_75t_SL g3641 ( 
.A1(n_3425),
.A2(n_3405),
.B(n_3461),
.C(n_3460),
.Y(n_3641)
);

INVx1_ASAP7_75t_L g3642 ( 
.A(n_3536),
.Y(n_3642)
);

INVx2_ASAP7_75t_L g3643 ( 
.A(n_3498),
.Y(n_3643)
);

INVx1_ASAP7_75t_L g3644 ( 
.A(n_3536),
.Y(n_3644)
);

INVx3_ASAP7_75t_L g3645 ( 
.A(n_3468),
.Y(n_3645)
);

INVx2_ASAP7_75t_L g3646 ( 
.A(n_3534),
.Y(n_3646)
);

INVx2_ASAP7_75t_L g3647 ( 
.A(n_3547),
.Y(n_3647)
);

NAND2xp5_ASAP7_75t_SL g3648 ( 
.A(n_3510),
.B(n_3419),
.Y(n_3648)
);

AND2x2_ASAP7_75t_L g3649 ( 
.A(n_3418),
.B(n_2937),
.Y(n_3649)
);

AND2x2_ASAP7_75t_L g3650 ( 
.A(n_3421),
.B(n_3423),
.Y(n_3650)
);

NOR2xp33_ASAP7_75t_L g3651 ( 
.A(n_3518),
.B(n_614),
.Y(n_3651)
);

INVx1_ASAP7_75t_L g3652 ( 
.A(n_3545),
.Y(n_3652)
);

AO32x2_ASAP7_75t_L g3653 ( 
.A1(n_3555),
.A2(n_3492),
.A3(n_3606),
.B1(n_3439),
.B2(n_3632),
.Y(n_3653)
);

O2A1O1Ixp33_ASAP7_75t_L g3654 ( 
.A1(n_3641),
.A2(n_3408),
.B(n_3436),
.C(n_3404),
.Y(n_3654)
);

OR2x2_ASAP7_75t_L g3655 ( 
.A(n_3563),
.B(n_3446),
.Y(n_3655)
);

A2O1A1Ixp33_ASAP7_75t_L g3656 ( 
.A1(n_3570),
.A2(n_3470),
.B(n_3413),
.C(n_3424),
.Y(n_3656)
);

BUFx3_ASAP7_75t_L g3657 ( 
.A(n_3620),
.Y(n_3657)
);

AOI22xp5_ASAP7_75t_L g3658 ( 
.A1(n_3601),
.A2(n_3422),
.B1(n_3538),
.B2(n_3441),
.Y(n_3658)
);

AND2x2_ASAP7_75t_SL g3659 ( 
.A(n_3639),
.B(n_3423),
.Y(n_3659)
);

INVx2_ASAP7_75t_SL g3660 ( 
.A(n_3579),
.Y(n_3660)
);

AND2x2_ASAP7_75t_L g3661 ( 
.A(n_3571),
.B(n_3488),
.Y(n_3661)
);

AND2x2_ASAP7_75t_L g3662 ( 
.A(n_3556),
.B(n_3471),
.Y(n_3662)
);

AND2x2_ASAP7_75t_L g3663 ( 
.A(n_3582),
.B(n_3546),
.Y(n_3663)
);

AOI221xp5_ASAP7_75t_L g3664 ( 
.A1(n_3614),
.A2(n_3452),
.B1(n_3489),
.B2(n_3482),
.C(n_3474),
.Y(n_3664)
);

AND2x2_ASAP7_75t_L g3665 ( 
.A(n_3589),
.B(n_3508),
.Y(n_3665)
);

OAI21x1_ASAP7_75t_L g3666 ( 
.A1(n_3591),
.A2(n_3448),
.B(n_3346),
.Y(n_3666)
);

OR2x2_ASAP7_75t_L g3667 ( 
.A(n_3572),
.B(n_3440),
.Y(n_3667)
);

A2O1A1Ixp33_ASAP7_75t_L g3668 ( 
.A1(n_3570),
.A2(n_3525),
.B(n_3270),
.C(n_3315),
.Y(n_3668)
);

OAI22xp5_ASAP7_75t_L g3669 ( 
.A1(n_3648),
.A2(n_3465),
.B1(n_3519),
.B2(n_3553),
.Y(n_3669)
);

AO32x2_ASAP7_75t_L g3670 ( 
.A1(n_3634),
.A2(n_3544),
.A3(n_3473),
.B1(n_3444),
.B2(n_3435),
.Y(n_3670)
);

AO32x2_ASAP7_75t_L g3671 ( 
.A1(n_3627),
.A2(n_3541),
.A3(n_3478),
.B1(n_3451),
.B2(n_3531),
.Y(n_3671)
);

AND2x2_ASAP7_75t_L g3672 ( 
.A(n_3597),
.B(n_3451),
.Y(n_3672)
);

O2A1O1Ixp33_ASAP7_75t_L g3673 ( 
.A1(n_3587),
.A2(n_3636),
.B(n_3605),
.C(n_3629),
.Y(n_3673)
);

A2O1A1Ixp33_ASAP7_75t_L g3674 ( 
.A1(n_3562),
.A2(n_3525),
.B(n_3311),
.C(n_3374),
.Y(n_3674)
);

A2O1A1Ixp33_ASAP7_75t_L g3675 ( 
.A1(n_3562),
.A2(n_3525),
.B(n_3241),
.C(n_3453),
.Y(n_3675)
);

AOI22xp5_ASAP7_75t_L g3676 ( 
.A1(n_3637),
.A2(n_3467),
.B1(n_3472),
.B2(n_3443),
.Y(n_3676)
);

OA21x2_ASAP7_75t_L g3677 ( 
.A1(n_3609),
.A2(n_3463),
.B(n_3326),
.Y(n_3677)
);

INVx3_ASAP7_75t_L g3678 ( 
.A(n_3633),
.Y(n_3678)
);

OR2x2_ASAP7_75t_L g3679 ( 
.A(n_3625),
.B(n_3238),
.Y(n_3679)
);

INVxp67_ASAP7_75t_L g3680 ( 
.A(n_3611),
.Y(n_3680)
);

AO21x2_ASAP7_75t_L g3681 ( 
.A1(n_3607),
.A2(n_3272),
.B(n_3239),
.Y(n_3681)
);

NAND2xp5_ASAP7_75t_L g3682 ( 
.A(n_3623),
.B(n_3262),
.Y(n_3682)
);

AND2x4_ASAP7_75t_L g3683 ( 
.A(n_3650),
.B(n_3546),
.Y(n_3683)
);

INVx2_ASAP7_75t_L g3684 ( 
.A(n_3558),
.Y(n_3684)
);

OR2x2_ASAP7_75t_L g3685 ( 
.A(n_3585),
.B(n_3263),
.Y(n_3685)
);

AO32x2_ASAP7_75t_L g3686 ( 
.A1(n_3584),
.A2(n_3297),
.A3(n_3295),
.B1(n_3153),
.B2(n_3412),
.Y(n_3686)
);

INVx3_ASAP7_75t_L g3687 ( 
.A(n_3600),
.Y(n_3687)
);

NOR2x1_ASAP7_75t_SL g3688 ( 
.A(n_3599),
.B(n_3427),
.Y(n_3688)
);

AOI221xp5_ASAP7_75t_L g3689 ( 
.A1(n_3624),
.A2(n_3383),
.B1(n_3354),
.B2(n_3365),
.C(n_3348),
.Y(n_3689)
);

AND2x2_ASAP7_75t_L g3690 ( 
.A(n_3617),
.B(n_3415),
.Y(n_3690)
);

AND2x2_ASAP7_75t_L g3691 ( 
.A(n_3619),
.B(n_3528),
.Y(n_3691)
);

INVx1_ASAP7_75t_L g3692 ( 
.A(n_3557),
.Y(n_3692)
);

AND2x4_ASAP7_75t_L g3693 ( 
.A(n_3600),
.B(n_3437),
.Y(n_3693)
);

A2O1A1Ixp33_ASAP7_75t_L g3694 ( 
.A1(n_3651),
.A2(n_3312),
.B(n_3318),
.C(n_3449),
.Y(n_3694)
);

NOR2x1_ASAP7_75t_R g3695 ( 
.A(n_3618),
.B(n_3454),
.Y(n_3695)
);

INVx2_ASAP7_75t_L g3696 ( 
.A(n_3561),
.Y(n_3696)
);

AOI221xp5_ASAP7_75t_L g3697 ( 
.A1(n_3586),
.A2(n_3366),
.B1(n_3334),
.B2(n_3459),
.C(n_3502),
.Y(n_3697)
);

NOR2xp33_ASAP7_75t_L g3698 ( 
.A(n_3581),
.B(n_614),
.Y(n_3698)
);

O2A1O1Ixp33_ASAP7_75t_L g3699 ( 
.A1(n_3622),
.A2(n_3313),
.B(n_3350),
.C(n_3233),
.Y(n_3699)
);

AND2x2_ASAP7_75t_SL g3700 ( 
.A(n_3616),
.B(n_3464),
.Y(n_3700)
);

OAI21xp5_ASAP7_75t_L g3701 ( 
.A1(n_3628),
.A2(n_3257),
.B(n_3242),
.Y(n_3701)
);

AOI21xp5_ASAP7_75t_L g3702 ( 
.A1(n_3580),
.A2(n_3588),
.B(n_3612),
.Y(n_3702)
);

OAI21xp5_ASAP7_75t_L g3703 ( 
.A1(n_3596),
.A2(n_3264),
.B(n_3259),
.Y(n_3703)
);

AO21x2_ASAP7_75t_L g3704 ( 
.A1(n_3559),
.A2(n_3307),
.B(n_3394),
.Y(n_3704)
);

NOR2xp33_ASAP7_75t_R g3705 ( 
.A(n_3564),
.B(n_3483),
.Y(n_3705)
);

AND2x2_ASAP7_75t_L g3706 ( 
.A(n_3565),
.B(n_2937),
.Y(n_3706)
);

BUFx6f_ASAP7_75t_L g3707 ( 
.A(n_3631),
.Y(n_3707)
);

AO32x1_ASAP7_75t_L g3708 ( 
.A1(n_3603),
.A2(n_3521),
.A3(n_3135),
.B1(n_3136),
.B2(n_3122),
.Y(n_3708)
);

INVx4_ASAP7_75t_L g3709 ( 
.A(n_3645),
.Y(n_3709)
);

AOI221xp5_ASAP7_75t_L g3710 ( 
.A1(n_3595),
.A2(n_3493),
.B1(n_3036),
.B2(n_3477),
.C(n_3396),
.Y(n_3710)
);

NOR2x1_ASAP7_75t_SL g3711 ( 
.A(n_3594),
.B(n_3646),
.Y(n_3711)
);

NOR2x1_ASAP7_75t_L g3712 ( 
.A(n_3657),
.B(n_3621),
.Y(n_3712)
);

AND2x2_ASAP7_75t_L g3713 ( 
.A(n_3663),
.B(n_3626),
.Y(n_3713)
);

INVx2_ASAP7_75t_L g3714 ( 
.A(n_3684),
.Y(n_3714)
);

AND2x4_ASAP7_75t_L g3715 ( 
.A(n_3683),
.B(n_3603),
.Y(n_3715)
);

INVx2_ASAP7_75t_L g3716 ( 
.A(n_3696),
.Y(n_3716)
);

AOI22xp33_ASAP7_75t_L g3717 ( 
.A1(n_3700),
.A2(n_3612),
.B1(n_3574),
.B2(n_3649),
.Y(n_3717)
);

NOR2xp33_ASAP7_75t_L g3718 ( 
.A(n_3658),
.B(n_3645),
.Y(n_3718)
);

AND2x2_ASAP7_75t_L g3719 ( 
.A(n_3680),
.B(n_3630),
.Y(n_3719)
);

OAI22xp5_ASAP7_75t_L g3720 ( 
.A1(n_3656),
.A2(n_3676),
.B1(n_3669),
.B2(n_3675),
.Y(n_3720)
);

INVx1_ASAP7_75t_L g3721 ( 
.A(n_3692),
.Y(n_3721)
);

AOI22xp5_ASAP7_75t_L g3722 ( 
.A1(n_3664),
.A2(n_3638),
.B1(n_3643),
.B2(n_3560),
.Y(n_3722)
);

AND2x4_ASAP7_75t_L g3723 ( 
.A(n_3711),
.B(n_3604),
.Y(n_3723)
);

NAND2xp5_ASAP7_75t_SL g3724 ( 
.A(n_3659),
.B(n_3647),
.Y(n_3724)
);

INVx2_ASAP7_75t_SL g3725 ( 
.A(n_3705),
.Y(n_3725)
);

NAND2xp5_ASAP7_75t_L g3726 ( 
.A(n_3706),
.B(n_3573),
.Y(n_3726)
);

INVx2_ASAP7_75t_L g3727 ( 
.A(n_3655),
.Y(n_3727)
);

NAND2xp5_ASAP7_75t_L g3728 ( 
.A(n_3682),
.B(n_3575),
.Y(n_3728)
);

INVx1_ASAP7_75t_L g3729 ( 
.A(n_3679),
.Y(n_3729)
);

INVx2_ASAP7_75t_L g3730 ( 
.A(n_3685),
.Y(n_3730)
);

INVx1_ASAP7_75t_L g3731 ( 
.A(n_3690),
.Y(n_3731)
);

HB1xp67_ASAP7_75t_L g3732 ( 
.A(n_3662),
.Y(n_3732)
);

INVx1_ASAP7_75t_L g3733 ( 
.A(n_3665),
.Y(n_3733)
);

INVx2_ASAP7_75t_SL g3734 ( 
.A(n_3660),
.Y(n_3734)
);

AND2x2_ASAP7_75t_L g3735 ( 
.A(n_3691),
.B(n_3583),
.Y(n_3735)
);

AND2x2_ASAP7_75t_L g3736 ( 
.A(n_3672),
.B(n_3642),
.Y(n_3736)
);

OR2x2_ASAP7_75t_L g3737 ( 
.A(n_3667),
.B(n_3566),
.Y(n_3737)
);

NAND2xp5_ASAP7_75t_L g3738 ( 
.A(n_3673),
.B(n_3644),
.Y(n_3738)
);

AND2x2_ASAP7_75t_L g3739 ( 
.A(n_3661),
.B(n_3644),
.Y(n_3739)
);

BUFx2_ASAP7_75t_L g3740 ( 
.A(n_3709),
.Y(n_3740)
);

INVx1_ASAP7_75t_L g3741 ( 
.A(n_3686),
.Y(n_3741)
);

OAI22xp5_ASAP7_75t_L g3742 ( 
.A1(n_3654),
.A2(n_3578),
.B1(n_3568),
.B2(n_3569),
.Y(n_3742)
);

INVx1_ASAP7_75t_L g3743 ( 
.A(n_3686),
.Y(n_3743)
);

HB1xp67_ASAP7_75t_L g3744 ( 
.A(n_3707),
.Y(n_3744)
);

INVx1_ASAP7_75t_L g3745 ( 
.A(n_3687),
.Y(n_3745)
);

INVx2_ASAP7_75t_L g3746 ( 
.A(n_3677),
.Y(n_3746)
);

AND2x2_ASAP7_75t_L g3747 ( 
.A(n_3671),
.B(n_3576),
.Y(n_3747)
);

INVx1_ASAP7_75t_L g3748 ( 
.A(n_3666),
.Y(n_3748)
);

INVx2_ASAP7_75t_L g3749 ( 
.A(n_3688),
.Y(n_3749)
);

INVx1_ASAP7_75t_L g3750 ( 
.A(n_3653),
.Y(n_3750)
);

AND2x2_ASAP7_75t_L g3751 ( 
.A(n_3693),
.B(n_3577),
.Y(n_3751)
);

NAND4xp25_ASAP7_75t_SL g3752 ( 
.A(n_3750),
.B(n_3670),
.C(n_3653),
.D(n_3702),
.Y(n_3752)
);

INVx3_ASAP7_75t_L g3753 ( 
.A(n_3723),
.Y(n_3753)
);

INVx2_ASAP7_75t_L g3754 ( 
.A(n_3730),
.Y(n_3754)
);

AND2x2_ASAP7_75t_L g3755 ( 
.A(n_3732),
.B(n_3670),
.Y(n_3755)
);

INVxp67_ASAP7_75t_L g3756 ( 
.A(n_3740),
.Y(n_3756)
);

AOI22xp5_ASAP7_75t_L g3757 ( 
.A1(n_3720),
.A2(n_3697),
.B1(n_3698),
.B2(n_3703),
.Y(n_3757)
);

AOI22xp33_ASAP7_75t_L g3758 ( 
.A1(n_3720),
.A2(n_3710),
.B1(n_3681),
.B2(n_3701),
.Y(n_3758)
);

AND2x2_ASAP7_75t_SL g3759 ( 
.A(n_3723),
.B(n_3678),
.Y(n_3759)
);

AOI21xp5_ASAP7_75t_SL g3760 ( 
.A1(n_3742),
.A2(n_3695),
.B(n_3674),
.Y(n_3760)
);

AOI221xp5_ASAP7_75t_L g3761 ( 
.A1(n_3741),
.A2(n_3699),
.B1(n_3694),
.B2(n_3689),
.C(n_3668),
.Y(n_3761)
);

NAND3xp33_ASAP7_75t_L g3762 ( 
.A(n_3743),
.B(n_3554),
.C(n_3635),
.Y(n_3762)
);

INVx2_ASAP7_75t_L g3763 ( 
.A(n_3714),
.Y(n_3763)
);

INVx1_ASAP7_75t_L g3764 ( 
.A(n_3729),
.Y(n_3764)
);

INVx5_ASAP7_75t_L g3765 ( 
.A(n_3725),
.Y(n_3765)
);

BUFx2_ASAP7_75t_L g3766 ( 
.A(n_3712),
.Y(n_3766)
);

AND2x2_ASAP7_75t_L g3767 ( 
.A(n_3736),
.B(n_3739),
.Y(n_3767)
);

AND2x2_ASAP7_75t_L g3768 ( 
.A(n_3713),
.B(n_3652),
.Y(n_3768)
);

INVx2_ASAP7_75t_L g3769 ( 
.A(n_3716),
.Y(n_3769)
);

INVx1_ASAP7_75t_SL g3770 ( 
.A(n_3744),
.Y(n_3770)
);

OAI221xp5_ASAP7_75t_L g3771 ( 
.A1(n_3718),
.A2(n_3515),
.B1(n_3289),
.B2(n_3288),
.C(n_3505),
.Y(n_3771)
);

AND2x2_ASAP7_75t_L g3772 ( 
.A(n_3727),
.B(n_3608),
.Y(n_3772)
);

NOR3xp33_ASAP7_75t_SL g3773 ( 
.A(n_3718),
.B(n_3349),
.C(n_2999),
.Y(n_3773)
);

AOI221xp5_ASAP7_75t_SL g3774 ( 
.A1(n_3717),
.A2(n_3747),
.B1(n_3738),
.B2(n_3749),
.C(n_3733),
.Y(n_3774)
);

AO21x2_ASAP7_75t_L g3775 ( 
.A1(n_3746),
.A2(n_3615),
.B(n_3567),
.Y(n_3775)
);

NAND2xp5_ASAP7_75t_L g3776 ( 
.A(n_3728),
.B(n_3590),
.Y(n_3776)
);

OAI33xp33_ASAP7_75t_L g3777 ( 
.A1(n_3738),
.A2(n_3592),
.A3(n_3593),
.B1(n_3590),
.B2(n_3602),
.B3(n_3598),
.Y(n_3777)
);

INVx3_ASAP7_75t_L g3778 ( 
.A(n_3715),
.Y(n_3778)
);

OAI221xp5_ASAP7_75t_L g3779 ( 
.A1(n_3717),
.A2(n_3007),
.B1(n_3058),
.B2(n_3003),
.C(n_2997),
.Y(n_3779)
);

NAND2xp5_ASAP7_75t_L g3780 ( 
.A(n_3728),
.B(n_3593),
.Y(n_3780)
);

INVx1_ASAP7_75t_SL g3781 ( 
.A(n_3744),
.Y(n_3781)
);

NOR3xp33_ASAP7_75t_L g3782 ( 
.A(n_3748),
.B(n_3745),
.C(n_3724),
.Y(n_3782)
);

INVx1_ASAP7_75t_L g3783 ( 
.A(n_3721),
.Y(n_3783)
);

AOI22xp33_ASAP7_75t_SL g3784 ( 
.A1(n_3734),
.A2(n_3704),
.B1(n_3610),
.B2(n_3613),
.Y(n_3784)
);

AND2x2_ASAP7_75t_L g3785 ( 
.A(n_3759),
.B(n_3751),
.Y(n_3785)
);

NOR2xp33_ASAP7_75t_L g3786 ( 
.A(n_3757),
.B(n_3731),
.Y(n_3786)
);

NOR2xp33_ASAP7_75t_L g3787 ( 
.A(n_3757),
.B(n_3722),
.Y(n_3787)
);

AND2x2_ASAP7_75t_L g3788 ( 
.A(n_3753),
.B(n_3719),
.Y(n_3788)
);

NOR2xp33_ASAP7_75t_L g3789 ( 
.A(n_3766),
.B(n_3735),
.Y(n_3789)
);

INVx2_ASAP7_75t_L g3790 ( 
.A(n_3754),
.Y(n_3790)
);

AND2x2_ASAP7_75t_L g3791 ( 
.A(n_3778),
.B(n_3755),
.Y(n_3791)
);

NAND2xp5_ASAP7_75t_L g3792 ( 
.A(n_3774),
.B(n_3726),
.Y(n_3792)
);

INVx1_ASAP7_75t_SL g3793 ( 
.A(n_3765),
.Y(n_3793)
);

INVx3_ASAP7_75t_L g3794 ( 
.A(n_3770),
.Y(n_3794)
);

INVxp67_ASAP7_75t_SL g3795 ( 
.A(n_3762),
.Y(n_3795)
);

NAND2xp5_ASAP7_75t_L g3796 ( 
.A(n_3774),
.B(n_3761),
.Y(n_3796)
);

NAND2xp5_ASAP7_75t_L g3797 ( 
.A(n_3764),
.B(n_3758),
.Y(n_3797)
);

NAND2xp5_ASAP7_75t_L g3798 ( 
.A(n_3796),
.B(n_3786),
.Y(n_3798)
);

AND2x2_ASAP7_75t_L g3799 ( 
.A(n_3791),
.B(n_3756),
.Y(n_3799)
);

INVx3_ASAP7_75t_L g3800 ( 
.A(n_3793),
.Y(n_3800)
);

AOI22xp5_ASAP7_75t_L g3801 ( 
.A1(n_3787),
.A2(n_3752),
.B1(n_3782),
.B2(n_3777),
.Y(n_3801)
);

AND2x4_ASAP7_75t_L g3802 ( 
.A(n_3785),
.B(n_3781),
.Y(n_3802)
);

AOI221xp5_ASAP7_75t_L g3803 ( 
.A1(n_3787),
.A2(n_3760),
.B1(n_3762),
.B2(n_3771),
.C(n_3783),
.Y(n_3803)
);

NAND2xp5_ASAP7_75t_L g3804 ( 
.A(n_3797),
.B(n_3792),
.Y(n_3804)
);

INVx2_ASAP7_75t_L g3805 ( 
.A(n_3794),
.Y(n_3805)
);

AND2x2_ASAP7_75t_L g3806 ( 
.A(n_3788),
.B(n_3768),
.Y(n_3806)
);

INVx1_ASAP7_75t_L g3807 ( 
.A(n_3790),
.Y(n_3807)
);

O2A1O1Ixp5_ASAP7_75t_R g3808 ( 
.A1(n_3795),
.A2(n_3776),
.B(n_3780),
.C(n_3784),
.Y(n_3808)
);

NAND2x1p5_ASAP7_75t_L g3809 ( 
.A(n_3789),
.B(n_3737),
.Y(n_3809)
);

AND2x2_ASAP7_75t_L g3810 ( 
.A(n_3795),
.B(n_3767),
.Y(n_3810)
);

NAND2x1p5_ASAP7_75t_L g3811 ( 
.A(n_3800),
.B(n_3772),
.Y(n_3811)
);

OAI222xp33_ASAP7_75t_L g3812 ( 
.A1(n_3801),
.A2(n_3763),
.B1(n_3769),
.B2(n_3779),
.C1(n_3773),
.C2(n_3602),
.Y(n_3812)
);

NOR2xp33_ASAP7_75t_L g3813 ( 
.A(n_3804),
.B(n_615),
.Y(n_3813)
);

NAND2xp5_ASAP7_75t_L g3814 ( 
.A(n_3810),
.B(n_3775),
.Y(n_3814)
);

NOR3xp33_ASAP7_75t_L g3815 ( 
.A(n_3803),
.B(n_3149),
.C(n_3071),
.Y(n_3815)
);

AO22x1_ASAP7_75t_L g3816 ( 
.A1(n_3808),
.A2(n_3708),
.B1(n_3598),
.B2(n_3640),
.Y(n_3816)
);

INVx1_ASAP7_75t_L g3817 ( 
.A(n_3799),
.Y(n_3817)
);

AND2x2_ASAP7_75t_L g3818 ( 
.A(n_3802),
.B(n_3640),
.Y(n_3818)
);

INVx1_ASAP7_75t_SL g3819 ( 
.A(n_3809),
.Y(n_3819)
);

INVx1_ASAP7_75t_SL g3820 ( 
.A(n_3805),
.Y(n_3820)
);

AND2x2_ASAP7_75t_L g3821 ( 
.A(n_3806),
.B(n_3243),
.Y(n_3821)
);

NAND2xp5_ASAP7_75t_L g3822 ( 
.A(n_3807),
.B(n_3200),
.Y(n_3822)
);

NAND2xp5_ASAP7_75t_L g3823 ( 
.A(n_3798),
.B(n_3251),
.Y(n_3823)
);

AOI22xp5_ASAP7_75t_L g3824 ( 
.A1(n_3819),
.A2(n_3322),
.B1(n_3336),
.B2(n_3327),
.Y(n_3824)
);

INVx1_ASAP7_75t_SL g3825 ( 
.A(n_3820),
.Y(n_3825)
);

OR2x6_ASAP7_75t_L g3826 ( 
.A(n_3811),
.B(n_3228),
.Y(n_3826)
);

NAND2xp5_ASAP7_75t_L g3827 ( 
.A(n_3817),
.B(n_616),
.Y(n_3827)
);

AOI222xp33_ASAP7_75t_L g3828 ( 
.A1(n_3812),
.A2(n_3110),
.B1(n_2852),
.B2(n_2785),
.C1(n_617),
.C2(n_618),
.Y(n_3828)
);

O2A1O1Ixp33_ASAP7_75t_L g3829 ( 
.A1(n_3813),
.A2(n_3082),
.B(n_3089),
.C(n_3080),
.Y(n_3829)
);

AOI21xp5_ASAP7_75t_L g3830 ( 
.A1(n_3823),
.A2(n_2852),
.B(n_2785),
.Y(n_3830)
);

AOI21xp5_ASAP7_75t_L g3831 ( 
.A1(n_3814),
.A2(n_2842),
.B(n_2823),
.Y(n_3831)
);

AOI211xp5_ASAP7_75t_L g3832 ( 
.A1(n_3825),
.A2(n_3815),
.B(n_3816),
.C(n_3818),
.Y(n_3832)
);

AND2x2_ASAP7_75t_L g3833 ( 
.A(n_3826),
.B(n_3821),
.Y(n_3833)
);

OR2x2_ASAP7_75t_L g3834 ( 
.A(n_3827),
.B(n_3822),
.Y(n_3834)
);

INVx1_ASAP7_75t_SL g3835 ( 
.A(n_3831),
.Y(n_3835)
);

OAI21xp5_ASAP7_75t_L g3836 ( 
.A1(n_3828),
.A2(n_620),
.B(n_621),
.Y(n_3836)
);

NOR4xp25_ASAP7_75t_L g3837 ( 
.A(n_3829),
.B(n_624),
.C(n_622),
.D(n_623),
.Y(n_3837)
);

OAI21xp5_ASAP7_75t_L g3838 ( 
.A1(n_3830),
.A2(n_3824),
.B(n_624),
.Y(n_3838)
);

INVx1_ASAP7_75t_SL g3839 ( 
.A(n_3825),
.Y(n_3839)
);

OAI221xp5_ASAP7_75t_L g3840 ( 
.A1(n_3837),
.A2(n_3832),
.B1(n_3838),
.B2(n_3836),
.C(n_3835),
.Y(n_3840)
);

AND2x2_ASAP7_75t_L g3841 ( 
.A(n_3833),
.B(n_628),
.Y(n_3841)
);

OAI22xp5_ASAP7_75t_L g3842 ( 
.A1(n_3834),
.A2(n_2864),
.B1(n_2895),
.B2(n_2849),
.Y(n_3842)
);

INVx1_ASAP7_75t_SL g3843 ( 
.A(n_3839),
.Y(n_3843)
);

NOR3xp33_ASAP7_75t_SL g3844 ( 
.A(n_3840),
.B(n_637),
.C(n_638),
.Y(n_3844)
);

AND2x2_ASAP7_75t_L g3845 ( 
.A(n_3841),
.B(n_638),
.Y(n_3845)
);

NOR2x1_ASAP7_75t_L g3846 ( 
.A(n_3842),
.B(n_641),
.Y(n_3846)
);

AND2x2_ASAP7_75t_L g3847 ( 
.A(n_3843),
.B(n_644),
.Y(n_3847)
);

INVx1_ASAP7_75t_L g3848 ( 
.A(n_3847),
.Y(n_3848)
);

OAI211xp5_ASAP7_75t_SL g3849 ( 
.A1(n_3844),
.A2(n_651),
.B(n_649),
.C(n_650),
.Y(n_3849)
);

INVx3_ASAP7_75t_SL g3850 ( 
.A(n_3845),
.Y(n_3850)
);

OAI222xp33_ASAP7_75t_L g3851 ( 
.A1(n_3846),
.A2(n_705),
.B1(n_707),
.B2(n_703),
.C1(n_704),
.C2(n_706),
.Y(n_3851)
);

AND2x2_ASAP7_75t_L g3852 ( 
.A(n_3850),
.B(n_708),
.Y(n_3852)
);

AOI221xp5_ASAP7_75t_SL g3853 ( 
.A1(n_3848),
.A2(n_712),
.B1(n_710),
.B2(n_711),
.C(n_713),
.Y(n_3853)
);

AOI22xp5_ASAP7_75t_L g3854 ( 
.A1(n_3849),
.A2(n_3113),
.B1(n_3069),
.B2(n_715),
.Y(n_3854)
);

XNOR2x1_ASAP7_75t_L g3855 ( 
.A(n_3851),
.B(n_717),
.Y(n_3855)
);

INVx1_ASAP7_75t_L g3856 ( 
.A(n_3852),
.Y(n_3856)
);

XOR2x2_ASAP7_75t_L g3857 ( 
.A(n_3855),
.B(n_719),
.Y(n_3857)
);

NAND4xp75_ASAP7_75t_L g3858 ( 
.A(n_3853),
.B(n_723),
.C(n_721),
.D(n_722),
.Y(n_3858)
);

INVx1_ASAP7_75t_L g3859 ( 
.A(n_3854),
.Y(n_3859)
);

INVx1_ASAP7_75t_L g3860 ( 
.A(n_3858),
.Y(n_3860)
);

NOR2x2_ASAP7_75t_L g3861 ( 
.A(n_3857),
.B(n_731),
.Y(n_3861)
);

NOR2x1_ASAP7_75t_L g3862 ( 
.A(n_3859),
.B(n_732),
.Y(n_3862)
);

AOI22xp5_ASAP7_75t_L g3863 ( 
.A1(n_3860),
.A2(n_3856),
.B1(n_734),
.B2(n_732),
.Y(n_3863)
);

OAI221xp5_ASAP7_75t_R g3864 ( 
.A1(n_3861),
.A2(n_735),
.B1(n_733),
.B2(n_734),
.C(n_736),
.Y(n_3864)
);

INVx1_ASAP7_75t_L g3865 ( 
.A(n_3862),
.Y(n_3865)
);

INVx2_ASAP7_75t_L g3866 ( 
.A(n_3865),
.Y(n_3866)
);

OAI22x1_ASAP7_75t_L g3867 ( 
.A1(n_3863),
.A2(n_740),
.B1(n_737),
.B2(n_738),
.Y(n_3867)
);

AO22x2_ASAP7_75t_L g3868 ( 
.A1(n_3864),
.A2(n_740),
.B1(n_737),
.B2(n_738),
.Y(n_3868)
);

INVx2_ASAP7_75t_L g3869 ( 
.A(n_3866),
.Y(n_3869)
);

AOI21xp5_ASAP7_75t_L g3870 ( 
.A1(n_3869),
.A2(n_3868),
.B(n_3867),
.Y(n_3870)
);

NAND2xp5_ASAP7_75t_SL g3871 ( 
.A(n_3870),
.B(n_742),
.Y(n_3871)
);

NOR3xp33_ASAP7_75t_L g3872 ( 
.A(n_3871),
.B(n_742),
.C(n_743),
.Y(n_3872)
);

NOR2xp33_ASAP7_75t_L g3873 ( 
.A(n_3871),
.B(n_744),
.Y(n_3873)
);

AO21x2_ASAP7_75t_L g3874 ( 
.A1(n_3873),
.A2(n_747),
.B(n_748),
.Y(n_3874)
);

OAI22xp33_ASAP7_75t_L g3875 ( 
.A1(n_3872),
.A2(n_749),
.B1(n_747),
.B2(n_748),
.Y(n_3875)
);

NOR2x1_ASAP7_75t_L g3876 ( 
.A(n_3874),
.B(n_3875),
.Y(n_3876)
);

OAI221xp5_ASAP7_75t_R g3877 ( 
.A1(n_3876),
.A2(n_756),
.B1(n_754),
.B2(n_755),
.C(n_757),
.Y(n_3877)
);

AOI211xp5_ASAP7_75t_L g3878 ( 
.A1(n_3877),
.A2(n_759),
.B(n_755),
.C(n_757),
.Y(n_3878)
);


endmodule