module fake_jpeg_18645_n_36 (n_3, n_2, n_1, n_0, n_4, n_5, n_36);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_36;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx1_ASAP7_75t_L g6 ( 
.A(n_1),
.Y(n_6)
);

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_0),
.Y(n_7)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_4),
.B(n_5),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_5),
.B(n_0),
.Y(n_10)
);

CKINVDCx16_ASAP7_75t_R g11 ( 
.A(n_4),
.Y(n_11)
);

INVx3_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx4_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx4_ASAP7_75t_SL g14 ( 
.A(n_12),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_14),
.B(n_18),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g15 ( 
.A1(n_12),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_15),
.A2(n_17),
.B1(n_11),
.B2(n_6),
.Y(n_22)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_16),
.B(n_6),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g17 ( 
.A(n_7),
.B(n_10),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_17),
.B(n_9),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_20),
.B(n_15),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_22),
.B(n_23),
.Y(n_25)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_22),
.B(n_17),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_24),
.B(n_26),
.Y(n_30)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_27),
.Y(n_28)
);

AO21x1_ASAP7_75t_L g29 ( 
.A1(n_25),
.A2(n_20),
.B(n_16),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_29),
.B(n_14),
.Y(n_32)
);

XOR2xp5_ASAP7_75t_L g31 ( 
.A(n_30),
.B(n_24),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_32),
.C(n_28),
.Y(n_34)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_32),
.Y(n_33)
);

AOI322xp5_ASAP7_75t_L g35 ( 
.A1(n_33),
.A2(n_34),
.A3(n_8),
.B1(n_29),
.B2(n_21),
.C1(n_18),
.C2(n_2),
.Y(n_35)
);

XOR2xp5_ASAP7_75t_L g36 ( 
.A(n_35),
.B(n_8),
.Y(n_36)
);


endmodule