module fake_jpeg_18912_n_231 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_231);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_231;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_2),
.B(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_0),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_43),
.Y(n_47)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_15),
.Y(n_40)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_27),
.Y(n_42)
);

OAI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_42),
.A2(n_23),
.B1(n_30),
.B2(n_28),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_0),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_41),
.A2(n_42),
.B1(n_40),
.B2(n_31),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_44),
.A2(n_56),
.B1(n_23),
.B2(n_19),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_43),
.A2(n_16),
.B1(n_27),
.B2(n_25),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_45),
.A2(n_20),
.B1(n_19),
.B2(n_16),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_25),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_38),
.A2(n_26),
.B1(n_30),
.B2(n_28),
.Y(n_56)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_58),
.Y(n_61)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_61),
.Y(n_104)
);

AO22x2_ASAP7_75t_L g62 ( 
.A1(n_57),
.A2(n_35),
.B1(n_39),
.B2(n_34),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_62),
.A2(n_83),
.B1(n_90),
.B2(n_24),
.Y(n_98)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_63),
.Y(n_97)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_64),
.Y(n_121)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_65),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_47),
.B(n_36),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_66),
.B(n_69),
.Y(n_96)
);

OAI21xp33_ASAP7_75t_SL g119 ( 
.A1(n_67),
.A2(n_75),
.B(n_3),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_51),
.B(n_37),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_68),
.B(n_74),
.Y(n_112)
);

OA22x2_ASAP7_75t_SL g70 ( 
.A1(n_45),
.A2(n_34),
.B1(n_33),
.B2(n_21),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_70),
.B(n_80),
.Y(n_107)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_71),
.B(n_72),
.Y(n_106)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_32),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_53),
.A2(n_16),
.B1(n_33),
.B2(n_22),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_21),
.Y(n_76)
);

FAx1_ASAP7_75t_SL g110 ( 
.A(n_76),
.B(n_78),
.CI(n_82),
.CON(n_110),
.SN(n_110)
);

A2O1A1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_47),
.A2(n_21),
.B(n_32),
.C(n_22),
.Y(n_78)
);

CKINVDCx12_ASAP7_75t_R g79 ( 
.A(n_55),
.Y(n_79)
);

INVx13_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_59),
.B(n_20),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_81),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_59),
.B(n_21),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_86),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_60),
.B(n_17),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_87),
.B(n_91),
.Y(n_113)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_52),
.A2(n_18),
.B1(n_17),
.B2(n_24),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_49),
.B(n_17),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

INVx13_ASAP7_75t_L g117 ( 
.A(n_92),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_93),
.Y(n_102)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_1),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_47),
.B(n_18),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_3),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_98),
.A2(n_89),
.B1(n_84),
.B2(n_85),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_95),
.A2(n_76),
.B1(n_70),
.B2(n_67),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_101),
.A2(n_75),
.B1(n_89),
.B2(n_86),
.Y(n_143)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_70),
.A2(n_24),
.B1(n_18),
.B2(n_4),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_108),
.A2(n_82),
.B1(n_93),
.B2(n_62),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_109),
.B(n_6),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_78),
.B(n_1),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_111),
.B(n_120),
.Y(n_130)
);

AOI22x1_ASAP7_75t_L g116 ( 
.A1(n_62),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_116)
);

OA22x2_ASAP7_75t_L g129 ( 
.A1(n_116),
.A2(n_119),
.B1(n_114),
.B2(n_111),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_118),
.A2(n_102),
.B1(n_110),
.B2(n_114),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_62),
.B(n_5),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_122),
.A2(n_126),
.B1(n_103),
.B2(n_77),
.Y(n_160)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_100),
.Y(n_123)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_123),
.Y(n_153)
);

AND2x2_ASAP7_75t_SL g124 ( 
.A(n_107),
.B(n_77),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_124),
.A2(n_129),
.B(n_135),
.Y(n_146)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_100),
.Y(n_125)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_125),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_107),
.A2(n_120),
.B1(n_101),
.B2(n_98),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_106),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_127),
.B(n_131),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_113),
.B(n_63),
.Y(n_128)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_128),
.Y(n_162)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_97),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_97),
.Y(n_132)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_132),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_133),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_104),
.Y(n_134)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_134),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_110),
.B(n_73),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_104),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_136),
.A2(n_117),
.B(n_99),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_137),
.B(n_139),
.Y(n_147)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_121),
.Y(n_138)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_138),
.Y(n_156)
);

NAND3xp33_ASAP7_75t_SL g139 ( 
.A(n_110),
.B(n_96),
.C(n_112),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_121),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_140),
.B(n_141),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_99),
.B(n_105),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_109),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_142),
.B(n_7),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_143),
.A2(n_144),
.B1(n_124),
.B2(n_135),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_126),
.B(n_118),
.C(n_102),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_145),
.B(n_157),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_148),
.A2(n_154),
.B1(n_158),
.B2(n_136),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_143),
.A2(n_116),
.B1(n_118),
.B2(n_115),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_133),
.B(n_116),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_124),
.A2(n_115),
.B1(n_103),
.B2(n_84),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_160),
.B(n_163),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_161),
.A2(n_146),
.B(n_158),
.Y(n_174)
);

A2O1A1Ixp33_ASAP7_75t_L g163 ( 
.A1(n_130),
.A2(n_129),
.B(n_135),
.C(n_122),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_164),
.B(n_140),
.Y(n_176)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_156),
.Y(n_165)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_165),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_156),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_166),
.B(n_173),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_168),
.A2(n_175),
.B1(n_152),
.B2(n_163),
.Y(n_186)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_149),
.Y(n_169)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_169),
.Y(n_187)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_149),
.Y(n_170)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_170),
.Y(n_190)
);

BUFx5_ASAP7_75t_L g171 ( 
.A(n_150),
.Y(n_171)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_171),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_151),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_174),
.B(n_176),
.Y(n_188)
);

A2O1A1Ixp33_ASAP7_75t_SL g175 ( 
.A1(n_148),
.A2(n_129),
.B(n_130),
.C(n_138),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_150),
.Y(n_177)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_177),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_151),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_178),
.B(n_180),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_145),
.A2(n_129),
.B1(n_125),
.B2(n_123),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_179),
.B(n_146),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_147),
.B(n_14),
.Y(n_180)
);

NOR3xp33_ASAP7_75t_SL g182 ( 
.A(n_175),
.B(n_155),
.C(n_147),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_182),
.B(n_154),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_183),
.B(n_191),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_186),
.B(n_175),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_167),
.B(n_157),
.C(n_162),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_189),
.B(n_179),
.C(n_174),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_167),
.B(n_152),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_194),
.B(n_183),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_195),
.B(n_196),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_182),
.B(n_171),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_181),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_197),
.B(n_199),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_188),
.A2(n_172),
.B(n_175),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_198),
.A2(n_204),
.B(n_161),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_189),
.B(n_168),
.C(n_172),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_201),
.A2(n_199),
.B1(n_202),
.B2(n_194),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_187),
.B(n_165),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_202),
.B(n_203),
.Y(n_209)
);

INVx13_ASAP7_75t_L g203 ( 
.A(n_185),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_192),
.B(n_177),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_201),
.A2(n_191),
.B1(n_186),
.B2(n_184),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_205),
.A2(n_212),
.B1(n_200),
.B2(n_170),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_207),
.B(n_200),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_210),
.B(n_211),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_198),
.A2(n_193),
.B(n_190),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_214),
.B(n_216),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_215),
.B(n_218),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_212),
.B(n_169),
.C(n_159),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_210),
.A2(n_206),
.B1(n_205),
.B2(n_208),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_217),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_209),
.B(n_153),
.C(n_164),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_213),
.A2(n_203),
.B(n_132),
.Y(n_220)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_220),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_221),
.Y(n_223)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_223),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_222),
.B(n_216),
.Y(n_225)
);

AOI322xp5_ASAP7_75t_L g227 ( 
.A1(n_225),
.A2(n_219),
.A3(n_213),
.B1(n_117),
.B2(n_131),
.C1(n_7),
.C2(n_10),
.Y(n_227)
);

AOI322xp5_ASAP7_75t_L g228 ( 
.A1(n_227),
.A2(n_224),
.A3(n_225),
.B1(n_9),
.B2(n_11),
.C1(n_7),
.C2(n_8),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_226),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_229),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_230),
.B(n_8),
.C(n_9),
.Y(n_231)
);


endmodule