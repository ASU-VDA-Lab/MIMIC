module fake_netlist_1_11472_n_37 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_37);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_37;
wire n_20;
wire n_36;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
BUFx6f_ASAP7_75t_L g14 ( .A(n_11), .Y(n_14) );
INVx3_ASAP7_75t_L g15 ( .A(n_0), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_5), .Y(n_16) );
INVx2_ASAP7_75t_L g17 ( .A(n_5), .Y(n_17) );
BUFx2_ASAP7_75t_L g18 ( .A(n_4), .Y(n_18) );
BUFx6f_ASAP7_75t_L g19 ( .A(n_8), .Y(n_19) );
INVx2_ASAP7_75t_L g20 ( .A(n_12), .Y(n_20) );
NAND2xp5_ASAP7_75t_L g21 ( .A(n_18), .B(n_0), .Y(n_21) );
BUFx8_ASAP7_75t_L g22 ( .A(n_18), .Y(n_22) );
AOI22xp5_ASAP7_75t_L g23 ( .A1(n_15), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_23) );
BUFx6f_ASAP7_75t_L g24 ( .A(n_21), .Y(n_24) );
AOI21x1_ASAP7_75t_L g25 ( .A1(n_23), .A2(n_20), .B(n_17), .Y(n_25) );
OR2x2_ASAP7_75t_L g26 ( .A(n_24), .B(n_22), .Y(n_26) );
OAI33xp33_ASAP7_75t_L g27 ( .A1(n_26), .A2(n_16), .A3(n_17), .B1(n_25), .B2(n_20), .B3(n_24), .Y(n_27) );
NAND2xp5_ASAP7_75t_L g28 ( .A(n_27), .B(n_24), .Y(n_28) );
NAND2xp5_ASAP7_75t_L g29 ( .A(n_27), .B(n_24), .Y(n_29) );
AOI22xp5_ASAP7_75t_L g30 ( .A1(n_28), .A2(n_29), .B1(n_15), .B2(n_19), .Y(n_30) );
NAND4xp75_ASAP7_75t_L g31 ( .A(n_28), .B(n_15), .C(n_2), .D(n_3), .Y(n_31) );
NOR2x1_ASAP7_75t_L g32 ( .A(n_31), .B(n_19), .Y(n_32) );
OR4x2_ASAP7_75t_L g33 ( .A(n_30), .B(n_1), .C(n_4), .D(n_6), .Y(n_33) );
XNOR2xp5_ASAP7_75t_L g34 ( .A(n_32), .B(n_6), .Y(n_34) );
AOI22x1_ASAP7_75t_L g35 ( .A1(n_33), .A2(n_14), .B1(n_19), .B2(n_9), .Y(n_35) );
AOI222xp33_ASAP7_75t_L g36 ( .A1(n_34), .A2(n_14), .B1(n_19), .B2(n_10), .C1(n_13), .C2(n_7), .Y(n_36) );
AOI22xp5_ASAP7_75t_L g37 ( .A1(n_36), .A2(n_34), .B1(n_14), .B2(n_35), .Y(n_37) );
endmodule