module fake_jpeg_10090_n_229 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_229);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_229;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx8_ASAP7_75t_SL g27 ( 
.A(n_10),
.Y(n_27)
);

INVx6_ASAP7_75t_SL g28 ( 
.A(n_5),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_14),
.B(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_31),
.B(n_32),
.Y(n_48)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_24),
.A2(n_20),
.B1(n_18),
.B2(n_23),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_34),
.A2(n_18),
.B1(n_20),
.B2(n_28),
.Y(n_50)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_35),
.B(n_37),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_14),
.B(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_15),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_38),
.B(n_1),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_14),
.B(n_0),
.Y(n_39)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_39),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_42),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_14),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_29),
.A2(n_24),
.B1(n_23),
.B2(n_18),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_43),
.A2(n_44),
.B1(n_50),
.B2(n_20),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_L g44 ( 
.A1(n_29),
.A2(n_24),
.B1(n_23),
.B2(n_28),
.Y(n_44)
);

CKINVDCx5p33_ASAP7_75t_R g45 ( 
.A(n_37),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_45),
.Y(n_69)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_53),
.Y(n_61)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_65),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_59),
.A2(n_26),
.B1(n_45),
.B2(n_17),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_60),
.Y(n_93)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_66),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_40),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_68),
.Y(n_81)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

AO22x2_ASAP7_75t_L g71 ( 
.A1(n_42),
.A2(n_38),
.B1(n_34),
.B2(n_35),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_71),
.A2(n_35),
.B1(n_48),
.B2(n_30),
.Y(n_88)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_72),
.A2(n_58),
.B1(n_74),
.B2(n_63),
.Y(n_84)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_74),
.Y(n_86)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_75),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_71),
.A2(n_29),
.B1(n_53),
.B2(n_40),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_76),
.A2(n_80),
.B1(n_82),
.B2(n_83),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_71),
.B(n_46),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_77),
.B(n_38),
.C(n_26),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_71),
.A2(n_41),
.B1(n_57),
.B2(n_55),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_62),
.A2(n_55),
.B1(n_52),
.B2(n_46),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_73),
.A2(n_52),
.B1(n_35),
.B2(n_32),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_84),
.A2(n_90),
.B1(n_72),
.B2(n_33),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_61),
.B(n_48),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_38),
.Y(n_105)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_87),
.B(n_91),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_88),
.A2(n_94),
.B1(n_56),
.B2(n_75),
.Y(n_100)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_68),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_65),
.A2(n_54),
.B1(n_33),
.B2(n_30),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_80),
.B(n_69),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_95),
.B(n_105),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_36),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_96),
.B(n_101),
.C(n_109),
.Y(n_126)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_99),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_100),
.A2(n_107),
.B1(n_108),
.B2(n_86),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_77),
.B(n_31),
.Y(n_101)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_102),
.Y(n_117)
);

A2O1A1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_77),
.A2(n_39),
.B(n_36),
.C(n_38),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_103),
.B(n_106),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_79),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_104),
.B(n_112),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_91),
.B(n_70),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_77),
.A2(n_33),
.B1(n_30),
.B2(n_56),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_85),
.A2(n_33),
.B1(n_56),
.B2(n_37),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_82),
.B(n_15),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_110),
.B(n_111),
.Y(n_119)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_79),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_83),
.B(n_15),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_113),
.B(n_86),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_109),
.B(n_87),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_114),
.A2(n_103),
.B(n_108),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_101),
.B(n_81),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_116),
.B(n_16),
.C(n_25),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_107),
.A2(n_81),
.B(n_94),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_118),
.A2(n_123),
.B(n_127),
.Y(n_140)
);

AND2x6_ASAP7_75t_L g120 ( 
.A(n_96),
.B(n_89),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_120),
.A2(n_131),
.B(n_95),
.Y(n_133)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_99),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_125),
.B(n_128),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_99),
.Y(n_128)
);

INVx13_ASAP7_75t_L g129 ( 
.A(n_102),
.Y(n_129)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_129),
.Y(n_144)
);

CKINVDCx14_ASAP7_75t_R g130 ( 
.A(n_97),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_130),
.B(n_97),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_104),
.A2(n_92),
.B(n_93),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_98),
.A2(n_89),
.B1(n_78),
.B2(n_93),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_132),
.A2(n_112),
.B1(n_111),
.B2(n_110),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_133),
.A2(n_138),
.B(n_146),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_116),
.B(n_98),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_134),
.B(n_135),
.C(n_141),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_126),
.B(n_105),
.Y(n_135)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_136),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_137),
.B(n_145),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_106),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_139),
.B(n_148),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_126),
.B(n_100),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_132),
.A2(n_78),
.B1(n_60),
.B2(n_22),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_142),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_120),
.B(n_10),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_143),
.B(n_118),
.Y(n_154)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_131),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_124),
.A2(n_25),
.B(n_22),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_115),
.B(n_14),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_149),
.B(n_119),
.C(n_124),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_127),
.A2(n_16),
.B1(n_21),
.B2(n_19),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_150),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_119),
.B(n_21),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_151),
.B(n_121),
.Y(n_167)
);

OR2x2_ASAP7_75t_L g152 ( 
.A(n_143),
.B(n_122),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_152),
.B(n_162),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_144),
.Y(n_153)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_153),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_154),
.B(n_166),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_SL g155 ( 
.A(n_138),
.B(n_114),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_155),
.B(n_140),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_147),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_151),
.B(n_125),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_163),
.B(n_165),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_136),
.B(n_128),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_167),
.B(n_144),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_135),
.B(n_114),
.C(n_117),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_134),
.C(n_141),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_169),
.B(n_170),
.C(n_172),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_159),
.B(n_133),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_159),
.B(n_140),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_173),
.B(n_154),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_160),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_174),
.B(n_177),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_168),
.B(n_149),
.C(n_139),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_175),
.B(n_181),
.C(n_182),
.Y(n_193)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_158),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_158),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_179),
.B(n_183),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_155),
.B(n_148),
.C(n_117),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_166),
.B(n_146),
.C(n_121),
.Y(n_182)
);

OR2x2_ASAP7_75t_L g184 ( 
.A(n_171),
.B(n_157),
.Y(n_184)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_184),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_180),
.B(n_156),
.Y(n_185)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_185),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_186),
.B(n_25),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_175),
.A2(n_161),
.B(n_164),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_189),
.B(n_190),
.C(n_191),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_181),
.A2(n_161),
.B(n_157),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_182),
.A2(n_152),
.B1(n_129),
.B2(n_150),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_173),
.A2(n_142),
.B(n_9),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_192),
.A2(n_7),
.B1(n_13),
.B2(n_3),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_170),
.B(n_25),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_194),
.B(n_176),
.C(n_25),
.Y(n_199)
);

A2O1A1Ixp33_ASAP7_75t_SL g197 ( 
.A1(n_184),
.A2(n_178),
.B(n_172),
.C(n_169),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_197),
.A2(n_203),
.B1(n_202),
.B2(n_4),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_199),
.B(n_7),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_193),
.B(n_8),
.C(n_13),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_200),
.B(n_205),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_201),
.B(n_19),
.Y(n_212)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_202),
.Y(n_209)
);

NOR3xp33_ASAP7_75t_L g204 ( 
.A(n_192),
.B(n_9),
.C(n_13),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_204),
.A2(n_11),
.B(n_12),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_193),
.B(n_7),
.C(n_12),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_198),
.A2(n_188),
.B1(n_195),
.B2(n_187),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_206),
.B(n_208),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_207),
.B(n_210),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_196),
.A2(n_187),
.B1(n_186),
.B2(n_194),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_211),
.B(n_212),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_208),
.B(n_197),
.C(n_21),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_214),
.B(n_219),
.Y(n_220)
);

OAI221xp5_ASAP7_75t_L g216 ( 
.A1(n_210),
.A2(n_197),
.B1(n_5),
.B2(n_6),
.C(n_11),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_216),
.A2(n_5),
.B(n_6),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_209),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_217),
.B(n_213),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_221),
.A2(n_223),
.B(n_220),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_222),
.B(n_215),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_218),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_224),
.B(n_225),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_226),
.A2(n_212),
.B1(n_1),
.B2(n_2),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_227),
.A2(n_1),
.B(n_2),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_2),
.Y(n_229)
);


endmodule