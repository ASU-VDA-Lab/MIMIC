module real_aes_1288_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_792;
wire n_386;
wire n_673;
wire n_635;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_545;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_815;
wire n_519;
wire n_638;
wire n_564;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_292;
wire n_539;
wire n_400;
wire n_626;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_502;
wire n_505;
wire n_434;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_785;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_L g515 ( .A(n_0), .B(n_212), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_1), .B(n_119), .Y(n_118) );
INVx1_ASAP7_75t_L g146 ( .A(n_2), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_3), .B(n_518), .Y(n_537) );
NAND2xp33_ASAP7_75t_SL g508 ( .A(n_4), .B(n_167), .Y(n_508) );
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_5), .B(n_180), .Y(n_203) );
INVx1_ASAP7_75t_L g500 ( .A(n_6), .Y(n_500) );
INVx1_ASAP7_75t_L g237 ( .A(n_7), .Y(n_237) );
CKINVDCx16_ASAP7_75t_R g119 ( .A(n_8), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g254 ( .A(n_9), .Y(n_254) );
AND2x2_ASAP7_75t_L g535 ( .A(n_10), .B(n_136), .Y(n_535) );
INVx2_ASAP7_75t_L g137 ( .A(n_11), .Y(n_137) );
CKINVDCx16_ASAP7_75t_R g112 ( .A(n_12), .Y(n_112) );
INVx1_ASAP7_75t_L g213 ( .A(n_13), .Y(n_213) );
AOI221x1_ASAP7_75t_L g503 ( .A1(n_14), .A2(n_169), .B1(n_504), .B2(n_506), .C(n_507), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g571 ( .A(n_15), .B(n_518), .Y(n_571) );
INVx1_ASAP7_75t_L g116 ( .A(n_16), .Y(n_116) );
INVx1_ASAP7_75t_L g210 ( .A(n_17), .Y(n_210) );
INVx1_ASAP7_75t_SL g158 ( .A(n_18), .Y(n_158) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_19), .B(n_161), .Y(n_183) );
AOI33xp33_ASAP7_75t_L g228 ( .A1(n_20), .A2(n_49), .A3(n_143), .B1(n_154), .B2(n_229), .B3(n_230), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_21), .A2(n_506), .B(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_22), .B(n_212), .Y(n_540) );
AOI221xp5_ASAP7_75t_SL g580 ( .A1(n_23), .A2(n_40), .B1(n_506), .B2(n_518), .C(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g247 ( .A(n_24), .Y(n_247) );
OR2x2_ASAP7_75t_L g138 ( .A(n_25), .B(n_89), .Y(n_138) );
OA21x2_ASAP7_75t_L g171 ( .A1(n_25), .A2(n_89), .B(n_137), .Y(n_171) );
INVxp67_ASAP7_75t_L g502 ( .A(n_26), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_27), .B(n_215), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g817 ( .A(n_28), .B(n_818), .Y(n_817) );
AND2x2_ASAP7_75t_L g529 ( .A(n_29), .B(n_135), .Y(n_529) );
CKINVDCx20_ASAP7_75t_R g787 ( .A(n_30), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_31), .B(n_141), .Y(n_140) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_32), .A2(n_506), .B(n_514), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_33), .B(n_215), .Y(n_582) );
AND2x2_ASAP7_75t_L g148 ( .A(n_34), .B(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g153 ( .A(n_34), .Y(n_153) );
AND2x2_ASAP7_75t_L g167 ( .A(n_34), .B(n_146), .Y(n_167) );
OR2x6_ASAP7_75t_L g114 ( .A(n_35), .B(n_115), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g249 ( .A(n_36), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_37), .B(n_141), .Y(n_274) );
AOI22xp5_ASAP7_75t_L g175 ( .A1(n_38), .A2(n_170), .B1(n_176), .B2(n_180), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_39), .B(n_185), .Y(n_184) );
AOI22xp5_ASAP7_75t_L g547 ( .A1(n_41), .A2(n_81), .B1(n_151), .B2(n_506), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_42), .B(n_161), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_43), .B(n_212), .Y(n_527) );
NAND2xp5_ASAP7_75t_SL g239 ( .A(n_44), .B(n_187), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_45), .B(n_161), .Y(n_238) );
CKINVDCx5p33_ASAP7_75t_R g179 ( .A(n_46), .Y(n_179) );
AND2x2_ASAP7_75t_L g519 ( .A(n_47), .B(n_135), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_48), .B(n_135), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_50), .B(n_161), .Y(n_278) );
CKINVDCx20_ASAP7_75t_R g426 ( .A(n_51), .Y(n_426) );
OAI22xp5_ASAP7_75t_L g814 ( .A1(n_51), .A2(n_61), .B1(n_426), .B2(n_815), .Y(n_814) );
INVx1_ASAP7_75t_L g144 ( .A(n_52), .Y(n_144) );
INVx1_ASAP7_75t_L g163 ( .A(n_52), .Y(n_163) );
AND2x2_ASAP7_75t_L g279 ( .A(n_53), .B(n_135), .Y(n_279) );
AOI221xp5_ASAP7_75t_L g235 ( .A1(n_54), .A2(n_74), .B1(n_141), .B2(n_151), .C(n_236), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_55), .B(n_141), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_56), .B(n_518), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_57), .B(n_170), .Y(n_256) );
AOI21xp5_ASAP7_75t_SL g192 ( .A1(n_58), .A2(n_151), .B(n_193), .Y(n_192) );
AND2x2_ASAP7_75t_L g556 ( .A(n_59), .B(n_135), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_60), .B(n_215), .Y(n_516) );
CKINVDCx20_ASAP7_75t_R g815 ( .A(n_61), .Y(n_815) );
INVx1_ASAP7_75t_L g206 ( .A(n_62), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_63), .B(n_212), .Y(n_554) );
AND2x2_ASAP7_75t_SL g576 ( .A(n_64), .B(n_136), .Y(n_576) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_65), .A2(n_506), .B(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g277 ( .A(n_66), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_67), .B(n_215), .Y(n_541) );
AND2x2_ASAP7_75t_SL g548 ( .A(n_68), .B(n_187), .Y(n_548) );
OAI22xp5_ASAP7_75t_L g783 ( .A1(n_69), .A2(n_100), .B1(n_784), .B2(n_785), .Y(n_783) );
CKINVDCx20_ASAP7_75t_R g784 ( .A(n_69), .Y(n_784) );
AOI21xp5_ASAP7_75t_L g275 ( .A1(n_70), .A2(n_151), .B(n_276), .Y(n_275) );
AOI221xp5_ASAP7_75t_L g101 ( .A1(n_71), .A2(n_102), .B1(n_120), .B2(n_793), .C(n_801), .Y(n_101) );
OAI22xp5_ASAP7_75t_L g812 ( .A1(n_71), .A2(n_813), .B1(n_814), .B2(n_816), .Y(n_812) );
CKINVDCx20_ASAP7_75t_R g813 ( .A(n_71), .Y(n_813) );
INVx1_ASAP7_75t_L g149 ( .A(n_72), .Y(n_149) );
INVx1_ASAP7_75t_L g165 ( .A(n_72), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_73), .B(n_141), .Y(n_231) );
AND2x2_ASAP7_75t_L g168 ( .A(n_75), .B(n_169), .Y(n_168) );
INVx1_ASAP7_75t_L g207 ( .A(n_76), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g150 ( .A1(n_77), .A2(n_151), .B(n_157), .Y(n_150) );
A2O1A1Ixp33_ASAP7_75t_L g181 ( .A1(n_78), .A2(n_151), .B(n_182), .C(n_186), .Y(n_181) );
AOI22xp5_ASAP7_75t_L g546 ( .A1(n_79), .A2(n_84), .B1(n_141), .B2(n_518), .Y(n_546) );
NAND2xp5_ASAP7_75t_SL g555 ( .A(n_80), .B(n_518), .Y(n_555) );
INVx1_ASAP7_75t_L g117 ( .A(n_82), .Y(n_117) );
AND2x2_ASAP7_75t_SL g190 ( .A(n_83), .B(n_169), .Y(n_190) );
AOI22xp5_ASAP7_75t_L g225 ( .A1(n_85), .A2(n_151), .B1(n_226), .B2(n_227), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_86), .B(n_212), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_87), .B(n_212), .Y(n_583) );
AOI21xp5_ASAP7_75t_L g551 ( .A1(n_88), .A2(n_506), .B(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g194 ( .A(n_90), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_91), .B(n_215), .Y(n_553) );
AND2x2_ASAP7_75t_L g232 ( .A(n_92), .B(n_169), .Y(n_232) );
A2O1A1Ixp33_ASAP7_75t_L g244 ( .A1(n_93), .A2(n_245), .B(n_246), .C(n_248), .Y(n_244) );
INVxp67_ASAP7_75t_L g505 ( .A(n_94), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_95), .B(n_518), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_96), .B(n_215), .Y(n_526) );
AOI21xp5_ASAP7_75t_L g572 ( .A1(n_97), .A2(n_506), .B(n_573), .Y(n_572) );
BUFx2_ASAP7_75t_SL g108 ( .A(n_98), .Y(n_108) );
BUFx2_ASAP7_75t_L g799 ( .A(n_98), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_99), .B(n_161), .Y(n_195) );
CKINVDCx20_ASAP7_75t_R g785 ( .A(n_100), .Y(n_785) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
AOI21xp5_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_109), .B(n_118), .Y(n_105) );
CKINVDCx11_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
CKINVDCx8_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
INVx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
BUFx2_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
BUFx2_ASAP7_75t_L g800 ( .A(n_111), .Y(n_800) );
BUFx3_ASAP7_75t_L g805 ( .A(n_111), .Y(n_805) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_112), .B(n_113), .Y(n_111) );
AND2x6_ASAP7_75t_SL g490 ( .A(n_112), .B(n_114), .Y(n_490) );
OR2x6_ASAP7_75t_SL g781 ( .A(n_112), .B(n_113), .Y(n_781) );
OR2x2_ASAP7_75t_L g789 ( .A(n_112), .B(n_114), .Y(n_789) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_114), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_116), .B(n_117), .Y(n_115) );
INVx2_ASAP7_75t_L g798 ( .A(n_118), .Y(n_798) );
OR2x2_ASAP7_75t_SL g821 ( .A(n_118), .B(n_799), .Y(n_821) );
NAND2xp5_ASAP7_75t_SL g120 ( .A(n_121), .B(n_790), .Y(n_120) );
AOI21xp33_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_782), .B(n_786), .Y(n_121) );
OAI22x1_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_489), .B1(n_491), .B2(n_779), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
OAI22xp5_ASAP7_75t_L g791 ( .A1(n_124), .A2(n_489), .B1(n_492), .B2(n_792), .Y(n_791) );
AND3x1_ASAP7_75t_L g124 ( .A(n_125), .B(n_483), .C(n_486), .Y(n_124) );
NAND5xp2_ASAP7_75t_L g125 ( .A(n_126), .B(n_383), .C(n_413), .D(n_427), .E(n_453), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
OAI21xp33_ASAP7_75t_L g483 ( .A1(n_127), .A2(n_426), .B(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g809 ( .A(n_127), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_128), .B(n_332), .Y(n_127) );
NOR3xp33_ASAP7_75t_SL g128 ( .A(n_129), .B(n_280), .C(n_314), .Y(n_128) );
A2O1A1Ixp33_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_197), .B(n_219), .C(n_258), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_131), .B(n_172), .Y(n_130) );
BUFx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_132), .B(n_270), .Y(n_335) );
AND2x2_ASAP7_75t_L g422 ( .A(n_132), .B(n_200), .Y(n_422) );
HB1xp67_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
OR2x2_ASAP7_75t_L g218 ( .A(n_133), .B(n_189), .Y(n_218) );
INVx1_ASAP7_75t_L g260 ( .A(n_133), .Y(n_260) );
INVx2_ASAP7_75t_L g265 ( .A(n_133), .Y(n_265) );
HB1xp67_ASAP7_75t_L g293 ( .A(n_133), .Y(n_293) );
INVx1_ASAP7_75t_L g307 ( .A(n_133), .Y(n_307) );
AND2x2_ASAP7_75t_L g311 ( .A(n_133), .B(n_202), .Y(n_311) );
AND2x2_ASAP7_75t_L g392 ( .A(n_133), .B(n_201), .Y(n_392) );
AO21x2_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_139), .B(n_168), .Y(n_133) );
AO21x2_ASAP7_75t_L g522 ( .A1(n_134), .A2(n_523), .B(n_529), .Y(n_522) );
AO21x2_ASAP7_75t_L g549 ( .A1(n_134), .A2(n_550), .B(n_556), .Y(n_549) );
AO21x2_ASAP7_75t_L g587 ( .A1(n_134), .A2(n_523), .B(n_529), .Y(n_587) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_135), .Y(n_134) );
OA21x2_ASAP7_75t_L g579 ( .A1(n_135), .A2(n_580), .B(n_584), .Y(n_579) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
AND2x2_ASAP7_75t_SL g136 ( .A(n_137), .B(n_138), .Y(n_136) );
AND2x4_ASAP7_75t_L g180 ( .A(n_137), .B(n_138), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_140), .B(n_150), .Y(n_139) );
INVx1_ASAP7_75t_L g257 ( .A(n_141), .Y(n_257) );
AOI22xp5_ASAP7_75t_L g498 ( .A1(n_141), .A2(n_151), .B1(n_499), .B2(n_501), .Y(n_498) );
AND2x4_ASAP7_75t_L g141 ( .A(n_142), .B(n_147), .Y(n_141) );
INVx1_ASAP7_75t_L g177 ( .A(n_142), .Y(n_177) );
AND2x2_ASAP7_75t_L g142 ( .A(n_143), .B(n_145), .Y(n_142) );
OR2x6_ASAP7_75t_L g159 ( .A(n_143), .B(n_155), .Y(n_159) );
INVxp33_ASAP7_75t_L g229 ( .A(n_143), .Y(n_229) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
AND2x2_ASAP7_75t_L g156 ( .A(n_144), .B(n_146), .Y(n_156) );
AND2x4_ASAP7_75t_L g215 ( .A(n_144), .B(n_164), .Y(n_215) );
HB1xp67_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx1_ASAP7_75t_L g178 ( .A(n_147), .Y(n_178) );
BUFx3_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
AND2x6_ASAP7_75t_L g506 ( .A(n_148), .B(n_156), .Y(n_506) );
INVx2_ASAP7_75t_L g155 ( .A(n_149), .Y(n_155) );
AND2x6_ASAP7_75t_L g212 ( .A(n_149), .B(n_162), .Y(n_212) );
INVxp67_ASAP7_75t_L g255 ( .A(n_151), .Y(n_255) );
AND2x4_ASAP7_75t_L g151 ( .A(n_152), .B(n_156), .Y(n_151) );
NOR2x1p5_ASAP7_75t_L g152 ( .A(n_153), .B(n_154), .Y(n_152) );
INVx1_ASAP7_75t_L g230 ( .A(n_154), .Y(n_230) );
INVx3_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
O2A1O1Ixp33_ASAP7_75t_SL g157 ( .A1(n_158), .A2(n_159), .B(n_160), .C(n_166), .Y(n_157) );
INVx2_ASAP7_75t_L g185 ( .A(n_159), .Y(n_185) );
O2A1O1Ixp33_ASAP7_75t_L g193 ( .A1(n_159), .A2(n_166), .B(n_194), .C(n_195), .Y(n_193) );
OAI22xp5_ASAP7_75t_L g205 ( .A1(n_159), .A2(n_206), .B1(n_207), .B2(n_208), .Y(n_205) );
O2A1O1Ixp33_ASAP7_75t_SL g236 ( .A1(n_159), .A2(n_166), .B(n_237), .C(n_238), .Y(n_236) );
INVxp67_ASAP7_75t_L g245 ( .A(n_159), .Y(n_245) );
O2A1O1Ixp33_ASAP7_75t_L g276 ( .A1(n_159), .A2(n_166), .B(n_277), .C(n_278), .Y(n_276) );
INVx1_ASAP7_75t_L g208 ( .A(n_161), .Y(n_208) );
AND2x4_ASAP7_75t_L g518 ( .A(n_161), .B(n_167), .Y(n_518) );
AND2x4_ASAP7_75t_L g161 ( .A(n_162), .B(n_164), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
AOI21xp5_ASAP7_75t_L g182 ( .A1(n_166), .A2(n_183), .B(n_184), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g216 ( .A(n_166), .B(n_180), .Y(n_216) );
INVx1_ASAP7_75t_L g226 ( .A(n_166), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_166), .A2(n_515), .B(n_516), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_166), .A2(n_526), .B(n_527), .Y(n_525) );
AOI21xp5_ASAP7_75t_L g539 ( .A1(n_166), .A2(n_540), .B(n_541), .Y(n_539) );
AOI21xp5_ASAP7_75t_L g552 ( .A1(n_166), .A2(n_553), .B(n_554), .Y(n_552) );
AOI21xp5_ASAP7_75t_L g573 ( .A1(n_166), .A2(n_574), .B(n_575), .Y(n_573) );
AOI21xp5_ASAP7_75t_L g581 ( .A1(n_166), .A2(n_582), .B(n_583), .Y(n_581) );
INVx5_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
HB1xp67_ASAP7_75t_L g248 ( .A(n_167), .Y(n_248) );
OAI22xp5_ASAP7_75t_L g243 ( .A1(n_169), .A2(n_244), .B1(n_249), .B2(n_250), .Y(n_243) );
INVx3_ASAP7_75t_L g250 ( .A(n_169), .Y(n_250) );
INVx4_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_170), .B(n_253), .Y(n_252) );
AOI21x1_ASAP7_75t_L g511 ( .A1(n_170), .A2(n_512), .B(n_519), .Y(n_511) );
INVx3_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
BUFx4f_ASAP7_75t_L g187 ( .A(n_171), .Y(n_187) );
AND2x4_ASAP7_75t_SL g172 ( .A(n_173), .B(n_188), .Y(n_172) );
HB1xp67_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx2_ASAP7_75t_L g217 ( .A(n_174), .Y(n_217) );
AND2x2_ASAP7_75t_L g261 ( .A(n_174), .B(n_202), .Y(n_261) );
AND2x2_ASAP7_75t_L g282 ( .A(n_174), .B(n_189), .Y(n_282) );
INVx1_ASAP7_75t_L g305 ( .A(n_174), .Y(n_305) );
AND2x4_ASAP7_75t_L g372 ( .A(n_174), .B(n_201), .Y(n_372) );
AND2x2_ASAP7_75t_L g174 ( .A(n_175), .B(n_181), .Y(n_174) );
NOR3xp33_ASAP7_75t_L g176 ( .A(n_177), .B(n_178), .C(n_179), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g191 ( .A1(n_180), .A2(n_192), .B(n_196), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_180), .B(n_500), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_180), .B(n_502), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_180), .B(n_505), .Y(n_504) );
NOR3xp33_ASAP7_75t_L g507 ( .A(n_180), .B(n_208), .C(n_508), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_180), .A2(n_537), .B(n_538), .Y(n_536) );
AO21x2_ASAP7_75t_L g223 ( .A1(n_186), .A2(n_224), .B(n_232), .Y(n_223) );
AO21x2_ASAP7_75t_L g287 ( .A1(n_186), .A2(n_224), .B(n_232), .Y(n_287) );
AOI21x1_ASAP7_75t_L g544 ( .A1(n_186), .A2(n_545), .B(n_548), .Y(n_544) );
INVx2_ASAP7_75t_SL g186 ( .A(n_187), .Y(n_186) );
OA21x2_ASAP7_75t_L g234 ( .A1(n_187), .A2(n_235), .B(n_239), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g570 ( .A1(n_187), .A2(n_571), .B(n_572), .Y(n_570) );
AND2x4_ASAP7_75t_L g388 ( .A(n_188), .B(n_305), .Y(n_388) );
OR2x2_ASAP7_75t_L g429 ( .A(n_188), .B(n_430), .Y(n_429) );
NOR2xp67_ASAP7_75t_SL g448 ( .A(n_188), .B(n_321), .Y(n_448) );
NOR2x1_ASAP7_75t_L g466 ( .A(n_188), .B(n_380), .Y(n_466) );
INVx4_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
NOR2x1_ASAP7_75t_SL g266 ( .A(n_189), .B(n_202), .Y(n_266) );
AND2x4_ASAP7_75t_L g304 ( .A(n_189), .B(n_305), .Y(n_304) );
BUFx6f_ASAP7_75t_L g310 ( .A(n_189), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_189), .B(n_264), .Y(n_342) );
INVx2_ASAP7_75t_L g356 ( .A(n_189), .Y(n_356) );
NAND2xp5_ASAP7_75t_SL g378 ( .A(n_189), .B(n_308), .Y(n_378) );
AND2x2_ASAP7_75t_L g470 ( .A(n_189), .B(n_328), .Y(n_470) );
OR2x6_ASAP7_75t_L g189 ( .A(n_190), .B(n_191), .Y(n_189) );
INVx1_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
NOR2x1_ASAP7_75t_L g198 ( .A(n_199), .B(n_218), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_200), .B(n_307), .Y(n_321) );
AND2x2_ASAP7_75t_SL g330 ( .A(n_200), .B(n_310), .Y(n_330) );
AND2x2_ASAP7_75t_L g200 ( .A(n_201), .B(n_217), .Y(n_200) );
INVx1_ASAP7_75t_L g308 ( .A(n_201), .Y(n_308) );
INVx3_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx2_ASAP7_75t_L g328 ( .A(n_202), .Y(n_328) );
AND2x4_ASAP7_75t_L g202 ( .A(n_203), .B(n_204), .Y(n_202) );
OAI21xp5_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_209), .B(n_216), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_208), .B(n_247), .Y(n_246) );
OAI22xp5_ASAP7_75t_L g209 ( .A1(n_210), .A2(n_211), .B1(n_213), .B2(n_214), .Y(n_209) );
INVxp67_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
INVxp67_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
INVx1_ASAP7_75t_L g361 ( .A(n_217), .Y(n_361) );
INVx2_ASAP7_75t_SL g406 ( .A(n_218), .Y(n_406) );
INVx1_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
AND2x2_ASAP7_75t_L g220 ( .A(n_221), .B(n_240), .Y(n_220) );
NAND2x1p5_ASAP7_75t_L g315 ( .A(n_221), .B(n_316), .Y(n_315) );
BUFx2_ASAP7_75t_L g352 ( .A(n_221), .Y(n_352) );
AND2x2_ASAP7_75t_L g476 ( .A(n_221), .B(n_301), .Y(n_476) );
AND2x2_ASAP7_75t_L g221 ( .A(n_222), .B(n_233), .Y(n_221) );
AND2x4_ASAP7_75t_L g289 ( .A(n_222), .B(n_271), .Y(n_289) );
INVx1_ASAP7_75t_L g300 ( .A(n_222), .Y(n_300) );
AND2x2_ASAP7_75t_L g331 ( .A(n_222), .B(n_286), .Y(n_331) );
INVx2_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_223), .B(n_234), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_223), .B(n_272), .Y(n_363) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_225), .B(n_231), .Y(n_224) );
INVx1_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
INVxp67_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
INVx2_ASAP7_75t_L g269 ( .A(n_234), .Y(n_269) );
AND2x4_ASAP7_75t_L g337 ( .A(n_234), .B(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g349 ( .A(n_234), .Y(n_349) );
INVx1_ASAP7_75t_L g391 ( .A(n_234), .Y(n_391) );
HB1xp67_ASAP7_75t_L g403 ( .A(n_234), .Y(n_403) );
AND2x2_ASAP7_75t_L g419 ( .A(n_234), .B(n_242), .Y(n_419) );
BUFx2_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
AND2x2_ASAP7_75t_L g366 ( .A(n_241), .B(n_324), .Y(n_366) );
INVx1_ASAP7_75t_SL g368 ( .A(n_241), .Y(n_368) );
AND2x2_ASAP7_75t_L g389 ( .A(n_241), .B(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
AND2x4_ASAP7_75t_L g268 ( .A(n_242), .B(n_269), .Y(n_268) );
INVx1_ASAP7_75t_L g296 ( .A(n_242), .Y(n_296) );
INVx2_ASAP7_75t_L g302 ( .A(n_242), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_242), .B(n_272), .Y(n_317) );
OR2x2_ASAP7_75t_L g242 ( .A(n_243), .B(n_251), .Y(n_242) );
AO21x2_ASAP7_75t_L g272 ( .A1(n_250), .A2(n_273), .B(n_279), .Y(n_272) );
AO21x2_ASAP7_75t_L g286 ( .A1(n_250), .A2(n_273), .B(n_279), .Y(n_286) );
OAI22xp5_ASAP7_75t_L g251 ( .A1(n_252), .A2(n_255), .B1(n_256), .B2(n_257), .Y(n_251) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
OAI21xp5_ASAP7_75t_L g258 ( .A1(n_259), .A2(n_262), .B(n_267), .Y(n_258) );
INVx1_ASAP7_75t_L g398 ( .A(n_259), .Y(n_398) );
AND2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_261), .Y(n_259) );
INVx2_ASAP7_75t_L g318 ( .A(n_261), .Y(n_318) );
AND2x2_ASAP7_75t_L g374 ( .A(n_261), .B(n_310), .Y(n_374) );
AND2x2_ASAP7_75t_L g262 ( .A(n_263), .B(n_266), .Y(n_262) );
INVx1_ASAP7_75t_L g288 ( .A(n_263), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_263), .B(n_304), .Y(n_350) );
NOR2xp33_ASAP7_75t_L g379 ( .A(n_263), .B(n_380), .Y(n_379) );
AND2x2_ASAP7_75t_L g395 ( .A(n_263), .B(n_388), .Y(n_395) );
AND2x2_ASAP7_75t_L g469 ( .A(n_263), .B(n_470), .Y(n_469) );
INVx3_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
HB1xp67_ASAP7_75t_L g457 ( .A(n_264), .Y(n_457) );
INVx2_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
HB1xp67_ASAP7_75t_L g377 ( .A(n_265), .Y(n_377) );
AND2x2_ASAP7_75t_L g290 ( .A(n_266), .B(n_291), .Y(n_290) );
OAI21xp33_ASAP7_75t_L g478 ( .A1(n_266), .A2(n_479), .B(n_481), .Y(n_478) );
AND2x2_ASAP7_75t_L g267 ( .A(n_268), .B(n_270), .Y(n_267) );
INVx3_ASAP7_75t_L g364 ( .A(n_268), .Y(n_364) );
NAND2x1_ASAP7_75t_SL g408 ( .A(n_268), .B(n_409), .Y(n_408) );
AND2x2_ASAP7_75t_L g411 ( .A(n_268), .B(n_289), .Y(n_411) );
AND2x2_ASAP7_75t_L g323 ( .A(n_270), .B(n_324), .Y(n_323) );
OR2x2_ASAP7_75t_L g460 ( .A(n_270), .B(n_461), .Y(n_460) );
AND2x2_ASAP7_75t_L g471 ( .A(n_270), .B(n_419), .Y(n_471) );
INVx3_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
NAND2x1p5_ASAP7_75t_L g347 ( .A(n_271), .B(n_348), .Y(n_347) );
INVx3_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g402 ( .A(n_272), .B(n_403), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
OAI21xp5_ASAP7_75t_SL g280 ( .A1(n_281), .A2(n_294), .B(n_297), .Y(n_280) );
AOI22xp5_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_283), .B1(n_289), .B2(n_290), .Y(n_281) );
HB1xp67_ASAP7_75t_L g339 ( .A(n_282), .Y(n_339) );
AND2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_288), .Y(n_283) );
AND2x2_ASAP7_75t_L g312 ( .A(n_284), .B(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g418 ( .A(n_284), .B(n_419), .Y(n_418) );
AOI22xp5_ASAP7_75t_L g436 ( .A1(n_284), .A2(n_437), .B1(n_438), .B2(n_439), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_284), .B(n_445), .Y(n_444) );
AND2x4_ASAP7_75t_L g284 ( .A(n_285), .B(n_287), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g301 ( .A(n_286), .B(n_302), .Y(n_301) );
NOR2xp67_ASAP7_75t_L g382 ( .A(n_286), .B(n_302), .Y(n_382) );
NOR2x1_ASAP7_75t_L g390 ( .A(n_286), .B(n_391), .Y(n_390) );
INVx2_ASAP7_75t_L g338 ( .A(n_287), .Y(n_338) );
AND2x2_ASAP7_75t_L g346 ( .A(n_287), .B(n_302), .Y(n_346) );
INVx1_ASAP7_75t_L g409 ( .A(n_287), .Y(n_409) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NAND2x1_ASAP7_75t_L g327 ( .A(n_292), .B(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g439 ( .A(n_295), .B(n_324), .Y(n_439) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx2_ASAP7_75t_L g313 ( .A(n_296), .Y(n_313) );
AND2x2_ASAP7_75t_L g336 ( .A(n_296), .B(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g424 ( .A(n_296), .B(n_331), .Y(n_424) );
AOI22xp5_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_303), .B1(n_309), .B2(n_312), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
OR2x2_ASAP7_75t_L g432 ( .A(n_299), .B(n_433), .Y(n_432) );
NAND2x1p5_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
AND2x2_ASAP7_75t_L g462 ( .A(n_302), .B(n_349), .Y(n_462) );
AND2x2_ASAP7_75t_SL g303 ( .A(n_304), .B(n_306), .Y(n_303) );
INVx2_ASAP7_75t_L g329 ( .A(n_304), .Y(n_329) );
OAI21xp33_ASAP7_75t_SL g475 ( .A1(n_304), .A2(n_476), .B(n_477), .Y(n_475) );
AND2x4_ASAP7_75t_SL g306 ( .A(n_307), .B(n_308), .Y(n_306) );
HB1xp67_ASAP7_75t_L g465 ( .A(n_307), .Y(n_465) );
AND2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
O2A1O1Ixp33_ASAP7_75t_SL g407 ( .A1(n_310), .A2(n_408), .B(n_410), .C(n_412), .Y(n_407) );
AND2x2_ASAP7_75t_SL g359 ( .A(n_311), .B(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g412 ( .A(n_311), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_311), .B(n_388), .Y(n_452) );
INVx1_ASAP7_75t_SL g319 ( .A(n_312), .Y(n_319) );
AND2x2_ASAP7_75t_L g400 ( .A(n_313), .B(n_337), .Y(n_400) );
INVx1_ASAP7_75t_L g445 ( .A(n_313), .Y(n_445) );
OAI221xp5_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_318), .B1(n_319), .B2(n_320), .C(n_322), .Y(n_314) );
HB1xp67_ASAP7_75t_L g434 ( .A(n_315), .Y(n_434) );
INVx2_ASAP7_75t_SL g316 ( .A(n_317), .Y(n_316) );
OR2x2_ASAP7_75t_L g482 ( .A(n_317), .B(n_325), .Y(n_482) );
OR2x2_ASAP7_75t_L g341 ( .A(n_318), .B(n_342), .Y(n_341) );
NOR2x1_ASAP7_75t_L g354 ( .A(n_318), .B(n_355), .Y(n_354) );
NOR2xp33_ASAP7_75t_L g441 ( .A(n_318), .B(n_442), .Y(n_441) );
OR2x2_ASAP7_75t_L g480 ( .A(n_318), .B(n_377), .Y(n_480) );
BUFx2_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
AOI32xp33_ASAP7_75t_L g322 ( .A1(n_323), .A2(n_326), .A3(n_329), .B1(n_330), .B2(n_331), .Y(n_322) );
INVx1_ASAP7_75t_L g343 ( .A(n_324), .Y(n_343) );
INVx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
NOR2xp33_ASAP7_75t_L g386 ( .A(n_326), .B(n_387), .Y(n_386) );
INVx2_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g438 ( .A(n_327), .Y(n_438) );
OAI22xp33_ASAP7_75t_SL g420 ( .A1(n_329), .A2(n_421), .B1(n_423), .B2(n_425), .Y(n_420) );
INVx1_ASAP7_75t_L g451 ( .A(n_330), .Y(n_451) );
AOI211x1_ASAP7_75t_L g332 ( .A1(n_333), .A2(n_339), .B(n_340), .C(n_357), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_334), .B(n_336), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_334), .B(n_419), .Y(n_425) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
AND2x4_ASAP7_75t_L g381 ( .A(n_337), .B(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g447 ( .A(n_337), .Y(n_447) );
OAI222xp33_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_343), .B1(n_344), .B2(n_350), .C1(n_351), .C2(n_353), .Y(n_340) );
INVxp67_ASAP7_75t_L g437 ( .A(n_341), .Y(n_437) );
OR2x2_ASAP7_75t_L g344 ( .A(n_345), .B(n_347), .Y(n_344) );
NOR2xp33_ASAP7_75t_L g477 ( .A(n_345), .B(n_430), .Y(n_477) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g393 ( .A(n_346), .B(n_390), .Y(n_393) );
INVx3_ASAP7_75t_L g433 ( .A(n_348), .Y(n_433) );
BUFx3_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g371 ( .A(n_356), .B(n_372), .Y(n_371) );
OAI221xp5_ASAP7_75t_L g357 ( .A1(n_358), .A2(n_362), .B1(n_365), .B2(n_370), .C(n_373), .Y(n_357) );
INVx1_ASAP7_75t_SL g358 ( .A(n_359), .Y(n_358) );
OAI21xp5_ASAP7_75t_L g415 ( .A1(n_359), .A2(n_416), .B(n_418), .Y(n_415) );
INVx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
OR2x2_ASAP7_75t_L g362 ( .A(n_363), .B(n_364), .Y(n_362) );
INVx1_ASAP7_75t_L g369 ( .A(n_363), .Y(n_369) );
OR2x2_ASAP7_75t_L g473 ( .A(n_364), .B(n_409), .Y(n_473) );
NOR2xp67_ASAP7_75t_L g365 ( .A(n_366), .B(n_367), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_367), .B(n_395), .Y(n_394) );
AND2x2_ASAP7_75t_L g367 ( .A(n_368), .B(n_369), .Y(n_367) );
OAI21xp5_ASAP7_75t_L g467 ( .A1(n_370), .A2(n_399), .B(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
OAI21xp5_ASAP7_75t_L g449 ( .A1(n_371), .A2(n_443), .B(n_450), .Y(n_449) );
INVx4_ASAP7_75t_L g380 ( .A(n_372), .Y(n_380) );
OAI31xp33_ASAP7_75t_SL g373 ( .A1(n_374), .A2(n_375), .A3(n_379), .B(n_381), .Y(n_373) );
INVx1_ASAP7_75t_L g431 ( .A(n_375), .Y(n_431) );
NOR2x1_ASAP7_75t_L g375 ( .A(n_376), .B(n_378), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx2_ASAP7_75t_L g405 ( .A(n_380), .Y(n_405) );
AND2x2_ASAP7_75t_L g383 ( .A(n_384), .B(n_396), .Y(n_383) );
NAND4xp25_ASAP7_75t_L g484 ( .A(n_384), .B(n_396), .C(n_415), .D(n_485), .Y(n_484) );
AND2x2_ASAP7_75t_L g384 ( .A(n_385), .B(n_394), .Y(n_384) );
AOI22xp5_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_389), .B1(n_392), .B2(n_393), .Y(n_385) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g456 ( .A(n_388), .B(n_457), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_389), .B(n_409), .Y(n_417) );
INVx1_ASAP7_75t_SL g430 ( .A(n_392), .Y(n_430) );
NOR2xp33_ASAP7_75t_L g396 ( .A(n_397), .B(n_407), .Y(n_396) );
OAI22xp5_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_399), .B1(n_401), .B2(n_404), .Y(n_397) );
INVx3_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVxp67_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
NAND2x1_ASAP7_75t_L g404 ( .A(n_405), .B(n_406), .Y(n_404) );
AOI22xp5_ASAP7_75t_L g468 ( .A1(n_406), .A2(n_469), .B1(n_471), .B2(n_472), .Y(n_468) );
INVx2_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
NOR3xp33_ASAP7_75t_L g413 ( .A(n_414), .B(n_420), .C(n_426), .Y(n_413) );
INVxp67_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g485 ( .A(n_420), .Y(n_485) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
OAI21xp33_ASAP7_75t_L g486 ( .A1(n_426), .A2(n_487), .B(n_488), .Y(n_486) );
INVxp33_ASAP7_75t_L g487 ( .A(n_427), .Y(n_487) );
AND2x2_ASAP7_75t_L g808 ( .A(n_427), .B(n_453), .Y(n_808) );
NOR2xp67_ASAP7_75t_L g427 ( .A(n_428), .B(n_435), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g428 ( .A1(n_429), .A2(n_431), .B1(n_432), .B2(n_434), .Y(n_428) );
OAI21xp5_ASAP7_75t_L g454 ( .A1(n_432), .A2(n_455), .B(n_458), .Y(n_454) );
INVx2_ASAP7_75t_L g442 ( .A(n_433), .Y(n_442) );
NAND3xp33_ASAP7_75t_SL g435 ( .A(n_436), .B(n_440), .C(n_449), .Y(n_435) );
AOI22xp5_ASAP7_75t_L g440 ( .A1(n_441), .A2(n_443), .B1(n_446), .B2(n_448), .Y(n_440) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_451), .B(n_452), .Y(n_450) );
INVxp33_ASAP7_75t_SL g488 ( .A(n_453), .Y(n_488) );
NOR3x1_ASAP7_75t_L g453 ( .A(n_454), .B(n_467), .C(n_474), .Y(n_453) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_459), .B(n_463), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_465), .B(n_466), .Y(n_464) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
NAND2xp5_ASAP7_75t_SL g474 ( .A(n_475), .B(n_478), .Y(n_474) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx1_ASAP7_75t_SL g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g810 ( .A(n_484), .Y(n_810) );
CKINVDCx11_ASAP7_75t_R g489 ( .A(n_490), .Y(n_489) );
INVx3_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
AND2x4_ASAP7_75t_L g492 ( .A(n_493), .B(n_656), .Y(n_492) );
NOR4xp25_ASAP7_75t_L g493 ( .A(n_494), .B(n_599), .C(n_638), .D(n_645), .Y(n_493) );
OAI221xp5_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_520), .B1(n_557), .B2(n_566), .C(n_585), .Y(n_494) );
OR2x2_ASAP7_75t_L g729 ( .A(n_495), .B(n_591), .Y(n_729) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
AND2x2_ASAP7_75t_L g644 ( .A(n_496), .B(n_569), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_496), .B(n_664), .Y(n_663) );
AND2x2_ASAP7_75t_SL g709 ( .A(n_496), .B(n_710), .Y(n_709) );
AND2x4_ASAP7_75t_L g496 ( .A(n_497), .B(n_509), .Y(n_496) );
AND2x4_ASAP7_75t_SL g568 ( .A(n_497), .B(n_569), .Y(n_568) );
INVx3_ASAP7_75t_L g590 ( .A(n_497), .Y(n_590) );
AND2x2_ASAP7_75t_L g625 ( .A(n_497), .B(n_598), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_497), .B(n_510), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_497), .B(n_592), .Y(n_677) );
OR2x2_ASAP7_75t_L g755 ( .A(n_497), .B(n_569), .Y(n_755) );
AND2x4_ASAP7_75t_L g497 ( .A(n_498), .B(n_503), .Y(n_497) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
AND2x2_ASAP7_75t_L g577 ( .A(n_510), .B(n_578), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_510), .B(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g603 ( .A(n_510), .Y(n_603) );
OR2x2_ASAP7_75t_L g608 ( .A(n_510), .B(n_592), .Y(n_608) );
AND2x2_ASAP7_75t_L g621 ( .A(n_510), .B(n_579), .Y(n_621) );
HB1xp67_ASAP7_75t_L g624 ( .A(n_510), .Y(n_624) );
INVx1_ASAP7_75t_L g636 ( .A(n_510), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_510), .B(n_590), .Y(n_701) );
INVx3_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_513), .B(n_517), .Y(n_512) );
NAND2xp5_ASAP7_75t_SL g520 ( .A(n_521), .B(n_530), .Y(n_520) );
HB1xp67_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
OR2x2_ASAP7_75t_L g565 ( .A(n_522), .B(n_549), .Y(n_565) );
AND2x4_ASAP7_75t_L g595 ( .A(n_522), .B(n_534), .Y(n_595) );
INVx2_ASAP7_75t_L g629 ( .A(n_522), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_522), .B(n_549), .Y(n_687) );
AND2x2_ASAP7_75t_L g734 ( .A(n_522), .B(n_563), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_524), .B(n_528), .Y(n_523) );
AOI222xp33_ASAP7_75t_L g722 ( .A1(n_530), .A2(n_594), .B1(n_637), .B2(n_697), .C1(n_723), .C2(n_725), .Y(n_722) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_532), .B(n_542), .Y(n_531) );
AND2x2_ASAP7_75t_L g641 ( .A(n_532), .B(n_561), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_532), .B(n_692), .Y(n_691) );
AND2x2_ASAP7_75t_L g770 ( .A(n_532), .B(n_610), .Y(n_770) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g600 ( .A1(n_533), .A2(n_601), .B(n_605), .Y(n_600) );
AND2x2_ASAP7_75t_L g681 ( .A(n_533), .B(n_564), .Y(n_681) );
OR2x2_ASAP7_75t_L g706 ( .A(n_533), .B(n_565), .Y(n_706) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx5_ASAP7_75t_L g560 ( .A(n_534), .Y(n_560) );
AND2x2_ASAP7_75t_L g647 ( .A(n_534), .B(n_629), .Y(n_647) );
AND2x2_ASAP7_75t_L g673 ( .A(n_534), .B(n_549), .Y(n_673) );
OR2x2_ASAP7_75t_L g676 ( .A(n_534), .B(n_563), .Y(n_676) );
HB1xp67_ASAP7_75t_L g694 ( .A(n_534), .Y(n_694) );
AND2x4_ASAP7_75t_SL g751 ( .A(n_534), .B(n_628), .Y(n_751) );
OR2x2_ASAP7_75t_L g760 ( .A(n_534), .B(n_587), .Y(n_760) );
OR2x6_ASAP7_75t_L g534 ( .A(n_535), .B(n_536), .Y(n_534) );
INVx1_ASAP7_75t_L g593 ( .A(n_542), .Y(n_593) );
AOI221xp5_ASAP7_75t_SL g711 ( .A1(n_542), .A2(n_595), .B1(n_712), .B2(n_714), .C(n_715), .Y(n_711) );
AND2x2_ASAP7_75t_L g542 ( .A(n_543), .B(n_549), .Y(n_542) );
OR2x2_ASAP7_75t_L g650 ( .A(n_543), .B(n_620), .Y(n_650) );
OR2x2_ASAP7_75t_L g660 ( .A(n_543), .B(n_661), .Y(n_660) );
OR2x2_ASAP7_75t_L g686 ( .A(n_543), .B(n_687), .Y(n_686) );
AND2x4_ASAP7_75t_L g692 ( .A(n_543), .B(n_611), .Y(n_692) );
NOR2xp33_ASAP7_75t_L g704 ( .A(n_543), .B(n_675), .Y(n_704) );
INVx2_ASAP7_75t_L g717 ( .A(n_543), .Y(n_717) );
NAND2xp5_ASAP7_75t_SL g738 ( .A(n_543), .B(n_595), .Y(n_738) );
AND2x2_ASAP7_75t_L g742 ( .A(n_543), .B(n_564), .Y(n_742) );
AND2x2_ASAP7_75t_L g750 ( .A(n_543), .B(n_751), .Y(n_750) );
BUFx6f_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx2_ASAP7_75t_L g563 ( .A(n_544), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_546), .B(n_547), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_549), .B(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g594 ( .A(n_549), .B(n_563), .Y(n_594) );
INVx2_ASAP7_75t_L g611 ( .A(n_549), .Y(n_611) );
AND2x4_ASAP7_75t_L g628 ( .A(n_549), .B(n_629), .Y(n_628) );
HB1xp67_ASAP7_75t_L g733 ( .A(n_549), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_551), .B(n_555), .Y(n_550) );
NOR2xp33_ASAP7_75t_L g557 ( .A(n_558), .B(n_561), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
OR2x2_ASAP7_75t_L g740 ( .A(n_559), .B(n_562), .Y(n_740) );
AND2x4_ASAP7_75t_L g586 ( .A(n_560), .B(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g627 ( .A(n_560), .B(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g654 ( .A(n_560), .B(n_594), .Y(n_654) );
AND2x2_ASAP7_75t_L g561 ( .A(n_562), .B(n_564), .Y(n_561) );
AND2x2_ASAP7_75t_L g758 ( .A(n_562), .B(n_759), .Y(n_758) );
BUFx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g610 ( .A(n_563), .B(n_611), .Y(n_610) );
OAI21xp5_ASAP7_75t_SL g630 ( .A1(n_564), .A2(n_631), .B(n_637), .Y(n_630) );
INVx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx1_ASAP7_75t_SL g566 ( .A(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_568), .B(n_577), .Y(n_567) );
INVx1_ASAP7_75t_SL g684 ( .A(n_568), .Y(n_684) );
AND2x2_ASAP7_75t_L g714 ( .A(n_568), .B(n_624), .Y(n_714) );
AND2x4_ASAP7_75t_L g725 ( .A(n_568), .B(n_726), .Y(n_725) );
OR2x2_ASAP7_75t_L g591 ( .A(n_569), .B(n_592), .Y(n_591) );
INVx2_ASAP7_75t_L g598 ( .A(n_569), .Y(n_598) );
AND2x4_ASAP7_75t_L g604 ( .A(n_569), .B(n_590), .Y(n_604) );
INVx2_ASAP7_75t_L g615 ( .A(n_569), .Y(n_615) );
INVx1_ASAP7_75t_L g664 ( .A(n_569), .Y(n_664) );
OR2x2_ASAP7_75t_L g685 ( .A(n_569), .B(n_669), .Y(n_685) );
OR2x2_ASAP7_75t_L g699 ( .A(n_569), .B(n_579), .Y(n_699) );
HB1xp67_ASAP7_75t_L g765 ( .A(n_569), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_569), .B(n_621), .Y(n_771) );
OR2x6_ASAP7_75t_L g569 ( .A(n_570), .B(n_576), .Y(n_569) );
INVx1_ASAP7_75t_L g616 ( .A(n_577), .Y(n_616) );
AND2x2_ASAP7_75t_L g749 ( .A(n_577), .B(n_615), .Y(n_749) );
AND2x2_ASAP7_75t_L g774 ( .A(n_577), .B(n_604), .Y(n_774) );
INVx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx2_ASAP7_75t_L g592 ( .A(n_579), .Y(n_592) );
BUFx3_ASAP7_75t_L g634 ( .A(n_579), .Y(n_634) );
HB1xp67_ASAP7_75t_L g661 ( .A(n_579), .Y(n_661) );
INVx1_ASAP7_75t_L g670 ( .A(n_579), .Y(n_670) );
AOI33xp33_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_588), .A3(n_593), .B1(n_594), .B2(n_595), .B3(n_596), .Y(n_585) );
AOI21x1_ASAP7_75t_SL g688 ( .A1(n_586), .A2(n_610), .B(n_672), .Y(n_688) );
INVx2_ASAP7_75t_L g718 ( .A(n_586), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_586), .B(n_717), .Y(n_724) );
AND2x2_ASAP7_75t_L g672 ( .A(n_587), .B(n_673), .Y(n_672) );
INVx1_ASAP7_75t_SL g588 ( .A(n_589), .Y(n_588) );
OR2x2_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
AND2x2_ASAP7_75t_L g635 ( .A(n_590), .B(n_636), .Y(n_635) );
INVx2_ASAP7_75t_L g736 ( .A(n_591), .Y(n_736) );
HB1xp67_ASAP7_75t_L g726 ( .A(n_592), .Y(n_726) );
OAI32xp33_ASAP7_75t_L g775 ( .A1(n_593), .A2(n_595), .A3(n_771), .B1(n_776), .B2(n_778), .Y(n_775) );
AND2x2_ASAP7_75t_L g693 ( .A(n_594), .B(n_694), .Y(n_693) );
INVx2_ASAP7_75t_SL g683 ( .A(n_595), .Y(n_683) );
AND2x2_ASAP7_75t_L g748 ( .A(n_595), .B(n_692), .Y(n_748) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
OAI221xp5_ASAP7_75t_L g599 ( .A1(n_600), .A2(n_609), .B1(n_612), .B2(n_626), .C(n_630), .Y(n_599) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_603), .B(n_604), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_603), .B(n_670), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_604), .B(n_607), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_604), .B(n_720), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_604), .B(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g653 ( .A(n_608), .Y(n_653) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
NOR3xp33_ASAP7_75t_L g612 ( .A(n_613), .B(n_617), .C(n_622), .Y(n_612) );
INVx1_ASAP7_75t_SL g613 ( .A(n_614), .Y(n_613) );
OAI22xp33_ASAP7_75t_L g715 ( .A1(n_614), .A2(n_676), .B1(n_716), .B2(n_719), .Y(n_715) );
OR2x2_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
INVx1_ASAP7_75t_L g619 ( .A(n_615), .Y(n_619) );
NOR2x1p5_ASAP7_75t_L g633 ( .A(n_615), .B(n_634), .Y(n_633) );
HB1xp67_ASAP7_75t_L g655 ( .A(n_615), .Y(n_655) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
OAI322xp33_ASAP7_75t_L g682 ( .A1(n_618), .A2(n_660), .A3(n_683), .B1(n_684), .B2(n_685), .C1(n_686), .C2(n_688), .Y(n_682) );
OR2x2_ASAP7_75t_L g618 ( .A(n_619), .B(n_620), .Y(n_618) );
A2O1A1Ixp33_ASAP7_75t_L g638 ( .A1(n_620), .A2(n_639), .B(n_640), .C(n_642), .Y(n_638) );
OR2x2_ASAP7_75t_L g730 ( .A(n_620), .B(n_684), .Y(n_730) );
INVx2_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g637 ( .A(n_621), .B(n_625), .Y(n_637) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_624), .B(n_625), .Y(n_623) );
INVx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g643 ( .A(n_627), .B(n_644), .Y(n_643) );
INVx3_ASAP7_75t_SL g675 ( .A(n_628), .Y(n_675) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_632), .B(n_696), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_633), .B(n_635), .Y(n_632) );
INVx1_ASAP7_75t_SL g679 ( .A(n_635), .Y(n_679) );
HB1xp67_ASAP7_75t_L g721 ( .A(n_636), .Y(n_721) );
OR2x6_ASAP7_75t_SL g776 ( .A(n_639), .B(n_777), .Y(n_776) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVxp67_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
AOI211xp5_ASAP7_75t_L g766 ( .A1(n_644), .A2(n_767), .B(n_768), .C(n_775), .Y(n_766) );
O2A1O1Ixp33_ASAP7_75t_SL g645 ( .A1(n_646), .A2(n_648), .B(n_651), .C(n_655), .Y(n_645) );
OAI211xp5_ASAP7_75t_SL g657 ( .A1(n_646), .A2(n_658), .B(n_665), .C(n_689), .Y(n_657) );
INVx2_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx3_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVxp67_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
AND2x2_ASAP7_75t_L g652 ( .A(n_653), .B(n_654), .Y(n_652) );
NOR3xp33_ASAP7_75t_L g656 ( .A(n_657), .B(n_702), .C(n_746), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_659), .B(n_662), .Y(n_658) );
INVx1_ASAP7_75t_SL g659 ( .A(n_660), .Y(n_659) );
HB1xp67_ASAP7_75t_L g753 ( .A(n_661), .Y(n_753) );
INVx1_ASAP7_75t_SL g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g708 ( .A(n_664), .Y(n_708) );
NOR3xp33_ASAP7_75t_SL g665 ( .A(n_666), .B(n_678), .C(n_682), .Y(n_665) );
OAI22xp5_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_671), .B1(n_674), .B2(n_677), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g710 ( .A(n_670), .Y(n_710) );
INVxp67_ASAP7_75t_SL g777 ( .A(n_670), .Y(n_777) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
OR2x2_ASAP7_75t_L g674 ( .A(n_675), .B(n_676), .Y(n_674) );
INVx1_ASAP7_75t_SL g763 ( .A(n_676), .Y(n_763) );
NOR2xp33_ASAP7_75t_L g678 ( .A(n_679), .B(n_680), .Y(n_678) );
OR2x2_ASAP7_75t_L g713 ( .A(n_679), .B(n_699), .Y(n_713) );
OR2x2_ASAP7_75t_L g764 ( .A(n_679), .B(n_765), .Y(n_764) );
INVx2_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g762 ( .A(n_687), .Y(n_762) );
OR2x2_ASAP7_75t_L g778 ( .A(n_687), .B(n_717), .Y(n_778) );
OAI21xp33_ASAP7_75t_L g689 ( .A1(n_690), .A2(n_693), .B(n_695), .Y(n_689) );
OAI31xp33_ASAP7_75t_L g703 ( .A1(n_690), .A2(n_704), .A3(n_705), .B(n_707), .Y(n_703) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
AND2x2_ASAP7_75t_L g697 ( .A(n_698), .B(n_700), .Y(n_697) );
INVx1_ASAP7_75t_SL g698 ( .A(n_699), .Y(n_698) );
AND2x4_ASAP7_75t_L g735 ( .A(n_700), .B(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
NAND4xp25_ASAP7_75t_SL g702 ( .A(n_703), .B(n_711), .C(n_722), .D(n_727), .Y(n_702) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
AND2x2_ASAP7_75t_L g707 ( .A(n_708), .B(n_709), .Y(n_707) );
HB1xp67_ASAP7_75t_L g745 ( .A(n_710), .Y(n_745) );
INVx1_ASAP7_75t_SL g712 ( .A(n_713), .Y(n_712) );
OR2x2_ASAP7_75t_L g716 ( .A(n_717), .B(n_718), .Y(n_716) );
INVxp67_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
AOI221xp5_ASAP7_75t_L g727 ( .A1(n_728), .A2(n_731), .B1(n_735), .B2(n_737), .C(n_739), .Y(n_727) );
NAND2xp33_ASAP7_75t_SL g728 ( .A(n_729), .B(n_730), .Y(n_728) );
INVx1_ASAP7_75t_L g772 ( .A(n_731), .Y(n_772) );
AND2x2_ASAP7_75t_SL g731 ( .A(n_732), .B(n_734), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
AOI21xp33_ASAP7_75t_L g739 ( .A1(n_740), .A2(n_741), .B(n_743), .Y(n_739) );
INVx1_ASAP7_75t_L g767 ( .A(n_741), .Y(n_767) );
INVx2_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
NAND2xp5_ASAP7_75t_SL g746 ( .A(n_747), .B(n_766), .Y(n_746) );
AOI221xp5_ASAP7_75t_L g747 ( .A1(n_748), .A2(n_749), .B1(n_750), .B2(n_752), .C(n_756), .Y(n_747) );
AND2x2_ASAP7_75t_L g752 ( .A(n_753), .B(n_754), .Y(n_752) );
INVx1_ASAP7_75t_SL g754 ( .A(n_755), .Y(n_754) );
AOI21xp33_ASAP7_75t_L g756 ( .A1(n_757), .A2(n_761), .B(n_764), .Y(n_756) );
INVxp33_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx1_ASAP7_75t_SL g759 ( .A(n_760), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_762), .B(n_763), .Y(n_761) );
OAI22xp5_ASAP7_75t_L g768 ( .A1(n_769), .A2(n_771), .B1(n_772), .B2(n_773), .Y(n_768) );
INVx1_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
CKINVDCx5p33_ASAP7_75t_R g779 ( .A(n_780), .Y(n_779) );
CKINVDCx20_ASAP7_75t_R g792 ( .A(n_780), .Y(n_792) );
CKINVDCx11_ASAP7_75t_R g780 ( .A(n_781), .Y(n_780) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_783), .B(n_791), .Y(n_790) );
NOR2xp33_ASAP7_75t_L g786 ( .A(n_787), .B(n_788), .Y(n_786) );
BUFx2_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
CKINVDCx20_ASAP7_75t_R g793 ( .A(n_794), .Y(n_793) );
INVx1_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
AND2x2_ASAP7_75t_L g795 ( .A(n_796), .B(n_800), .Y(n_795) );
INVxp67_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
NAND2xp5_ASAP7_75t_SL g797 ( .A(n_798), .B(n_799), .Y(n_797) );
INVx1_ASAP7_75t_SL g818 ( .A(n_800), .Y(n_818) );
AOI21xp33_ASAP7_75t_L g801 ( .A1(n_802), .A2(n_817), .B(n_819), .Y(n_801) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_803), .B(n_806), .Y(n_802) );
CKINVDCx11_ASAP7_75t_R g803 ( .A(n_804), .Y(n_803) );
CKINVDCx20_ASAP7_75t_R g804 ( .A(n_805), .Y(n_804) );
XNOR2xp5_ASAP7_75t_L g806 ( .A(n_807), .B(n_811), .Y(n_806) );
NAND3x1_ASAP7_75t_L g807 ( .A(n_808), .B(n_809), .C(n_810), .Y(n_807) );
CKINVDCx5p33_ASAP7_75t_R g811 ( .A(n_812), .Y(n_811) );
INVx1_ASAP7_75t_L g816 ( .A(n_814), .Y(n_816) );
INVx2_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
INVx1_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
endmodule