module real_aes_16451_n_376 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_374, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_376);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_374;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_376;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_1797;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_1903;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1929;
wire n_1737;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_1888;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_1972;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1730;
wire n_1744;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1936;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1873;
wire n_1835;
wire n_1871;
wire n_1468;
wire n_1713;
wire n_1967;
wire n_1920;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_1859;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1845;
wire n_1415;
wire n_1160;
wire n_1849;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1805;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1441;
wire n_1225;
wire n_875;
wire n_1199;
wire n_951;
wire n_1382;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1833;
wire n_1477;
wire n_1944;
wire n_595;
wire n_1893;
wire n_1960;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1959;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_1809;
wire n_682;
wire n_1745;
wire n_1820;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_1883;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1981;
wire n_1196;
wire n_1013;
wire n_1905;
wire n_808;
wire n_1694;
wire n_1639;
wire n_1224;
wire n_1872;
wire n_688;
wire n_1042;
wire n_1588;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_1966;
wire n_1346;
wire n_552;
wire n_1383;
wire n_1890;
wire n_1675;
wire n_1954;
wire n_590;
wire n_1293;
wire n_1880;
wire n_432;
wire n_1882;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_1865;
wire n_805;
wire n_1600;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1583;
wire n_1284;
wire n_1987;
wire n_859;
wire n_1465;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_1658;
wire n_1866;
wire n_954;
wire n_702;
wire n_1874;
wire n_1007;
wire n_1906;
wire n_1926;
wire n_898;
wire n_562;
wire n_1897;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1632;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1768;
wire n_1243;
wire n_1846;
wire n_1003;
wire n_749;
wire n_1870;
wire n_914;
wire n_1837;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1813;
wire n_1978;
wire n_1628;
wire n_1587;
wire n_1821;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_1397;
wire n_765;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1825;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1956;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_1940;
wire n_1666;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_1814;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1510;
wire n_1495;
wire n_1727;
wire n_712;
wire n_1921;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1648;
wire n_1914;
wire n_440;
wire n_1945;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_1787;
wire n_424;
wire n_877;
wire n_802;
wire n_1876;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1979;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1828;
wire n_1860;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1973;
wire n_1561;
wire n_635;
wire n_792;
wire n_1542;
wire n_1392;
wire n_665;
wire n_667;
wire n_991;
wire n_1712;
wire n_1556;
wire n_1004;
wire n_580;
wire n_1417;
wire n_1370;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_1951;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_1606;
wire n_1129;
wire n_1760;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_1852;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1830;
wire n_1594;
wire n_1864;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1991;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_1499;
wire n_399;
wire n_700;
wire n_948;
wire n_1269;
wire n_677;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1839;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1881;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1884;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1946;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_1879;
wire n_746;
wire n_1614;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_1853;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_1977;
wire n_1930;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1985;
wire n_1812;
wire n_1769;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_1971;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_1854;
wire n_617;
wire n_602;
wire n_1404;
wire n_402;
wire n_733;
wire n_676;
wire n_658;
wire n_1856;
wire n_531;
wire n_1848;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_1145;
wire n_645;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_777;
wire n_985;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_1907;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_1857;
wire n_1984;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_1234;
wire n_1915;
wire n_622;
wire n_1634;
wire n_1353;
wire n_1002;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_1862;
wire n_1965;
wire n_850;
wire n_720;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_1699;
wire n_1794;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_1970;
wire n_526;
wire n_1513;
wire n_1983;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_1934;
wire n_809;
wire n_1532;
wire n_679;
wire n_520;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1784;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1474;
wire n_1032;
wire n_721;
wire n_1431;
wire n_1806;
wire n_1829;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_1976;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_1524;
wire n_762;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1807;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1910;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1957;
wire n_1184;
wire n_583;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1961;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_1904;
wire n_450;
wire n_1578;
wire n_473;
wire n_1779;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1908;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_1840;
wire n_968;
wire n_710;
wire n_1040;
wire n_1185;
wire n_1102;
wire n_661;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1451;
wire n_1069;
wire n_842;
wire n_1788;
wire n_1938;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1816;
wire n_1952;
wire n_1811;
wire n_1066;
wire n_1917;
wire n_1377;
wire n_800;
wire n_1170;
wire n_1175;
wire n_778;
wire n_522;
wire n_1475;
wire n_1928;
wire n_977;
wire n_943;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_1980;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1932;
wire n_1707;
wire n_856;
wire n_594;
wire n_1146;
wire n_1685;
wire n_1810;
wire n_1435;
wire n_1800;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_1990;
wire n_427;
wire n_1540;
wire n_519;
wire n_1878;
wire n_1116;
wire n_709;
wire n_1834;
wire n_388;
wire n_1913;
wire n_1899;
wire n_816;
wire n_1470;
wire n_625;
wire n_953;
wire n_1565;
wire n_1953;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_584;
wire n_896;
wire n_1817;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1638;
wire n_1072;
wire n_1663;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1923;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1850;
wire n_1332;
wire n_1927;
wire n_1263;
wire n_1411;
wire n_1922;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1827;
wire n_1726;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1949;
wire n_1029;
wire n_1989;
wire n_1207;
wire n_1555;
wire n_1962;
wire n_664;
wire n_1017;
wire n_1942;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_1939;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1869;
wire n_1259;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_1671;
wire n_502;
wire n_434;
wire n_769;
wire n_1455;
wire n_1212;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1895;
wire n_1670;
wire n_1941;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1986;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_1948;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1886;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_1832;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_1605;
wire n_1592;
wire n_1802;
wire n_1855;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1774;
wire n_1785;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1838;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_1863;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_1191;
wire n_705;
wire n_1206;
wire n_1824;
wire n_1933;
wire n_1270;
wire n_1988;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_1761;
wire n_863;
wire n_525;
wire n_1226;
wire n_1617;
wire n_1790;
wire n_644;
wire n_1150;
wire n_1861;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_1143;
wire n_929;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_1457;
wire n_465;
wire n_719;
wire n_1343;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1799;
wire n_640;
wire n_1176;
wire n_1691;
wire n_1721;
wire n_1931;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_1964;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1844;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1937;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_1841;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_987;
wire n_1596;
wire n_1982;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_1822;
wire n_718;
wire n_1955;
wire n_669;
wire n_1091;
wire n_423;
wire n_1969;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_1777;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1819;
wire n_1887;
wire n_1674;
wire n_491;
wire n_1294;
wire n_1902;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_1889;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_1896;
wire n_767;
wire n_889;
wire n_1398;
wire n_1911;
wire n_379;
wire n_1847;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1912;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1654;
wire n_1099;
wire n_626;
wire n_539;
wire n_1919;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1541;
wire n_1272;
wire n_408;
wire n_1754;
wire n_892;
wire n_578;
wire n_938;
wire n_774;
wire n_1049;
wire n_466;
wire n_559;
wire n_1277;
wire n_1584;
wire n_1950;
wire n_984;
wire n_726;
wire n_517;
wire n_931;
wire n_780;
wire n_1851;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_1916;
wire n_532;
wire n_1025;
wire n_1875;
wire n_1826;
wire n_1836;
wire n_1909;
wire n_924;
wire n_1264;
wire n_1858;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1901;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1943;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1318;
wire n_1290;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_1818;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1974;
wire n_1547;
wire n_1823;
wire n_1867;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1891;
wire n_1267;
wire n_790;
wire n_1262;
wire n_1843;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1885;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_1992;
wire n_1963;
wire n_1958;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1925;
wire n_1801;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_1968;
wire n_430;
wire n_1252;
wire n_1647;
wire n_1132;
wire n_1947;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1894;
wire n_1296;
wire n_1484;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_1808;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_1481;
wire n_1430;
wire n_907;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_1877;
wire n_1900;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1842;
wire n_1536;
wire n_1746;
wire n_1898;
wire n_1711;
wire n_482;
wire n_633;
wire n_1892;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_1573;
wire n_1130;
wire n_1918;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_1831;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_1372;
wire n_698;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1815;
wire n_1924;
wire n_1412;
wire n_1868;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1975;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_1352;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_703;
wire n_1369;
wire n_1097;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1935;
wire n_1645;
wire n_429;
INVx1_ASAP7_75t_L g413 ( .A(n_0), .Y(n_413) );
INVx1_ASAP7_75t_L g798 ( .A(n_1), .Y(n_798) );
INVx1_ASAP7_75t_L g1627 ( .A(n_2), .Y(n_1627) );
OAI211xp5_ASAP7_75t_L g1653 ( .A1(n_2), .A2(n_1654), .B(n_1655), .C(n_1659), .Y(n_1653) );
NOR2xp33_ASAP7_75t_L g445 ( .A(n_3), .B(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g471 ( .A(n_3), .Y(n_471) );
AND2x2_ASAP7_75t_L g797 ( .A(n_3), .B(n_281), .Y(n_797) );
AND2x2_ASAP7_75t_L g811 ( .A(n_3), .B(n_501), .Y(n_811) );
OAI211xp5_ASAP7_75t_SL g477 ( .A1(n_4), .A2(n_478), .B(n_481), .C(n_487), .Y(n_477) );
INVx1_ASAP7_75t_L g538 ( .A(n_4), .Y(n_538) );
INVx1_ASAP7_75t_L g1142 ( .A(n_5), .Y(n_1142) );
OAI22xp5_ASAP7_75t_L g799 ( .A1(n_6), .A2(n_292), .B1(n_800), .B2(n_804), .Y(n_799) );
OAI211xp5_ASAP7_75t_L g808 ( .A1(n_6), .A2(n_809), .B(n_812), .C(n_819), .Y(n_808) );
INVx1_ASAP7_75t_L g1386 ( .A(n_7), .Y(n_1386) );
OAI22xp5_ASAP7_75t_L g1513 ( .A1(n_8), .A2(n_170), .B1(n_644), .B2(n_1514), .Y(n_1513) );
OAI22xp5_ASAP7_75t_L g1526 ( .A1(n_8), .A2(n_170), .B1(n_622), .B2(n_1377), .Y(n_1526) );
OAI22xp33_ASAP7_75t_L g975 ( .A1(n_9), .A2(n_310), .B1(n_693), .B2(n_908), .Y(n_975) );
OAI22xp33_ASAP7_75t_L g981 ( .A1(n_9), .A2(n_310), .B1(n_982), .B2(n_983), .Y(n_981) );
OAI22xp33_ASAP7_75t_L g1515 ( .A1(n_10), .A2(n_303), .B1(n_641), .B2(n_642), .Y(n_1515) );
OAI22xp33_ASAP7_75t_L g1521 ( .A1(n_10), .A2(n_303), .B1(n_633), .B2(n_902), .Y(n_1521) );
AOI22xp33_ASAP7_75t_L g711 ( .A1(n_11), .A2(n_84), .B1(n_706), .B2(n_707), .Y(n_711) );
AOI22xp33_ASAP7_75t_L g743 ( .A1(n_11), .A2(n_250), .B1(n_724), .B2(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g1074 ( .A(n_12), .Y(n_1074) );
AOI22xp33_ASAP7_75t_L g1384 ( .A1(n_13), .A2(n_90), .B1(n_686), .B2(n_773), .Y(n_1384) );
AOI221xp5_ASAP7_75t_L g1401 ( .A1(n_13), .A2(n_24), .B1(n_826), .B2(n_1402), .C(n_1404), .Y(n_1401) );
INVx1_ASAP7_75t_L g560 ( .A(n_14), .Y(n_560) );
OAI22xp5_ASAP7_75t_L g1098 ( .A1(n_15), .A2(n_52), .B1(n_1036), .B2(n_1099), .Y(n_1098) );
OAI22xp5_ASAP7_75t_L g1107 ( .A1(n_15), .A2(n_52), .B1(n_642), .B2(n_1108), .Y(n_1107) );
INVx1_ASAP7_75t_L g1568 ( .A(n_16), .Y(n_1568) );
AOI22xp33_ASAP7_75t_L g776 ( .A1(n_17), .A2(n_325), .B1(n_706), .B2(n_777), .Y(n_776) );
AOI22xp33_ASAP7_75t_L g825 ( .A1(n_17), .A2(n_369), .B1(n_826), .B2(n_827), .Y(n_825) );
AOI22xp33_ASAP7_75t_L g1645 ( .A1(n_18), .A2(n_199), .B1(n_771), .B2(n_1646), .Y(n_1645) );
INVx1_ASAP7_75t_L g1656 ( .A(n_18), .Y(n_1656) );
AOI22xp33_ASAP7_75t_L g1276 ( .A1(n_19), .A2(n_33), .B1(n_715), .B2(n_1248), .Y(n_1276) );
INVx1_ASAP7_75t_L g1316 ( .A(n_19), .Y(n_1316) );
INVx1_ASAP7_75t_L g859 ( .A(n_20), .Y(n_859) );
INVx1_ASAP7_75t_L g928 ( .A(n_21), .Y(n_928) );
INVx1_ASAP7_75t_L g1030 ( .A(n_22), .Y(n_1030) );
OAI22xp33_ASAP7_75t_L g1980 ( .A1(n_23), .A2(n_186), .B1(n_901), .B2(n_902), .Y(n_1980) );
OAI22xp33_ASAP7_75t_L g1982 ( .A1(n_23), .A2(n_186), .B1(n_641), .B2(n_1167), .Y(n_1982) );
AOI22xp33_ASAP7_75t_SL g1393 ( .A1(n_24), .A2(n_266), .B1(n_704), .B2(n_715), .Y(n_1393) );
INVx2_ASAP7_75t_L g394 ( .A(n_25), .Y(n_394) );
AOI22xp5_ASAP7_75t_L g1726 ( .A1(n_26), .A2(n_29), .B1(n_1690), .B2(n_1698), .Y(n_1726) );
AOI22xp33_ASAP7_75t_L g1603 ( .A1(n_27), .A2(n_374), .B1(n_846), .B2(n_1604), .Y(n_1603) );
INVx1_ASAP7_75t_L g1612 ( .A(n_27), .Y(n_1612) );
OAI22xp33_ASAP7_75t_L g888 ( .A1(n_28), .A2(n_314), .B1(n_508), .B2(n_641), .Y(n_888) );
OAI22xp5_ASAP7_75t_L g900 ( .A1(n_28), .A2(n_314), .B1(n_901), .B2(n_902), .Y(n_900) );
INVx1_ASAP7_75t_L g1492 ( .A(n_30), .Y(n_1492) );
INVx1_ASAP7_75t_L g1926 ( .A(n_31), .Y(n_1926) );
INVx1_ASAP7_75t_L g425 ( .A(n_32), .Y(n_425) );
AOI221xp5_ASAP7_75t_L g1293 ( .A1(n_33), .A2(n_51), .B1(n_846), .B2(n_1294), .C(n_1296), .Y(n_1293) );
INVx1_ASAP7_75t_L g1003 ( .A(n_34), .Y(n_1003) );
INVx1_ASAP7_75t_L g1390 ( .A(n_35), .Y(n_1390) );
INVx1_ASAP7_75t_L g584 ( .A(n_36), .Y(n_584) );
OAI22xp5_ASAP7_75t_L g1158 ( .A1(n_37), .A2(n_318), .B1(n_540), .B2(n_633), .Y(n_1158) );
OAI22xp5_ASAP7_75t_L g1168 ( .A1(n_37), .A2(n_347), .B1(n_644), .B2(n_646), .Y(n_1168) );
INVx1_ASAP7_75t_L g677 ( .A(n_38), .Y(n_677) );
OA222x2_ASAP7_75t_L g1184 ( .A1(n_39), .A2(n_95), .B1(n_276), .B2(n_1185), .C1(n_1187), .C2(n_1193), .Y(n_1184) );
INVx1_ASAP7_75t_L g1245 ( .A(n_39), .Y(n_1245) );
HB1xp67_ASAP7_75t_L g1677 ( .A(n_40), .Y(n_1677) );
AND2x2_ASAP7_75t_L g1691 ( .A(n_40), .B(n_1675), .Y(n_1691) );
AOI22xp33_ASAP7_75t_L g1771 ( .A1(n_41), .A2(n_228), .B1(n_1698), .B2(n_1722), .Y(n_1771) );
INVx1_ASAP7_75t_L g1448 ( .A(n_42), .Y(n_1448) );
AOI22xp33_ASAP7_75t_L g1340 ( .A1(n_43), .A2(n_352), .B1(n_671), .B2(n_745), .Y(n_1340) );
INVxp67_ASAP7_75t_SL g1358 ( .A(n_43), .Y(n_1358) );
AOI22xp33_ASAP7_75t_L g1592 ( .A1(n_44), .A2(n_236), .B1(n_728), .B2(n_1593), .Y(n_1592) );
AOI22xp33_ASAP7_75t_L g1618 ( .A1(n_44), .A2(n_296), .B1(n_780), .B2(n_1619), .Y(n_1618) );
AOI22xp33_ASAP7_75t_L g1277 ( .A1(n_45), .A2(n_247), .B1(n_706), .B2(n_1246), .Y(n_1277) );
INVx1_ASAP7_75t_L g1299 ( .A(n_45), .Y(n_1299) );
INVx1_ASAP7_75t_L g1574 ( .A(n_46), .Y(n_1574) );
INVx1_ASAP7_75t_L g1075 ( .A(n_47), .Y(n_1075) );
INVx1_ASAP7_75t_L g869 ( .A(n_48), .Y(n_869) );
OAI22xp5_ASAP7_75t_L g1032 ( .A1(n_49), .A2(n_300), .B1(n_639), .B2(n_642), .Y(n_1032) );
OAI22xp5_ASAP7_75t_L g1039 ( .A1(n_49), .A2(n_212), .B1(n_633), .B2(n_693), .Y(n_1039) );
OAI22xp33_ASAP7_75t_L g965 ( .A1(n_50), .A2(n_211), .B1(n_966), .B2(n_968), .Y(n_965) );
OAI22xp33_ASAP7_75t_L g984 ( .A1(n_50), .A2(n_211), .B1(n_508), .B2(n_641), .Y(n_984) );
AOI22xp33_ASAP7_75t_SL g1282 ( .A1(n_51), .A2(n_344), .B1(n_715), .B2(n_1283), .Y(n_1282) );
INVxp67_ASAP7_75t_SL g1389 ( .A(n_53), .Y(n_1389) );
OAI22xp5_ASAP7_75t_L g1409 ( .A1(n_53), .A2(n_198), .B1(n_450), .B2(n_1410), .Y(n_1409) );
AOI22xp33_ASAP7_75t_SL g1042 ( .A1(n_54), .A2(n_145), .B1(n_1043), .B2(n_1044), .Y(n_1042) );
AOI22xp33_ASAP7_75t_SL g1062 ( .A1(n_54), .A2(n_280), .B1(n_1056), .B2(n_1063), .Y(n_1062) );
INVx1_ASAP7_75t_L g576 ( .A(n_55), .Y(n_576) );
INVx1_ASAP7_75t_L g1958 ( .A(n_56), .Y(n_1958) );
INVx1_ASAP7_75t_L g1917 ( .A(n_57), .Y(n_1917) );
INVx1_ASAP7_75t_L g923 ( .A(n_58), .Y(n_923) );
OAI211xp5_ASAP7_75t_L g889 ( .A1(n_59), .A2(n_653), .B(n_890), .C(n_891), .Y(n_889) );
INVx1_ASAP7_75t_L g906 ( .A(n_59), .Y(n_906) );
CKINVDCx5p33_ASAP7_75t_R g1211 ( .A(n_60), .Y(n_1211) );
INVx1_ASAP7_75t_L g1397 ( .A(n_61), .Y(n_1397) );
INVx1_ASAP7_75t_L g1136 ( .A(n_62), .Y(n_1136) );
INVx1_ASAP7_75t_L g1639 ( .A(n_63), .Y(n_1639) );
AOI21xp33_ASAP7_75t_L g1660 ( .A1(n_63), .A2(n_843), .B(n_1050), .Y(n_1660) );
AOI22xp33_ASAP7_75t_SL g1345 ( .A1(n_64), .A2(n_291), .B1(n_671), .B2(n_1346), .Y(n_1345) );
AOI22xp33_ASAP7_75t_L g1359 ( .A1(n_64), .A2(n_270), .B1(n_1063), .B2(n_1237), .Y(n_1359) );
INVx1_ASAP7_75t_L g1977 ( .A(n_65), .Y(n_1977) );
AOI22xp5_ASAP7_75t_L g1720 ( .A1(n_66), .A2(n_245), .B1(n_1690), .B2(n_1695), .Y(n_1720) );
CKINVDCx5p33_ASAP7_75t_R g1388 ( .A(n_67), .Y(n_1388) );
INVx1_ASAP7_75t_L g1420 ( .A(n_68), .Y(n_1420) );
AOI22xp5_ASAP7_75t_L g1706 ( .A1(n_68), .A2(n_363), .B1(n_1698), .B2(n_1707), .Y(n_1706) );
BUFx6f_ASAP7_75t_L g454 ( .A(n_69), .Y(n_454) );
AOI22xp33_ASAP7_75t_L g1278 ( .A1(n_70), .A2(n_85), .B1(n_1279), .B2(n_1281), .Y(n_1278) );
INVx1_ASAP7_75t_L g1298 ( .A(n_70), .Y(n_1298) );
INVx1_ASAP7_75t_L g1954 ( .A(n_71), .Y(n_1954) );
OAI22xp33_ASAP7_75t_SL g1335 ( .A1(n_72), .A2(n_279), .B1(n_607), .B2(n_1000), .Y(n_1335) );
INVx1_ASAP7_75t_L g1372 ( .A(n_72), .Y(n_1372) );
AOI22xp33_ASAP7_75t_L g1476 ( .A1(n_73), .A2(n_122), .B1(n_1191), .B2(n_1213), .Y(n_1476) );
AOI22xp33_ASAP7_75t_L g1501 ( .A1(n_73), .A2(n_256), .B1(n_706), .B2(n_707), .Y(n_1501) );
INVx1_ASAP7_75t_L g1635 ( .A(n_74), .Y(n_1635) );
OAI22xp5_ASAP7_75t_L g1650 ( .A1(n_74), .A2(n_337), .B1(n_1651), .B2(n_1652), .Y(n_1650) );
XNOR2xp5_ASAP7_75t_L g554 ( .A(n_75), .B(n_555), .Y(n_554) );
INVx1_ASAP7_75t_L g1452 ( .A(n_76), .Y(n_1452) );
INVx1_ASAP7_75t_L g1531 ( .A(n_77), .Y(n_1531) );
CKINVDCx5p33_ASAP7_75t_R g1269 ( .A(n_78), .Y(n_1269) );
XOR2x2_ASAP7_75t_L g1468 ( .A(n_79), .B(n_1469), .Y(n_1468) );
AOI22xp5_ASAP7_75t_L g1721 ( .A1(n_80), .A2(n_343), .B1(n_1698), .B2(n_1722), .Y(n_1721) );
INVx1_ASAP7_75t_L g862 ( .A(n_81), .Y(n_862) );
AOI22xp5_ASAP7_75t_L g1730 ( .A1(n_82), .A2(n_144), .B1(n_1690), .B2(n_1695), .Y(n_1730) );
AOI21xp33_ASAP7_75t_L g1602 ( .A1(n_83), .A2(n_732), .B(n_1339), .Y(n_1602) );
AOI22xp33_ASAP7_75t_L g1613 ( .A1(n_83), .A2(n_236), .B1(n_1248), .B2(n_1614), .Y(n_1613) );
AOI22xp33_ASAP7_75t_SL g730 ( .A1(n_84), .A2(n_118), .B1(n_731), .B2(n_734), .Y(n_730) );
INVx1_ASAP7_75t_L g1320 ( .A(n_85), .Y(n_1320) );
OAI211xp5_ASAP7_75t_L g1902 ( .A1(n_86), .A2(n_527), .B(n_1137), .C(n_1903), .Y(n_1902) );
INVx1_ASAP7_75t_L g1910 ( .A(n_86), .Y(n_1910) );
INVx1_ASAP7_75t_L g631 ( .A(n_87), .Y(n_631) );
OAI211xp5_ASAP7_75t_L g649 ( .A1(n_87), .A2(n_650), .B(n_653), .C(n_654), .Y(n_649) );
INVx1_ASAP7_75t_L g948 ( .A(n_88), .Y(n_948) );
OAI211xp5_ASAP7_75t_L g952 ( .A1(n_88), .A2(n_625), .B(n_904), .C(n_953), .Y(n_952) );
OAI22xp33_ASAP7_75t_L g757 ( .A1(n_89), .A2(n_332), .B1(n_758), .B2(n_764), .Y(n_757) );
INVx1_ASAP7_75t_L g813 ( .A(n_89), .Y(n_813) );
INVx1_ASAP7_75t_L g1419 ( .A(n_90), .Y(n_1419) );
INVx1_ASAP7_75t_L g1139 ( .A(n_91), .Y(n_1139) );
INVx1_ASAP7_75t_L g1925 ( .A(n_92), .Y(n_1925) );
INVx1_ASAP7_75t_L g921 ( .A(n_93), .Y(n_921) );
CKINVDCx5p33_ASAP7_75t_R g1585 ( .A(n_94), .Y(n_1585) );
OAI221xp5_ASAP7_75t_L g1230 ( .A1(n_95), .A2(n_223), .B1(n_1231), .B2(n_1233), .C(n_1235), .Y(n_1230) );
OAI22xp5_ASAP7_75t_L g1307 ( .A1(n_96), .A2(n_329), .B1(n_450), .B2(n_457), .Y(n_1307) );
INVx1_ASAP7_75t_L g1322 ( .A(n_96), .Y(n_1322) );
INVx1_ASAP7_75t_L g1201 ( .A(n_97), .Y(n_1201) );
AOI22xp33_ASAP7_75t_L g1261 ( .A1(n_97), .A2(n_159), .B1(n_709), .B2(n_780), .Y(n_1261) );
INVx1_ASAP7_75t_L g1923 ( .A(n_98), .Y(n_1923) );
XOR2x2_ASAP7_75t_L g1424 ( .A(n_99), .B(n_1425), .Y(n_1424) );
INVx1_ASAP7_75t_L g1005 ( .A(n_100), .Y(n_1005) );
OAI22xp5_ASAP7_75t_L g894 ( .A1(n_101), .A2(n_196), .B1(n_895), .B2(n_896), .Y(n_894) );
OAI22xp33_ASAP7_75t_L g907 ( .A1(n_101), .A2(n_196), .B1(n_621), .B2(n_908), .Y(n_907) );
INVx1_ASAP7_75t_L g396 ( .A(n_102), .Y(n_396) );
INVx1_ASAP7_75t_L g491 ( .A(n_103), .Y(n_491) );
INVx1_ASAP7_75t_L g676 ( .A(n_104), .Y(n_676) );
AOI22xp5_ASAP7_75t_L g1711 ( .A1(n_105), .A2(n_371), .B1(n_1690), .B2(n_1695), .Y(n_1711) );
AOI22xp33_ASAP7_75t_SL g714 ( .A1(n_106), .A2(n_193), .B1(n_715), .B2(n_717), .Y(n_714) );
AOI22xp33_ASAP7_75t_L g723 ( .A1(n_106), .A2(n_253), .B1(n_724), .B2(n_726), .Y(n_723) );
INVx1_ASAP7_75t_L g1429 ( .A(n_107), .Y(n_1429) );
XOR2x2_ASAP7_75t_L g1119 ( .A(n_108), .B(n_1120), .Y(n_1119) );
INVx1_ASAP7_75t_L g573 ( .A(n_109), .Y(n_573) );
XNOR2xp5_ASAP7_75t_L g911 ( .A(n_110), .B(n_912), .Y(n_911) );
CKINVDCx5p33_ASAP7_75t_R g1396 ( .A(n_111), .Y(n_1396) );
INVx1_ASAP7_75t_L g1905 ( .A(n_112), .Y(n_1905) );
OAI211xp5_ASAP7_75t_L g1908 ( .A1(n_112), .A2(n_481), .B(n_1449), .C(n_1909), .Y(n_1908) );
AOI22xp33_ASAP7_75t_SL g779 ( .A1(n_113), .A2(n_282), .B1(n_718), .B2(n_780), .Y(n_779) );
AOI221xp5_ASAP7_75t_L g820 ( .A1(n_113), .A2(n_335), .B1(n_821), .B2(n_823), .C(n_824), .Y(n_820) );
AOI22xp33_ASAP7_75t_L g1392 ( .A1(n_114), .A2(n_348), .B1(n_707), .B2(n_1279), .Y(n_1392) );
AOI221xp5_ASAP7_75t_L g1416 ( .A1(n_114), .A2(n_242), .B1(n_671), .B2(n_846), .C(n_1417), .Y(n_1416) );
OAI211xp5_ASAP7_75t_L g1516 ( .A1(n_115), .A2(n_481), .B(n_1156), .C(n_1517), .Y(n_1516) );
INVx1_ASAP7_75t_L g1525 ( .A(n_115), .Y(n_1525) );
AOI22xp5_ASAP7_75t_SL g1712 ( .A1(n_116), .A2(n_252), .B1(n_1698), .B2(n_1707), .Y(n_1712) );
INVx1_ASAP7_75t_L g1955 ( .A(n_117), .Y(n_1955) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_118), .A2(n_250), .B1(n_706), .B2(n_707), .Y(n_705) );
INVx1_ASAP7_75t_L g1325 ( .A(n_119), .Y(n_1325) );
INVx1_ASAP7_75t_L g1922 ( .A(n_120), .Y(n_1922) );
INVx1_ASAP7_75t_L g892 ( .A(n_121), .Y(n_892) );
AOI22xp33_ASAP7_75t_L g1502 ( .A1(n_122), .A2(n_143), .B1(n_570), .B2(n_1281), .Y(n_1502) );
INVx1_ASAP7_75t_L g1644 ( .A(n_123), .Y(n_1644) );
AOI22xp33_ASAP7_75t_L g1658 ( .A1(n_123), .A2(n_283), .B1(n_671), .B2(n_745), .Y(n_1658) );
CKINVDCx5p33_ASAP7_75t_R g1584 ( .A(n_124), .Y(n_1584) );
INVx1_ASAP7_75t_L g1675 ( .A(n_125), .Y(n_1675) );
INVx1_ASAP7_75t_L g568 ( .A(n_126), .Y(n_568) );
XOR2x2_ASAP7_75t_L g962 ( .A(n_127), .B(n_963), .Y(n_962) );
OAI22xp5_ASAP7_75t_L g1493 ( .A1(n_128), .A2(n_194), .B1(n_1324), .B2(n_1494), .Y(n_1493) );
INVx1_ASAP7_75t_L g1126 ( .A(n_129), .Y(n_1126) );
OAI211xp5_ASAP7_75t_L g1427 ( .A1(n_130), .A2(n_481), .B(n_1353), .C(n_1428), .Y(n_1427) );
INVx1_ASAP7_75t_L g1437 ( .A(n_130), .Y(n_1437) );
OAI22xp5_ASAP7_75t_L g949 ( .A1(n_131), .A2(n_180), .B1(n_895), .B2(n_896), .Y(n_949) );
OAI22xp33_ASAP7_75t_L g956 ( .A1(n_131), .A2(n_180), .B1(n_621), .B2(n_957), .Y(n_956) );
INVx1_ASAP7_75t_L g1519 ( .A(n_132), .Y(n_1519) );
OAI211xp5_ASAP7_75t_L g1522 ( .A1(n_132), .A2(n_625), .B(n_1523), .C(n_1524), .Y(n_1522) );
INVxp67_ASAP7_75t_SL g1487 ( .A(n_133), .Y(n_1487) );
AOI22xp33_ASAP7_75t_L g1503 ( .A1(n_133), .A2(n_305), .B1(n_773), .B2(n_1283), .Y(n_1503) );
AOI22xp5_ASAP7_75t_L g1714 ( .A1(n_134), .A2(n_351), .B1(n_1695), .B2(n_1707), .Y(n_1714) );
OAI22xp5_ASAP7_75t_L g1334 ( .A1(n_135), .A2(n_175), .B1(n_1076), .B2(n_1202), .Y(n_1334) );
NOR2xp33_ASAP7_75t_L g1376 ( .A(n_135), .B(n_1377), .Y(n_1376) );
INVx1_ASAP7_75t_L g439 ( .A(n_136), .Y(n_439) );
CKINVDCx5p33_ASAP7_75t_R g1289 ( .A(n_137), .Y(n_1289) );
INVx1_ASAP7_75t_L g428 ( .A(n_138), .Y(n_428) );
INVx1_ASAP7_75t_L g436 ( .A(n_139), .Y(n_436) );
OAI22xp5_ASAP7_75t_L g498 ( .A1(n_140), .A2(n_155), .B1(n_499), .B2(n_502), .Y(n_498) );
OAI22xp33_ASAP7_75t_L g539 ( .A1(n_140), .A2(n_155), .B1(n_540), .B2(n_543), .Y(n_539) );
INVx1_ASAP7_75t_L g864 ( .A(n_141), .Y(n_864) );
INVx1_ASAP7_75t_L g1455 ( .A(n_142), .Y(n_1455) );
AOI221xp5_ASAP7_75t_L g1488 ( .A1(n_143), .A2(n_256), .B1(n_843), .B2(n_1050), .C(n_1489), .Y(n_1488) );
AOI22xp33_ASAP7_75t_L g1053 ( .A1(n_145), .A2(n_258), .B1(n_717), .B2(n_1054), .Y(n_1053) );
AOI22xp33_ASAP7_75t_L g774 ( .A1(n_146), .A2(n_369), .B1(n_706), .B2(n_775), .Y(n_774) );
AOI21xp33_ASAP7_75t_L g840 ( .A1(n_146), .A2(n_841), .B(n_843), .Y(n_840) );
INVx1_ASAP7_75t_L g999 ( .A(n_147), .Y(n_999) );
INVx1_ASAP7_75t_L g497 ( .A(n_148), .Y(n_497) );
OAI211xp5_ASAP7_75t_L g523 ( .A1(n_148), .A2(n_524), .B(n_527), .C(n_531), .Y(n_523) );
OAI22xp5_ASAP7_75t_L g1163 ( .A1(n_149), .A2(n_347), .B1(n_622), .B2(n_1164), .Y(n_1163) );
OAI22xp33_ASAP7_75t_L g1166 ( .A1(n_149), .A2(n_318), .B1(n_641), .B2(n_1167), .Y(n_1166) );
INVx1_ASAP7_75t_L g404 ( .A(n_150), .Y(n_404) );
AOI22xp33_ASAP7_75t_SL g1641 ( .A1(n_151), .A2(n_306), .B1(n_686), .B2(n_1056), .Y(n_1641) );
AOI21xp33_ASAP7_75t_L g1657 ( .A1(n_151), .A2(n_841), .B(n_1339), .Y(n_1657) );
INVx1_ASAP7_75t_L g1904 ( .A(n_152), .Y(n_1904) );
INVx1_ASAP7_75t_L g1957 ( .A(n_153), .Y(n_1957) );
INVx1_ASAP7_75t_L g674 ( .A(n_154), .Y(n_674) );
INVx1_ASAP7_75t_L g947 ( .A(n_156), .Y(n_947) );
INVx1_ASAP7_75t_L g1104 ( .A(n_157), .Y(n_1104) );
OAI211xp5_ASAP7_75t_L g1110 ( .A1(n_157), .A2(n_1111), .B(n_1112), .C(n_1114), .Y(n_1110) );
OAI211xp5_ASAP7_75t_L g1972 ( .A1(n_158), .A2(n_625), .B(n_1973), .C(n_1976), .Y(n_1972) );
INVx1_ASAP7_75t_L g1986 ( .A(n_158), .Y(n_1986) );
AOI22xp33_ASAP7_75t_L g1212 ( .A1(n_159), .A2(n_207), .B1(n_1191), .B2(n_1213), .Y(n_1212) );
INVx1_ASAP7_75t_L g917 ( .A(n_160), .Y(n_917) );
AOI221xp5_ASAP7_75t_L g1474 ( .A1(n_161), .A2(n_305), .B1(n_823), .B2(n_824), .C(n_1475), .Y(n_1474) );
AOI22xp33_ASAP7_75t_L g1498 ( .A1(n_161), .A2(n_261), .B1(n_704), .B2(n_1499), .Y(n_1498) );
OAI22xp5_ASAP7_75t_L g1431 ( .A1(n_162), .A2(n_358), .B1(n_895), .B2(n_896), .Y(n_1431) );
OAI22xp5_ASAP7_75t_L g1434 ( .A1(n_162), .A2(n_358), .B1(n_543), .B2(n_1377), .Y(n_1434) );
INVx1_ASAP7_75t_L g1965 ( .A(n_163), .Y(n_1965) );
OAI22xp5_ASAP7_75t_L g1218 ( .A1(n_164), .A2(n_223), .B1(n_802), .B2(n_1219), .Y(n_1218) );
INVx1_ASAP7_75t_L g1247 ( .A(n_164), .Y(n_1247) );
INVx1_ASAP7_75t_L g1920 ( .A(n_165), .Y(n_1920) );
INVx1_ASAP7_75t_L g1082 ( .A(n_166), .Y(n_1082) );
OAI22xp33_ASAP7_75t_L g1432 ( .A1(n_167), .A2(n_214), .B1(n_506), .B2(n_1167), .Y(n_1432) );
OAI22xp33_ASAP7_75t_L g1438 ( .A1(n_167), .A2(n_214), .B1(n_518), .B2(n_635), .Y(n_1438) );
OAI22xp33_ASAP7_75t_L g505 ( .A1(n_168), .A2(n_272), .B1(n_506), .B2(n_508), .Y(n_505) );
OAI22xp33_ASAP7_75t_L g517 ( .A1(n_168), .A2(n_272), .B1(n_518), .B2(n_519), .Y(n_517) );
INVx1_ASAP7_75t_L g786 ( .A(n_169), .Y(n_786) );
OAI221xp5_ASAP7_75t_L g829 ( .A1(n_169), .A2(n_226), .B1(n_830), .B2(n_834), .C(n_838), .Y(n_829) );
OAI22xp33_ASAP7_75t_L g1906 ( .A1(n_171), .A2(n_190), .B1(n_635), .B2(n_1099), .Y(n_1906) );
OAI22xp33_ASAP7_75t_L g1912 ( .A1(n_171), .A2(n_190), .B1(n_506), .B2(n_1167), .Y(n_1912) );
OAI221xp5_ASAP7_75t_L g1349 ( .A1(n_172), .A2(n_355), .B1(n_1350), .B2(n_1352), .C(n_1353), .Y(n_1349) );
INVx1_ASAP7_75t_L g1369 ( .A(n_172), .Y(n_1369) );
INVx1_ASAP7_75t_L g1337 ( .A(n_173), .Y(n_1337) );
AOI22xp33_ASAP7_75t_L g1364 ( .A1(n_173), .A2(n_291), .B1(n_718), .B2(n_1237), .Y(n_1364) );
CKINVDCx5p33_ASAP7_75t_R g1342 ( .A(n_174), .Y(n_1342) );
INVx1_ASAP7_75t_L g1371 ( .A(n_175), .Y(n_1371) );
INVx1_ASAP7_75t_L g974 ( .A(n_176), .Y(n_974) );
OAI211xp5_ASAP7_75t_L g977 ( .A1(n_176), .A2(n_652), .B(n_978), .C(n_979), .Y(n_977) );
INVx1_ASAP7_75t_L g1029 ( .A(n_177), .Y(n_1029) );
OAI211xp5_ASAP7_75t_L g1037 ( .A1(n_177), .A2(n_625), .B(n_873), .C(n_1038), .Y(n_1037) );
OAI211xp5_ASAP7_75t_L g1159 ( .A1(n_178), .A2(n_527), .B(n_873), .C(n_1160), .Y(n_1159) );
INVx1_ASAP7_75t_L g1172 ( .A(n_178), .Y(n_1172) );
OAI22xp33_ASAP7_75t_L g632 ( .A1(n_179), .A2(n_285), .B1(n_633), .B2(n_635), .Y(n_632) );
OAI22xp5_ASAP7_75t_L g638 ( .A1(n_179), .A2(n_285), .B1(n_639), .B2(n_642), .Y(n_638) );
INVx1_ASAP7_75t_L g1518 ( .A(n_181), .Y(n_1518) );
INVx1_ASAP7_75t_L g564 ( .A(n_182), .Y(n_564) );
INVx1_ASAP7_75t_L g996 ( .A(n_183), .Y(n_996) );
INVx1_ASAP7_75t_L g580 ( .A(n_184), .Y(n_580) );
INVx1_ASAP7_75t_L g1962 ( .A(n_185), .Y(n_1962) );
OAI22xp33_ASAP7_75t_L g620 ( .A1(n_187), .A2(n_221), .B1(n_621), .B2(n_622), .Y(n_620) );
OAI22xp33_ASAP7_75t_L g643 ( .A1(n_187), .A2(n_221), .B1(n_644), .B2(n_646), .Y(n_643) );
INVx1_ASAP7_75t_L g872 ( .A(n_188), .Y(n_872) );
INVx1_ASAP7_75t_L g931 ( .A(n_189), .Y(n_931) );
XNOR2xp5_ASAP7_75t_L g664 ( .A(n_191), .B(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g1001 ( .A(n_192), .Y(n_1001) );
AOI22xp33_ASAP7_75t_SL g739 ( .A1(n_193), .A2(n_331), .B1(n_731), .B2(n_740), .Y(n_739) );
OAI211xp5_ASAP7_75t_L g1471 ( .A1(n_194), .A2(n_1472), .B(n_1473), .C(n_1477), .Y(n_1471) );
AOI221xp5_ASAP7_75t_L g1588 ( .A1(n_195), .A2(n_361), .B1(n_1199), .B2(n_1589), .C(n_1591), .Y(n_1588) );
AOI22xp33_ASAP7_75t_L g1617 ( .A1(n_195), .A2(n_374), .B1(n_777), .B2(n_927), .Y(n_1617) );
XOR2x2_ASAP7_75t_L g1069 ( .A(n_197), .B(n_1070), .Y(n_1069) );
INVxp67_ASAP7_75t_SL g1399 ( .A(n_198), .Y(n_1399) );
AOI22xp33_ASAP7_75t_L g1661 ( .A1(n_199), .A2(n_306), .B1(n_671), .B2(n_745), .Y(n_1661) );
CKINVDCx5p33_ASAP7_75t_R g1208 ( .A(n_200), .Y(n_1208) );
INVx1_ASAP7_75t_L g1919 ( .A(n_201), .Y(n_1919) );
INVx1_ASAP7_75t_L g1103 ( .A(n_202), .Y(n_1103) );
INVx1_ASAP7_75t_L g1086 ( .A(n_203), .Y(n_1086) );
INVx1_ASAP7_75t_L g1328 ( .A(n_204), .Y(n_1328) );
INVx1_ASAP7_75t_L g1768 ( .A(n_205), .Y(n_1768) );
INVx1_ASAP7_75t_L g679 ( .A(n_206), .Y(n_679) );
OAI22xp5_ASAP7_75t_L g688 ( .A1(n_206), .A2(n_323), .B1(n_689), .B2(n_690), .Y(n_688) );
INVx1_ASAP7_75t_L g1257 ( .A(n_207), .Y(n_1257) );
XNOR2xp5_ASAP7_75t_L g852 ( .A(n_208), .B(n_853), .Y(n_852) );
AOI22xp5_ASAP7_75t_SL g1729 ( .A1(n_208), .A2(n_218), .B1(n_1698), .B2(n_1707), .Y(n_1729) );
INVx1_ASAP7_75t_L g930 ( .A(n_209), .Y(n_930) );
INVx1_ASAP7_75t_L g1451 ( .A(n_210), .Y(n_1451) );
INVx1_ASAP7_75t_L g1027 ( .A(n_212), .Y(n_1027) );
INVx1_ASAP7_75t_L g1430 ( .A(n_213), .Y(n_1430) );
OAI211xp5_ASAP7_75t_L g1435 ( .A1(n_213), .A2(n_524), .B(n_527), .C(n_1436), .Y(n_1435) );
OAI22xp33_ASAP7_75t_L g1979 ( .A1(n_215), .A2(n_364), .B1(n_540), .B2(n_622), .Y(n_1979) );
OAI22xp33_ASAP7_75t_L g1983 ( .A1(n_215), .A2(n_364), .B1(n_644), .B2(n_646), .Y(n_1983) );
INVx1_ASAP7_75t_L g990 ( .A(n_216), .Y(n_990) );
AOI221x1_ASAP7_75t_SL g1195 ( .A1(n_217), .A2(n_288), .B1(n_1196), .B2(n_1198), .C(n_1200), .Y(n_1195) );
AOI21xp33_ASAP7_75t_L g1259 ( .A1(n_217), .A2(n_767), .B(n_1260), .Y(n_1259) );
INVx1_ASAP7_75t_L g1478 ( .A(n_219), .Y(n_1478) );
OAI22xp33_ASAP7_75t_L g1507 ( .A1(n_219), .A2(n_333), .B1(n_764), .B2(n_1508), .Y(n_1507) );
OAI221xp5_ASAP7_75t_L g1481 ( .A1(n_220), .A2(n_289), .B1(n_1482), .B2(n_1483), .C(n_1485), .Y(n_1481) );
INVx1_ASAP7_75t_L g1505 ( .A(n_220), .Y(n_1505) );
INVx2_ASAP7_75t_L g1693 ( .A(n_222), .Y(n_1693) );
AND2x2_ASAP7_75t_L g1696 ( .A(n_222), .B(n_1694), .Y(n_1696) );
AND2x2_ASAP7_75t_L g1701 ( .A(n_222), .B(n_326), .Y(n_1701) );
OAI22xp33_ASAP7_75t_L g1105 ( .A1(n_224), .A2(n_287), .B1(n_543), .B2(n_693), .Y(n_1105) );
OAI22xp33_ASAP7_75t_L g1116 ( .A1(n_224), .A2(n_287), .B1(n_895), .B2(n_1117), .Y(n_1116) );
AOI22xp5_ASAP7_75t_SL g1725 ( .A1(n_225), .A2(n_286), .B1(n_1695), .B2(n_1700), .Y(n_1725) );
INVx1_ASAP7_75t_L g782 ( .A(n_226), .Y(n_782) );
INVx1_ASAP7_75t_L g1031 ( .A(n_227), .Y(n_1031) );
AOI22xp5_ASAP7_75t_L g1697 ( .A1(n_229), .A2(n_349), .B1(n_1698), .B2(n_1700), .Y(n_1697) );
INVx1_ASAP7_75t_L g973 ( .A(n_230), .Y(n_973) );
INVx1_ASAP7_75t_L g1161 ( .A(n_231), .Y(n_1161) );
OAI22xp5_ASAP7_75t_L g1565 ( .A1(n_232), .A2(n_1566), .B1(n_1620), .B2(n_1621), .Y(n_1565) );
INVxp67_ASAP7_75t_L g1621 ( .A(n_232), .Y(n_1621) );
AOI22xp5_ASAP7_75t_L g1705 ( .A1(n_233), .A2(n_290), .B1(n_1690), .B2(n_1695), .Y(n_1705) );
CKINVDCx5p33_ASAP7_75t_R g1203 ( .A(n_234), .Y(n_1203) );
AOI22xp33_ASAP7_75t_L g1045 ( .A1(n_235), .A2(n_360), .B1(n_724), .B2(n_740), .Y(n_1045) );
AOI22xp33_ASAP7_75t_L g1058 ( .A1(n_235), .A2(n_241), .B1(n_1059), .B2(n_1061), .Y(n_1058) );
XOR2x2_ASAP7_75t_L g1509 ( .A(n_237), .B(n_1510), .Y(n_1509) );
INVx1_ASAP7_75t_L g857 ( .A(n_238), .Y(n_857) );
AOI22xp5_ASAP7_75t_L g1715 ( .A1(n_239), .A2(n_307), .B1(n_1690), .B2(n_1698), .Y(n_1715) );
OAI221xp5_ASAP7_75t_SL g1580 ( .A1(n_240), .A2(n_320), .B1(n_1581), .B2(n_1582), .C(n_1583), .Y(n_1580) );
INVx1_ASAP7_75t_L g1598 ( .A(n_240), .Y(n_1598) );
AOI22xp33_ASAP7_75t_SL g1051 ( .A1(n_241), .A2(n_357), .B1(n_724), .B2(n_744), .Y(n_1051) );
AOI22xp33_ASAP7_75t_L g1383 ( .A1(n_242), .A2(n_336), .B1(n_570), .B2(n_1281), .Y(n_1383) );
INVx1_ASAP7_75t_L g1079 ( .A(n_243), .Y(n_1079) );
INVx1_ASAP7_75t_L g1143 ( .A(n_244), .Y(n_1143) );
OAI22xp5_ASAP7_75t_L g1901 ( .A1(n_246), .A2(n_263), .B1(n_622), .B2(n_693), .Y(n_1901) );
OAI22xp5_ASAP7_75t_L g1911 ( .A1(n_246), .A2(n_263), .B1(n_895), .B2(n_896), .Y(n_1911) );
INVx1_ASAP7_75t_L g1318 ( .A(n_247), .Y(n_1318) );
INVx1_ASAP7_75t_L g1080 ( .A(n_248), .Y(n_1080) );
INVx2_ASAP7_75t_L g393 ( .A(n_249), .Y(n_393) );
INVx1_ASAP7_75t_L g433 ( .A(n_249), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_249), .B(n_394), .Y(n_763) );
XNOR2xp5_ASAP7_75t_L g746 ( .A(n_251), .B(n_747), .Y(n_746) );
AOI22xp33_ASAP7_75t_SL g699 ( .A1(n_253), .A2(n_331), .B1(n_700), .B2(n_704), .Y(n_699) );
OAI22xp33_ASAP7_75t_L g944 ( .A1(n_254), .A2(n_284), .B1(n_508), .B2(n_641), .Y(n_944) );
OAI22xp5_ASAP7_75t_L g951 ( .A1(n_254), .A2(n_284), .B1(n_635), .B2(n_901), .Y(n_951) );
BUFx3_ASAP7_75t_L g401 ( .A(n_255), .Y(n_401) );
INVx1_ASAP7_75t_L g1571 ( .A(n_257), .Y(n_1571) );
AOI22xp33_ASAP7_75t_SL g1048 ( .A1(n_258), .A2(n_280), .B1(n_734), .B2(n_1049), .Y(n_1048) );
INVx1_ASAP7_75t_L g1088 ( .A(n_259), .Y(n_1088) );
INVx1_ASAP7_75t_L g1978 ( .A(n_260), .Y(n_1978) );
OAI211xp5_ASAP7_75t_L g1984 ( .A1(n_260), .A2(n_650), .B(n_653), .C(n_1985), .Y(n_1984) );
INVxp67_ASAP7_75t_SL g1486 ( .A(n_261), .Y(n_1486) );
INVx1_ASAP7_75t_L g867 ( .A(n_262), .Y(n_867) );
AOI22xp5_ASAP7_75t_L g1689 ( .A1(n_264), .A2(n_302), .B1(n_1690), .B2(n_1695), .Y(n_1689) );
OA22x2_ASAP7_75t_L g1898 ( .A1(n_264), .A2(n_1899), .B1(n_1935), .B2(n_1936), .Y(n_1898) );
INVxp67_ASAP7_75t_L g1936 ( .A(n_264), .Y(n_1936) );
AOI22xp33_ASAP7_75t_L g1943 ( .A1(n_264), .A2(n_1944), .B1(n_1947), .B2(n_1987), .Y(n_1943) );
AOI22xp33_ASAP7_75t_L g770 ( .A1(n_265), .A2(n_335), .B1(n_704), .B2(n_771), .Y(n_770) );
AOI22xp33_ASAP7_75t_L g845 ( .A1(n_265), .A2(n_282), .B1(n_826), .B2(n_846), .Y(n_845) );
INVx1_ASAP7_75t_L g1418 ( .A(n_266), .Y(n_1418) );
INVx1_ASAP7_75t_L g1444 ( .A(n_267), .Y(n_1444) );
INVx1_ASAP7_75t_L g893 ( .A(n_268), .Y(n_893) );
OAI211xp5_ASAP7_75t_SL g903 ( .A1(n_268), .A2(n_527), .B(n_904), .C(n_905), .Y(n_903) );
INVx1_ASAP7_75t_L g988 ( .A(n_269), .Y(n_988) );
AOI21xp33_ASAP7_75t_L g1338 ( .A1(n_270), .A2(n_732), .B(n_1339), .Y(n_1338) );
XNOR2xp5_ASAP7_75t_L g1948 ( .A(n_271), .B(n_1949), .Y(n_1948) );
INVx1_ASAP7_75t_L g1132 ( .A(n_273), .Y(n_1132) );
INVx1_ASAP7_75t_L g1534 ( .A(n_274), .Y(n_1534) );
INVx1_ASAP7_75t_L g993 ( .A(n_275), .Y(n_993) );
INVx1_ASAP7_75t_L g1236 ( .A(n_276), .Y(n_1236) );
INVx1_ASAP7_75t_L g1631 ( .A(n_277), .Y(n_1631) );
INVx1_ASAP7_75t_L g583 ( .A(n_278), .Y(n_583) );
INVx1_ASAP7_75t_L g1375 ( .A(n_279), .Y(n_1375) );
BUFx3_ASAP7_75t_L g446 ( .A(n_281), .Y(n_446) );
INVx1_ASAP7_75t_L g501 ( .A(n_281), .Y(n_501) );
INVx1_ASAP7_75t_L g1640 ( .A(n_283), .Y(n_1640) );
XNOR2xp5_ASAP7_75t_L g383 ( .A(n_286), .B(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g1256 ( .A(n_288), .Y(n_1256) );
INVx1_ASAP7_75t_L g1506 ( .A(n_289), .Y(n_1506) );
INVx1_ASAP7_75t_L g1182 ( .A(n_293), .Y(n_1182) );
INVx1_ASAP7_75t_L g419 ( .A(n_294), .Y(n_419) );
INVx1_ASAP7_75t_L g1542 ( .A(n_295), .Y(n_1542) );
INVx1_ASAP7_75t_L g1601 ( .A(n_296), .Y(n_1601) );
INVx1_ASAP7_75t_L g1129 ( .A(n_297), .Y(n_1129) );
INVx1_ASAP7_75t_L g925 ( .A(n_298), .Y(n_925) );
INVx1_ASAP7_75t_L g1447 ( .A(n_299), .Y(n_1447) );
OAI22xp5_ASAP7_75t_L g1035 ( .A1(n_300), .A2(n_375), .B1(n_543), .B2(n_1036), .Y(n_1035) );
INVx1_ASAP7_75t_L g1541 ( .A(n_301), .Y(n_1541) );
CKINVDCx5p33_ASAP7_75t_R g1291 ( .A(n_304), .Y(n_1291) );
INVx1_ASAP7_75t_L g1538 ( .A(n_308), .Y(n_1538) );
INVx1_ASAP7_75t_L g403 ( .A(n_309), .Y(n_403) );
INVx1_ASAP7_75t_L g410 ( .A(n_309), .Y(n_410) );
OAI22xp5_ASAP7_75t_L g1622 ( .A1(n_311), .A2(n_1623), .B1(n_1624), .B2(n_1666), .Y(n_1622) );
INVxp67_ASAP7_75t_L g1666 ( .A(n_311), .Y(n_1666) );
INVx1_ASAP7_75t_L g1548 ( .A(n_312), .Y(n_1548) );
INVx1_ASAP7_75t_L g1960 ( .A(n_313), .Y(n_1960) );
INVxp67_ASAP7_75t_SL g1628 ( .A(n_315), .Y(n_1628) );
OAI221xp5_ASAP7_75t_L g1663 ( .A1(n_315), .A2(n_362), .B1(n_796), .B2(n_1484), .C(n_1664), .Y(n_1663) );
INVx1_ASAP7_75t_L g1131 ( .A(n_316), .Y(n_1131) );
OAI211xp5_ASAP7_75t_L g945 ( .A1(n_317), .A2(n_653), .B(n_890), .C(n_946), .Y(n_945) );
INVx1_ASAP7_75t_L g955 ( .A(n_317), .Y(n_955) );
INVx1_ASAP7_75t_L g629 ( .A(n_319), .Y(n_629) );
INVx1_ASAP7_75t_L g1607 ( .A(n_320), .Y(n_1607) );
CKINVDCx5p33_ASAP7_75t_R g1632 ( .A(n_321), .Y(n_1632) );
INVx1_ASAP7_75t_L g1084 ( .A(n_322), .Y(n_1084) );
INVx1_ASAP7_75t_L g681 ( .A(n_323), .Y(n_681) );
CKINVDCx5p33_ASAP7_75t_R g1285 ( .A(n_324), .Y(n_1285) );
INVxp67_ASAP7_75t_SL g839 ( .A(n_325), .Y(n_839) );
INVx1_ASAP7_75t_L g1694 ( .A(n_326), .Y(n_1694) );
AND2x2_ASAP7_75t_L g1699 ( .A(n_326), .B(n_1693), .Y(n_1699) );
OAI211xp5_ASAP7_75t_SL g623 ( .A1(n_327), .A2(n_624), .B(n_625), .C(n_626), .Y(n_623) );
INVx1_ASAP7_75t_L g658 ( .A(n_327), .Y(n_658) );
INVx1_ASAP7_75t_L g682 ( .A(n_328), .Y(n_682) );
INVx1_ASAP7_75t_L g1272 ( .A(n_329), .Y(n_1272) );
OAI211xp5_ASAP7_75t_L g1101 ( .A1(n_330), .A2(n_527), .B(n_971), .C(n_1102), .Y(n_1101) );
INVx1_ASAP7_75t_L g1115 ( .A(n_330), .Y(n_1115) );
INVx1_ASAP7_75t_L g816 ( .A(n_332), .Y(n_816) );
INVx1_ASAP7_75t_L g1479 ( .A(n_333), .Y(n_1479) );
INVx1_ASAP7_75t_L g1442 ( .A(n_334), .Y(n_1442) );
INVx1_ASAP7_75t_L g1406 ( .A(n_336), .Y(n_1406) );
INVx1_ASAP7_75t_L g1636 ( .A(n_337), .Y(n_1636) );
INVx1_ASAP7_75t_L g1348 ( .A(n_338), .Y(n_1348) );
INVx1_ASAP7_75t_L g918 ( .A(n_339), .Y(n_918) );
INVx1_ASAP7_75t_L g1770 ( .A(n_340), .Y(n_1770) );
CKINVDCx5p33_ASAP7_75t_R g1643 ( .A(n_341), .Y(n_1643) );
INVx1_ASAP7_75t_L g1547 ( .A(n_342), .Y(n_1547) );
OAI22xp5_ASAP7_75t_L g1020 ( .A1(n_343), .A2(n_1021), .B1(n_1064), .B2(n_1065), .Y(n_1020) );
INVxp67_ASAP7_75t_SL g1065 ( .A(n_343), .Y(n_1065) );
AOI211xp5_ASAP7_75t_SL g1314 ( .A1(n_344), .A2(n_680), .B(n_1315), .C(n_1317), .Y(n_1314) );
AOI21xp5_ASAP7_75t_SL g1343 ( .A1(n_345), .A2(n_732), .B(n_1344), .Y(n_1343) );
INVx1_ASAP7_75t_L g1357 ( .A(n_345), .Y(n_1357) );
INVx1_ASAP7_75t_L g875 ( .A(n_346), .Y(n_875) );
INVx1_ASAP7_75t_L g1405 ( .A(n_348), .Y(n_1405) );
INVx1_ASAP7_75t_L g1964 ( .A(n_350), .Y(n_1964) );
INVxp67_ASAP7_75t_L g1363 ( .A(n_352), .Y(n_1363) );
OAI211xp5_ASAP7_75t_L g969 ( .A1(n_353), .A2(n_527), .B(n_970), .C(n_972), .Y(n_969) );
INVx1_ASAP7_75t_L g980 ( .A(n_353), .Y(n_980) );
INVx1_ASAP7_75t_L g1916 ( .A(n_354), .Y(n_1916) );
INVxp67_ASAP7_75t_SL g1374 ( .A(n_355), .Y(n_1374) );
BUFx6f_ASAP7_75t_L g453 ( .A(n_356), .Y(n_453) );
AOI22xp33_ASAP7_75t_SL g1055 ( .A1(n_357), .A2(n_360), .B1(n_707), .B2(n_1056), .Y(n_1055) );
CKINVDCx5p33_ASAP7_75t_R g1223 ( .A(n_359), .Y(n_1223) );
INVx1_ASAP7_75t_L g1611 ( .A(n_361), .Y(n_1611) );
INVx1_ASAP7_75t_L g1630 ( .A(n_362), .Y(n_1630) );
INVx1_ASAP7_75t_L g669 ( .A(n_365), .Y(n_669) );
INVx1_ASAP7_75t_L g1454 ( .A(n_366), .Y(n_1454) );
INVx1_ASAP7_75t_L g1539 ( .A(n_367), .Y(n_1539) );
INVx1_ASAP7_75t_L g1162 ( .A(n_368), .Y(n_1162) );
OAI211xp5_ASAP7_75t_L g1169 ( .A1(n_368), .A2(n_653), .B(n_890), .C(n_1170), .Y(n_1169) );
INVx1_ASAP7_75t_L g391 ( .A(n_370), .Y(n_391) );
INVx2_ASAP7_75t_L g431 ( .A(n_370), .Y(n_431) );
INVx1_ASAP7_75t_L g589 ( .A(n_370), .Y(n_589) );
CKINVDCx5p33_ASAP7_75t_R g1226 ( .A(n_372), .Y(n_1226) );
CKINVDCx5p33_ASAP7_75t_R g1274 ( .A(n_373), .Y(n_1274) );
INVx1_ASAP7_75t_L g1025 ( .A(n_375), .Y(n_1025) );
AOI21xp5_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_1668), .B(n_1681), .Y(n_376) );
XNOR2xp5_ASAP7_75t_L g377 ( .A(n_378), .B(n_1175), .Y(n_377) );
OAI22xp5_ASAP7_75t_L g378 ( .A1(n_379), .A2(n_380), .B1(n_660), .B2(n_1174), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AOI22xp5_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_382), .B1(n_552), .B2(n_553), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
HB1xp67_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
NAND3xp33_ASAP7_75t_L g384 ( .A(n_385), .B(n_476), .C(n_516), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g385 ( .A(n_386), .B(n_440), .Y(n_385) );
OAI33xp33_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_395), .A3(n_412), .B1(n_424), .B2(n_429), .B3(n_435), .Y(n_386) );
OAI33xp33_ASAP7_75t_L g1456 ( .A1(n_387), .A2(n_429), .A3(n_1457), .B1(n_1458), .B2(n_1460), .B3(n_1462), .Y(n_1456) );
OAI33xp33_ASAP7_75t_L g1927 ( .A1(n_387), .A2(n_585), .A3(n_1928), .B1(n_1932), .B2(n_1933), .B3(n_1934), .Y(n_1927) );
BUFx2_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
BUFx4f_ASAP7_75t_L g558 ( .A(n_388), .Y(n_558) );
BUFx8_ASAP7_75t_L g915 ( .A(n_388), .Y(n_915) );
BUFx4f_ASAP7_75t_L g1124 ( .A(n_388), .Y(n_1124) );
OR2x2_ASAP7_75t_L g388 ( .A(n_389), .B(n_392), .Y(n_388) );
AND2x2_ASAP7_75t_SL g469 ( .A(n_389), .B(n_470), .Y(n_469) );
HB1xp67_ASAP7_75t_L g551 ( .A(n_389), .Y(n_551) );
INVx1_ASAP7_75t_L g611 ( .A(n_389), .Y(n_611) );
OR2x2_ASAP7_75t_L g762 ( .A(n_389), .B(n_763), .Y(n_762) );
INVx2_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
BUFx2_ASAP7_75t_L g515 ( .A(n_390), .Y(n_515) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
BUFx2_ASAP7_75t_L g1260 ( .A(n_392), .Y(n_1260) );
NAND2xp33_ASAP7_75t_SL g392 ( .A(n_393), .B(n_394), .Y(n_392) );
HB1xp67_ASAP7_75t_L g549 ( .A(n_393), .Y(n_549) );
AND3x4_ASAP7_75t_L g697 ( .A(n_393), .B(n_534), .C(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g756 ( .A(n_393), .Y(n_756) );
INVx3_ASAP7_75t_L g434 ( .A(n_394), .Y(n_434) );
BUFx3_ASAP7_75t_L g534 ( .A(n_394), .Y(n_534) );
OAI22xp33_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_397), .B1(n_404), .B2(n_405), .Y(n_395) );
OAI22xp33_ASAP7_75t_L g447 ( .A1(n_396), .A2(n_436), .B1(n_448), .B2(n_455), .Y(n_447) );
OAI22xp33_ASAP7_75t_L g871 ( .A1(n_397), .A2(n_872), .B1(n_873), .B2(n_875), .Y(n_871) );
BUFx4f_ASAP7_75t_SL g397 ( .A(n_398), .Y(n_397) );
OAI22xp33_ASAP7_75t_L g435 ( .A1(n_398), .A2(n_436), .B1(n_437), .B2(n_439), .Y(n_435) );
OAI22xp33_ASAP7_75t_L g1090 ( .A1(n_398), .A2(n_1074), .B1(n_1082), .B2(n_1091), .Y(n_1090) );
OAI22xp33_ASAP7_75t_L g1094 ( .A1(n_398), .A2(n_405), .B1(n_1075), .B2(n_1084), .Y(n_1094) );
OAI22xp33_ASAP7_75t_L g1457 ( .A1(n_398), .A2(n_971), .B1(n_1442), .B2(n_1451), .Y(n_1457) );
OAI22xp33_ASAP7_75t_L g1462 ( .A1(n_398), .A2(n_566), .B1(n_1444), .B2(n_1452), .Y(n_1462) );
INVx3_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx2_ASAP7_75t_SL g759 ( .A(n_399), .Y(n_759) );
INVx2_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
OR2x4_ASAP7_75t_L g518 ( .A(n_400), .B(n_434), .Y(n_518) );
OR2x4_ASAP7_75t_L g542 ( .A(n_400), .B(n_521), .Y(n_542) );
BUFx3_ASAP7_75t_L g563 ( .A(n_400), .Y(n_563) );
BUFx3_ASAP7_75t_L g858 ( .A(n_400), .Y(n_858) );
BUFx4f_ASAP7_75t_L g1128 ( .A(n_400), .Y(n_1128) );
OR2x2_ASAP7_75t_L g400 ( .A(n_401), .B(n_402), .Y(n_400) );
BUFx6f_ASAP7_75t_L g411 ( .A(n_401), .Y(n_411) );
INVx2_ASAP7_75t_L g418 ( .A(n_401), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_401), .B(n_410), .Y(n_423) );
AND2x4_ASAP7_75t_L g529 ( .A(n_401), .B(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g703 ( .A(n_402), .Y(n_703) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVxp67_ASAP7_75t_L g417 ( .A(n_403), .Y(n_417) );
OAI22xp5_ASAP7_75t_L g467 ( .A1(n_404), .A2(n_439), .B1(n_461), .B2(n_464), .Y(n_467) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVxp67_ASAP7_75t_L g624 ( .A(n_406), .Y(n_624) );
INVx1_ASAP7_75t_L g1931 ( .A(n_406), .Y(n_1931) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g1975 ( .A(n_407), .Y(n_1975) );
BUFx2_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
BUFx6f_ASAP7_75t_L g438 ( .A(n_408), .Y(n_438) );
BUFx3_ASAP7_75t_L g566 ( .A(n_408), .Y(n_566) );
NAND2x1p5_ASAP7_75t_L g408 ( .A(n_409), .B(n_411), .Y(n_408) );
BUFx2_ASAP7_75t_L g537 ( .A(n_409), .Y(n_537) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx2_ASAP7_75t_L g530 ( .A(n_410), .Y(n_530) );
BUFx2_ASAP7_75t_L g535 ( .A(n_411), .Y(n_535) );
AND2x4_ASAP7_75t_L g709 ( .A(n_411), .B(n_710), .Y(n_709) );
INVx2_ASAP7_75t_L g785 ( .A(n_411), .Y(n_785) );
OAI22xp5_ASAP7_75t_L g412 ( .A1(n_413), .A2(n_414), .B1(n_419), .B2(n_420), .Y(n_412) );
OAI22xp5_ASAP7_75t_L g460 ( .A1(n_413), .A2(n_425), .B1(n_461), .B2(n_464), .Y(n_460) );
OAI22xp5_ASAP7_75t_L g424 ( .A1(n_414), .A2(n_425), .B1(n_426), .B2(n_428), .Y(n_424) );
INVx2_ASAP7_75t_L g1054 ( .A(n_414), .Y(n_1054) );
OAI22xp5_ASAP7_75t_L g1458 ( .A1(n_414), .A2(n_1447), .B1(n_1454), .B2(n_1459), .Y(n_1458) );
OAI221xp5_ASAP7_75t_L g1642 ( .A1(n_414), .A2(n_420), .B1(n_1643), .B2(n_1644), .C(n_1645), .Y(n_1642) );
BUFx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g927 ( .A(n_415), .Y(n_927) );
INVx3_ASAP7_75t_L g1362 ( .A(n_415), .Y(n_1362) );
INVx2_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
BUFx6f_ASAP7_75t_L g522 ( .A(n_416), .Y(n_522) );
BUFx6f_ASAP7_75t_L g572 ( .A(n_416), .Y(n_572) );
BUFx8_ASAP7_75t_L g767 ( .A(n_416), .Y(n_767) );
AND2x4_ASAP7_75t_L g416 ( .A(n_417), .B(n_418), .Y(n_416) );
AND2x4_ASAP7_75t_L g702 ( .A(n_418), .B(n_703), .Y(n_702) );
OAI22xp5_ASAP7_75t_L g472 ( .A1(n_419), .A2(n_428), .B1(n_473), .B2(n_475), .Y(n_472) );
OAI22xp5_ASAP7_75t_L g1092 ( .A1(n_420), .A2(n_1079), .B1(n_1086), .B2(n_1093), .Y(n_1092) );
OAI22xp5_ASAP7_75t_L g1460 ( .A1(n_420), .A2(n_1448), .B1(n_1455), .B2(n_1461), .Y(n_1460) );
OAI22xp5_ASAP7_75t_L g1557 ( .A1(n_420), .A2(n_1539), .B1(n_1548), .B2(n_1558), .Y(n_1557) );
INVx3_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx3_ASAP7_75t_L g581 ( .A(n_421), .Y(n_581) );
CKINVDCx8_ASAP7_75t_R g865 ( .A(n_421), .Y(n_865) );
INVx1_ASAP7_75t_L g1459 ( .A(n_421), .Y(n_1459) );
INVx3_ASAP7_75t_L g1556 ( .A(n_421), .Y(n_1556) );
BUFx6f_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g427 ( .A(n_422), .Y(n_427) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
BUFx2_ASAP7_75t_L g546 ( .A(n_423), .Y(n_546) );
BUFx3_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
OR2x2_ASAP7_75t_L g794 ( .A(n_427), .B(n_762), .Y(n_794) );
INVx1_ASAP7_75t_L g778 ( .A(n_429), .Y(n_778) );
OAI33xp33_ASAP7_75t_L g1089 ( .A1(n_429), .A2(n_915), .A3(n_1090), .B1(n_1092), .B2(n_1094), .B3(n_1095), .Y(n_1089) );
OR2x6_ASAP7_75t_L g429 ( .A(n_430), .B(n_432), .Y(n_429) );
AND2x4_ASAP7_75t_L g444 ( .A(n_430), .B(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g1263 ( .A(n_430), .Y(n_1263) );
BUFx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g698 ( .A(n_431), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g1217 ( .A(n_431), .B(n_797), .Y(n_1217) );
INVx3_ASAP7_75t_L g1254 ( .A(n_432), .Y(n_1254) );
NAND2x1p5_ASAP7_75t_L g432 ( .A(n_433), .B(n_434), .Y(n_432) );
NAND3x1_ASAP7_75t_L g587 ( .A(n_433), .B(n_434), .C(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g521 ( .A(n_434), .Y(n_521) );
AND2x4_ASAP7_75t_L g528 ( .A(n_434), .B(n_529), .Y(n_528) );
OR2x6_ASAP7_75t_L g545 ( .A(n_434), .B(n_546), .Y(n_545) );
AND2x4_ASAP7_75t_L g755 ( .A(n_434), .B(n_756), .Y(n_755) );
HB1xp67_ASAP7_75t_L g860 ( .A(n_437), .Y(n_860) );
INVx1_ASAP7_75t_L g1138 ( .A(n_437), .Y(n_1138) );
OAI22xp33_ASAP7_75t_L g1934 ( .A1(n_437), .A2(n_1917), .B1(n_1923), .B2(n_1929), .Y(n_1934) );
BUFx6f_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx4_ASAP7_75t_L g526 ( .A(n_438), .Y(n_526) );
OR2x2_ASAP7_75t_L g801 ( .A(n_438), .B(n_762), .Y(n_801) );
INVx3_ASAP7_75t_L g874 ( .A(n_438), .Y(n_874) );
OAI33xp33_ASAP7_75t_L g440 ( .A1(n_441), .A2(n_447), .A3(n_460), .B1(n_467), .B2(n_468), .B3(n_472), .Y(n_440) );
OAI33xp33_ASAP7_75t_L g986 ( .A1(n_441), .A2(n_987), .A3(n_992), .B1(n_997), .B2(n_1002), .B3(n_1006), .Y(n_986) );
OAI33xp33_ASAP7_75t_L g1072 ( .A1(n_441), .A2(n_1006), .A3(n_1073), .B1(n_1078), .B2(n_1081), .B3(n_1085), .Y(n_1072) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx2_ASAP7_75t_SL g442 ( .A(n_443), .Y(n_442) );
INVx2_ASAP7_75t_SL g1046 ( .A(n_443), .Y(n_1046) );
INVx4_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g591 ( .A(n_444), .Y(n_591) );
INVx2_ASAP7_75t_L g722 ( .A(n_444), .Y(n_722) );
INVx2_ASAP7_75t_L g1145 ( .A(n_444), .Y(n_1145) );
INVx1_ASAP7_75t_L g1205 ( .A(n_444), .Y(n_1205) );
INVx2_ASAP7_75t_L g1445 ( .A(n_444), .Y(n_1445) );
AND2x4_ASAP7_75t_L g470 ( .A(n_446), .B(n_471), .Y(n_470) );
INVx2_ASAP7_75t_L g484 ( .A(n_446), .Y(n_484) );
BUFx2_ASAP7_75t_L g489 ( .A(n_446), .Y(n_489) );
AND2x4_ASAP7_75t_L g494 ( .A(n_446), .B(n_495), .Y(n_494) );
OAI221xp5_ASAP7_75t_L g1485 ( .A1(n_448), .A2(n_475), .B1(n_1486), .B2(n_1487), .C(n_1488), .Y(n_1485) );
OAI22xp5_ASAP7_75t_L g1924 ( .A1(n_448), .A2(n_1004), .B1(n_1925), .B2(n_1926), .Y(n_1924) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_SL g449 ( .A(n_450), .Y(n_449) );
OR2x6_ASAP7_75t_L g506 ( .A(n_450), .B(n_507), .Y(n_506) );
BUFx3_ASAP7_75t_L g989 ( .A(n_450), .Y(n_989) );
BUFx3_ASAP7_75t_L g1202 ( .A(n_450), .Y(n_1202) );
BUFx6f_ASAP7_75t_L g1443 ( .A(n_450), .Y(n_1443) );
INVx3_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx2_ASAP7_75t_L g474 ( .A(n_451), .Y(n_474) );
BUFx4f_ASAP7_75t_L g595 ( .A(n_451), .Y(n_595) );
INVx3_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
OR2x2_ASAP7_75t_L g452 ( .A(n_453), .B(n_454), .Y(n_452) );
INVx2_ASAP7_75t_L g459 ( .A(n_453), .Y(n_459) );
INVx2_ASAP7_75t_L g463 ( .A(n_453), .Y(n_463) );
NAND2x1_ASAP7_75t_L g466 ( .A(n_453), .B(n_454), .Y(n_466) );
AND2x2_ASAP7_75t_L g486 ( .A(n_453), .B(n_454), .Y(n_486) );
INVx1_ASAP7_75t_L g496 ( .A(n_453), .Y(n_496) );
AND2x2_ASAP7_75t_L g510 ( .A(n_453), .B(n_511), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_454), .B(n_459), .Y(n_458) );
OR2x2_ASAP7_75t_L g462 ( .A(n_454), .B(n_463), .Y(n_462) );
BUFx2_ASAP7_75t_L g490 ( .A(n_454), .Y(n_490) );
INVx2_ASAP7_75t_L g511 ( .A(n_454), .Y(n_511) );
INVx1_ASAP7_75t_L g673 ( .A(n_454), .Y(n_673) );
AND2x2_ASAP7_75t_L g729 ( .A(n_454), .B(n_459), .Y(n_729) );
OAI22xp5_ASAP7_75t_L g1317 ( .A1(n_455), .A2(n_1318), .B1(n_1319), .B2(n_1320), .Y(n_1317) );
OAI22xp33_ASAP7_75t_L g1441 ( .A1(n_455), .A2(n_1442), .B1(n_1443), .B2(n_1444), .Y(n_1441) );
INVx2_ASAP7_75t_L g1536 ( .A(n_455), .Y(n_1536) );
INVx4_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
BUFx6f_ASAP7_75t_L g597 ( .A(n_456), .Y(n_597) );
INVx1_ASAP7_75t_L g618 ( .A(n_456), .Y(n_618) );
INVx1_ASAP7_75t_L g936 ( .A(n_456), .Y(n_936) );
INVx2_ASAP7_75t_L g991 ( .A(n_456), .Y(n_991) );
INVx2_ASAP7_75t_L g1077 ( .A(n_456), .Y(n_1077) );
INVx2_ASAP7_75t_SL g1150 ( .A(n_456), .Y(n_1150) );
INVx2_ASAP7_75t_L g1410 ( .A(n_456), .Y(n_1410) );
INVx8_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
BUFx2_ASAP7_75t_L g475 ( .A(n_457), .Y(n_475) );
OR2x2_ASAP7_75t_L g504 ( .A(n_457), .B(n_489), .Y(n_504) );
BUFx6f_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
OAI22xp5_ASAP7_75t_SL g1446 ( .A1(n_461), .A2(n_1447), .B1(n_1448), .B2(n_1449), .Y(n_1446) );
BUFx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx2_ASAP7_75t_L g602 ( .A(n_462), .Y(n_602) );
BUFx3_ASAP7_75t_L g607 ( .A(n_462), .Y(n_607) );
BUFx2_ASAP7_75t_L g941 ( .A(n_462), .Y(n_941) );
INVx1_ASAP7_75t_L g1210 ( .A(n_462), .Y(n_1210) );
AND2x2_ASAP7_75t_L g672 ( .A(n_463), .B(n_673), .Y(n_672) );
HB1xp67_ASAP7_75t_L g1312 ( .A(n_463), .Y(n_1312) );
BUFx2_ASAP7_75t_L g890 ( .A(n_464), .Y(n_890) );
OAI211xp5_ASAP7_75t_L g1655 ( .A1(n_464), .A2(n_1656), .B(n_1657), .C(n_1658), .Y(n_1655) );
OAI211xp5_ASAP7_75t_SL g1659 ( .A1(n_464), .A2(n_1643), .B(n_1660), .C(n_1661), .Y(n_1659) );
BUFx3_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx2_ASAP7_75t_SL g604 ( .A(n_465), .Y(n_604) );
BUFx2_ASAP7_75t_SL g885 ( .A(n_465), .Y(n_885) );
OR2x2_ASAP7_75t_L g1193 ( .A(n_465), .B(n_1190), .Y(n_1193) );
NAND2xp5_ASAP7_75t_L g1309 ( .A(n_465), .B(n_1310), .Y(n_1309) );
NAND2xp5_ASAP7_75t_L g1412 ( .A(n_465), .B(n_1413), .Y(n_1412) );
BUFx3_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
BUFx6f_ASAP7_75t_L g480 ( .A(n_466), .Y(n_480) );
OAI33xp33_ASAP7_75t_L g1440 ( .A1(n_468), .A2(n_1441), .A3(n_1445), .B1(n_1446), .B2(n_1450), .B3(n_1453), .Y(n_1440) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
AND2x4_ASAP7_75t_L g609 ( .A(n_470), .B(n_610), .Y(n_609) );
INVx1_ASAP7_75t_SL g824 ( .A(n_470), .Y(n_824) );
OAI21xp33_ASAP7_75t_L g1315 ( .A1(n_470), .A2(n_607), .B(n_1316), .Y(n_1315) );
INVx4_ASAP7_75t_L g1339 ( .A(n_470), .Y(n_1339) );
OAI221xp5_ASAP7_75t_L g1417 ( .A1(n_470), .A2(n_480), .B1(n_607), .B2(n_1418), .C(n_1419), .Y(n_1417) );
NAND2xp5_ASAP7_75t_L g1545 ( .A(n_470), .B(n_610), .Y(n_1545) );
INVx1_ASAP7_75t_L g513 ( .A(n_471), .Y(n_513) );
AND2x4_ASAP7_75t_L g844 ( .A(n_471), .B(n_484), .Y(n_844) );
OAI22xp5_ASAP7_75t_L g1002 ( .A1(n_473), .A2(n_1003), .B1(n_1004), .B2(n_1005), .Y(n_1002) );
OAI22xp33_ASAP7_75t_L g1073 ( .A1(n_473), .A2(n_1074), .B1(n_1075), .B2(n_1076), .Y(n_1073) );
OAI22xp33_ASAP7_75t_L g1453 ( .A1(n_473), .A2(n_1004), .B1(n_1454), .B2(n_1455), .Y(n_1453) );
BUFx4f_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
OR2x6_ASAP7_75t_L g499 ( .A(n_474), .B(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g616 ( .A(n_474), .Y(n_616) );
OR2x6_ASAP7_75t_L g641 ( .A(n_474), .B(n_507), .Y(n_641) );
OAI31xp33_ASAP7_75t_L g476 ( .A1(n_477), .A2(n_498), .A3(n_505), .B(n_512), .Y(n_476) );
OAI211xp5_ASAP7_75t_SL g838 ( .A1(n_478), .A2(n_839), .B(n_840), .C(n_845), .Y(n_838) );
OAI22xp5_ASAP7_75t_L g1450 ( .A1(n_478), .A2(n_998), .B1(n_1451), .B2(n_1452), .Y(n_1450) );
INVx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g1156 ( .A(n_479), .Y(n_1156) );
INVx2_ASAP7_75t_L g1297 ( .A(n_479), .Y(n_1297) );
INVx1_ASAP7_75t_L g1449 ( .A(n_479), .Y(n_1449) );
INVx4_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
BUFx4f_ASAP7_75t_L g652 ( .A(n_480), .Y(n_652) );
BUFx4f_ASAP7_75t_L g1000 ( .A(n_480), .Y(n_1000) );
BUFx4f_ASAP7_75t_L g1111 ( .A(n_480), .Y(n_1111) );
BUFx4f_ASAP7_75t_L g1153 ( .A(n_480), .Y(n_1153) );
OR2x6_ASAP7_75t_L g1214 ( .A(n_480), .B(n_1215), .Y(n_1214) );
BUFx6f_ASAP7_75t_L g1353 ( .A(n_480), .Y(n_1353) );
NAND4xp25_ASAP7_75t_L g667 ( .A(n_481), .B(n_668), .C(n_675), .D(n_678), .Y(n_667) );
NAND3xp33_ASAP7_75t_L g1023 ( .A(n_481), .B(n_1024), .C(n_1028), .Y(n_1023) );
INVx3_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g653 ( .A(n_482), .Y(n_653) );
INVx1_ASAP7_75t_L g978 ( .A(n_482), .Y(n_978) );
AND2x2_ASAP7_75t_L g482 ( .A(n_483), .B(n_485), .Y(n_482) );
AND2x2_ASAP7_75t_L g1113 ( .A(n_483), .B(n_742), .Y(n_1113) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVxp67_ASAP7_75t_L g507 ( .A(n_484), .Y(n_507) );
BUFx3_ASAP7_75t_L g680 ( .A(n_485), .Y(n_680) );
BUFx3_ASAP7_75t_L g823 ( .A(n_485), .Y(n_823) );
AND2x6_ASAP7_75t_L g828 ( .A(n_485), .B(n_797), .Y(n_828) );
AND2x4_ASAP7_75t_SL g833 ( .A(n_485), .B(n_811), .Y(n_833) );
BUFx6f_ASAP7_75t_L g1199 ( .A(n_485), .Y(n_1199) );
INVx1_ASAP7_75t_L g1490 ( .A(n_485), .Y(n_1490) );
BUFx6f_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g738 ( .A(n_486), .Y(n_738) );
AOI22xp33_ASAP7_75t_L g487 ( .A1(n_488), .A2(n_491), .B1(n_492), .B2(n_497), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g891 ( .A1(n_488), .A2(n_657), .B1(n_892), .B2(n_893), .Y(n_891) );
AOI22xp33_ASAP7_75t_L g979 ( .A1(n_488), .A2(n_657), .B1(n_973), .B2(n_980), .Y(n_979) );
AOI222xp33_ASAP7_75t_L g1028 ( .A1(n_488), .A2(n_492), .B1(n_823), .B2(n_1029), .C1(n_1030), .C2(n_1031), .Y(n_1028) );
AOI22xp33_ASAP7_75t_L g1909 ( .A1(n_488), .A2(n_492), .B1(n_1904), .B2(n_1910), .Y(n_1909) );
AND2x2_ASAP7_75t_L g488 ( .A(n_489), .B(n_490), .Y(n_488) );
AND2x4_ASAP7_75t_L g656 ( .A(n_489), .B(n_490), .Y(n_656) );
AND2x2_ASAP7_75t_L g670 ( .A(n_489), .B(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g836 ( .A(n_490), .Y(n_836) );
INVx1_ASAP7_75t_L g1221 ( .A(n_490), .Y(n_1221) );
AOI22xp33_ASAP7_75t_L g1310 ( .A1(n_490), .A2(n_1269), .B1(n_1289), .B2(n_1311), .Y(n_1310) );
BUFx2_ASAP7_75t_L g1414 ( .A(n_490), .Y(n_1414) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_491), .A2(n_532), .B1(n_536), .B2(n_538), .Y(n_531) );
AOI222xp33_ASAP7_75t_L g678 ( .A1(n_492), .A2(n_656), .B1(n_679), .B2(n_680), .C1(n_681), .C2(n_682), .Y(n_678) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx2_ASAP7_75t_L g657 ( .A(n_493), .Y(n_657) );
INVx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g946 ( .A1(n_494), .A2(n_656), .B1(n_947), .B2(n_948), .Y(n_946) );
AOI22xp33_ASAP7_75t_L g1114 ( .A1(n_494), .A2(n_656), .B1(n_1103), .B2(n_1115), .Y(n_1114) );
BUFx3_ASAP7_75t_L g1171 ( .A(n_494), .Y(n_1171) );
AOI22xp33_ASAP7_75t_L g1428 ( .A1(n_494), .A2(n_656), .B1(n_1429), .B2(n_1430), .Y(n_1428) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_495), .B(n_797), .Y(n_803) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g645 ( .A(n_499), .Y(n_645) );
BUFx6f_ASAP7_75t_L g895 ( .A(n_499), .Y(n_895) );
BUFx2_ASAP7_75t_L g982 ( .A(n_499), .Y(n_982) );
AND2x4_ASAP7_75t_L g509 ( .A(n_500), .B(n_510), .Y(n_509) );
HB1xp67_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx2_ASAP7_75t_L g1026 ( .A(n_502), .Y(n_1026) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g668 ( .A1(n_503), .A2(n_669), .B1(n_670), .B2(n_674), .Y(n_668) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
BUFx2_ASAP7_75t_L g648 ( .A(n_504), .Y(n_648) );
INVx2_ASAP7_75t_L g897 ( .A(n_504), .Y(n_897) );
INVx1_ASAP7_75t_L g1109 ( .A(n_506), .Y(n_1109) );
INVx4_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx3_ASAP7_75t_SL g642 ( .A(n_509), .Y(n_642) );
AOI22xp33_ASAP7_75t_L g675 ( .A1(n_509), .A2(n_640), .B1(n_676), .B2(n_677), .Y(n_675) );
CKINVDCx16_ASAP7_75t_R g1167 ( .A(n_509), .Y(n_1167) );
BUFx6f_ASAP7_75t_L g733 ( .A(n_510), .Y(n_733) );
BUFx3_ASAP7_75t_L g822 ( .A(n_510), .Y(n_822) );
INVx2_ASAP7_75t_L g842 ( .A(n_510), .Y(n_842) );
BUFx2_ASAP7_75t_SL g659 ( .A(n_512), .Y(n_659) );
AOI22xp5_ASAP7_75t_L g666 ( .A1(n_512), .A2(n_667), .B1(n_683), .B2(n_684), .Y(n_666) );
BUFx3_ASAP7_75t_L g898 ( .A(n_512), .Y(n_898) );
BUFx2_ASAP7_75t_L g1033 ( .A(n_512), .Y(n_1033) );
INVx1_ASAP7_75t_L g1511 ( .A(n_512), .Y(n_1511) );
AND2x4_ASAP7_75t_L g512 ( .A(n_513), .B(n_514), .Y(n_512) );
INVx1_ASAP7_75t_L g1680 ( .A(n_513), .Y(n_1680) );
NOR2xp33_ASAP7_75t_L g1942 ( .A(n_513), .B(n_1672), .Y(n_1942) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
OR2x2_ASAP7_75t_L g802 ( .A(n_515), .B(n_803), .Y(n_802) );
INVxp67_ASAP7_75t_L g806 ( .A(n_515), .Y(n_806) );
INVx1_ASAP7_75t_L g1225 ( .A(n_515), .Y(n_1225) );
OAI31xp33_ASAP7_75t_L g516 ( .A1(n_517), .A2(n_523), .A3(n_539), .B(n_547), .Y(n_516) );
INVx2_ASAP7_75t_SL g634 ( .A(n_518), .Y(n_634) );
HB1xp67_ASAP7_75t_L g901 ( .A(n_518), .Y(n_901) );
INVx2_ASAP7_75t_SL g967 ( .A(n_518), .Y(n_967) );
INVx1_ASAP7_75t_L g1100 ( .A(n_518), .Y(n_1100) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g635 ( .A(n_520), .Y(n_635) );
AOI22xp33_ASAP7_75t_L g694 ( .A1(n_520), .A2(n_634), .B1(n_676), .B2(n_677), .Y(n_694) );
INVx1_ASAP7_75t_L g902 ( .A(n_520), .Y(n_902) );
INVx2_ASAP7_75t_L g968 ( .A(n_520), .Y(n_968) );
INVxp67_ASAP7_75t_L g1036 ( .A(n_520), .Y(n_1036) );
INVx1_ASAP7_75t_L g1164 ( .A(n_520), .Y(n_1164) );
AOI22xp33_ASAP7_75t_L g1626 ( .A1(n_520), .A2(n_544), .B1(n_1627), .B2(n_1628), .Y(n_1626) );
AND2x4_ASAP7_75t_L g520 ( .A(n_521), .B(n_522), .Y(n_520) );
BUFx6f_ASAP7_75t_L g706 ( .A(n_522), .Y(n_706) );
INVx1_ASAP7_75t_L g868 ( .A(n_522), .Y(n_868) );
BUFx6f_ASAP7_75t_L g1012 ( .A(n_522), .Y(n_1012) );
INVx2_ASAP7_75t_L g1096 ( .A(n_522), .Y(n_1096) );
HB1xp67_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
OAI221xp5_ASAP7_75t_L g1253 ( .A1(n_525), .A2(n_858), .B1(n_1203), .B2(n_1211), .C(n_1254), .Y(n_1253) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx2_ASAP7_75t_L g904 ( .A(n_526), .Y(n_904) );
INVx1_ASAP7_75t_L g1009 ( .A(n_526), .Y(n_1009) );
INVx1_ASAP7_75t_L g1091 ( .A(n_526), .Y(n_1091) );
INVx1_ASAP7_75t_L g1523 ( .A(n_526), .Y(n_1523) );
CKINVDCx8_ASAP7_75t_R g527 ( .A(n_528), .Y(n_527) );
CKINVDCx8_ASAP7_75t_R g625 ( .A(n_528), .Y(n_625) );
AOI211xp5_ASAP7_75t_L g685 ( .A1(n_528), .A2(n_682), .B(n_686), .C(n_688), .Y(n_685) );
OAI31xp33_ASAP7_75t_L g1366 ( .A1(n_528), .A2(n_1367), .A3(n_1376), .B(n_1378), .Y(n_1366) );
INVx2_ASAP7_75t_L g687 ( .A(n_529), .Y(n_687) );
BUFx2_ASAP7_75t_L g704 ( .A(n_529), .Y(n_704) );
BUFx2_ASAP7_75t_L g718 ( .A(n_529), .Y(n_718) );
BUFx2_ASAP7_75t_L g752 ( .A(n_529), .Y(n_752) );
BUFx3_ASAP7_75t_L g1238 ( .A(n_529), .Y(n_1238) );
BUFx2_ASAP7_75t_L g1248 ( .A(n_529), .Y(n_1248) );
BUFx2_ASAP7_75t_L g1633 ( .A(n_529), .Y(n_1633) );
INVx1_ASAP7_75t_L g710 ( .A(n_530), .Y(n_710) );
INVx1_ASAP7_75t_L g689 ( .A(n_532), .Y(n_689) );
AOI22xp33_ASAP7_75t_L g1102 ( .A1(n_532), .A2(n_536), .B1(n_1103), .B2(n_1104), .Y(n_1102) );
AOI22xp33_ASAP7_75t_L g1160 ( .A1(n_532), .A2(n_536), .B1(n_1161), .B2(n_1162), .Y(n_1160) );
AOI22xp5_ASAP7_75t_L g1373 ( .A1(n_532), .A2(n_536), .B1(n_1374), .B2(n_1375), .Y(n_1373) );
AOI22xp33_ASAP7_75t_L g1436 ( .A1(n_532), .A2(n_536), .B1(n_1429), .B2(n_1437), .Y(n_1436) );
AOI22xp33_ASAP7_75t_L g1903 ( .A1(n_532), .A2(n_536), .B1(n_1904), .B2(n_1905), .Y(n_1903) );
AND2x4_ASAP7_75t_L g532 ( .A(n_533), .B(n_535), .Y(n_532) );
AND2x4_ASAP7_75t_L g536 ( .A(n_533), .B(n_537), .Y(n_536) );
AND2x2_ASAP7_75t_L g628 ( .A(n_533), .B(n_535), .Y(n_628) );
A2O1A1Ixp33_ASAP7_75t_L g1367 ( .A1(n_533), .A2(n_1368), .B(n_1370), .C(n_1373), .Y(n_1367) );
INVx3_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
BUFx6f_ASAP7_75t_L g630 ( .A(n_536), .Y(n_630) );
INVx1_ASAP7_75t_L g690 ( .A(n_536), .Y(n_690) );
AOI22xp33_ASAP7_75t_SL g972 ( .A1(n_536), .A2(n_954), .B1(n_973), .B2(n_974), .Y(n_972) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g1634 ( .A1(n_541), .A2(n_634), .B1(n_1635), .B2(n_1636), .Y(n_1634) );
INVx2_ASAP7_75t_SL g541 ( .A(n_542), .Y(n_541) );
BUFx2_ASAP7_75t_L g621 ( .A(n_542), .Y(n_621) );
BUFx3_ASAP7_75t_L g693 ( .A(n_542), .Y(n_693) );
BUFx2_ASAP7_75t_L g1377 ( .A(n_542), .Y(n_1377) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_544), .A2(n_669), .B1(n_674), .B2(n_692), .Y(n_691) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
BUFx3_ASAP7_75t_L g622 ( .A(n_545), .Y(n_622) );
INVx1_ASAP7_75t_L g909 ( .A(n_545), .Y(n_909) );
INVx1_ASAP7_75t_L g958 ( .A(n_545), .Y(n_958) );
BUFx3_ASAP7_75t_L g574 ( .A(n_546), .Y(n_574) );
INVx1_ASAP7_75t_L g1015 ( .A(n_546), .Y(n_1015) );
OAI31xp33_ASAP7_75t_L g1097 ( .A1(n_547), .A2(n_1098), .A3(n_1101), .B(n_1105), .Y(n_1097) );
OAI31xp33_ASAP7_75t_L g1433 ( .A1(n_547), .A2(n_1434), .A3(n_1435), .B(n_1438), .Y(n_1433) );
AND2x2_ASAP7_75t_L g547 ( .A(n_548), .B(n_550), .Y(n_547) );
AND2x2_ASAP7_75t_L g636 ( .A(n_548), .B(n_550), .Y(n_636) );
AND2x4_ASAP7_75t_L g683 ( .A(n_548), .B(n_550), .Y(n_683) );
AND2x2_ASAP7_75t_SL g910 ( .A(n_548), .B(n_550), .Y(n_910) );
AND2x2_ASAP7_75t_L g1378 ( .A(n_548), .B(n_550), .Y(n_1378) );
INVx1_ASAP7_75t_SL g548 ( .A(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
HB1xp67_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
AND3x1_ASAP7_75t_L g555 ( .A(n_556), .B(n_619), .C(n_637), .Y(n_555) );
NOR2xp33_ASAP7_75t_L g556 ( .A(n_557), .B(n_590), .Y(n_556) );
OAI33xp33_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_559), .A3(n_567), .B1(n_575), .B2(n_582), .B3(n_585), .Y(n_557) );
OAI33xp33_ASAP7_75t_L g855 ( .A1(n_558), .A2(n_856), .A3(n_861), .B1(n_866), .B2(n_870), .B3(n_871), .Y(n_855) );
OAI33xp33_ASAP7_75t_L g1549 ( .A1(n_558), .A2(n_585), .A3(n_1550), .B1(n_1555), .B2(n_1557), .B3(n_1560), .Y(n_1549) );
OAI211xp5_ASAP7_75t_SL g1609 ( .A1(n_558), .A2(n_750), .B(n_1610), .C(n_1616), .Y(n_1609) );
OAI33xp33_ASAP7_75t_L g1952 ( .A1(n_558), .A2(n_585), .A3(n_1953), .B1(n_1956), .B2(n_1959), .B3(n_1963), .Y(n_1952) );
OAI22xp33_ASAP7_75t_L g559 ( .A1(n_560), .A2(n_561), .B1(n_564), .B2(n_565), .Y(n_559) );
OAI22xp33_ASAP7_75t_L g592 ( .A1(n_560), .A2(n_583), .B1(n_593), .B2(n_596), .Y(n_592) );
OAI22xp33_ASAP7_75t_L g582 ( .A1(n_561), .A2(n_565), .B1(n_583), .B2(n_584), .Y(n_582) );
OAI22xp33_ASAP7_75t_L g1008 ( .A1(n_561), .A2(n_988), .B1(n_999), .B2(n_1009), .Y(n_1008) );
OAI22xp33_ASAP7_75t_L g1019 ( .A1(n_561), .A2(n_904), .B1(n_990), .B2(n_1001), .Y(n_1019) );
OAI22xp33_ASAP7_75t_L g1953 ( .A1(n_561), .A2(n_565), .B1(n_1954), .B2(n_1955), .Y(n_1953) );
OAI22xp33_ASAP7_75t_L g1963 ( .A1(n_561), .A2(n_1553), .B1(n_1964), .B2(n_1965), .Y(n_1963) );
INVx2_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g1930 ( .A(n_563), .Y(n_1930) );
OAI22xp33_ASAP7_75t_L g605 ( .A1(n_564), .A2(n_584), .B1(n_603), .B2(n_606), .Y(n_605) );
OAI22xp33_ASAP7_75t_L g1125 ( .A1(n_565), .A2(n_1126), .B1(n_1127), .B2(n_1129), .Y(n_1125) );
OAI22xp33_ASAP7_75t_L g1560 ( .A1(n_565), .A2(n_1534), .B1(n_1542), .B2(n_1561), .Y(n_1560) );
BUFx6f_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
HB1xp67_ASAP7_75t_L g919 ( .A(n_566), .Y(n_919) );
HB1xp67_ASAP7_75t_L g932 ( .A(n_566), .Y(n_932) );
INVx2_ASAP7_75t_L g1554 ( .A(n_566), .Y(n_1554) );
OAI22xp5_ASAP7_75t_L g567 ( .A1(n_568), .A2(n_569), .B1(n_573), .B2(n_574), .Y(n_567) );
OAI22xp5_ASAP7_75t_L g598 ( .A1(n_568), .A2(n_576), .B1(n_599), .B2(n_603), .Y(n_598) );
OAI22xp5_ASAP7_75t_L g1956 ( .A1(n_569), .A2(n_574), .B1(n_1957), .B2(n_1958), .Y(n_1956) );
INVx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx8_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
BUFx3_ASAP7_75t_L g922 ( .A(n_571), .Y(n_922) );
OAI22xp5_ASAP7_75t_L g1016 ( .A1(n_571), .A2(n_996), .B1(n_1005), .B2(n_1013), .Y(n_1016) );
INVx5_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx3_ASAP7_75t_L g579 ( .A(n_572), .Y(n_579) );
INVx2_ASAP7_75t_SL g863 ( .A(n_572), .Y(n_863) );
INVx2_ASAP7_75t_SL g1280 ( .A(n_572), .Y(n_1280) );
AOI22xp33_ASAP7_75t_L g1370 ( .A1(n_572), .A2(n_715), .B1(n_1371), .B2(n_1372), .Y(n_1370) );
HB1xp67_ASAP7_75t_L g1559 ( .A(n_572), .Y(n_1559) );
OAI22xp5_ASAP7_75t_L g612 ( .A1(n_573), .A2(n_580), .B1(n_613), .B2(n_617), .Y(n_612) );
OAI22xp5_ASAP7_75t_L g924 ( .A1(n_574), .A2(n_925), .B1(n_926), .B2(n_928), .Y(n_924) );
OAI22xp5_ASAP7_75t_L g1933 ( .A1(n_574), .A2(n_1361), .B1(n_1920), .B2(n_1926), .Y(n_1933) );
OAI22xp5_ASAP7_75t_L g575 ( .A1(n_576), .A2(n_577), .B1(n_580), .B2(n_581), .Y(n_575) );
OAI22xp33_ASAP7_75t_SL g1130 ( .A1(n_577), .A2(n_1131), .B1(n_1132), .B2(n_1133), .Y(n_1130) );
INVx2_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g1242 ( .A1(n_578), .A2(n_1223), .B1(n_1226), .B2(n_1243), .Y(n_1242) );
INVx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
OAI22xp5_ASAP7_75t_L g866 ( .A1(n_581), .A2(n_867), .B1(n_868), .B2(n_869), .Y(n_866) );
OAI22xp5_ASAP7_75t_L g1140 ( .A1(n_581), .A2(n_1141), .B1(n_1142), .B2(n_1143), .Y(n_1140) );
OAI22xp5_ASAP7_75t_L g1959 ( .A1(n_581), .A2(n_1960), .B1(n_1961), .B2(n_1962), .Y(n_1959) );
OAI33xp33_ASAP7_75t_L g1122 ( .A1(n_585), .A2(n_1123), .A3(n_1125), .B1(n_1130), .B2(n_1134), .B3(n_1140), .Y(n_1122) );
OAI22xp5_ASAP7_75t_L g1637 ( .A1(n_585), .A2(n_1123), .B1(n_1638), .B2(n_1642), .Y(n_1637) );
INVx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
CKINVDCx5p33_ASAP7_75t_R g870 ( .A(n_586), .Y(n_870) );
NAND3xp33_ASAP7_75t_L g1057 ( .A(n_586), .B(n_1058), .C(n_1062), .Y(n_1057) );
INVx2_ASAP7_75t_L g1365 ( .A(n_586), .Y(n_1365) );
NAND3xp33_ASAP7_75t_L g1616 ( .A(n_586), .B(n_1617), .C(n_1618), .Y(n_1616) );
INVx3_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx3_ASAP7_75t_L g713 ( .A(n_587), .Y(n_713) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g754 ( .A(n_589), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g1190 ( .A(n_589), .B(n_811), .Y(n_1190) );
OAI33xp33_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_592), .A3(n_598), .B1(n_605), .B2(n_608), .B3(n_612), .Y(n_590) );
OAI33xp33_ASAP7_75t_L g1966 ( .A1(n_591), .A2(n_608), .A3(n_1967), .B1(n_1968), .B2(n_1969), .B3(n_1970), .Y(n_1966) );
OAI22xp5_ASAP7_75t_L g942 ( .A1(n_593), .A2(n_596), .B1(n_923), .B2(n_928), .Y(n_942) );
OAI22xp33_ASAP7_75t_L g1967 ( .A1(n_593), .A2(n_596), .B1(n_1954), .B2(n_1964), .Y(n_1967) );
INVx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx2_ASAP7_75t_L g935 ( .A(n_594), .Y(n_935) );
INVx3_ASAP7_75t_L g1087 ( .A(n_594), .Y(n_1087) );
INVx2_ASAP7_75t_SL g1147 ( .A(n_594), .Y(n_1147) );
BUFx6f_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx3_ASAP7_75t_L g880 ( .A(n_595), .Y(n_880) );
INVx4_ASAP7_75t_L g1319 ( .A(n_595), .Y(n_1319) );
OAI22xp5_ASAP7_75t_L g877 ( .A1(n_596), .A2(n_857), .B1(n_872), .B2(n_878), .Y(n_877) );
OAI22xp5_ASAP7_75t_L g886 ( .A1(n_596), .A2(n_864), .B1(n_869), .B2(n_880), .Y(n_886) );
INVx6_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx5_ASAP7_75t_L g1004 ( .A(n_597), .Y(n_1004) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
OAI221xp5_ASAP7_75t_L g1404 ( .A1(n_601), .A2(n_844), .B1(n_1297), .B2(n_1405), .C(n_1406), .Y(n_1404) );
OAI22xp5_ASAP7_75t_L g1537 ( .A1(n_601), .A2(n_1111), .B1(n_1538), .B2(n_1539), .Y(n_1537) );
OAI22xp5_ASAP7_75t_L g1540 ( .A1(n_601), .A2(n_603), .B1(n_1541), .B2(n_1542), .Y(n_1540) );
INVx2_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
BUFx2_ASAP7_75t_L g883 ( .A(n_602), .Y(n_883) );
INVx2_ASAP7_75t_L g1300 ( .A(n_602), .Y(n_1300) );
OAI22xp5_ASAP7_75t_L g881 ( .A1(n_603), .A2(n_862), .B1(n_867), .B2(n_882), .Y(n_881) );
OAI22xp5_ASAP7_75t_L g937 ( .A1(n_603), .A2(n_882), .B1(n_921), .B2(n_925), .Y(n_937) );
OAI22xp5_ASAP7_75t_L g1078 ( .A1(n_603), .A2(n_998), .B1(n_1079), .B2(n_1080), .Y(n_1078) );
OAI211xp5_ASAP7_75t_L g1600 ( .A1(n_603), .A2(n_1601), .B(n_1602), .C(n_1603), .Y(n_1600) );
OAI22xp5_ASAP7_75t_L g1918 ( .A1(n_603), .A2(n_1209), .B1(n_1919), .B2(n_1920), .Y(n_1918) );
OAI22xp5_ASAP7_75t_L g1969 ( .A1(n_603), .A2(n_1152), .B1(n_1955), .B2(n_1965), .Y(n_1969) );
INVx5_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
HB1xp67_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx2_ASAP7_75t_L g995 ( .A(n_607), .Y(n_995) );
OAI22xp5_ASAP7_75t_L g1968 ( .A1(n_607), .A2(n_1153), .B1(n_1957), .B2(n_1960), .Y(n_1968) );
OAI33xp33_ASAP7_75t_L g876 ( .A1(n_608), .A2(n_721), .A3(n_877), .B1(n_881), .B2(n_884), .B3(n_886), .Y(n_876) );
OAI33xp33_ASAP7_75t_L g933 ( .A1(n_608), .A2(n_721), .A3(n_934), .B1(n_937), .B2(n_938), .B3(n_942), .Y(n_933) );
OAI33xp33_ASAP7_75t_L g1144 ( .A1(n_608), .A2(n_1145), .A3(n_1146), .B1(n_1151), .B2(n_1154), .B3(n_1155), .Y(n_1144) );
INVx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
AOI33xp33_ASAP7_75t_L g719 ( .A1(n_609), .A2(n_720), .A3(n_723), .B1(n_730), .B2(n_739), .B3(n_743), .Y(n_719) );
CKINVDCx5p33_ASAP7_75t_R g1006 ( .A(n_609), .Y(n_1006) );
NAND3xp33_ASAP7_75t_L g1047 ( .A(n_609), .B(n_1048), .C(n_1051), .Y(n_1047) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
OAI22xp33_ASAP7_75t_L g1155 ( .A1(n_613), .A2(n_1132), .B1(n_1139), .B2(n_1156), .Y(n_1155) );
OAI22xp33_ASAP7_75t_L g1970 ( .A1(n_613), .A2(n_1004), .B1(n_1958), .B2(n_1962), .Y(n_1970) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
BUFx3_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
OAI31xp33_ASAP7_75t_L g619 ( .A1(n_620), .A2(n_623), .A3(n_632), .B(n_636), .Y(n_619) );
NAND4xp25_ASAP7_75t_L g1625 ( .A(n_625), .B(n_1626), .C(n_1629), .D(n_1634), .Y(n_1625) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_627), .A2(n_629), .B1(n_630), .B2(n_631), .Y(n_626) );
AOI22xp33_ASAP7_75t_L g905 ( .A1(n_627), .A2(n_630), .B1(n_892), .B2(n_906), .Y(n_905) );
AOI22xp33_ASAP7_75t_L g1038 ( .A1(n_627), .A2(n_630), .B1(n_1030), .B2(n_1031), .Y(n_1038) );
AOI22xp33_ASAP7_75t_L g1524 ( .A1(n_627), .A2(n_630), .B1(n_1518), .B2(n_1525), .Y(n_1524) );
AOI22xp33_ASAP7_75t_L g1976 ( .A1(n_627), .A2(n_630), .B1(n_1977), .B2(n_1978), .Y(n_1976) );
BUFx3_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
BUFx3_ASAP7_75t_L g954 ( .A(n_628), .Y(n_954) );
AOI22xp33_ASAP7_75t_L g654 ( .A1(n_629), .A2(n_655), .B1(n_657), .B2(n_658), .Y(n_654) );
AOI22xp33_ASAP7_75t_L g953 ( .A1(n_630), .A2(n_947), .B1(n_954), .B2(n_955), .Y(n_953) );
AOI222xp33_ASAP7_75t_L g1629 ( .A1(n_630), .A2(n_954), .B1(n_1630), .B2(n_1631), .C1(n_1632), .C2(n_1633), .Y(n_1629) );
INVx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
OAI31xp33_ASAP7_75t_SL g637 ( .A1(n_638), .A2(n_643), .A3(n_649), .B(n_659), .Y(n_637) );
INVxp67_ASAP7_75t_SL g639 ( .A(n_640), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g1679 ( .A(n_640), .B(n_1680), .Y(n_1679) );
AND2x4_ASAP7_75t_SL g1941 ( .A(n_640), .B(n_1942), .Y(n_1941) );
INVx3_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx2_ASAP7_75t_SL g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
OAI22xp5_ASAP7_75t_L g992 ( .A1(n_652), .A2(n_993), .B1(n_994), .B2(n_996), .Y(n_992) );
OAI22xp5_ASAP7_75t_L g1081 ( .A1(n_652), .A2(n_1082), .B1(n_1083), .B2(n_1084), .Y(n_1081) );
OAI22xp5_ASAP7_75t_L g1921 ( .A1(n_652), .A2(n_1209), .B1(n_1922), .B2(n_1923), .Y(n_1921) );
AOI22xp33_ASAP7_75t_L g1170 ( .A1(n_655), .A2(n_1161), .B1(n_1171), .B2(n_1172), .Y(n_1170) );
AOI22xp33_ASAP7_75t_L g1517 ( .A1(n_655), .A2(n_1171), .B1(n_1518), .B2(n_1519), .Y(n_1517) );
AOI22xp33_ASAP7_75t_L g1985 ( .A1(n_655), .A2(n_657), .B1(n_1977), .B2(n_1986), .Y(n_1985) );
BUFx3_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
OAI31xp33_ASAP7_75t_L g943 ( .A1(n_659), .A2(n_944), .A3(n_945), .B(n_949), .Y(n_943) );
OAI31xp33_ASAP7_75t_L g976 ( .A1(n_659), .A2(n_977), .A3(n_981), .B(n_984), .Y(n_976) );
OAI31xp33_ASAP7_75t_L g1165 ( .A1(n_659), .A2(n_1166), .A3(n_1168), .B(n_1169), .Y(n_1165) );
OAI31xp33_ASAP7_75t_L g1426 ( .A1(n_659), .A2(n_1427), .A3(n_1431), .B(n_1432), .Y(n_1426) );
OAI31xp33_ASAP7_75t_L g1907 ( .A1(n_659), .A2(n_1908), .A3(n_1911), .B(n_1912), .Y(n_1907) );
OAI31xp33_ASAP7_75t_L g1981 ( .A1(n_659), .A2(n_1982), .A3(n_1983), .B(n_1984), .Y(n_1981) );
INVx1_ASAP7_75t_L g1174 ( .A(n_660), .Y(n_1174) );
XNOR2xp5_ASAP7_75t_L g660 ( .A(n_661), .B(n_960), .Y(n_660) );
AOI22xp33_ASAP7_75t_SL g661 ( .A1(n_662), .A2(n_663), .B1(n_851), .B2(n_959), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
XNOR2x1_ASAP7_75t_L g663 ( .A(n_664), .B(n_746), .Y(n_663) );
NAND3x1_ASAP7_75t_L g665 ( .A(n_666), .B(n_695), .C(n_719), .Y(n_665) );
AOI22xp5_ASAP7_75t_L g1024 ( .A1(n_670), .A2(n_1025), .B1(n_1026), .B2(n_1027), .Y(n_1024) );
BUFx6f_ASAP7_75t_L g826 ( .A(n_671), .Y(n_826) );
INVx3_ASAP7_75t_L g1295 ( .A(n_671), .Y(n_1295) );
A2O1A1Ixp33_ASAP7_75t_L g1308 ( .A1(n_671), .A2(n_1274), .B(n_1309), .C(n_1313), .Y(n_1308) );
A2O1A1Ixp33_ASAP7_75t_L g1411 ( .A1(n_671), .A2(n_1390), .B(n_1412), .C(n_1415), .Y(n_1411) );
BUFx6f_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx3_ASAP7_75t_L g725 ( .A(n_672), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_672), .B(n_797), .Y(n_796) );
AND2x2_ASAP7_75t_L g815 ( .A(n_672), .B(n_811), .Y(n_815) );
OAI31xp33_ASAP7_75t_L g964 ( .A1(n_683), .A2(n_965), .A3(n_969), .B(n_975), .Y(n_964) );
OAI31xp33_ASAP7_75t_L g1034 ( .A1(n_683), .A2(n_1035), .A3(n_1037), .B(n_1039), .Y(n_1034) );
CKINVDCx14_ASAP7_75t_R g1527 ( .A(n_683), .Y(n_1527) );
AOI211xp5_ASAP7_75t_L g1624 ( .A1(n_683), .A2(n_1625), .B(n_1637), .C(n_1648), .Y(n_1624) );
OAI31xp33_ASAP7_75t_L g1900 ( .A1(n_683), .A2(n_1901), .A3(n_1902), .B(n_1906), .Y(n_1900) );
OAI31xp33_ASAP7_75t_L g1971 ( .A1(n_683), .A2(n_1972), .A3(n_1979), .B(n_1980), .Y(n_1971) );
NAND3xp33_ASAP7_75t_L g684 ( .A(n_685), .B(n_691), .C(n_694), .Y(n_684) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx2_ASAP7_75t_L g1063 ( .A(n_687), .Y(n_1063) );
INVx1_ASAP7_75t_L g1283 ( .A(n_687), .Y(n_1283) );
INVx2_ASAP7_75t_L g1619 ( .A(n_687), .Y(n_1619) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
AOI33xp33_ASAP7_75t_L g695 ( .A1(n_696), .A2(n_699), .A3(n_705), .B1(n_711), .B2(n_712), .B3(n_714), .Y(n_695) );
NAND3xp33_ASAP7_75t_L g1052 ( .A(n_696), .B(n_1053), .C(n_1055), .Y(n_1052) );
BUFx3_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
AOI33xp33_ASAP7_75t_L g769 ( .A1(n_697), .A2(n_770), .A3(n_774), .B1(n_776), .B2(n_778), .B3(n_779), .Y(n_769) );
AOI33xp33_ASAP7_75t_L g1275 ( .A1(n_697), .A2(n_778), .A3(n_1276), .B1(n_1277), .B2(n_1278), .B3(n_1282), .Y(n_1275) );
NAND3xp33_ASAP7_75t_L g1382 ( .A(n_697), .B(n_1383), .C(n_1384), .Y(n_1382) );
AOI33xp33_ASAP7_75t_L g1497 ( .A1(n_697), .A2(n_778), .A3(n_1498), .B1(n_1501), .B2(n_1502), .B3(n_1503), .Y(n_1497) );
INVx1_ASAP7_75t_L g850 ( .A(n_698), .Y(n_850) );
BUFx2_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g1615 ( .A(n_701), .Y(n_1615) );
BUFx3_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx8_ASAP7_75t_L g716 ( .A(n_702), .Y(n_716) );
BUFx3_ASAP7_75t_L g773 ( .A(n_702), .Y(n_773) );
NAND2x1p5_ASAP7_75t_L g805 ( .A(n_702), .B(n_755), .Y(n_805) );
HB1xp67_ASAP7_75t_L g1243 ( .A(n_702), .Y(n_1243) );
INVx1_ASAP7_75t_L g1093 ( .A(n_706), .Y(n_1093) );
INVx2_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx2_ASAP7_75t_R g775 ( .A(n_708), .Y(n_775) );
INVx1_ASAP7_75t_L g1061 ( .A(n_708), .Y(n_1061) );
INVx5_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
BUFx12f_ASAP7_75t_L g777 ( .A(n_709), .Y(n_777) );
BUFx3_ASAP7_75t_L g1246 ( .A(n_709), .Y(n_1246) );
BUFx3_ASAP7_75t_L g1281 ( .A(n_709), .Y(n_1281) );
INVx1_ASAP7_75t_L g790 ( .A(n_710), .Y(n_790) );
BUFx2_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
BUFx2_ASAP7_75t_L g1018 ( .A(n_713), .Y(n_1018) );
INVx8_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx3_ASAP7_75t_L g780 ( .A(n_716), .Y(n_780) );
CKINVDCx5p33_ASAP7_75t_R g1237 ( .A(n_716), .Y(n_1237) );
INVx2_ASAP7_75t_L g1271 ( .A(n_716), .Y(n_1271) );
HB1xp67_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
BUFx6f_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx2_ASAP7_75t_L g1213 ( .A(n_725), .Y(n_1213) );
INVx2_ASAP7_75t_L g1593 ( .A(n_725), .Y(n_1593) );
INVx2_ASAP7_75t_SL g1596 ( .A(n_725), .Y(n_1596) );
INVx1_ASAP7_75t_L g1604 ( .A(n_725), .Y(n_1604) );
INVx1_ASAP7_75t_SL g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_SL g727 ( .A(n_728), .Y(n_727) );
BUFx3_ASAP7_75t_L g1044 ( .A(n_728), .Y(n_1044) );
BUFx3_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
BUFx6f_ASAP7_75t_L g745 ( .A(n_729), .Y(n_745) );
BUFx3_ASAP7_75t_L g846 ( .A(n_729), .Y(n_846) );
INVx2_ASAP7_75t_L g1192 ( .A(n_729), .Y(n_1192) );
BUFx3_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
BUFx6f_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
AND2x4_ASAP7_75t_L g818 ( .A(n_733), .B(n_811), .Y(n_818) );
AND2x2_ASAP7_75t_L g1228 ( .A(n_733), .B(n_811), .Y(n_1228) );
INVx2_ASAP7_75t_L g1306 ( .A(n_733), .Y(n_1306) );
INVx1_ASAP7_75t_L g1590 ( .A(n_733), .Y(n_1590) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
AOI221xp5_ASAP7_75t_L g1597 ( .A1(n_736), .A2(n_1311), .B1(n_1351), .B2(n_1585), .C(n_1598), .Y(n_1597) );
INVx2_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
BUFx2_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g742 ( .A(n_738), .Y(n_742) );
INVx2_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
BUFx2_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
AND2x4_ASAP7_75t_L g810 ( .A(n_745), .B(n_811), .Y(n_810) );
HB1xp67_ASAP7_75t_L g827 ( .A(n_745), .Y(n_827) );
INVx1_ASAP7_75t_L g1403 ( .A(n_745), .Y(n_1403) );
AND3x1_ASAP7_75t_L g747 ( .A(n_748), .B(n_791), .C(n_807), .Y(n_747) );
NOR3xp33_ASAP7_75t_L g748 ( .A(n_749), .B(n_757), .C(n_768), .Y(n_748) );
NOR3xp33_ASAP7_75t_L g1495 ( .A(n_749), .B(n_1496), .C(n_1507), .Y(n_1495) );
INVx2_ASAP7_75t_SL g749 ( .A(n_750), .Y(n_749) );
INVx3_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
AOI221xp5_ASAP7_75t_L g1287 ( .A1(n_751), .A2(n_1288), .B1(n_1289), .B2(n_1290), .C(n_1291), .Y(n_1287) );
AOI221xp5_ASAP7_75t_L g1395 ( .A1(n_751), .A2(n_1288), .B1(n_1290), .B2(n_1396), .C(n_1397), .Y(n_1395) );
AND2x4_ASAP7_75t_L g751 ( .A(n_752), .B(n_753), .Y(n_751) );
AND2x2_ASAP7_75t_L g783 ( .A(n_753), .B(n_784), .Y(n_783) );
AND2x4_ASAP7_75t_L g787 ( .A(n_753), .B(n_788), .Y(n_787) );
AND2x4_ASAP7_75t_SL g1288 ( .A(n_753), .B(n_784), .Y(n_1288) );
AND2x4_ASAP7_75t_SL g1290 ( .A(n_753), .B(n_788), .Y(n_1290) );
AND2x4_ASAP7_75t_L g753 ( .A(n_754), .B(n_755), .Y(n_753) );
OR2x2_ASAP7_75t_L g795 ( .A(n_754), .B(n_796), .Y(n_795) );
AND2x6_ASAP7_75t_L g1232 ( .A(n_755), .B(n_784), .Y(n_1232) );
AND2x2_ASAP7_75t_L g1234 ( .A(n_755), .B(n_790), .Y(n_1234) );
INVx1_ASAP7_75t_L g1240 ( .A(n_755), .Y(n_1240) );
NAND2xp5_ASAP7_75t_L g1572 ( .A(n_758), .B(n_1573), .Y(n_1572) );
OR2x6_ASAP7_75t_L g758 ( .A(n_759), .B(n_760), .Y(n_758) );
OR2x2_ASAP7_75t_L g1508 ( .A(n_759), .B(n_760), .Y(n_1508) );
INVx2_ASAP7_75t_SL g1562 ( .A(n_759), .Y(n_1562) );
INVxp67_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
AND2x2_ASAP7_75t_L g1577 ( .A(n_761), .B(n_1362), .Y(n_1577) );
INVx1_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVx1_ASAP7_75t_L g766 ( .A(n_762), .Y(n_766) );
INVx1_ASAP7_75t_L g1251 ( .A(n_763), .Y(n_1251) );
INVx2_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g1284 ( .A(n_765), .B(n_1285), .Y(n_1284) );
NAND2xp5_ASAP7_75t_L g1385 ( .A(n_765), .B(n_1386), .Y(n_1385) );
AND2x4_ASAP7_75t_L g765 ( .A(n_766), .B(n_767), .Y(n_765) );
AND2x4_ASAP7_75t_L g1270 ( .A(n_766), .B(n_1271), .Y(n_1270) );
INVx3_ASAP7_75t_L g1060 ( .A(n_767), .Y(n_1060) );
INVx2_ASAP7_75t_SL g1461 ( .A(n_767), .Y(n_1461) );
INVx3_ASAP7_75t_L g1961 ( .A(n_767), .Y(n_1961) );
NAND2xp5_ASAP7_75t_SL g768 ( .A(n_769), .B(n_781), .Y(n_768) );
INVx1_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
BUFx3_ASAP7_75t_L g1056 ( .A(n_773), .Y(n_1056) );
INVx2_ASAP7_75t_SL g1500 ( .A(n_773), .Y(n_1500) );
AOI22xp33_ASAP7_75t_L g1368 ( .A1(n_777), .A2(n_1238), .B1(n_1348), .B2(n_1369), .Y(n_1368) );
NAND3xp33_ASAP7_75t_L g1391 ( .A(n_778), .B(n_1392), .C(n_1393), .Y(n_1391) );
AOI22xp33_ASAP7_75t_L g781 ( .A1(n_782), .A2(n_783), .B1(n_786), .B2(n_787), .Y(n_781) );
AOI22xp33_ASAP7_75t_L g1504 ( .A1(n_783), .A2(n_787), .B1(n_1505), .B2(n_1506), .Y(n_1504) );
INVx3_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
INVx2_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
AOI21xp33_ASAP7_75t_L g791 ( .A1(n_792), .A2(n_798), .B(n_799), .Y(n_791) );
AOI21xp33_ASAP7_75t_SL g1491 ( .A1(n_792), .A2(n_1492), .B(n_1493), .Y(n_1491) );
INVx8_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
AND2x4_ASAP7_75t_L g793 ( .A(n_794), .B(n_795), .Y(n_793) );
INVx1_ASAP7_75t_L g1273 ( .A(n_794), .Y(n_1273) );
INVx1_ASAP7_75t_L g1186 ( .A(n_795), .Y(n_1186) );
INVx1_ASAP7_75t_L g837 ( .A(n_797), .Y(n_837) );
HB1xp67_ASAP7_75t_L g1313 ( .A(n_797), .Y(n_1313) );
AND2x4_ASAP7_75t_L g800 ( .A(n_801), .B(n_802), .Y(n_800) );
INVx2_ASAP7_75t_L g1268 ( .A(n_801), .Y(n_1268) );
AND2x4_ASAP7_75t_L g1494 ( .A(n_801), .B(n_802), .Y(n_1494) );
INVx1_ASAP7_75t_L g1665 ( .A(n_803), .Y(n_1665) );
OR2x2_ASAP7_75t_L g804 ( .A(n_805), .B(n_806), .Y(n_804) );
OR2x6_ASAP7_75t_L g1324 ( .A(n_805), .B(n_806), .Y(n_1324) );
OAI21xp5_ASAP7_75t_SL g807 ( .A1(n_808), .A2(n_829), .B(n_847), .Y(n_807) );
INVx3_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
INVx2_ASAP7_75t_SL g1472 ( .A(n_810), .Y(n_1472) );
BUFx2_ASAP7_75t_L g1303 ( .A(n_811), .Y(n_1303) );
AND2x2_ASAP7_75t_L g1606 ( .A(n_811), .B(n_1191), .Y(n_1606) );
AOI22xp33_ASAP7_75t_L g812 ( .A1(n_813), .A2(n_814), .B1(n_816), .B2(n_817), .Y(n_812) );
AOI22xp33_ASAP7_75t_L g1477 ( .A1(n_814), .A2(n_1478), .B1(n_1479), .B2(n_1480), .Y(n_1477) );
INVx1_ASAP7_75t_L g1651 ( .A(n_814), .Y(n_1651) );
BUFx6f_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
AND2x4_ASAP7_75t_L g1224 ( .A(n_815), .B(n_1225), .Y(n_1224) );
BUFx6f_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
HB1xp67_ASAP7_75t_L g1480 ( .A(n_818), .Y(n_1480) );
INVx1_ASAP7_75t_L g1654 ( .A(n_818), .Y(n_1654) );
AOI21xp5_ASAP7_75t_L g819 ( .A1(n_820), .A2(n_825), .B(n_828), .Y(n_819) );
HB1xp67_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
BUFx2_ASAP7_75t_L g1043 ( .A(n_822), .Y(n_1043) );
A2O1A1Ixp33_ASAP7_75t_SL g1347 ( .A1(n_826), .A2(n_1313), .B(n_1348), .C(n_1349), .Y(n_1347) );
AOI21xp5_ASAP7_75t_SL g1473 ( .A1(n_828), .A2(n_1474), .B(n_1476), .Y(n_1473) );
AOI211xp5_ASAP7_75t_SL g1662 ( .A1(n_828), .A2(n_1608), .B(n_1631), .C(n_1663), .Y(n_1662) );
INVx2_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
INVx1_ASAP7_75t_L g1482 ( .A(n_831), .Y(n_1482) );
INVx4_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
INVx2_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
BUFx3_ASAP7_75t_L g1608 ( .A(n_833), .Y(n_1608) );
INVx2_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
INVx2_ASAP7_75t_L g1484 ( .A(n_835), .Y(n_1484) );
NOR2x1_ASAP7_75t_L g835 ( .A(n_836), .B(n_837), .Y(n_835) );
INVx1_ASAP7_75t_L g1351 ( .A(n_836), .Y(n_1351) );
INVx1_ASAP7_75t_L g1415 ( .A(n_837), .Y(n_1415) );
INVx2_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
INVx2_ASAP7_75t_L g1050 ( .A(n_842), .Y(n_1050) );
INVx3_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
OAI221xp5_ASAP7_75t_L g1296 ( .A1(n_844), .A2(n_1297), .B1(n_1298), .B2(n_1299), .C(n_1300), .Y(n_1296) );
INVx1_ASAP7_75t_L g1344 ( .A(n_844), .Y(n_1344) );
INVx2_ASAP7_75t_L g1591 ( .A(n_844), .Y(n_1591) );
OAI21xp33_ASAP7_75t_L g1470 ( .A1(n_847), .A2(n_1471), .B(n_1481), .Y(n_1470) );
INVx1_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
AOI21xp33_ASAP7_75t_L g1648 ( .A1(n_848), .A2(n_1649), .B(n_1662), .Y(n_1648) );
INVx1_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
BUFx2_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
OAI31xp33_ASAP7_75t_L g1292 ( .A1(n_850), .A2(n_1293), .A3(n_1301), .B(n_1314), .Y(n_1292) );
HB1xp67_ASAP7_75t_L g1331 ( .A(n_850), .Y(n_1331) );
OAI31xp33_ASAP7_75t_L g1400 ( .A1(n_850), .A2(n_1401), .A3(n_1407), .B(n_1416), .Y(n_1400) );
INVx1_ASAP7_75t_L g959 ( .A(n_851), .Y(n_959) );
XOR2x2_ASAP7_75t_L g851 ( .A(n_852), .B(n_911), .Y(n_851) );
AND3x1_ASAP7_75t_L g853 ( .A(n_854), .B(n_887), .C(n_899), .Y(n_853) );
NOR2xp33_ASAP7_75t_L g854 ( .A(n_855), .B(n_876), .Y(n_854) );
OAI22xp33_ASAP7_75t_L g856 ( .A1(n_857), .A2(n_858), .B1(n_859), .B2(n_860), .Y(n_856) );
OAI22xp33_ASAP7_75t_L g916 ( .A1(n_858), .A2(n_917), .B1(n_918), .B2(n_919), .Y(n_916) );
OAI22xp33_ASAP7_75t_L g929 ( .A1(n_858), .A2(n_930), .B1(n_931), .B2(n_932), .Y(n_929) );
OAI22xp5_ASAP7_75t_L g884 ( .A1(n_859), .A2(n_875), .B1(n_882), .B2(n_885), .Y(n_884) );
OAI22xp5_ASAP7_75t_L g861 ( .A1(n_862), .A2(n_863), .B1(n_864), .B2(n_865), .Y(n_861) );
OAI22xp5_ASAP7_75t_L g920 ( .A1(n_865), .A2(n_921), .B1(n_922), .B2(n_923), .Y(n_920) );
OAI22xp5_ASAP7_75t_L g1095 ( .A1(n_865), .A2(n_1080), .B1(n_1088), .B2(n_1096), .Y(n_1095) );
OAI22xp5_ASAP7_75t_L g1255 ( .A1(n_865), .A2(n_1011), .B1(n_1256), .B2(n_1257), .Y(n_1255) );
OAI221xp5_ASAP7_75t_L g1355 ( .A1(n_865), .A2(n_1356), .B1(n_1357), .B2(n_1358), .C(n_1359), .Y(n_1355) );
OAI221xp5_ASAP7_75t_L g1360 ( .A1(n_865), .A2(n_1342), .B1(n_1361), .B2(n_1363), .C(n_1364), .Y(n_1360) );
OAI221xp5_ASAP7_75t_L g1638 ( .A1(n_865), .A2(n_1135), .B1(n_1639), .B2(n_1640), .C(n_1641), .Y(n_1638) );
OAI22xp33_ASAP7_75t_L g1932 ( .A1(n_865), .A2(n_1356), .B1(n_1919), .B2(n_1925), .Y(n_1932) );
OAI33xp33_ASAP7_75t_L g914 ( .A1(n_870), .A2(n_915), .A3(n_916), .B1(n_920), .B2(n_924), .B3(n_929), .Y(n_914) );
INVx2_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
INVx2_ASAP7_75t_L g971 ( .A(n_874), .Y(n_971) );
INVx2_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
INVx2_ASAP7_75t_SL g879 ( .A(n_880), .Y(n_879) );
INVx4_ASAP7_75t_L g882 ( .A(n_883), .Y(n_882) );
OAI22xp5_ASAP7_75t_L g938 ( .A1(n_885), .A2(n_918), .B1(n_931), .B2(n_939), .Y(n_938) );
OAI31xp33_ASAP7_75t_L g887 ( .A1(n_888), .A2(n_889), .A3(n_894), .B(n_898), .Y(n_887) );
INVx2_ASAP7_75t_L g896 ( .A(n_897), .Y(n_896) );
INVx1_ASAP7_75t_L g983 ( .A(n_897), .Y(n_983) );
INVx1_ASAP7_75t_L g1117 ( .A(n_897), .Y(n_1117) );
OAI31xp33_ASAP7_75t_L g899 ( .A1(n_900), .A2(n_903), .A3(n_907), .B(n_910), .Y(n_899) );
INVx1_ASAP7_75t_L g908 ( .A(n_909), .Y(n_908) );
OAI31xp33_ASAP7_75t_L g950 ( .A1(n_910), .A2(n_951), .A3(n_952), .B(n_956), .Y(n_950) );
OAI31xp33_ASAP7_75t_SL g1157 ( .A1(n_910), .A2(n_1158), .A3(n_1159), .B(n_1163), .Y(n_1157) );
AND3x1_ASAP7_75t_L g912 ( .A(n_913), .B(n_943), .C(n_950), .Y(n_912) );
NOR2xp33_ASAP7_75t_L g913 ( .A(n_914), .B(n_933), .Y(n_913) );
OAI33xp33_ASAP7_75t_L g1007 ( .A1(n_915), .A2(n_1008), .A3(n_1010), .B1(n_1016), .B2(n_1017), .B3(n_1019), .Y(n_1007) );
OAI22xp33_ASAP7_75t_L g934 ( .A1(n_917), .A2(n_930), .B1(n_935), .B2(n_936), .Y(n_934) );
INVx1_ASAP7_75t_L g926 ( .A(n_927), .Y(n_926) );
INVx1_ASAP7_75t_L g1135 ( .A(n_927), .Y(n_1135) );
INVx2_ASAP7_75t_L g939 ( .A(n_940), .Y(n_939) );
INVx4_ASAP7_75t_L g998 ( .A(n_940), .Y(n_998) );
INVx2_ASAP7_75t_L g1083 ( .A(n_940), .Y(n_1083) );
INVx2_ASAP7_75t_L g1152 ( .A(n_940), .Y(n_1152) );
INVx4_ASAP7_75t_L g940 ( .A(n_941), .Y(n_940) );
INVx1_ASAP7_75t_L g957 ( .A(n_958), .Y(n_957) );
XOR2xp5_ASAP7_75t_L g960 ( .A(n_961), .B(n_1068), .Y(n_960) );
OAI22xp5_ASAP7_75t_L g961 ( .A1(n_962), .A2(n_1020), .B1(n_1066), .B2(n_1067), .Y(n_961) );
INVx1_ASAP7_75t_L g1066 ( .A(n_962), .Y(n_1066) );
NAND3xp33_ASAP7_75t_L g963 ( .A(n_964), .B(n_976), .C(n_985), .Y(n_963) );
INVx2_ASAP7_75t_SL g966 ( .A(n_967), .Y(n_966) );
HB1xp67_ASAP7_75t_L g970 ( .A(n_971), .Y(n_970) );
OAI211xp5_ASAP7_75t_L g1258 ( .A1(n_971), .A2(n_1208), .B(n_1259), .C(n_1261), .Y(n_1258) );
NOR2xp33_ASAP7_75t_L g985 ( .A(n_986), .B(n_1007), .Y(n_985) );
OAI22xp33_ASAP7_75t_L g987 ( .A1(n_988), .A2(n_989), .B1(n_990), .B2(n_991), .Y(n_987) );
OAI22xp5_ASAP7_75t_L g1085 ( .A1(n_991), .A2(n_1086), .B1(n_1087), .B2(n_1088), .Y(n_1085) );
OAI22xp5_ASAP7_75t_L g1010 ( .A1(n_993), .A2(n_1003), .B1(n_1011), .B2(n_1013), .Y(n_1010) );
OAI22xp5_ASAP7_75t_L g1154 ( .A1(n_994), .A2(n_1129), .B1(n_1143), .B2(n_1148), .Y(n_1154) );
INVx3_ASAP7_75t_L g994 ( .A(n_995), .Y(n_994) );
OAI22xp5_ASAP7_75t_L g997 ( .A1(n_998), .A2(n_999), .B1(n_1000), .B2(n_1001), .Y(n_997) );
OAI221xp5_ASAP7_75t_L g1207 ( .A1(n_1000), .A2(n_1208), .B1(n_1209), .B2(n_1211), .C(n_1212), .Y(n_1207) );
OAI211xp5_ASAP7_75t_SL g1336 ( .A1(n_1000), .A2(n_1337), .B(n_1338), .C(n_1340), .Y(n_1336) );
OAI211xp5_ASAP7_75t_SL g1341 ( .A1(n_1000), .A2(n_1342), .B(n_1343), .C(n_1345), .Y(n_1341) );
OAI22xp33_ASAP7_75t_L g1915 ( .A1(n_1004), .A2(n_1087), .B1(n_1916), .B2(n_1917), .Y(n_1915) );
OAI21xp5_ASAP7_75t_L g1206 ( .A1(n_1006), .A2(n_1207), .B(n_1214), .Y(n_1206) );
OAI33xp33_ASAP7_75t_L g1914 ( .A1(n_1006), .A2(n_1445), .A3(n_1915), .B1(n_1918), .B2(n_1921), .B3(n_1924), .Y(n_1914) );
INVx2_ASAP7_75t_L g1011 ( .A(n_1012), .Y(n_1011) );
INVx2_ASAP7_75t_SL g1356 ( .A(n_1012), .Y(n_1356) );
OAI221xp5_ASAP7_75t_L g1610 ( .A1(n_1013), .A2(n_1096), .B1(n_1611), .B2(n_1612), .C(n_1613), .Y(n_1610) );
INVx3_ASAP7_75t_L g1013 ( .A(n_1014), .Y(n_1013) );
BUFx2_ASAP7_75t_L g1014 ( .A(n_1015), .Y(n_1014) );
INVx1_ASAP7_75t_L g1133 ( .A(n_1015), .Y(n_1133) );
INVx1_ASAP7_75t_L g1017 ( .A(n_1018), .Y(n_1017) );
INVx2_ASAP7_75t_L g1067 ( .A(n_1020), .Y(n_1067) );
INVx1_ASAP7_75t_L g1064 ( .A(n_1021), .Y(n_1064) );
NAND3xp33_ASAP7_75t_L g1021 ( .A(n_1022), .B(n_1034), .C(n_1040), .Y(n_1021) );
OAI21xp5_ASAP7_75t_L g1022 ( .A1(n_1023), .A2(n_1032), .B(n_1033), .Y(n_1022) );
INVx2_ASAP7_75t_L g1514 ( .A(n_1026), .Y(n_1514) );
OAI31xp33_ASAP7_75t_SL g1106 ( .A1(n_1033), .A2(n_1107), .A3(n_1110), .B(n_1116), .Y(n_1106) );
AND4x1_ASAP7_75t_L g1040 ( .A(n_1041), .B(n_1047), .C(n_1052), .D(n_1057), .Y(n_1040) );
NAND3xp33_ASAP7_75t_L g1041 ( .A(n_1042), .B(n_1045), .C(n_1046), .Y(n_1041) );
HB1xp67_ASAP7_75t_L g1049 ( .A(n_1050), .Y(n_1049) );
INVx2_ASAP7_75t_L g1197 ( .A(n_1050), .Y(n_1197) );
INVx1_ASAP7_75t_L g1059 ( .A(n_1060), .Y(n_1059) );
OAI22xp5_ASAP7_75t_L g1068 ( .A1(n_1069), .A2(n_1118), .B1(n_1119), .B2(n_1173), .Y(n_1068) );
INVx2_ASAP7_75t_SL g1173 ( .A(n_1069), .Y(n_1173) );
NAND3xp33_ASAP7_75t_L g1070 ( .A(n_1071), .B(n_1097), .C(n_1106), .Y(n_1070) );
NOR2xp33_ASAP7_75t_L g1071 ( .A(n_1072), .B(n_1089), .Y(n_1071) );
OAI22xp5_ASAP7_75t_L g1200 ( .A1(n_1076), .A2(n_1201), .B1(n_1202), .B2(n_1203), .Y(n_1200) );
BUFx6f_ASAP7_75t_L g1076 ( .A(n_1077), .Y(n_1076) );
INVx1_ASAP7_75t_L g1099 ( .A(n_1100), .Y(n_1099) );
INVx1_ASAP7_75t_L g1108 ( .A(n_1109), .Y(n_1108) );
INVx2_ASAP7_75t_L g1112 ( .A(n_1113), .Y(n_1112) );
INVx2_ASAP7_75t_SL g1118 ( .A(n_1119), .Y(n_1118) );
NAND3xp33_ASAP7_75t_L g1120 ( .A(n_1121), .B(n_1157), .C(n_1165), .Y(n_1120) );
NOR2xp33_ASAP7_75t_SL g1121 ( .A(n_1122), .B(n_1144), .Y(n_1121) );
OAI22xp33_ASAP7_75t_L g1354 ( .A1(n_1123), .A2(n_1355), .B1(n_1360), .B2(n_1365), .Y(n_1354) );
BUFx3_ASAP7_75t_L g1123 ( .A(n_1124), .Y(n_1123) );
OAI22xp5_ASAP7_75t_L g1146 ( .A1(n_1126), .A2(n_1142), .B1(n_1147), .B2(n_1148), .Y(n_1146) );
HB1xp67_ASAP7_75t_L g1127 ( .A(n_1128), .Y(n_1127) );
HB1xp67_ASAP7_75t_L g1141 ( .A(n_1128), .Y(n_1141) );
INVx1_ASAP7_75t_L g1552 ( .A(n_1128), .Y(n_1552) );
OAI22xp5_ASAP7_75t_L g1151 ( .A1(n_1131), .A2(n_1136), .B1(n_1152), .B2(n_1153), .Y(n_1151) );
OAI22xp5_ASAP7_75t_L g1134 ( .A1(n_1135), .A2(n_1136), .B1(n_1137), .B2(n_1139), .Y(n_1134) );
OAI22xp5_ASAP7_75t_L g1555 ( .A1(n_1135), .A2(n_1538), .B1(n_1547), .B2(n_1556), .Y(n_1555) );
INVx2_ASAP7_75t_SL g1137 ( .A(n_1138), .Y(n_1137) );
INVx1_ASAP7_75t_L g1148 ( .A(n_1149), .Y(n_1148) );
INVx1_ASAP7_75t_L g1149 ( .A(n_1150), .Y(n_1149) );
OAI22xp5_ASAP7_75t_SL g1175 ( .A1(n_1176), .A2(n_1464), .B1(n_1465), .B2(n_1667), .Y(n_1175) );
AOI22xp33_ASAP7_75t_L g1176 ( .A1(n_1177), .A2(n_1422), .B1(n_1423), .B2(n_1463), .Y(n_1176) );
INVx3_ASAP7_75t_SL g1463 ( .A(n_1177), .Y(n_1463) );
AOI22xp33_ASAP7_75t_L g1667 ( .A1(n_1177), .A2(n_1422), .B1(n_1423), .B2(n_1463), .Y(n_1667) );
BUFx3_ASAP7_75t_L g1177 ( .A(n_1178), .Y(n_1177) );
OA22x2_ASAP7_75t_L g1178 ( .A1(n_1179), .A2(n_1180), .B1(n_1326), .B2(n_1421), .Y(n_1178) );
INVx1_ASAP7_75t_L g1179 ( .A(n_1180), .Y(n_1179) );
XOR2xp5_ASAP7_75t_L g1180 ( .A(n_1181), .B(n_1264), .Y(n_1180) );
XNOR2x1_ASAP7_75t_L g1181 ( .A(n_1182), .B(n_1183), .Y(n_1181) );
NAND4xp75_ASAP7_75t_L g1183 ( .A(n_1184), .B(n_1194), .C(n_1222), .D(n_1229), .Y(n_1183) );
INVx1_ASAP7_75t_L g1185 ( .A(n_1186), .Y(n_1185) );
INVx1_ASAP7_75t_L g1187 ( .A(n_1188), .Y(n_1187) );
AND2x4_ASAP7_75t_L g1188 ( .A(n_1189), .B(n_1191), .Y(n_1188) );
INVx1_ASAP7_75t_L g1189 ( .A(n_1190), .Y(n_1189) );
INVx3_ASAP7_75t_L g1191 ( .A(n_1192), .Y(n_1191) );
INVx1_ASAP7_75t_L g1346 ( .A(n_1192), .Y(n_1346) );
AOI211x1_ASAP7_75t_L g1194 ( .A1(n_1195), .A2(n_1204), .B(n_1206), .C(n_1218), .Y(n_1194) );
INVx2_ASAP7_75t_L g1196 ( .A(n_1197), .Y(n_1196) );
INVx2_ASAP7_75t_L g1475 ( .A(n_1197), .Y(n_1475) );
BUFx2_ASAP7_75t_L g1198 ( .A(n_1199), .Y(n_1198) );
AOI221xp5_ASAP7_75t_L g1304 ( .A1(n_1199), .A2(n_1285), .B1(n_1291), .B2(n_1305), .C(n_1307), .Y(n_1304) );
AOI221xp5_ASAP7_75t_L g1408 ( .A1(n_1199), .A2(n_1305), .B1(n_1386), .B2(n_1397), .C(n_1409), .Y(n_1408) );
INVx1_ASAP7_75t_L g1533 ( .A(n_1202), .Y(n_1533) );
INVx1_ASAP7_75t_L g1204 ( .A(n_1205), .Y(n_1204) );
INVx2_ASAP7_75t_L g1209 ( .A(n_1210), .Y(n_1209) );
INVx1_ASAP7_75t_L g1215 ( .A(n_1216), .Y(n_1215) );
NAND2x2_ASAP7_75t_L g1219 ( .A(n_1216), .B(n_1220), .Y(n_1219) );
INVx2_ASAP7_75t_L g1216 ( .A(n_1217), .Y(n_1216) );
INVx2_ASAP7_75t_SL g1220 ( .A(n_1221), .Y(n_1220) );
AOI22xp5_ASAP7_75t_L g1222 ( .A1(n_1223), .A2(n_1224), .B1(n_1226), .B2(n_1227), .Y(n_1222) );
INVx3_ASAP7_75t_L g1573 ( .A(n_1224), .Y(n_1573) );
AND2x4_ASAP7_75t_L g1227 ( .A(n_1225), .B(n_1228), .Y(n_1227) );
INVx2_ASAP7_75t_L g1578 ( .A(n_1227), .Y(n_1578) );
OAI31xp67_ASAP7_75t_L g1229 ( .A1(n_1230), .A2(n_1241), .A3(n_1252), .B(n_1262), .Y(n_1229) );
INVx4_ASAP7_75t_L g1231 ( .A(n_1232), .Y(n_1231) );
INVx2_ASAP7_75t_L g1233 ( .A(n_1234), .Y(n_1233) );
A2O1A1Ixp33_ASAP7_75t_L g1235 ( .A1(n_1236), .A2(n_1237), .B(n_1238), .C(n_1239), .Y(n_1235) );
INVx1_ASAP7_75t_L g1239 ( .A(n_1240), .Y(n_1239) );
AOI21xp33_ASAP7_75t_L g1241 ( .A1(n_1242), .A2(n_1244), .B(n_1249), .Y(n_1241) );
AOI22xp33_ASAP7_75t_L g1244 ( .A1(n_1245), .A2(n_1246), .B1(n_1247), .B2(n_1248), .Y(n_1244) );
INVx1_ASAP7_75t_L g1249 ( .A(n_1250), .Y(n_1249) );
HB1xp67_ASAP7_75t_L g1250 ( .A(n_1251), .Y(n_1250) );
OAI21xp5_ASAP7_75t_SL g1252 ( .A1(n_1253), .A2(n_1255), .B(n_1258), .Y(n_1252) );
AOI31xp33_ASAP7_75t_L g1586 ( .A1(n_1262), .A2(n_1587), .A3(n_1600), .B(n_1605), .Y(n_1586) );
BUFx2_ASAP7_75t_L g1262 ( .A(n_1263), .Y(n_1262) );
XNOR2x1_ASAP7_75t_L g1264 ( .A(n_1265), .B(n_1325), .Y(n_1264) );
OR2x2_ASAP7_75t_L g1265 ( .A(n_1266), .B(n_1286), .Y(n_1265) );
NAND3xp33_ASAP7_75t_L g1266 ( .A(n_1267), .B(n_1275), .C(n_1284), .Y(n_1266) );
AOI222xp33_ASAP7_75t_L g1267 ( .A1(n_1268), .A2(n_1269), .B1(n_1270), .B2(n_1272), .C1(n_1273), .C2(n_1274), .Y(n_1267) );
AOI222xp33_ASAP7_75t_L g1387 ( .A1(n_1268), .A2(n_1270), .B1(n_1273), .B2(n_1388), .C1(n_1389), .C2(n_1390), .Y(n_1387) );
AOI22xp5_ASAP7_75t_L g1583 ( .A1(n_1268), .A2(n_1273), .B1(n_1584), .B2(n_1585), .Y(n_1583) );
INVx2_ASAP7_75t_L g1279 ( .A(n_1280), .Y(n_1279) );
NAND3xp33_ASAP7_75t_SL g1286 ( .A(n_1287), .B(n_1292), .C(n_1321), .Y(n_1286) );
INVx1_ASAP7_75t_L g1581 ( .A(n_1288), .Y(n_1581) );
INVx1_ASAP7_75t_L g1582 ( .A(n_1290), .Y(n_1582) );
INVx1_ASAP7_75t_L g1294 ( .A(n_1295), .Y(n_1294) );
OAI21xp33_ASAP7_75t_L g1301 ( .A1(n_1302), .A2(n_1304), .B(n_1308), .Y(n_1301) );
OAI21xp5_ASAP7_75t_SL g1407 ( .A1(n_1302), .A2(n_1408), .B(n_1411), .Y(n_1407) );
INVxp67_ASAP7_75t_L g1302 ( .A(n_1303), .Y(n_1302) );
OAI21xp5_ASAP7_75t_L g1333 ( .A1(n_1303), .A2(n_1334), .B(n_1335), .Y(n_1333) );
INVx2_ASAP7_75t_L g1305 ( .A(n_1306), .Y(n_1305) );
INVx1_ASAP7_75t_L g1352 ( .A(n_1311), .Y(n_1352) );
AOI22xp5_ASAP7_75t_L g1413 ( .A1(n_1311), .A2(n_1388), .B1(n_1396), .B2(n_1414), .Y(n_1413) );
INVx1_ASAP7_75t_L g1311 ( .A(n_1312), .Y(n_1311) );
INVx1_ASAP7_75t_L g1599 ( .A(n_1313), .Y(n_1599) );
NAND2xp5_ASAP7_75t_L g1321 ( .A(n_1322), .B(n_1323), .Y(n_1321) );
NAND2xp5_ASAP7_75t_L g1398 ( .A(n_1323), .B(n_1399), .Y(n_1398) );
INVx5_ASAP7_75t_L g1323 ( .A(n_1324), .Y(n_1323) );
INVx3_ASAP7_75t_L g1569 ( .A(n_1324), .Y(n_1569) );
XNOR2xp5_ASAP7_75t_L g1326 ( .A(n_1327), .B(n_1379), .Y(n_1326) );
XOR2xp5_ASAP7_75t_L g1421 ( .A(n_1327), .B(n_1379), .Y(n_1421) );
XNOR2x1_ASAP7_75t_L g1327 ( .A(n_1328), .B(n_1329), .Y(n_1327) );
AND2x2_ASAP7_75t_L g1329 ( .A(n_1330), .B(n_1366), .Y(n_1329) );
AOI21xp5_ASAP7_75t_L g1330 ( .A1(n_1331), .A2(n_1332), .B(n_1354), .Y(n_1330) );
NAND4xp25_ASAP7_75t_L g1332 ( .A(n_1333), .B(n_1336), .C(n_1341), .D(n_1347), .Y(n_1332) );
INVx1_ASAP7_75t_L g1350 ( .A(n_1351), .Y(n_1350) );
INVx2_ASAP7_75t_L g1361 ( .A(n_1362), .Y(n_1361) );
XNOR2x1_ASAP7_75t_L g1379 ( .A(n_1380), .B(n_1420), .Y(n_1379) );
OR2x2_ASAP7_75t_L g1380 ( .A(n_1381), .B(n_1394), .Y(n_1380) );
NAND4xp25_ASAP7_75t_SL g1381 ( .A(n_1382), .B(n_1385), .C(n_1387), .D(n_1391), .Y(n_1381) );
NAND3xp33_ASAP7_75t_SL g1394 ( .A(n_1395), .B(n_1398), .C(n_1400), .Y(n_1394) );
INVx1_ASAP7_75t_L g1402 ( .A(n_1403), .Y(n_1402) );
INVx1_ASAP7_75t_L g1422 ( .A(n_1423), .Y(n_1422) );
INVx1_ASAP7_75t_L g1423 ( .A(n_1424), .Y(n_1423) );
NAND3xp33_ASAP7_75t_L g1425 ( .A(n_1426), .B(n_1433), .C(n_1439), .Y(n_1425) );
NOR2xp33_ASAP7_75t_SL g1439 ( .A(n_1440), .B(n_1456), .Y(n_1439) );
OAI33xp33_ASAP7_75t_L g1529 ( .A1(n_1445), .A2(n_1530), .A3(n_1537), .B1(n_1540), .B2(n_1543), .B3(n_1546), .Y(n_1529) );
INVx2_ASAP7_75t_SL g1464 ( .A(n_1465), .Y(n_1464) );
AO22x1_ASAP7_75t_L g1465 ( .A1(n_1466), .A2(n_1467), .B1(n_1563), .B2(n_1564), .Y(n_1465) );
INVx1_ASAP7_75t_L g1466 ( .A(n_1467), .Y(n_1466) );
XNOR2xp5_ASAP7_75t_L g1467 ( .A(n_1468), .B(n_1509), .Y(n_1467) );
NAND3xp33_ASAP7_75t_L g1469 ( .A(n_1470), .B(n_1491), .C(n_1495), .Y(n_1469) );
BUFx2_ASAP7_75t_L g1483 ( .A(n_1484), .Y(n_1483) );
INVx1_ASAP7_75t_L g1489 ( .A(n_1490), .Y(n_1489) );
NAND2xp5_ASAP7_75t_SL g1496 ( .A(n_1497), .B(n_1504), .Y(n_1496) );
INVx2_ASAP7_75t_L g1499 ( .A(n_1500), .Y(n_1499) );
OAI221xp5_ASAP7_75t_L g1510 ( .A1(n_1511), .A2(n_1512), .B1(n_1520), .B2(n_1527), .C(n_1528), .Y(n_1510) );
NOR3xp33_ASAP7_75t_L g1512 ( .A(n_1513), .B(n_1515), .C(n_1516), .Y(n_1512) );
NOR3xp33_ASAP7_75t_L g1520 ( .A(n_1521), .B(n_1522), .C(n_1526), .Y(n_1520) );
NOR2xp33_ASAP7_75t_L g1528 ( .A(n_1529), .B(n_1549), .Y(n_1528) );
OAI22xp5_ASAP7_75t_L g1530 ( .A1(n_1531), .A2(n_1532), .B1(n_1534), .B2(n_1535), .Y(n_1530) );
OAI22xp33_ASAP7_75t_L g1550 ( .A1(n_1531), .A2(n_1541), .B1(n_1551), .B2(n_1553), .Y(n_1550) );
OAI22xp5_ASAP7_75t_L g1546 ( .A1(n_1532), .A2(n_1535), .B1(n_1547), .B2(n_1548), .Y(n_1546) );
INVx2_ASAP7_75t_L g1532 ( .A(n_1533), .Y(n_1532) );
INVx2_ASAP7_75t_L g1535 ( .A(n_1536), .Y(n_1535) );
INVx2_ASAP7_75t_L g1543 ( .A(n_1544), .Y(n_1543) );
INVx1_ASAP7_75t_L g1544 ( .A(n_1545), .Y(n_1544) );
INVx2_ASAP7_75t_L g1551 ( .A(n_1552), .Y(n_1551) );
INVx2_ASAP7_75t_L g1553 ( .A(n_1554), .Y(n_1553) );
INVx1_ASAP7_75t_L g1558 ( .A(n_1559), .Y(n_1558) );
INVx1_ASAP7_75t_L g1561 ( .A(n_1562), .Y(n_1561) );
INVx2_ASAP7_75t_L g1563 ( .A(n_1564), .Y(n_1563) );
XOR2x2_ASAP7_75t_L g1564 ( .A(n_1565), .B(n_1622), .Y(n_1564) );
INVx1_ASAP7_75t_L g1620 ( .A(n_1566), .Y(n_1620) );
NAND3xp33_ASAP7_75t_L g1566 ( .A(n_1567), .B(n_1570), .C(n_1579), .Y(n_1566) );
NAND2xp5_ASAP7_75t_L g1567 ( .A(n_1568), .B(n_1569), .Y(n_1567) );
AOI22xp33_ASAP7_75t_L g1605 ( .A1(n_1568), .A2(n_1606), .B1(n_1607), .B2(n_1608), .Y(n_1605) );
AOI22xp33_ASAP7_75t_L g1570 ( .A1(n_1571), .A2(n_1572), .B1(n_1574), .B2(n_1575), .Y(n_1570) );
NAND2x1_ASAP7_75t_L g1575 ( .A(n_1576), .B(n_1578), .Y(n_1575) );
INVx2_ASAP7_75t_SL g1576 ( .A(n_1577), .Y(n_1576) );
NOR3xp33_ASAP7_75t_SL g1579 ( .A(n_1580), .B(n_1586), .C(n_1609), .Y(n_1579) );
NAND2xp5_ASAP7_75t_L g1595 ( .A(n_1584), .B(n_1596), .Y(n_1595) );
AOI21xp5_ASAP7_75t_L g1587 ( .A1(n_1588), .A2(n_1592), .B(n_1594), .Y(n_1587) );
INVx2_ASAP7_75t_SL g1589 ( .A(n_1590), .Y(n_1589) );
AOI21xp5_ASAP7_75t_L g1594 ( .A1(n_1595), .A2(n_1597), .B(n_1599), .Y(n_1594) );
INVx2_ASAP7_75t_L g1652 ( .A(n_1606), .Y(n_1652) );
INVx1_ASAP7_75t_L g1614 ( .A(n_1615), .Y(n_1614) );
INVx1_ASAP7_75t_L g1623 ( .A(n_1624), .Y(n_1623) );
NAND2xp5_ASAP7_75t_L g1664 ( .A(n_1632), .B(n_1665), .Y(n_1664) );
INVx1_ASAP7_75t_L g1647 ( .A(n_1633), .Y(n_1647) );
INVx1_ASAP7_75t_L g1646 ( .A(n_1647), .Y(n_1646) );
NOR2xp33_ASAP7_75t_L g1649 ( .A(n_1650), .B(n_1653), .Y(n_1649) );
BUFx2_ASAP7_75t_L g1668 ( .A(n_1669), .Y(n_1668) );
BUFx4f_ASAP7_75t_L g1669 ( .A(n_1670), .Y(n_1669) );
INVx3_ASAP7_75t_L g1670 ( .A(n_1671), .Y(n_1670) );
OR2x2_ASAP7_75t_L g1671 ( .A(n_1672), .B(n_1678), .Y(n_1671) );
INVx1_ASAP7_75t_L g1672 ( .A(n_1673), .Y(n_1672) );
NOR2xp33_ASAP7_75t_L g1673 ( .A(n_1674), .B(n_1676), .Y(n_1673) );
NOR2xp33_ASAP7_75t_L g1946 ( .A(n_1674), .B(n_1677), .Y(n_1946) );
INVx1_ASAP7_75t_L g1989 ( .A(n_1674), .Y(n_1989) );
HB1xp67_ASAP7_75t_L g1674 ( .A(n_1675), .Y(n_1674) );
INVx1_ASAP7_75t_L g1676 ( .A(n_1677), .Y(n_1676) );
NOR2xp33_ASAP7_75t_L g1992 ( .A(n_1677), .B(n_1989), .Y(n_1992) );
INVx1_ASAP7_75t_L g1678 ( .A(n_1679), .Y(n_1678) );
OAI221xp5_ASAP7_75t_L g1681 ( .A1(n_1682), .A2(n_1896), .B1(n_1898), .B2(n_1937), .C(n_1943), .Y(n_1681) );
AOI21xp5_ASAP7_75t_L g1682 ( .A1(n_1683), .A2(n_1822), .B(n_1870), .Y(n_1682) );
NAND5xp2_ASAP7_75t_L g1683 ( .A(n_1684), .B(n_1772), .C(n_1788), .D(n_1801), .E(n_1814), .Y(n_1683) );
AOI211xp5_ASAP7_75t_L g1684 ( .A1(n_1685), .A2(n_1716), .B(n_1731), .C(n_1756), .Y(n_1684) );
AND2x2_ASAP7_75t_L g1685 ( .A(n_1686), .B(n_1702), .Y(n_1685) );
AND2x2_ASAP7_75t_L g1848 ( .A(n_1686), .B(n_1783), .Y(n_1848) );
CKINVDCx5p33_ASAP7_75t_R g1686 ( .A(n_1687), .Y(n_1686) );
OR2x2_ASAP7_75t_L g1774 ( .A(n_1687), .B(n_1740), .Y(n_1774) );
AND2x2_ASAP7_75t_L g1782 ( .A(n_1687), .B(n_1783), .Y(n_1782) );
AOI322xp5_ASAP7_75t_L g1801 ( .A1(n_1687), .A2(n_1758), .A3(n_1802), .B1(n_1806), .B2(n_1807), .C1(n_1811), .C2(n_1812), .Y(n_1801) );
NAND2xp5_ASAP7_75t_L g1840 ( .A(n_1687), .B(n_1841), .Y(n_1840) );
NAND2xp5_ASAP7_75t_L g1857 ( .A(n_1687), .B(n_1858), .Y(n_1857) );
NAND2xp5_ASAP7_75t_L g1886 ( .A(n_1687), .B(n_1748), .Y(n_1886) );
O2A1O1Ixp33_ASAP7_75t_SL g1892 ( .A1(n_1687), .A2(n_1742), .B(n_1757), .C(n_1842), .Y(n_1892) );
INVx4_ASAP7_75t_L g1687 ( .A(n_1688), .Y(n_1687) );
INVx4_ASAP7_75t_L g1738 ( .A(n_1688), .Y(n_1738) );
NAND2xp5_ASAP7_75t_SL g1747 ( .A(n_1688), .B(n_1704), .Y(n_1747) );
AND2x2_ASAP7_75t_L g1775 ( .A(n_1688), .B(n_1776), .Y(n_1775) );
NOR2xp33_ASAP7_75t_L g1791 ( .A(n_1688), .B(n_1723), .Y(n_1791) );
OR2x2_ASAP7_75t_L g1810 ( .A(n_1688), .B(n_1704), .Y(n_1810) );
NOR2xp33_ASAP7_75t_L g1811 ( .A(n_1688), .B(n_1709), .Y(n_1811) );
NAND2xp5_ASAP7_75t_L g1837 ( .A(n_1688), .B(n_1817), .Y(n_1837) );
AND2x2_ASAP7_75t_L g1869 ( .A(n_1688), .B(n_1777), .Y(n_1869) );
AOI321xp33_ASAP7_75t_R g1881 ( .A1(n_1688), .A2(n_1716), .A3(n_1775), .B1(n_1787), .B2(n_1806), .C(n_1882), .Y(n_1881) );
AND2x4_ASAP7_75t_SL g1688 ( .A(n_1689), .B(n_1697), .Y(n_1688) );
AND2x4_ASAP7_75t_L g1690 ( .A(n_1691), .B(n_1692), .Y(n_1690) );
AND2x6_ASAP7_75t_L g1695 ( .A(n_1691), .B(n_1696), .Y(n_1695) );
AND2x6_ASAP7_75t_L g1698 ( .A(n_1691), .B(n_1699), .Y(n_1698) );
AND2x2_ASAP7_75t_L g1700 ( .A(n_1691), .B(n_1701), .Y(n_1700) );
AND2x2_ASAP7_75t_L g1707 ( .A(n_1691), .B(n_1701), .Y(n_1707) );
AND2x2_ASAP7_75t_L g1722 ( .A(n_1691), .B(n_1701), .Y(n_1722) );
NAND2xp5_ASAP7_75t_L g1767 ( .A(n_1691), .B(n_1692), .Y(n_1767) );
HB1xp67_ASAP7_75t_L g1990 ( .A(n_1692), .Y(n_1990) );
AND2x2_ASAP7_75t_L g1692 ( .A(n_1693), .B(n_1694), .Y(n_1692) );
INVx2_ASAP7_75t_L g1769 ( .A(n_1695), .Y(n_1769) );
AOI221xp5_ASAP7_75t_L g1890 ( .A1(n_1702), .A2(n_1832), .B1(n_1855), .B2(n_1891), .C(n_1892), .Y(n_1890) );
AND2x2_ASAP7_75t_L g1702 ( .A(n_1703), .B(n_1708), .Y(n_1702) );
OR2x2_ASAP7_75t_L g1752 ( .A(n_1703), .B(n_1709), .Y(n_1752) );
AND2x2_ASAP7_75t_L g1776 ( .A(n_1703), .B(n_1777), .Y(n_1776) );
OR2x2_ASAP7_75t_L g1842 ( .A(n_1703), .B(n_1742), .Y(n_1842) );
AND2x2_ASAP7_75t_L g1872 ( .A(n_1703), .B(n_1821), .Y(n_1872) );
INVx1_ASAP7_75t_L g1703 ( .A(n_1704), .Y(n_1703) );
NAND2xp5_ASAP7_75t_L g1790 ( .A(n_1704), .B(n_1713), .Y(n_1790) );
OR2x2_ASAP7_75t_L g1794 ( .A(n_1704), .B(n_1710), .Y(n_1794) );
AND2x2_ASAP7_75t_L g1796 ( .A(n_1704), .B(n_1748), .Y(n_1796) );
AND2x2_ASAP7_75t_L g1799 ( .A(n_1704), .B(n_1800), .Y(n_1799) );
AND2x2_ASAP7_75t_L g1853 ( .A(n_1704), .B(n_1778), .Y(n_1853) );
OR2x2_ASAP7_75t_L g1889 ( .A(n_1704), .B(n_1778), .Y(n_1889) );
AND2x2_ASAP7_75t_L g1704 ( .A(n_1705), .B(n_1706), .Y(n_1704) );
AND2x2_ASAP7_75t_L g1741 ( .A(n_1705), .B(n_1706), .Y(n_1741) );
NAND2xp5_ASAP7_75t_L g1781 ( .A(n_1708), .B(n_1782), .Y(n_1781) );
NAND3xp33_ASAP7_75t_L g1835 ( .A(n_1708), .B(n_1827), .C(n_1836), .Y(n_1835) );
NAND2xp5_ASAP7_75t_L g1849 ( .A(n_1708), .B(n_1834), .Y(n_1849) );
AND2x2_ASAP7_75t_L g1880 ( .A(n_1708), .B(n_1746), .Y(n_1880) );
INVx1_ASAP7_75t_L g1708 ( .A(n_1709), .Y(n_1708) );
OR2x2_ASAP7_75t_L g1830 ( .A(n_1709), .B(n_1810), .Y(n_1830) );
OR2x2_ASAP7_75t_L g1709 ( .A(n_1710), .B(n_1713), .Y(n_1709) );
NAND2xp5_ASAP7_75t_L g1742 ( .A(n_1710), .B(n_1743), .Y(n_1742) );
AND2x2_ASAP7_75t_L g1748 ( .A(n_1710), .B(n_1713), .Y(n_1748) );
INVx2_ASAP7_75t_L g1778 ( .A(n_1710), .Y(n_1778) );
NAND2x1p5_ASAP7_75t_L g1710 ( .A(n_1711), .B(n_1712), .Y(n_1710) );
INVx1_ASAP7_75t_L g1743 ( .A(n_1713), .Y(n_1743) );
AND2x2_ASAP7_75t_L g1777 ( .A(n_1713), .B(n_1778), .Y(n_1777) );
INVx1_ASAP7_75t_L g1800 ( .A(n_1713), .Y(n_1800) );
OR2x2_ASAP7_75t_L g1859 ( .A(n_1713), .B(n_1741), .Y(n_1859) );
AND2x2_ASAP7_75t_L g1713 ( .A(n_1714), .B(n_1715), .Y(n_1713) );
AOI221xp5_ASAP7_75t_L g1871 ( .A1(n_1716), .A2(n_1761), .B1(n_1872), .B2(n_1873), .C(n_1874), .Y(n_1871) );
INVx1_ASAP7_75t_L g1716 ( .A(n_1717), .Y(n_1716) );
OR2x2_ASAP7_75t_L g1717 ( .A(n_1718), .B(n_1723), .Y(n_1717) );
AOI221xp5_ASAP7_75t_L g1772 ( .A1(n_1718), .A2(n_1758), .B1(n_1773), .B2(n_1775), .C(n_1779), .Y(n_1772) );
AOI221xp5_ASAP7_75t_L g1788 ( .A1(n_1718), .A2(n_1789), .B1(n_1791), .B2(n_1792), .C(n_1797), .Y(n_1788) );
OAI322xp33_ASAP7_75t_L g1846 ( .A1(n_1718), .A2(n_1741), .A3(n_1847), .B1(n_1849), .B2(n_1850), .C1(n_1851), .C2(n_1852), .Y(n_1846) );
AND2x2_ASAP7_75t_L g1868 ( .A(n_1718), .B(n_1834), .Y(n_1868) );
INVx1_ASAP7_75t_L g1718 ( .A(n_1719), .Y(n_1718) );
INVx3_ASAP7_75t_L g1734 ( .A(n_1719), .Y(n_1734) );
AND2x2_ASAP7_75t_L g1750 ( .A(n_1719), .B(n_1751), .Y(n_1750) );
AND2x2_ASAP7_75t_L g1786 ( .A(n_1719), .B(n_1727), .Y(n_1786) );
OR2x2_ASAP7_75t_L g1818 ( .A(n_1719), .B(n_1727), .Y(n_1818) );
AND2x2_ASAP7_75t_L g1719 ( .A(n_1720), .B(n_1721), .Y(n_1719) );
AOI21xp33_ASAP7_75t_L g1895 ( .A1(n_1723), .A2(n_1774), .B(n_1795), .Y(n_1895) );
OR2x2_ASAP7_75t_L g1723 ( .A(n_1724), .B(n_1727), .Y(n_1723) );
INVx1_ASAP7_75t_L g1739 ( .A(n_1724), .Y(n_1739) );
INVx1_ASAP7_75t_L g1755 ( .A(n_1724), .Y(n_1755) );
NAND2xp5_ASAP7_75t_L g1724 ( .A(n_1725), .B(n_1726), .Y(n_1724) );
A2O1A1Ixp33_ASAP7_75t_L g1744 ( .A1(n_1727), .A2(n_1745), .B(n_1749), .C(n_1753), .Y(n_1744) );
INVx1_ASAP7_75t_L g1751 ( .A(n_1727), .Y(n_1751) );
AND2x2_ASAP7_75t_L g1758 ( .A(n_1727), .B(n_1734), .Y(n_1758) );
OR2x2_ASAP7_75t_L g1784 ( .A(n_1727), .B(n_1755), .Y(n_1784) );
OAI22xp5_ASAP7_75t_L g1792 ( .A1(n_1727), .A2(n_1793), .B1(n_1794), .B2(n_1795), .Y(n_1792) );
AND2x2_ASAP7_75t_L g1806 ( .A(n_1727), .B(n_1739), .Y(n_1806) );
INVx2_ASAP7_75t_L g1827 ( .A(n_1727), .Y(n_1827) );
INVx2_ASAP7_75t_L g1727 ( .A(n_1728), .Y(n_1727) );
OR2x2_ASAP7_75t_L g1820 ( .A(n_1728), .B(n_1755), .Y(n_1820) );
NAND2xp5_ASAP7_75t_L g1728 ( .A(n_1729), .B(n_1730), .Y(n_1728) );
NAND2xp5_ASAP7_75t_L g1731 ( .A(n_1732), .B(n_1744), .Y(n_1731) );
NAND2xp5_ASAP7_75t_L g1732 ( .A(n_1733), .B(n_1735), .Y(n_1732) );
CKINVDCx14_ASAP7_75t_R g1733 ( .A(n_1734), .Y(n_1733) );
NAND2xp5_ASAP7_75t_L g1813 ( .A(n_1734), .B(n_1739), .Y(n_1813) );
OR2x2_ASAP7_75t_L g1845 ( .A(n_1734), .B(n_1754), .Y(n_1845) );
OR2x2_ASAP7_75t_L g1850 ( .A(n_1734), .B(n_1739), .Y(n_1850) );
OR2x2_ASAP7_75t_L g1851 ( .A(n_1734), .B(n_1784), .Y(n_1851) );
AND2x2_ASAP7_75t_L g1855 ( .A(n_1734), .B(n_1783), .Y(n_1855) );
O2A1O1Ixp33_ASAP7_75t_SL g1874 ( .A1(n_1734), .A2(n_1805), .B(n_1875), .C(n_1877), .Y(n_1874) );
OR2x2_ASAP7_75t_L g1888 ( .A(n_1734), .B(n_1820), .Y(n_1888) );
A2O1A1Ixp33_ASAP7_75t_R g1893 ( .A1(n_1734), .A2(n_1848), .B(n_1894), .C(n_1895), .Y(n_1893) );
AOI221xp5_ASAP7_75t_L g1823 ( .A1(n_1735), .A2(n_1758), .B1(n_1784), .B2(n_1824), .C(n_1829), .Y(n_1823) );
NOR2xp33_ASAP7_75t_L g1735 ( .A(n_1736), .B(n_1740), .Y(n_1735) );
INVx1_ASAP7_75t_L g1736 ( .A(n_1737), .Y(n_1736) );
OAI21xp33_ASAP7_75t_L g1785 ( .A1(n_1737), .A2(n_1786), .B(n_1787), .Y(n_1785) );
AND2x2_ASAP7_75t_L g1737 ( .A(n_1738), .B(n_1739), .Y(n_1737) );
AND2x2_ASAP7_75t_L g1761 ( .A(n_1738), .B(n_1762), .Y(n_1761) );
NOR2x1_ASAP7_75t_L g1821 ( .A(n_1738), .B(n_1804), .Y(n_1821) );
NAND2x1_ASAP7_75t_L g1825 ( .A(n_1738), .B(n_1796), .Y(n_1825) );
CKINVDCx5p33_ASAP7_75t_R g1834 ( .A(n_1738), .Y(n_1834) );
NOR2xp33_ASAP7_75t_L g1876 ( .A(n_1738), .B(n_1751), .Y(n_1876) );
INVx2_ASAP7_75t_L g1817 ( .A(n_1739), .Y(n_1817) );
AND2x2_ASAP7_75t_L g1833 ( .A(n_1739), .B(n_1834), .Y(n_1833) );
NAND2xp5_ASAP7_75t_L g1789 ( .A(n_1740), .B(n_1790), .Y(n_1789) );
OR2x2_ASAP7_75t_L g1740 ( .A(n_1741), .B(n_1742), .Y(n_1740) );
AND2x2_ASAP7_75t_L g1787 ( .A(n_1741), .B(n_1777), .Y(n_1787) );
OR2x2_ASAP7_75t_L g1803 ( .A(n_1741), .B(n_1804), .Y(n_1803) );
AOI321xp33_ASAP7_75t_L g1865 ( .A1(n_1741), .A2(n_1763), .A3(n_1812), .B1(n_1866), .B2(n_1868), .C(n_1869), .Y(n_1865) );
OAI221xp5_ASAP7_75t_L g1756 ( .A1(n_1742), .A2(n_1757), .B1(n_1759), .B2(n_1760), .C(n_1763), .Y(n_1756) );
INVx1_ASAP7_75t_L g1762 ( .A(n_1742), .Y(n_1762) );
NAND2xp5_ASAP7_75t_L g1866 ( .A(n_1742), .B(n_1867), .Y(n_1866) );
INVx1_ASAP7_75t_L g1780 ( .A(n_1745), .Y(n_1780) );
AND2x2_ASAP7_75t_L g1745 ( .A(n_1746), .B(n_1748), .Y(n_1745) );
INVx1_ASAP7_75t_L g1746 ( .A(n_1747), .Y(n_1746) );
INVx1_ASAP7_75t_L g1804 ( .A(n_1748), .Y(n_1804) );
NAND2xp5_ASAP7_75t_L g1808 ( .A(n_1748), .B(n_1809), .Y(n_1808) );
OAI31xp33_ASAP7_75t_L g1814 ( .A1(n_1749), .A2(n_1815), .A3(n_1819), .B(n_1821), .Y(n_1814) );
NOR2xp33_ASAP7_75t_L g1749 ( .A(n_1750), .B(n_1752), .Y(n_1749) );
INVx1_ASAP7_75t_L g1759 ( .A(n_1750), .Y(n_1759) );
AOI221xp5_ASAP7_75t_L g1854 ( .A1(n_1750), .A2(n_1855), .B1(n_1856), .B2(n_1860), .C(n_1861), .Y(n_1854) );
OAI22xp5_ASAP7_75t_L g1824 ( .A1(n_1751), .A2(n_1825), .B1(n_1826), .B2(n_1828), .Y(n_1824) );
INVx1_ASAP7_75t_L g1864 ( .A(n_1752), .Y(n_1864) );
OAI211xp5_ASAP7_75t_L g1779 ( .A1(n_1753), .A2(n_1780), .B(n_1781), .C(n_1785), .Y(n_1779) );
INVx1_ASAP7_75t_L g1753 ( .A(n_1754), .Y(n_1753) );
NAND2xp5_ASAP7_75t_L g1757 ( .A(n_1754), .B(n_1758), .Y(n_1757) );
INVx1_ASAP7_75t_L g1754 ( .A(n_1755), .Y(n_1754) );
NOR2xp33_ASAP7_75t_L g1878 ( .A(n_1755), .B(n_1879), .Y(n_1878) );
A2O1A1Ixp33_ASAP7_75t_L g1883 ( .A1(n_1755), .A2(n_1786), .B(n_1821), .C(n_1843), .Y(n_1883) );
AND2x2_ASAP7_75t_L g1891 ( .A(n_1758), .B(n_1833), .Y(n_1891) );
INVx1_ASAP7_75t_L g1760 ( .A(n_1761), .Y(n_1760) );
INVx2_ASAP7_75t_L g1763 ( .A(n_1764), .Y(n_1763) );
INVx1_ASAP7_75t_L g1764 ( .A(n_1765), .Y(n_1764) );
INVx1_ASAP7_75t_L g1765 ( .A(n_1766), .Y(n_1765) );
OAI221xp5_ASAP7_75t_L g1766 ( .A1(n_1767), .A2(n_1768), .B1(n_1769), .B2(n_1770), .C(n_1771), .Y(n_1766) );
CKINVDCx5p33_ASAP7_75t_R g1897 ( .A(n_1767), .Y(n_1897) );
INVx1_ASAP7_75t_L g1773 ( .A(n_1774), .Y(n_1773) );
NAND2xp5_ASAP7_75t_L g1828 ( .A(n_1777), .B(n_1809), .Y(n_1828) );
INVx1_ASAP7_75t_L g1867 ( .A(n_1777), .Y(n_1867) );
INVx1_ASAP7_75t_L g1793 ( .A(n_1782), .Y(n_1793) );
NAND2xp5_ASAP7_75t_L g1798 ( .A(n_1782), .B(n_1799), .Y(n_1798) );
CKINVDCx5p33_ASAP7_75t_R g1783 ( .A(n_1784), .Y(n_1783) );
INVx1_ASAP7_75t_L g1894 ( .A(n_1790), .Y(n_1894) );
INVx1_ASAP7_75t_L g1832 ( .A(n_1794), .Y(n_1832) );
INVx1_ASAP7_75t_L g1795 ( .A(n_1796), .Y(n_1795) );
INVxp67_ASAP7_75t_L g1797 ( .A(n_1798), .Y(n_1797) );
INVx1_ASAP7_75t_L g1805 ( .A(n_1799), .Y(n_1805) );
NAND2xp5_ASAP7_75t_SL g1802 ( .A(n_1803), .B(n_1805), .Y(n_1802) );
INVx1_ASAP7_75t_L g1860 ( .A(n_1803), .Y(n_1860) );
INVx1_ASAP7_75t_L g1807 ( .A(n_1808), .Y(n_1807) );
OAI211xp5_ASAP7_75t_L g1884 ( .A1(n_1809), .A2(n_1885), .B(n_1887), .C(n_1889), .Y(n_1884) );
INVx1_ASAP7_75t_L g1809 ( .A(n_1810), .Y(n_1809) );
INVx1_ASAP7_75t_L g1812 ( .A(n_1813), .Y(n_1812) );
INVx1_ASAP7_75t_L g1815 ( .A(n_1816), .Y(n_1815) );
OR2x2_ASAP7_75t_L g1816 ( .A(n_1817), .B(n_1818), .Y(n_1816) );
CKINVDCx5p33_ASAP7_75t_R g1819 ( .A(n_1820), .Y(n_1819) );
OAI211xp5_ASAP7_75t_L g1829 ( .A1(n_1820), .A2(n_1830), .B(n_1831), .C(n_1835), .Y(n_1829) );
NAND4xp25_ASAP7_75t_L g1822 ( .A(n_1823), .B(n_1838), .C(n_1854), .D(n_1865), .Y(n_1822) );
NAND3xp33_ASAP7_75t_L g1831 ( .A(n_1826), .B(n_1832), .C(n_1833), .Y(n_1831) );
INVx1_ASAP7_75t_L g1826 ( .A(n_1827), .Y(n_1826) );
INVx1_ASAP7_75t_L g1843 ( .A(n_1830), .Y(n_1843) );
INVx1_ASAP7_75t_L g1836 ( .A(n_1837), .Y(n_1836) );
O2A1O1Ixp33_ASAP7_75t_L g1838 ( .A1(n_1839), .A2(n_1843), .B(n_1844), .C(n_1846), .Y(n_1838) );
INVxp67_ASAP7_75t_L g1839 ( .A(n_1840), .Y(n_1839) );
INVx1_ASAP7_75t_L g1841 ( .A(n_1842), .Y(n_1841) );
INVx1_ASAP7_75t_L g1844 ( .A(n_1845), .Y(n_1844) );
INVx1_ASAP7_75t_L g1847 ( .A(n_1848), .Y(n_1847) );
INVx1_ASAP7_75t_L g1863 ( .A(n_1850), .Y(n_1863) );
INVx1_ASAP7_75t_L g1873 ( .A(n_1851), .Y(n_1873) );
CKINVDCx14_ASAP7_75t_R g1852 ( .A(n_1853), .Y(n_1852) );
INVx1_ASAP7_75t_L g1856 ( .A(n_1857), .Y(n_1856) );
INVxp67_ASAP7_75t_L g1858 ( .A(n_1859), .Y(n_1858) );
INVx1_ASAP7_75t_L g1861 ( .A(n_1862), .Y(n_1861) );
NAND2xp5_ASAP7_75t_L g1862 ( .A(n_1863), .B(n_1864), .Y(n_1862) );
NAND4xp25_ASAP7_75t_L g1870 ( .A(n_1871), .B(n_1881), .C(n_1890), .D(n_1893), .Y(n_1870) );
INVx1_ASAP7_75t_L g1875 ( .A(n_1876), .Y(n_1875) );
INVx1_ASAP7_75t_L g1877 ( .A(n_1878), .Y(n_1877) );
INVx1_ASAP7_75t_L g1879 ( .A(n_1880), .Y(n_1879) );
NAND2xp5_ASAP7_75t_SL g1882 ( .A(n_1883), .B(n_1884), .Y(n_1882) );
INVxp67_ASAP7_75t_SL g1885 ( .A(n_1886), .Y(n_1885) );
INVx1_ASAP7_75t_L g1887 ( .A(n_1888), .Y(n_1887) );
CKINVDCx20_ASAP7_75t_R g1896 ( .A(n_1897), .Y(n_1896) );
INVx1_ASAP7_75t_L g1935 ( .A(n_1899), .Y(n_1935) );
NAND3xp33_ASAP7_75t_L g1899 ( .A(n_1900), .B(n_1907), .C(n_1913), .Y(n_1899) );
NOR2xp33_ASAP7_75t_L g1913 ( .A(n_1914), .B(n_1927), .Y(n_1913) );
OAI22xp33_ASAP7_75t_L g1928 ( .A1(n_1916), .A2(n_1922), .B1(n_1929), .B2(n_1931), .Y(n_1928) );
INVx2_ASAP7_75t_L g1929 ( .A(n_1930), .Y(n_1929) );
CKINVDCx20_ASAP7_75t_R g1937 ( .A(n_1938), .Y(n_1937) );
CKINVDCx20_ASAP7_75t_R g1938 ( .A(n_1939), .Y(n_1938) );
INVx3_ASAP7_75t_L g1939 ( .A(n_1940), .Y(n_1939) );
BUFx3_ASAP7_75t_L g1940 ( .A(n_1941), .Y(n_1940) );
HB1xp67_ASAP7_75t_L g1944 ( .A(n_1945), .Y(n_1944) );
BUFx3_ASAP7_75t_L g1945 ( .A(n_1946), .Y(n_1945) );
INVxp33_ASAP7_75t_SL g1947 ( .A(n_1948), .Y(n_1947) );
HB1xp67_ASAP7_75t_L g1949 ( .A(n_1950), .Y(n_1949) );
AND3x1_ASAP7_75t_L g1950 ( .A(n_1951), .B(n_1971), .C(n_1981), .Y(n_1950) );
NOR2xp33_ASAP7_75t_L g1951 ( .A(n_1952), .B(n_1966), .Y(n_1951) );
HB1xp67_ASAP7_75t_L g1973 ( .A(n_1974), .Y(n_1973) );
INVxp67_ASAP7_75t_SL g1974 ( .A(n_1975), .Y(n_1974) );
HB1xp67_ASAP7_75t_L g1987 ( .A(n_1988), .Y(n_1987) );
OAI21xp5_ASAP7_75t_L g1988 ( .A1(n_1989), .A2(n_1990), .B(n_1991), .Y(n_1988) );
INVx1_ASAP7_75t_L g1991 ( .A(n_1992), .Y(n_1991) );
endmodule