module fake_jpeg_31533_n_133 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_133);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_133;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

BUFx10_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_21),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_41),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_5),
.B(n_26),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_42),
.Y(n_56)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_55),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_55),
.Y(n_58)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_0),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_60),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_1),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_2),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_64),
.Y(n_67)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_59),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_68),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_62),
.A2(n_52),
.B1(n_51),
.B2(n_43),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_69),
.A2(n_43),
.B1(n_48),
.B2(n_49),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_64),
.A2(n_52),
.B1(n_51),
.B2(n_46),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_71),
.A2(n_56),
.B1(n_47),
.B2(n_54),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_53),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_73),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_46),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_45),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_2),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_46),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_68),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_79),
.A2(n_85),
.B1(n_88),
.B2(n_91),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_77),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_80),
.B(n_83),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_73),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_87),
.Y(n_97)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_71),
.A2(n_40),
.B1(n_20),
.B2(n_22),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_75),
.A2(n_3),
.B(n_4),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_6),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_67),
.A2(n_19),
.B1(n_37),
.B2(n_36),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_90),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_78),
.A2(n_17),
.B1(n_35),
.B2(n_34),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_70),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_92),
.A2(n_93),
.B(n_76),
.Y(n_96)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_84),
.A2(n_76),
.B(n_68),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_94),
.A2(n_108),
.B(n_109),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_82),
.B(n_81),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_99),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_SL g98 ( 
.A(n_89),
.B(n_16),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_SL g118 ( 
.A(n_98),
.B(n_102),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_100),
.B(n_104),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_79),
.B(n_23),
.Y(n_102)
);

AND2x6_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_18),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_90),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_105),
.A2(n_15),
.B1(n_25),
.B2(n_28),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_87),
.A2(n_7),
.B(n_8),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_107),
.Y(n_112)
);

HAxp5_ASAP7_75t_SL g108 ( 
.A(n_86),
.B(n_9),
.CON(n_108),
.SN(n_108)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_27),
.Y(n_109)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_106),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_110),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_103),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_111),
.B(n_113),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_101),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_116),
.A2(n_97),
.B(n_108),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_120),
.A2(n_119),
.B1(n_115),
.B2(n_114),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_114),
.A2(n_119),
.B(n_117),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_121),
.A2(n_94),
.B(n_98),
.Y(n_127)
);

BUFx24_ASAP7_75t_SL g123 ( 
.A(n_112),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g126 ( 
.A(n_123),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_125),
.A2(n_127),
.B1(n_124),
.B2(n_118),
.Y(n_128)
);

AOI322xp5_ASAP7_75t_L g129 ( 
.A1(n_128),
.A2(n_118),
.A3(n_104),
.B1(n_102),
.B2(n_126),
.C1(n_110),
.C2(n_122),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_129),
.A2(n_29),
.B(n_30),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_130),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_131),
.A2(n_31),
.B(n_32),
.Y(n_132)
);

FAx1_ASAP7_75t_SL g133 ( 
.A(n_132),
.B(n_38),
.CI(n_130),
.CON(n_133),
.SN(n_133)
);


endmodule