module real_jpeg_7993_n_12 (n_252, n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_252;
input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_215;
wire n_166;
wire n_221;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_164;
wire n_48;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_198;
wire n_203;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_193;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_187;
wire n_97;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_244;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

BUFx24_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g19 ( 
.A1(n_1),
.A2(n_11),
.B1(n_20),
.B2(n_21),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_1),
.A2(n_20),
.B1(n_24),
.B2(n_25),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_1),
.A2(n_20),
.B1(n_40),
.B2(n_41),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_1),
.A2(n_20),
.B1(n_55),
.B2(n_56),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_2),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_23)
);

INVx2_ASAP7_75t_SL g26 ( 
.A(n_2),
.Y(n_26)
);

AOI21xp33_ASAP7_75t_L g193 ( 
.A1(n_2),
.A2(n_10),
.B(n_25),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_3),
.A2(n_40),
.B1(n_41),
.B2(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_3),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_3),
.A2(n_55),
.B1(n_56),
.B2(n_63),
.Y(n_78)
);

BUFx10_ASAP7_75t_L g83 ( 
.A(n_4),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_5),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_6),
.A2(n_55),
.B1(n_56),
.B2(n_59),
.Y(n_54)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_6),
.Y(n_59)
);

A2O1A1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_6),
.A2(n_40),
.B(n_54),
.C(n_61),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_6),
.B(n_40),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_6),
.A2(n_10),
.B(n_56),
.Y(n_135)
);

BUFx6f_ASAP7_75t_SL g39 ( 
.A(n_7),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_9),
.A2(n_24),
.B1(n_25),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_9),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_9),
.A2(n_37),
.B1(n_40),
.B2(n_41),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_9),
.A2(n_37),
.B1(n_55),
.B2(n_56),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_10),
.A2(n_11),
.B1(n_21),
.B2(n_29),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_10),
.A2(n_24),
.B1(n_25),
.B2(n_29),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_10),
.A2(n_29),
.B1(n_40),
.B2(n_41),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_10),
.A2(n_29),
.B1(n_55),
.B2(n_56),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_10),
.B(n_74),
.Y(n_153)
);

O2A1O1Ixp33_ASAP7_75t_L g163 ( 
.A1(n_10),
.A2(n_24),
.B(n_39),
.C(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_10),
.B(n_22),
.Y(n_175)
);

INVx2_ASAP7_75t_SL g21 ( 
.A(n_11),
.Y(n_21)
);

A2O1A1Ixp33_ASAP7_75t_L g30 ( 
.A1(n_11),
.A2(n_23),
.B(n_26),
.C(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_11),
.B(n_26),
.Y(n_31)
);

A2O1A1Ixp33_ASAP7_75t_L g192 ( 
.A1(n_11),
.A2(n_26),
.B(n_29),
.C(n_193),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_116),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_114),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_93),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_15),
.B(n_93),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g15 ( 
.A1(n_16),
.A2(n_75),
.B1(n_76),
.B2(n_92),
.Y(n_15)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_16),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_66),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_32),
.B1(n_33),
.B2(n_65),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_18),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_18),
.A2(n_65),
.B1(n_184),
.B2(n_185),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_18),
.B(n_107),
.C(n_186),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_18),
.A2(n_65),
.B1(n_219),
.B2(n_220),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_18),
.B(n_217),
.C(n_219),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_22),
.B(n_27),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_19),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_23),
.B(n_30),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_23),
.A2(n_28),
.B1(n_30),
.B2(n_106),
.Y(n_105)
);

A2O1A1Ixp33_ASAP7_75t_L g48 ( 
.A1(n_24),
.A2(n_38),
.B(n_39),
.C(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_24),
.B(n_39),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_30),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_28),
.Y(n_90)
);

A2O1A1Ixp33_ASAP7_75t_L g134 ( 
.A1(n_29),
.A2(n_41),
.B(n_59),
.C(n_135),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_29),
.B(n_82),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_29),
.B(n_54),
.Y(n_143)
);

OAI21xp33_ASAP7_75t_L g164 ( 
.A1(n_29),
.A2(n_40),
.B(n_44),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_33),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_34),
.A2(n_50),
.B1(n_51),
.B2(n_64),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_34),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_38),
.B(n_45),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_40),
.B1(n_41),
.B2(n_44),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_39),
.Y(n_44)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_46),
.A2(n_71),
.B(n_74),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_48),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_47),
.B(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_52),
.B(n_62),
.Y(n_51)
);

INVxp33_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_53),
.B(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_60),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_54),
.A2(n_60),
.B1(n_62),
.B2(n_68),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_54),
.A2(n_68),
.B(n_86),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_54),
.A2(n_60),
.B1(n_88),
.B2(n_103),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_54),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_55),
.B(n_141),
.Y(n_140)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_56),
.B(n_82),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx24_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_60),
.B(n_88),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_66),
.A2(n_67),
.B(n_69),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_69),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_69),
.A2(n_70),
.B1(n_172),
.B2(n_173),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_69),
.A2(n_70),
.B1(n_104),
.B2(n_105),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_70),
.B(n_124),
.C(n_175),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_70),
.B(n_104),
.C(n_209),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_72),
.B1(n_73),
.B2(n_74),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_72),
.B(n_74),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_84),
.B(n_89),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_85),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_77),
.A2(n_89),
.B1(n_112),
.B2(n_113),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_77),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_77),
.A2(n_85),
.B1(n_112),
.B2(n_237),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_79),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_79),
.B(n_128),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_80),
.B(n_83),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_80),
.A2(n_83),
.B1(n_99),
.B2(n_100),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_81),
.B(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_81),
.A2(n_82),
.B1(n_126),
.B2(n_128),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_82),
.A2(n_204),
.B(n_205),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_83),
.A2(n_125),
.B(n_127),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_SL g110 ( 
.A(n_84),
.B(n_111),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_85),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_87),
.A2(n_131),
.B(n_132),
.Y(n_130)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_88),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_89),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_91),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_108),
.C(n_109),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_94),
.A2(n_95),
.B1(n_242),
.B2(n_243),
.Y(n_241)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_104),
.C(n_107),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_96),
.A2(n_97),
.B1(n_233),
.B2(n_234),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_101),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_98),
.A2(n_101),
.B1(n_102),
.B2(n_215),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_98),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_99),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_101),
.A2(n_102),
.B1(n_152),
.B2(n_153),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_101),
.A2(n_102),
.B1(n_177),
.B2(n_178),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_102),
.B(n_144),
.C(n_152),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_102),
.B(n_171),
.C(n_178),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_103),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_104),
.A2(n_105),
.B1(n_107),
.B2(n_161),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_107),
.A2(n_130),
.B1(n_136),
.B2(n_161),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_107),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_107),
.B(n_130),
.C(n_166),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_107),
.A2(n_161),
.B1(n_186),
.B2(n_188),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_108),
.A2(n_109),
.B1(n_110),
.B2(n_244),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_108),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

AOI321xp33_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_226),
.A3(n_239),
.B1(n_245),
.B2(n_250),
.C(n_252),
.Y(n_116)
);

NOR3xp33_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_198),
.C(n_223),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_180),
.B(n_197),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_168),
.B(n_179),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_156),
.B(n_167),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_122),
.A2(n_147),
.B(n_155),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_137),
.B(n_146),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_129),
.Y(n_123)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_124),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_124),
.B(n_129),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_124),
.A2(n_139),
.B1(n_174),
.B2(n_175),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_127),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_133),
.B1(n_134),
.B2(n_136),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_130),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_130),
.B(n_134),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_130),
.A2(n_136),
.B1(n_202),
.B2(n_203),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_136),
.B(n_203),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_142),
.B(n_145),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_144),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_143),
.B(n_144),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_144),
.A2(n_150),
.B1(n_151),
.B2(n_154),
.Y(n_149)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_144),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_144),
.A2(n_154),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_144),
.B(n_191),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_149),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_148),
.B(n_149),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_157),
.B(n_158),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_159),
.A2(n_160),
.B1(n_162),
.B2(n_166),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_162),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_165),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_163),
.B(n_165),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_169),
.B(n_170),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_176),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_177),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_181),
.B(n_182),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_189),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_183),
.B(n_190),
.C(n_196),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_186),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_194),
.B1(n_195),
.B2(n_196),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_190),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_194),
.Y(n_196)
);

CKINVDCx14_ASAP7_75t_R g198 ( 
.A(n_199),
.Y(n_198)
);

AOI21xp33_ASAP7_75t_L g246 ( 
.A1(n_199),
.A2(n_247),
.B(n_248),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_210),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_200),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_200),
.B(n_210),
.Y(n_248)
);

FAx1_ASAP7_75t_SL g200 ( 
.A(n_201),
.B(n_206),
.CI(n_207),
.CON(n_200),
.SN(n_200)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_203),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_212),
.B1(n_213),
.B2(n_222),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_211),
.Y(n_222)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_216),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_214),
.B(n_216),
.C(n_222),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_224),
.B(n_225),
.Y(n_247)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_227),
.A2(n_246),
.B(n_249),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_228),
.B(n_229),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_238),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_231),
.A2(n_232),
.B1(n_235),
.B2(n_236),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_231),
.B(n_236),
.C(n_238),
.Y(n_240)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_234),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_240),
.B(n_241),
.Y(n_250)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);


endmodule