module fake_jpeg_11258_n_204 (n_13, n_21, n_53, n_33, n_54, n_1, n_45, n_10, n_23, n_27, n_55, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_204);

input n_13;
input n_21;
input n_53;
input n_33;
input n_54;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_55;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_204;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g56 ( 
.A(n_55),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_52),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_20),
.Y(n_59)
);

BUFx4f_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_34),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_7),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_6),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_9),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_14),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_28),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_46),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_11),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_26),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_24),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_7),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_1),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_8),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_48),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_33),
.Y(n_79)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_12),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_35),
.Y(n_82)
);

BUFx10_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_15),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_37),
.Y(n_85)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_83),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_83),
.Y(n_88)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_62),
.B(n_0),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_89),
.B(n_92),
.Y(n_99)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_83),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_93),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_57),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_94),
.B(n_84),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_95),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_92),
.A2(n_90),
.B1(n_86),
.B2(n_88),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_96),
.A2(n_100),
.B1(n_82),
.B2(n_73),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_92),
.A2(n_81),
.B1(n_71),
.B2(n_75),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_101),
.B(n_102),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_63),
.C(n_64),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_87),
.A2(n_75),
.B1(n_56),
.B2(n_68),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_103),
.A2(n_111),
.B1(n_84),
.B2(n_93),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_89),
.B(n_67),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_109),
.B(n_110),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_94),
.B(n_66),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_95),
.A2(n_71),
.B1(n_81),
.B2(n_82),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_107),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_112),
.B(n_113),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_99),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_114),
.Y(n_154)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_106),
.Y(n_115)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_115),
.Y(n_134)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_105),
.Y(n_116)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_116),
.Y(n_140)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_104),
.Y(n_117)
);

INVx3_ASAP7_75t_SL g138 ( 
.A(n_117),
.Y(n_138)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_105),
.Y(n_118)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_118),
.Y(n_146)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_97),
.Y(n_119)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_119),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_121),
.A2(n_128),
.B1(n_60),
.B2(n_1),
.Y(n_136)
);

A2O1A1Ixp33_ASAP7_75t_L g122 ( 
.A1(n_103),
.A2(n_77),
.B(n_70),
.C(n_74),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_122),
.B(n_132),
.Y(n_135)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_104),
.Y(n_123)
);

INVx2_ASAP7_75t_SL g139 ( 
.A(n_123),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_96),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_124),
.B(n_130),
.Y(n_137)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_108),
.Y(n_125)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_125),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_100),
.A2(n_81),
.B1(n_82),
.B2(n_73),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_126),
.A2(n_131),
.B1(n_133),
.B2(n_4),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_98),
.A2(n_59),
.B1(n_85),
.B2(n_79),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_98),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_129),
.Y(n_145)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_108),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_111),
.A2(n_61),
.B1(n_69),
.B2(n_72),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_109),
.B(n_94),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_111),
.A2(n_78),
.B1(n_60),
.B2(n_2),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_136),
.A2(n_155),
.B1(n_11),
.B2(n_12),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_127),
.B(n_0),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_141),
.B(n_143),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_120),
.B(n_2),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_131),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_144),
.B(n_151),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_129),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_147),
.Y(n_172)
);

BUFx5_ASAP7_75t_L g148 ( 
.A(n_117),
.Y(n_148)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_148),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_114),
.A2(n_3),
.B(n_4),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_150),
.A2(n_13),
.B(n_14),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_133),
.B(n_3),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_152),
.A2(n_5),
.B1(n_9),
.B2(n_10),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_126),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_155)
);

AO21x1_ASAP7_75t_L g184 ( 
.A1(n_156),
.A2(n_162),
.B(n_165),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_142),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_157),
.B(n_160),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_149),
.B(n_54),
.C(n_30),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_159),
.B(n_163),
.Y(n_185)
);

OR2x2_ASAP7_75t_L g160 ( 
.A(n_135),
.B(n_10),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_137),
.B(n_32),
.C(n_47),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_146),
.B(n_134),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_164),
.B(n_166),
.Y(n_178)
);

INVxp33_ASAP7_75t_L g165 ( 
.A(n_138),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_140),
.B(n_13),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_154),
.A2(n_139),
.B1(n_138),
.B2(n_155),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_167),
.B(n_169),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_168),
.B(n_170),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_154),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_169)
);

OR2x2_ASAP7_75t_L g170 ( 
.A(n_153),
.B(n_19),
.Y(n_170)
);

OA21x2_ASAP7_75t_L g173 ( 
.A1(n_150),
.A2(n_21),
.B(n_23),
.Y(n_173)
);

AO22x1_ASAP7_75t_SL g175 ( 
.A1(n_173),
.A2(n_27),
.B1(n_29),
.B2(n_31),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_158),
.Y(n_174)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_174),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_175),
.Y(n_188)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_161),
.Y(n_176)
);

NAND3xp33_ASAP7_75t_L g190 ( 
.A(n_176),
.B(n_181),
.C(n_183),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_171),
.B(n_139),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_177),
.B(n_160),
.C(n_170),
.Y(n_186)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_172),
.Y(n_181)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_172),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_186),
.B(n_189),
.Y(n_195)
);

BUFx24_ASAP7_75t_SL g189 ( 
.A(n_179),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_184),
.A2(n_182),
.B1(n_173),
.B2(n_165),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_191),
.A2(n_182),
.B1(n_180),
.B2(n_175),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_178),
.B(n_159),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_192),
.B(n_185),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_193),
.B(n_194),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_196),
.A2(n_188),
.B(n_195),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_197),
.A2(n_190),
.B(n_194),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_198),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_199),
.A2(n_187),
.B(n_38),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_200),
.B(n_147),
.C(n_145),
.Y(n_201)
);

OAI311xp33_ASAP7_75t_L g202 ( 
.A1(n_201),
.A2(n_36),
.A3(n_39),
.B1(n_40),
.C1(n_41),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_202),
.B(n_43),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_203),
.B(n_45),
.Y(n_204)
);


endmodule