module fake_jpeg_312_n_148 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_148);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_148;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx6_ASAP7_75t_SL g41 ( 
.A(n_22),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_23),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_35),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_34),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_0),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_0),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_55),
.Y(n_58)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_57),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_53),
.A2(n_48),
.B1(n_44),
.B2(n_46),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_60),
.A2(n_48),
.B1(n_50),
.B2(n_38),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_61),
.B(n_63),
.Y(n_76)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_37),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_37),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_66),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_38),
.Y(n_66)
);

INVxp33_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_69),
.Y(n_97)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_70),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_64),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_71),
.B(n_77),
.Y(n_92)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_75),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_68),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_82),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_45),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_60),
.A2(n_50),
.B1(n_42),
.B2(n_47),
.Y(n_81)
);

OA21x2_ASAP7_75t_L g86 ( 
.A1(n_81),
.A2(n_49),
.B(n_45),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_83),
.B(n_40),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_80),
.B(n_42),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_85),
.B(n_91),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_86),
.Y(n_101)
);

AND2x2_ASAP7_75t_SL g87 ( 
.A(n_72),
.B(n_45),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_87),
.Y(n_114)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_89),
.Y(n_103)
);

A2O1A1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_76),
.A2(n_51),
.B(n_43),
.C(n_3),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_69),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_95),
.Y(n_99)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_82),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_96),
.A2(n_14),
.B1(n_36),
.B2(n_32),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_81),
.C(n_79),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_18),
.C(n_30),
.Y(n_123)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_98),
.Y(n_104)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_104),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_92),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_105),
.B(n_107),
.Y(n_122)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_97),
.Y(n_106)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_106),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_85),
.B(n_40),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_108),
.B(n_112),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_86),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_109),
.A2(n_110),
.B1(n_113),
.B2(n_6),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_89),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_97),
.Y(n_111)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_111),
.Y(n_117)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_94),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_113)
);

AO22x1_ASAP7_75t_SL g118 ( 
.A1(n_109),
.A2(n_84),
.B1(n_88),
.B2(n_95),
.Y(n_118)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_118),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_119),
.B(n_124),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_114),
.A2(n_20),
.B(n_31),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_123),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_114),
.A2(n_16),
.B(n_29),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_99),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_125),
.B(n_126),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_8),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_103),
.B(n_8),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_SL g128 ( 
.A(n_127),
.B(n_108),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_128),
.B(n_132),
.Y(n_135)
);

AOI321xp33_ASAP7_75t_L g132 ( 
.A1(n_120),
.A2(n_101),
.A3(n_102),
.B1(n_9),
.B2(n_10),
.C(n_13),
.Y(n_132)
);

A2O1A1O1Ixp25_ASAP7_75t_L g133 ( 
.A1(n_122),
.A2(n_104),
.B(n_25),
.C(n_11),
.D(n_12),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_133),
.B(n_123),
.Y(n_138)
);

INVx1_ASAP7_75t_SL g136 ( 
.A(n_129),
.Y(n_136)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_136),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_131),
.A2(n_119),
.B1(n_118),
.B2(n_115),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_137),
.B(n_138),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_117),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_134),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_135),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_139),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_144),
.B(n_130),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_145),
.A2(n_131),
.B(n_136),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_146),
.A2(n_116),
.B(n_118),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_26),
.Y(n_148)
);


endmodule