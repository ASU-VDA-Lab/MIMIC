module fake_jpeg_299_n_672 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_672);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_672;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_145;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_16),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_12),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx6_ASAP7_75t_SL g38 ( 
.A(n_16),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx24_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_17),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_5),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_5),
.Y(n_44)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_15),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_4),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_13),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_56),
.Y(n_59)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_59),
.Y(n_136)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_56),
.Y(n_60)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_60),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_61),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_23),
.B(n_9),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_62),
.B(n_95),
.Y(n_137)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_63),
.Y(n_149)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_64),
.Y(n_158)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g211 ( 
.A(n_65),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_66),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_29),
.B(n_9),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_67),
.B(n_72),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_68),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_69),
.Y(n_181)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_70),
.Y(n_161)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_71),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_29),
.B(n_9),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_33),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_73),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_74),
.Y(n_186)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_38),
.Y(n_75)
);

INVx2_ASAP7_75t_SL g213 ( 
.A(n_75),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_50),
.B(n_9),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_76),
.B(n_80),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_33),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_77),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_78),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_79),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_8),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_81),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_82),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

INVx8_ASAP7_75t_L g148 ( 
.A(n_83),
.Y(n_148)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_34),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_84),
.Y(n_196)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_85),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

INVx8_ASAP7_75t_L g162 ( 
.A(n_86),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_22),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_87),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_22),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_88),
.Y(n_221)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_22),
.Y(n_89)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_89),
.Y(n_166)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_40),
.Y(n_90)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_90),
.Y(n_134)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_23),
.Y(n_91)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_91),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_35),
.A2(n_8),
.B1(n_18),
.B2(n_16),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_92),
.A2(n_25),
.B1(n_42),
.B2(n_51),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_35),
.B(n_8),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_93),
.B(n_99),
.Y(n_224)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_35),
.Y(n_94)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_94),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_30),
.B(n_58),
.Y(n_95)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_22),
.Y(n_96)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_96),
.Y(n_173)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_31),
.Y(n_97)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_97),
.Y(n_176)
);

BUFx12_ASAP7_75t_L g98 ( 
.A(n_45),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g143 ( 
.A(n_98),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_27),
.B(n_8),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_22),
.Y(n_100)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_100),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_22),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g189 ( 
.A(n_101),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_31),
.Y(n_102)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_102),
.Y(n_179)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_34),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g155 ( 
.A(n_103),
.Y(n_155)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_31),
.Y(n_104)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_104),
.Y(n_193)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_31),
.Y(n_105)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_105),
.Y(n_195)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_34),
.Y(n_106)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_106),
.Y(n_182)
);

INVx13_ASAP7_75t_L g107 ( 
.A(n_45),
.Y(n_107)
);

BUFx8_ASAP7_75t_L g194 ( 
.A(n_107),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_57),
.Y(n_108)
);

INVx5_ASAP7_75t_L g180 ( 
.A(n_108),
.Y(n_180)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

INVx5_ASAP7_75t_L g187 ( 
.A(n_109),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_34),
.Y(n_110)
);

INVx5_ASAP7_75t_L g188 ( 
.A(n_110),
.Y(n_188)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_57),
.Y(n_111)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_111),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_27),
.B(n_10),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_112),
.B(n_114),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_57),
.Y(n_113)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_113),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_27),
.B(n_10),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_57),
.Y(n_115)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_115),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_21),
.Y(n_116)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_116),
.Y(n_171)
);

AOI21xp33_ASAP7_75t_L g117 ( 
.A1(n_21),
.A2(n_19),
.B(n_18),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_117),
.B(n_120),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_57),
.Y(n_118)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_118),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_21),
.Y(n_119)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_119),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_30),
.B(n_16),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_32),
.Y(n_121)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_121),
.Y(n_163)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_32),
.Y(n_122)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_122),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_28),
.B(n_15),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_123),
.B(n_51),
.Y(n_135)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_32),
.Y(n_124)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_124),
.Y(n_169)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_43),
.Y(n_125)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_125),
.Y(n_210)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_43),
.Y(n_126)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_126),
.Y(n_223)
);

BUFx5_ASAP7_75t_L g127 ( 
.A(n_40),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_127),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_43),
.Y(n_128)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_128),
.Y(n_226)
);

INVx11_ASAP7_75t_L g129 ( 
.A(n_40),
.Y(n_129)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_129),
.Y(n_200)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_45),
.Y(n_130)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_130),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_28),
.B(n_15),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_131),
.B(n_14),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_75),
.A2(n_36),
.B1(n_41),
.B2(n_39),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_132),
.A2(n_147),
.B1(n_150),
.B2(n_151),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_135),
.B(n_141),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_62),
.A2(n_36),
.B1(n_41),
.B2(n_39),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_138),
.A2(n_164),
.B1(n_184),
.B2(n_216),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_145),
.B(n_3),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_129),
.A2(n_36),
.B1(n_41),
.B2(n_39),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_65),
.A2(n_28),
.B1(n_58),
.B2(n_44),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_70),
.A2(n_58),
.B1(n_44),
.B2(n_42),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_71),
.A2(n_44),
.B1(n_42),
.B2(n_25),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_154),
.A2(n_174),
.B1(n_40),
.B2(n_53),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_156),
.A2(n_160),
.B1(n_177),
.B2(n_199),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_85),
.A2(n_51),
.B1(n_25),
.B2(n_55),
.Y(n_157)
);

OR2x2_ASAP7_75t_L g233 ( 
.A(n_157),
.B(n_26),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_89),
.B(n_20),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_159),
.B(n_172),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_61),
.A2(n_20),
.B1(n_54),
.B2(n_48),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_73),
.A2(n_20),
.B1(n_54),
.B2(n_48),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_96),
.B(n_54),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_110),
.A2(n_40),
.B1(n_46),
.B2(n_48),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_66),
.A2(n_55),
.B1(n_26),
.B2(n_47),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_116),
.B(n_47),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_178),
.B(n_204),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_74),
.A2(n_78),
.B1(n_79),
.B2(n_82),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_128),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_185),
.Y(n_232)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_119),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_197),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_68),
.A2(n_55),
.B1(n_26),
.B2(n_47),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_111),
.B(n_46),
.Y(n_204)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_130),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_206),
.B(n_208),
.Y(n_258)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_103),
.Y(n_207)
);

INVxp67_ASAP7_75t_SL g272 ( 
.A(n_207),
.Y(n_272)
);

NOR3xp33_ASAP7_75t_L g208 ( 
.A(n_107),
.B(n_46),
.C(n_37),
.Y(n_208)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_106),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_212),
.B(n_215),
.Y(n_267)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_103),
.Y(n_214)
);

INVx4_ASAP7_75t_SL g231 ( 
.A(n_214),
.Y(n_231)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_102),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_L g216 ( 
.A1(n_77),
.A2(n_86),
.B1(n_83),
.B2(n_69),
.Y(n_216)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_84),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_218),
.B(n_219),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_109),
.B(n_118),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_87),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_220),
.B(n_225),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_113),
.B(n_37),
.Y(n_225)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_88),
.Y(n_229)
);

INVx2_ASAP7_75t_SL g302 ( 
.A(n_229),
.Y(n_302)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_226),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g369 ( 
.A(n_230),
.Y(n_369)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_233),
.Y(n_319)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_142),
.Y(n_235)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_235),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_228),
.A2(n_108),
.B1(n_101),
.B2(n_37),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g366 ( 
.A1(n_236),
.A2(n_251),
.B(n_283),
.Y(n_366)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_227),
.Y(n_237)
);

BUFx2_ASAP7_75t_L g331 ( 
.A(n_237),
.Y(n_331)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_211),
.Y(n_238)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_238),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_211),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g354 ( 
.A(n_239),
.Y(n_354)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_194),
.Y(n_240)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_240),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_SL g362 ( 
.A1(n_241),
.A2(n_250),
.B1(n_254),
.B2(n_262),
.Y(n_362)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_164),
.Y(n_242)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_242),
.Y(n_351)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_209),
.Y(n_243)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_243),
.Y(n_358)
);

OAI22xp33_ASAP7_75t_L g244 ( 
.A1(n_154),
.A2(n_40),
.B1(n_53),
.B2(n_45),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_244),
.A2(n_246),
.B1(n_295),
.B2(n_133),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_L g245 ( 
.A1(n_210),
.A2(n_53),
.B1(n_14),
.B2(n_13),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_245),
.A2(n_259),
.B1(n_285),
.B2(n_298),
.Y(n_327)
);

OAI22xp33_ASAP7_75t_L g246 ( 
.A1(n_151),
.A2(n_53),
.B1(n_98),
.B2(n_2),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_136),
.Y(n_247)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_247),
.Y(n_334)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_139),
.Y(n_249)
);

INVx3_ASAP7_75t_L g332 ( 
.A(n_249),
.Y(n_332)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_223),
.A2(n_98),
.B1(n_14),
.B2(n_13),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_224),
.A2(n_14),
.B1(n_13),
.B2(n_11),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_183),
.Y(n_252)
);

INVx3_ASAP7_75t_L g350 ( 
.A(n_252),
.Y(n_350)
);

CKINVDCx14_ASAP7_75t_R g253 ( 
.A(n_194),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_253),
.B(n_263),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_163),
.A2(n_11),
.B1(n_1),
.B2(n_2),
.Y(n_254)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_194),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_256),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_217),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_169),
.Y(n_260)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_260),
.Y(n_371)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_161),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_261),
.B(n_265),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_171),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_161),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_153),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_264),
.B(n_275),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_208),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_182),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_266),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_171),
.B(n_7),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_268),
.Y(n_329)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_176),
.Y(n_269)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_269),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_135),
.B(n_3),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_271),
.B(n_283),
.Y(n_316)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_193),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_273),
.Y(n_337)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_195),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_274),
.Y(n_355)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_179),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_144),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_277),
.B(n_280),
.Y(n_333)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_166),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_278),
.Y(n_361)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_149),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_279),
.Y(n_372)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_158),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_153),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_281),
.B(n_284),
.Y(n_335)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_173),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_282),
.B(n_287),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_137),
.B(n_3),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_L g285 ( 
.A1(n_184),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_285)
);

BUFx12f_ASAP7_75t_L g286 ( 
.A(n_191),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_286),
.B(n_288),
.Y(n_345)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_201),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_180),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_213),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_289),
.B(n_300),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_222),
.B(n_4),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_290),
.B(n_299),
.Y(n_317)
);

AND2x2_ASAP7_75t_SL g291 ( 
.A(n_167),
.B(n_4),
.Y(n_291)
);

MAJx2_ASAP7_75t_L g359 ( 
.A(n_291),
.B(n_296),
.C(n_168),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_187),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_292),
.B(n_293),
.Y(n_349)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_202),
.Y(n_293)
);

OAI22xp33_ASAP7_75t_L g295 ( 
.A1(n_150),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_295)
);

AND2x2_ASAP7_75t_SL g296 ( 
.A(n_201),
.B(n_6),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_188),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_297),
.B(n_301),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_216),
.A2(n_7),
.B1(n_190),
.B2(n_192),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_203),
.B(n_132),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_213),
.B(n_152),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_165),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g346 ( 
.A(n_304),
.B(n_271),
.Y(n_346)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_143),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_305),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_155),
.B(n_175),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_306),
.B(n_205),
.C(n_221),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_146),
.B(n_143),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_307),
.B(n_189),
.Y(n_341)
);

INVx4_ASAP7_75t_L g308 ( 
.A(n_143),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_308),
.Y(n_336)
);

AOI22xp33_ASAP7_75t_L g309 ( 
.A1(n_183),
.A2(n_190),
.B1(n_186),
.B2(n_192),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_309),
.A2(n_148),
.B1(n_162),
.B2(n_189),
.Y(n_360)
);

AOI22xp33_ASAP7_75t_SL g310 ( 
.A1(n_155),
.A2(n_134),
.B1(n_196),
.B2(n_200),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_310),
.A2(n_312),
.B1(n_314),
.B2(n_240),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_174),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_311),
.Y(n_365)
);

AOI22xp33_ASAP7_75t_SL g312 ( 
.A1(n_134),
.A2(n_196),
.B1(n_198),
.B2(n_165),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_198),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_313),
.B(n_289),
.Y(n_342)
);

INVx5_ASAP7_75t_L g314 ( 
.A(n_133),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_315),
.B(n_360),
.Y(n_396)
);

AOI22xp33_ASAP7_75t_L g325 ( 
.A1(n_242),
.A2(n_186),
.B1(n_170),
.B2(n_181),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_325),
.A2(n_330),
.B1(n_357),
.B2(n_363),
.Y(n_384)
);

AOI22xp33_ASAP7_75t_L g330 ( 
.A1(n_294),
.A2(n_140),
.B1(n_181),
.B2(n_170),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_299),
.A2(n_147),
.B(n_221),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g416 ( 
.A1(n_339),
.A2(n_364),
.B(n_237),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_255),
.B(n_140),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_340),
.B(n_374),
.C(n_375),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_341),
.B(n_329),
.Y(n_424)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_342),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_343),
.B(n_347),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_SL g381 ( 
.A(n_346),
.B(n_267),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_291),
.B(n_146),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_348),
.B(n_370),
.Y(n_400)
);

O2A1O1Ixp33_ASAP7_75t_L g353 ( 
.A1(n_311),
.A2(n_265),
.B(n_233),
.C(n_234),
.Y(n_353)
);

A2O1A1Ixp33_ASAP7_75t_SL g380 ( 
.A1(n_353),
.A2(n_300),
.B(n_287),
.C(n_277),
.Y(n_380)
);

AOI22xp33_ASAP7_75t_SL g379 ( 
.A1(n_356),
.A2(n_360),
.B1(n_256),
.B2(n_263),
.Y(n_379)
);

AOI22xp33_ASAP7_75t_L g357 ( 
.A1(n_294),
.A2(n_168),
.B1(n_205),
.B2(n_148),
.Y(n_357)
);

MAJx2_ASAP7_75t_L g402 ( 
.A(n_359),
.B(n_302),
.C(n_238),
.Y(n_402)
);

AOI22xp33_ASAP7_75t_L g363 ( 
.A1(n_258),
.A2(n_162),
.B1(n_189),
.B2(n_248),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_L g364 ( 
.A1(n_233),
.A2(n_259),
.B(n_257),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_366),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g367 ( 
.A1(n_248),
.A2(n_298),
.B1(n_236),
.B2(n_306),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_367),
.A2(n_376),
.B1(n_268),
.B2(n_284),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_295),
.A2(n_246),
.B1(n_303),
.B2(n_244),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_368),
.A2(n_232),
.B1(n_314),
.B2(n_302),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_291),
.B(n_296),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_290),
.B(n_276),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_235),
.B(n_260),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_296),
.A2(n_251),
.B1(n_307),
.B2(n_268),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_344),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_377),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_378),
.B(n_385),
.Y(n_453)
);

AOI22xp33_ASAP7_75t_SL g460 ( 
.A1(n_379),
.A2(n_380),
.B1(n_414),
.B2(n_336),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_381),
.B(n_404),
.Y(n_431)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_344),
.Y(n_382)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_382),
.Y(n_428)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_371),
.Y(n_383)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_383),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_L g385 ( 
.A1(n_319),
.A2(n_297),
.B(n_270),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_317),
.A2(n_230),
.B1(n_243),
.B2(n_292),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_386),
.A2(n_392),
.B1(n_396),
.B2(n_401),
.Y(n_426)
);

INVx3_ASAP7_75t_L g387 ( 
.A(n_323),
.Y(n_387)
);

INVx3_ASAP7_75t_L g437 ( 
.A(n_387),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_367),
.A2(n_317),
.B1(n_319),
.B2(n_339),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_388),
.A2(n_421),
.B1(n_315),
.B2(n_320),
.Y(n_440)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_371),
.Y(n_390)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_390),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_330),
.A2(n_232),
.B1(n_288),
.B2(n_274),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_326),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_393),
.B(n_405),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_SL g394 ( 
.A1(n_353),
.A2(n_300),
.B(n_264),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g439 ( 
.A1(n_394),
.A2(n_397),
.B(n_412),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_364),
.B(n_278),
.Y(n_395)
);

NAND3xp33_ASAP7_75t_L g448 ( 
.A(n_395),
.B(n_347),
.C(n_322),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_L g397 ( 
.A1(n_353),
.A2(n_270),
.B(n_282),
.Y(n_397)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_331),
.Y(n_399)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_399),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_402),
.B(n_423),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_340),
.B(n_269),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_403),
.B(n_413),
.C(n_419),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_SL g404 ( 
.A(n_335),
.B(n_273),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_326),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_365),
.A2(n_302),
.B1(n_261),
.B2(n_275),
.Y(n_406)
);

OA22x2_ASAP7_75t_L g456 ( 
.A1(n_406),
.A2(n_356),
.B1(n_380),
.B2(n_323),
.Y(n_456)
);

AOI21xp33_ASAP7_75t_L g407 ( 
.A1(n_370),
.A2(n_281),
.B(n_247),
.Y(n_407)
);

XOR2x1_ASAP7_75t_SL g444 ( 
.A(n_407),
.B(n_415),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_359),
.B(n_280),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_408),
.B(n_411),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_347),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_409),
.B(n_369),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_357),
.A2(n_249),
.B1(n_279),
.B2(n_252),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_410),
.A2(n_351),
.B1(n_327),
.B2(n_369),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_359),
.B(n_293),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_365),
.A2(n_308),
.B(n_305),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_343),
.B(n_272),
.C(n_301),
.Y(n_413)
);

AOI22xp33_ASAP7_75t_SL g414 ( 
.A1(n_320),
.A2(n_313),
.B1(n_231),
.B2(n_286),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_347),
.B(n_320),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_416),
.B(n_425),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_375),
.B(n_231),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_417),
.B(n_424),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_SL g418 ( 
.A1(n_320),
.A2(n_231),
.B(n_286),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g457 ( 
.A1(n_418),
.A2(n_322),
.B(n_345),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_374),
.B(n_252),
.C(n_286),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_333),
.Y(n_420)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_420),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_327),
.A2(n_351),
.B1(n_376),
.B2(n_368),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_333),
.Y(n_422)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_422),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_348),
.B(n_341),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_404),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_427),
.B(n_445),
.Y(n_490)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_430),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_421),
.A2(n_388),
.B1(n_396),
.B2(n_378),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g475 ( 
.A1(n_432),
.A2(n_454),
.B1(n_458),
.B2(n_466),
.Y(n_475)
);

AOI211xp5_ASAP7_75t_L g435 ( 
.A1(n_391),
.A2(n_346),
.B(n_335),
.C(n_366),
.Y(n_435)
);

OAI21xp33_ASAP7_75t_L g480 ( 
.A1(n_435),
.A2(n_448),
.B(n_452),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_398),
.B(n_316),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_436),
.B(n_442),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_440),
.A2(n_384),
.B1(n_420),
.B2(n_422),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_398),
.B(n_316),
.Y(n_442)
);

CKINVDCx16_ASAP7_75t_R g445 ( 
.A(n_386),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_403),
.B(n_423),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_450),
.B(n_451),
.C(n_463),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_408),
.B(n_352),
.C(n_342),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_396),
.A2(n_349),
.B1(n_352),
.B2(n_345),
.Y(n_454)
);

INVxp67_ASAP7_75t_L g484 ( 
.A(n_456),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_SL g469 ( 
.A1(n_457),
.A2(n_460),
.B(n_394),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_396),
.A2(n_349),
.B1(n_362),
.B2(n_369),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_382),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_461),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_411),
.B(n_338),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_383),
.Y(n_464)
);

CKINVDCx16_ASAP7_75t_R g489 ( 
.A(n_464),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_400),
.B(n_373),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_465),
.B(n_385),
.C(n_402),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_401),
.A2(n_373),
.B1(n_358),
.B2(n_350),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_SL g534 ( 
.A1(n_469),
.A2(n_470),
.B(n_471),
.Y(n_534)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_439),
.A2(n_397),
.B(n_416),
.Y(n_470)
);

OAI21xp5_ASAP7_75t_L g471 ( 
.A1(n_439),
.A2(n_394),
.B(n_380),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_438),
.Y(n_472)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_472),
.Y(n_512)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_438),
.Y(n_473)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_473),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_L g508 ( 
.A1(n_474),
.A2(n_481),
.B1(n_482),
.B2(n_492),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_459),
.B(n_425),
.Y(n_476)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_476),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_459),
.B(n_417),
.Y(n_477)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_477),
.Y(n_528)
);

OAI21xp5_ASAP7_75t_SL g478 ( 
.A1(n_453),
.A2(n_412),
.B(n_380),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_L g509 ( 
.A1(n_478),
.A2(n_495),
.B(n_497),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_462),
.B(n_389),
.Y(n_479)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_479),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_L g481 ( 
.A1(n_432),
.A2(n_384),
.B1(n_400),
.B2(n_413),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_L g482 ( 
.A1(n_426),
.A2(n_419),
.B1(n_380),
.B2(n_415),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_436),
.B(n_402),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g533 ( 
.A(n_485),
.B(n_483),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_431),
.B(n_381),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_486),
.B(n_494),
.Y(n_514)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_441),
.Y(n_487)
);

INVxp67_ASAP7_75t_L g523 ( 
.A(n_487),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g526 ( 
.A(n_491),
.B(n_444),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_440),
.A2(n_395),
.B1(n_424),
.B2(n_415),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_441),
.Y(n_493)
);

INVxp67_ASAP7_75t_L g527 ( 
.A(n_493),
.Y(n_527)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_428),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_453),
.A2(n_415),
.B1(n_380),
.B2(n_407),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_462),
.B(n_377),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_496),
.B(n_501),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_453),
.A2(n_392),
.B1(n_390),
.B2(n_410),
.Y(n_497)
);

A2O1A1Ixp33_ASAP7_75t_L g498 ( 
.A1(n_433),
.A2(n_418),
.B(n_338),
.C(n_336),
.Y(n_498)
);

OAI21xp5_ASAP7_75t_L g511 ( 
.A1(n_498),
.A2(n_502),
.B(n_505),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_426),
.A2(n_387),
.B1(n_350),
.B2(n_399),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_SL g542 ( 
.A1(n_499),
.A2(n_350),
.B1(n_332),
.B2(n_331),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_450),
.B(n_358),
.C(n_338),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_500),
.B(n_429),
.C(n_443),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_465),
.B(n_338),
.Y(n_501)
);

OAI21xp5_ASAP7_75t_L g502 ( 
.A1(n_454),
.A2(n_406),
.B(n_328),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_449),
.B(n_337),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_503),
.B(n_504),
.Y(n_519)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_434),
.Y(n_504)
);

OAI21xp5_ASAP7_75t_L g505 ( 
.A1(n_457),
.A2(n_328),
.B(n_361),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_506),
.B(n_507),
.C(n_526),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_483),
.B(n_429),
.C(n_443),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_496),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_510),
.B(n_530),
.Y(n_551)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_475),
.A2(n_458),
.B1(n_435),
.B2(n_446),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_L g555 ( 
.A1(n_516),
.A2(n_518),
.B1(n_524),
.B2(n_529),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_486),
.B(n_442),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_SL g564 ( 
.A(n_517),
.B(n_525),
.Y(n_564)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_475),
.A2(n_446),
.B1(n_430),
.B2(n_447),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_SL g520 ( 
.A(n_485),
.B(n_463),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_SL g547 ( 
.A(n_520),
.B(n_533),
.Y(n_547)
);

OAI21xp5_ASAP7_75t_L g521 ( 
.A1(n_470),
.A2(n_447),
.B(n_444),
.Y(n_521)
);

OAI21xp5_ASAP7_75t_SL g569 ( 
.A1(n_521),
.A2(n_473),
.B(n_472),
.Y(n_569)
);

AOI22xp5_ASAP7_75t_L g524 ( 
.A1(n_474),
.A2(n_466),
.B1(n_456),
.B2(n_451),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_489),
.B(n_324),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_L g529 ( 
.A1(n_481),
.A2(n_456),
.B1(n_434),
.B2(n_437),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g530 ( 
.A(n_479),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g531 ( 
.A(n_468),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_531),
.B(n_532),
.Y(n_546)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_468),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_476),
.B(n_455),
.Y(n_535)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_535),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_483),
.B(n_456),
.C(n_355),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_536),
.B(n_488),
.C(n_500),
.Y(n_553)
);

CKINVDCx16_ASAP7_75t_R g537 ( 
.A(n_490),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_537),
.B(n_489),
.Y(n_566)
);

XOR2x2_ASAP7_75t_L g538 ( 
.A(n_495),
.B(n_437),
.Y(n_538)
);

XNOR2x1_ASAP7_75t_L g570 ( 
.A(n_538),
.B(n_487),
.Y(n_570)
);

XOR2xp5_ASAP7_75t_L g539 ( 
.A(n_488),
.B(n_455),
.Y(n_539)
);

XOR2xp5_ASAP7_75t_L g552 ( 
.A(n_539),
.B(n_500),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g540 ( 
.A(n_503),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_540),
.B(n_477),
.Y(n_550)
);

AOI22xp5_ASAP7_75t_L g548 ( 
.A1(n_542),
.A2(n_467),
.B1(n_504),
.B2(n_494),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_SL g545 ( 
.A1(n_518),
.A2(n_484),
.B1(n_492),
.B2(n_490),
.Y(n_545)
);

AOI22xp5_ASAP7_75t_L g587 ( 
.A1(n_545),
.A2(n_560),
.B1(n_511),
.B2(n_541),
.Y(n_587)
);

OAI22xp5_ASAP7_75t_L g584 ( 
.A1(n_548),
.A2(n_557),
.B1(n_558),
.B2(n_562),
.Y(n_584)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_514),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_549),
.B(n_556),
.Y(n_583)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_550),
.Y(n_575)
);

XOR2xp5_ASAP7_75t_L g598 ( 
.A(n_552),
.B(n_565),
.Y(n_598)
);

XNOR2xp5_ASAP7_75t_L g577 ( 
.A(n_553),
.B(n_561),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_539),
.B(n_488),
.C(n_491),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_554),
.B(n_559),
.C(n_571),
.Y(n_574)
);

OAI21xp33_ASAP7_75t_SL g556 ( 
.A1(n_534),
.A2(n_469),
.B(n_478),
.Y(n_556)
);

CKINVDCx20_ASAP7_75t_R g557 ( 
.A(n_514),
.Y(n_557)
);

AOI22xp5_ASAP7_75t_L g558 ( 
.A1(n_529),
.A2(n_467),
.B1(n_482),
.B2(n_480),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_507),
.B(n_506),
.C(n_533),
.Y(n_559)
);

OAI22xp5_ASAP7_75t_SL g560 ( 
.A1(n_516),
.A2(n_497),
.B1(n_471),
.B2(n_502),
.Y(n_560)
);

XNOR2xp5_ASAP7_75t_L g561 ( 
.A(n_526),
.B(n_491),
.Y(n_561)
);

AOI22xp5_ASAP7_75t_L g562 ( 
.A1(n_508),
.A2(n_498),
.B1(n_505),
.B2(n_499),
.Y(n_562)
);

HB1xp67_ASAP7_75t_L g563 ( 
.A(n_519),
.Y(n_563)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_563),
.Y(n_578)
);

XOR2xp5_ASAP7_75t_L g565 ( 
.A(n_520),
.B(n_498),
.Y(n_565)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_566),
.Y(n_593)
);

XNOR2xp5_ASAP7_75t_L g567 ( 
.A(n_521),
.B(n_501),
.Y(n_567)
);

XNOR2xp5_ASAP7_75t_L g592 ( 
.A(n_567),
.B(n_568),
.Y(n_592)
);

XOR2xp5_ASAP7_75t_L g568 ( 
.A(n_536),
.B(n_493),
.Y(n_568)
);

XOR2xp5_ASAP7_75t_SL g588 ( 
.A(n_569),
.B(n_570),
.Y(n_588)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_528),
.B(n_354),
.C(n_321),
.Y(n_571)
);

XNOR2xp5_ASAP7_75t_L g572 ( 
.A(n_524),
.B(n_372),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g580 ( 
.A(n_572),
.B(n_523),
.C(n_527),
.Y(n_580)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_519),
.Y(n_573)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_573),
.Y(n_596)
);

AOI21xp5_ASAP7_75t_L g576 ( 
.A1(n_570),
.A2(n_534),
.B(n_511),
.Y(n_576)
);

INVxp33_ASAP7_75t_L g602 ( 
.A(n_576),
.Y(n_602)
);

AOI22xp5_ASAP7_75t_SL g579 ( 
.A1(n_560),
.A2(n_540),
.B1(n_530),
.B2(n_528),
.Y(n_579)
);

OAI22xp5_ASAP7_75t_SL g604 ( 
.A1(n_579),
.A2(n_587),
.B1(n_551),
.B2(n_548),
.Y(n_604)
);

XNOR2xp5_ASAP7_75t_L g600 ( 
.A(n_580),
.B(n_567),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_546),
.B(n_523),
.Y(n_581)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_581),
.Y(n_611)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_559),
.B(n_538),
.C(n_509),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_582),
.B(n_586),
.Y(n_615)
);

OAI22xp5_ASAP7_75t_SL g585 ( 
.A1(n_558),
.A2(n_522),
.B1(n_510),
.B2(n_541),
.Y(n_585)
);

AOI22xp5_ASAP7_75t_L g601 ( 
.A1(n_585),
.A2(n_544),
.B1(n_545),
.B2(n_562),
.Y(n_601)
);

MAJIxp5_ASAP7_75t_L g586 ( 
.A(n_554),
.B(n_538),
.C(n_509),
.Y(n_586)
);

CKINVDCx16_ASAP7_75t_R g589 ( 
.A(n_546),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_589),
.B(n_550),
.Y(n_603)
);

MAJIxp5_ASAP7_75t_L g590 ( 
.A(n_552),
.B(n_535),
.C(n_515),
.Y(n_590)
);

MAJIxp5_ASAP7_75t_L g610 ( 
.A(n_590),
.B(n_594),
.C(n_597),
.Y(n_610)
);

INVx1_ASAP7_75t_SL g591 ( 
.A(n_571),
.Y(n_591)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_591),
.Y(n_612)
);

MAJIxp5_ASAP7_75t_L g594 ( 
.A(n_543),
.B(n_553),
.C(n_568),
.Y(n_594)
);

OAI22xp5_ASAP7_75t_L g595 ( 
.A1(n_555),
.A2(n_522),
.B1(n_532),
.B2(n_531),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_595),
.B(n_542),
.Y(n_617)
);

MAJIxp5_ASAP7_75t_L g597 ( 
.A(n_543),
.B(n_515),
.C(n_527),
.Y(n_597)
);

XNOR2x1_ASAP7_75t_SL g599 ( 
.A(n_587),
.B(n_565),
.Y(n_599)
);

OAI21xp33_ASAP7_75t_SL g623 ( 
.A1(n_599),
.A2(n_617),
.B(n_601),
.Y(n_623)
);

HB1xp67_ASAP7_75t_L g619 ( 
.A(n_600),
.Y(n_619)
);

OAI22xp5_ASAP7_75t_SL g634 ( 
.A1(n_601),
.A2(n_588),
.B1(n_592),
.B2(n_323),
.Y(n_634)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_603),
.Y(n_621)
);

INVxp67_ASAP7_75t_L g620 ( 
.A(n_604),
.Y(n_620)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_581),
.Y(n_605)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_605),
.Y(n_627)
);

XOR2xp5_ASAP7_75t_L g606 ( 
.A(n_598),
.B(n_572),
.Y(n_606)
);

MAJIxp5_ASAP7_75t_L g628 ( 
.A(n_606),
.B(n_613),
.C(n_614),
.Y(n_628)
);

OAI22xp5_ASAP7_75t_SL g607 ( 
.A1(n_579),
.A2(n_569),
.B1(n_512),
.B2(n_513),
.Y(n_607)
);

AOI22xp5_ASAP7_75t_L g635 ( 
.A1(n_607),
.A2(n_592),
.B1(n_332),
.B2(n_354),
.Y(n_635)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_578),
.Y(n_608)
);

INVxp67_ASAP7_75t_SL g624 ( 
.A(n_608),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_597),
.B(n_564),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_SL g625 ( 
.A(n_609),
.B(n_616),
.Y(n_625)
);

MAJIxp5_ASAP7_75t_L g613 ( 
.A(n_594),
.B(n_561),
.C(n_547),
.Y(n_613)
);

MAJIxp5_ASAP7_75t_L g614 ( 
.A(n_574),
.B(n_547),
.C(n_513),
.Y(n_614)
);

XNOR2xp5_ASAP7_75t_L g616 ( 
.A(n_574),
.B(n_512),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_SL g618 ( 
.A(n_593),
.B(n_334),
.Y(n_618)
);

NOR2x1_ASAP7_75t_L g626 ( 
.A(n_618),
.B(n_596),
.Y(n_626)
);

AOI22xp5_ASAP7_75t_L g622 ( 
.A1(n_604),
.A2(n_585),
.B1(n_584),
.B2(n_575),
.Y(n_622)
);

OAI22xp5_ASAP7_75t_SL g642 ( 
.A1(n_622),
.A2(n_630),
.B1(n_633),
.B2(n_635),
.Y(n_642)
);

AOI22xp5_ASAP7_75t_L g640 ( 
.A1(n_623),
.A2(n_634),
.B1(n_602),
.B2(n_611),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_626),
.B(n_629),
.Y(n_646)
);

OAI21xp5_ASAP7_75t_SL g629 ( 
.A1(n_602),
.A2(n_583),
.B(n_576),
.Y(n_629)
);

AOI22xp5_ASAP7_75t_L g630 ( 
.A1(n_607),
.A2(n_591),
.B1(n_582),
.B2(n_586),
.Y(n_630)
);

MAJIxp5_ASAP7_75t_L g631 ( 
.A(n_616),
.B(n_577),
.C(n_590),
.Y(n_631)
);

MAJIxp5_ASAP7_75t_L g647 ( 
.A(n_631),
.B(n_632),
.C(n_332),
.Y(n_647)
);

MAJIxp5_ASAP7_75t_L g632 ( 
.A(n_610),
.B(n_577),
.C(n_598),
.Y(n_632)
);

FAx1_ASAP7_75t_SL g633 ( 
.A(n_599),
.B(n_588),
.CI(n_580),
.CON(n_633),
.SN(n_633)
);

NOR2xp67_ASAP7_75t_L g636 ( 
.A(n_621),
.B(n_610),
.Y(n_636)
);

OAI21x1_ASAP7_75t_L g656 ( 
.A1(n_636),
.A2(n_645),
.B(n_646),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_625),
.B(n_612),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_637),
.B(n_638),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_SL g638 ( 
.A(n_631),
.B(n_614),
.Y(n_638)
);

XOR2xp5_ASAP7_75t_L g639 ( 
.A(n_630),
.B(n_600),
.Y(n_639)
);

MAJIxp5_ASAP7_75t_L g653 ( 
.A(n_639),
.B(n_645),
.C(n_628),
.Y(n_653)
);

INVxp67_ASAP7_75t_SL g655 ( 
.A(n_640),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_SL g641 ( 
.A(n_628),
.B(n_615),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_641),
.B(n_643),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_620),
.B(n_608),
.Y(n_643)
);

OAI22xp5_ASAP7_75t_SL g644 ( 
.A1(n_620),
.A2(n_605),
.B1(n_617),
.B2(n_606),
.Y(n_644)
);

INVxp33_ASAP7_75t_L g649 ( 
.A(n_644),
.Y(n_649)
);

XOR2xp5_ASAP7_75t_L g645 ( 
.A(n_629),
.B(n_613),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_SL g650 ( 
.A(n_647),
.B(n_648),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_619),
.B(n_331),
.Y(n_648)
);

OAI21xp5_ASAP7_75t_SL g652 ( 
.A1(n_646),
.A2(n_622),
.B(n_627),
.Y(n_652)
);

OAI21xp5_ASAP7_75t_SL g659 ( 
.A1(n_652),
.A2(n_657),
.B(n_640),
.Y(n_659)
);

XOR2xp5_ASAP7_75t_L g663 ( 
.A(n_653),
.B(n_642),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_656),
.B(n_639),
.Y(n_660)
);

AOI21xp5_ASAP7_75t_L g657 ( 
.A1(n_647),
.A2(n_632),
.B(n_635),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_651),
.B(n_626),
.Y(n_658)
);

OAI21xp5_ASAP7_75t_L g665 ( 
.A1(n_658),
.A2(n_659),
.B(n_660),
.Y(n_665)
);

O2A1O1Ixp33_ASAP7_75t_SL g661 ( 
.A1(n_655),
.A2(n_633),
.B(n_642),
.C(n_624),
.Y(n_661)
);

OAI21xp5_ASAP7_75t_SL g664 ( 
.A1(n_661),
.A2(n_662),
.B(n_663),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_654),
.B(n_644),
.Y(n_662)
);

OAI21xp5_ASAP7_75t_SL g666 ( 
.A1(n_658),
.A2(n_649),
.B(n_655),
.Y(n_666)
);

AOI21xp5_ASAP7_75t_L g668 ( 
.A1(n_666),
.A2(n_633),
.B(n_318),
.Y(n_668)
);

MAJIxp5_ASAP7_75t_L g667 ( 
.A(n_665),
.B(n_634),
.C(n_650),
.Y(n_667)
);

MAJIxp5_ASAP7_75t_L g669 ( 
.A(n_667),
.B(n_668),
.C(n_664),
.Y(n_669)
);

BUFx24_ASAP7_75t_SL g670 ( 
.A(n_669),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_670),
.B(n_334),
.Y(n_671)
);

XNOR2xp5_ASAP7_75t_L g672 ( 
.A(n_671),
.B(n_318),
.Y(n_672)
);


endmodule