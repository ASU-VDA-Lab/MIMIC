module fake_jpeg_26843_n_134 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_134);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_134;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_7),
.B(n_6),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_28),
.B(n_17),
.Y(n_43)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_13),
.B(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_20),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

CKINVDCx6p67_ASAP7_75t_R g37 ( 
.A(n_32),
.Y(n_37)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_35),
.B(n_43),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_23),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_23),
.Y(n_50)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_26),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_25),
.C(n_22),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_32),
.Y(n_58)
);

A2O1A1Ixp33_ASAP7_75t_L g45 ( 
.A1(n_44),
.A2(n_31),
.B(n_14),
.C(n_12),
.Y(n_45)
);

A2O1A1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_45),
.A2(n_56),
.B(n_15),
.C(n_14),
.Y(n_71)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_47),
.Y(n_64)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_51),
.Y(n_67)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_52),
.Y(n_60)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_33),
.Y(n_62)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_27),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g56 ( 
.A1(n_36),
.A2(n_38),
.B(n_29),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_34),
.A2(n_24),
.B1(n_21),
.B2(n_20),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_18),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_32),
.Y(n_66)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_59),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_62),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_19),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_63),
.B(n_72),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_66),
.A2(n_71),
.B(n_74),
.Y(n_78)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_70),
.Y(n_87)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_38),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_19),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_36),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_73),
.A2(n_24),
.B1(n_21),
.B2(n_17),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_58),
.B(n_30),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_54),
.Y(n_89)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_76),
.A2(n_60),
.B(n_61),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_77),
.B(n_15),
.Y(n_94)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_79),
.B(n_80),
.Y(n_92)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_68),
.A2(n_33),
.B1(n_45),
.B2(n_40),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_82),
.A2(n_84),
.B1(n_69),
.B2(n_61),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_45),
.C(n_30),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_85),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_71),
.A2(n_33),
.B1(n_40),
.B2(n_49),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_67),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_66),
.A2(n_47),
.B1(n_46),
.B2(n_48),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_90),
.A2(n_75),
.B1(n_76),
.B2(n_74),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_91),
.A2(n_95),
.B1(n_102),
.B2(n_42),
.Y(n_107)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_85),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_94),
.Y(n_111)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_90),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_96),
.A2(n_98),
.B(n_99),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_78),
.A2(n_74),
.B(n_64),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_78),
.A2(n_64),
.B(n_67),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_100),
.B(n_101),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_83),
.A2(n_86),
.B1(n_81),
.B2(n_89),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_97),
.B(n_98),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_103),
.B(n_106),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_97),
.B(n_86),
.C(n_80),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_107),
.B(n_110),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_101),
.B(n_79),
.C(n_88),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_108),
.B(n_109),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_32),
.C(n_26),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_100),
.B(n_12),
.Y(n_110)
);

OA21x2_ASAP7_75t_L g113 ( 
.A1(n_105),
.A2(n_96),
.B(n_91),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_113),
.B(n_109),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_106),
.A2(n_99),
.B(n_92),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_114),
.B(n_116),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_104),
.A2(n_0),
.B(n_1),
.Y(n_116)
);

AOI221xp5_ASAP7_75t_L g118 ( 
.A1(n_111),
.A2(n_22),
.B1(n_10),
.B2(n_9),
.C(n_18),
.Y(n_118)
);

NOR2xp67_ASAP7_75t_SL g120 ( 
.A(n_118),
.B(n_10),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_119),
.B(n_120),
.Y(n_127)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_113),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_121),
.B(n_115),
.C(n_108),
.Y(n_124)
);

NAND2xp33_ASAP7_75t_SL g122 ( 
.A(n_112),
.B(n_103),
.Y(n_122)
);

MAJx2_ASAP7_75t_L g125 ( 
.A(n_122),
.B(n_117),
.C(n_22),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_124),
.B(n_126),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_125),
.B(n_122),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_123),
.B(n_53),
.C(n_52),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_128),
.B(n_51),
.C(n_2),
.Y(n_131)
);

AOI322xp5_ASAP7_75t_L g129 ( 
.A1(n_127),
.A2(n_51),
.A3(n_52),
.B1(n_2),
.B2(n_3),
.C1(n_4),
.C2(n_0),
.Y(n_129)
);

OAI21x1_ASAP7_75t_L g132 ( 
.A1(n_129),
.A2(n_1),
.B(n_3),
.Y(n_132)
);

OAI221xp5_ASAP7_75t_L g133 ( 
.A1(n_131),
.A2(n_132),
.B1(n_130),
.B2(n_6),
.C(n_7),
.Y(n_133)
);

AOI221xp5_ASAP7_75t_L g134 ( 
.A1(n_133),
.A2(n_3),
.B1(n_7),
.B2(n_8),
.C(n_128),
.Y(n_134)
);


endmodule