module fake_jpeg_31115_n_328 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_328);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_328;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx5_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx4f_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_2),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_26),
.B(n_28),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_45),
.B(n_53),
.Y(n_83)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_46),
.Y(n_102)
);

INVx6_ASAP7_75t_SL g47 ( 
.A(n_22),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_47),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_22),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_48),
.B(n_58),
.Y(n_74)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_26),
.B(n_18),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_51),
.B(n_37),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_21),
.B(n_15),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_52),
.B(n_56),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_28),
.B(n_0),
.Y(n_53)
);

BUFx10_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_54),
.Y(n_97)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_21),
.B(n_33),
.Y(n_56)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_65),
.Y(n_79)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_30),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

BUFx8_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

NAND3xp33_ASAP7_75t_L g65 ( 
.A(n_36),
.B(n_1),
.C(n_2),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_66),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_33),
.B(n_14),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_67),
.B(n_69),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_70),
.Y(n_105)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_71),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_47),
.A2(n_41),
.B1(n_38),
.B2(n_24),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_72),
.A2(n_81),
.B1(n_98),
.B2(n_101),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_75),
.B(n_96),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_51),
.B(n_37),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_80),
.B(n_92),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_66),
.A2(n_39),
.B1(n_32),
.B2(n_22),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_54),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_93),
.B(n_95),
.Y(n_128)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_61),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_70),
.B(n_36),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_55),
.A2(n_71),
.B1(n_63),
.B2(n_68),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_60),
.B(n_42),
.Y(n_100)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_100),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_63),
.A2(n_39),
.B1(n_25),
.B2(n_40),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_68),
.B(n_39),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_103),
.B(n_54),
.Y(n_125)
);

CKINVDCx12_ASAP7_75t_R g104 ( 
.A(n_64),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_104),
.Y(n_145)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_59),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_106),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_48),
.B(n_42),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_107),
.B(n_109),
.Y(n_151)
);

AND2x2_ASAP7_75t_SL g109 ( 
.A(n_50),
.B(n_1),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_62),
.A2(n_25),
.B1(n_38),
.B2(n_23),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_110),
.A2(n_40),
.B1(n_27),
.B2(n_29),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_54),
.Y(n_111)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_111),
.B(n_64),
.Y(n_132)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_44),
.Y(n_112)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_112),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_57),
.A2(n_25),
.B1(n_31),
.B2(n_29),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_113),
.A2(n_58),
.B1(n_2),
.B2(n_3),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_74),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_114),
.B(n_126),
.Y(n_154)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_87),
.Y(n_115)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_115),
.Y(n_183)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_99),
.Y(n_116)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_116),
.Y(n_152)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_87),
.Y(n_117)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_117),
.Y(n_153)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_73),
.Y(n_118)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_118),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_119),
.A2(n_123),
.B1(n_150),
.B2(n_142),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_72),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_120),
.B(n_121),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_113),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_76),
.A2(n_69),
.B1(n_20),
.B2(n_31),
.Y(n_123)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_78),
.Y(n_124)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_124),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_125),
.B(n_146),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_97),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_109),
.B(n_27),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_131),
.B(n_139),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_132),
.B(n_138),
.Y(n_170)
);

O2A1O1Ixp33_ASAP7_75t_L g135 ( 
.A1(n_103),
.A2(n_64),
.B(n_46),
.C(n_69),
.Y(n_135)
);

OR2x2_ASAP7_75t_L g175 ( 
.A(n_135),
.B(n_136),
.Y(n_175)
);

OR2x4_ASAP7_75t_L g136 ( 
.A(n_109),
.B(n_69),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_137),
.A2(n_82),
.B(n_10),
.Y(n_160)
);

A2O1A1Ixp33_ASAP7_75t_L g138 ( 
.A1(n_79),
.A2(n_83),
.B(n_94),
.C(n_85),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_99),
.B(n_1),
.Y(n_139)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_73),
.Y(n_140)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_140),
.Y(n_177)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_97),
.Y(n_141)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_141),
.Y(n_180)
);

O2A1O1Ixp33_ASAP7_75t_L g142 ( 
.A1(n_108),
.A2(n_58),
.B(n_5),
.C(n_6),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_142),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_77),
.A2(n_58),
.B1(n_5),
.B2(n_6),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_143),
.A2(n_144),
.B1(n_81),
.B2(n_108),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_77),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_105),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_105),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_147),
.B(n_90),
.Y(n_158)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_91),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_148),
.B(n_13),
.Y(n_173)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_78),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_149),
.A2(n_82),
.B1(n_102),
.B2(n_86),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_90),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_155),
.B(n_149),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_156),
.Y(n_187)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_158),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_121),
.A2(n_120),
.B1(n_125),
.B2(n_119),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_159),
.B(n_162),
.Y(n_185)
);

HAxp5_ASAP7_75t_SL g188 ( 
.A(n_160),
.B(n_167),
.CON(n_188),
.SN(n_188)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_130),
.A2(n_89),
.B1(n_88),
.B2(n_86),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_136),
.A2(n_85),
.B(n_88),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_163),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_151),
.A2(n_89),
.B1(n_91),
.B2(n_84),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_164),
.A2(n_181),
.B1(n_182),
.B2(n_148),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_151),
.B(n_102),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_165),
.B(n_171),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_139),
.B(n_102),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_166),
.B(n_172),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_131),
.A2(n_84),
.B(n_11),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_167),
.A2(n_115),
.B(n_117),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_127),
.B(n_9),
.C(n_12),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_133),
.B(n_12),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_173),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_132),
.A2(n_14),
.B1(n_135),
.B2(n_129),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_176),
.B(n_178),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_129),
.A2(n_14),
.B1(n_147),
.B2(n_146),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_134),
.B(n_128),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_179),
.B(n_138),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_122),
.A2(n_134),
.B1(n_116),
.B2(n_124),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_186),
.A2(n_188),
.B(n_157),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_190),
.A2(n_197),
.B1(n_206),
.B2(n_208),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_179),
.B(n_141),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_193),
.B(n_195),
.Y(n_227)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_152),
.Y(n_194)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_194),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_154),
.B(n_166),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_170),
.B(n_145),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_196),
.B(n_211),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_168),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_201),
.B(n_202),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_176),
.Y(n_202)
);

INVx13_ASAP7_75t_L g203 ( 
.A(n_183),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_203),
.Y(n_223)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_158),
.Y(n_204)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_204),
.Y(n_220)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_180),
.Y(n_205)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_205),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_178),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_206),
.Y(n_229)
);

INVx13_ASAP7_75t_L g207 ( 
.A(n_183),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_207),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_182),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_208),
.B(n_212),
.Y(n_234)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_180),
.Y(n_209)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_209),
.Y(n_230)
);

CKINVDCx11_ASAP7_75t_R g210 ( 
.A(n_184),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_210),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_163),
.B(n_118),
.Y(n_211)
);

INVxp67_ASAP7_75t_SL g213 ( 
.A(n_159),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_213),
.B(n_214),
.Y(n_237)
);

INVx13_ASAP7_75t_L g214 ( 
.A(n_153),
.Y(n_214)
);

INVx13_ASAP7_75t_L g215 ( 
.A(n_153),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_215),
.B(n_194),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_211),
.A2(n_175),
.B(n_161),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_216),
.A2(n_217),
.B(n_225),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_187),
.A2(n_175),
.B(n_161),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_185),
.A2(n_160),
.B1(n_161),
.B2(n_162),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_218),
.B(n_221),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_185),
.A2(n_157),
.B1(n_155),
.B2(n_164),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_198),
.B(n_165),
.C(n_172),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_226),
.B(n_236),
.C(n_192),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_186),
.A2(n_171),
.B(n_169),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_228),
.A2(n_238),
.B(n_191),
.Y(n_254)
);

OAI32xp33_ASAP7_75t_L g233 ( 
.A1(n_213),
.A2(n_174),
.A3(n_169),
.B1(n_177),
.B2(n_152),
.Y(n_233)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_233),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_198),
.B(n_177),
.C(n_174),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_186),
.A2(n_140),
.B(n_189),
.Y(n_238)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_239),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_200),
.A2(n_188),
.B(n_197),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_240),
.B(n_202),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_241),
.B(n_190),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_220),
.B(n_193),
.Y(n_243)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_243),
.Y(n_264)
);

XNOR2x1_ASAP7_75t_L g244 ( 
.A(n_236),
.B(n_192),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_244),
.B(n_217),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_245),
.A2(n_254),
.B(n_255),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_220),
.B(n_227),
.Y(n_246)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_246),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_247),
.B(n_249),
.C(n_258),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_236),
.B(n_195),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_224),
.Y(n_250)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_250),
.Y(n_270)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_224),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_251),
.Y(n_274)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_230),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_253),
.B(n_256),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_231),
.B(n_212),
.Y(n_256)
);

OA21x2_ASAP7_75t_SL g257 ( 
.A1(n_232),
.A2(n_210),
.B(n_200),
.Y(n_257)
);

NOR3xp33_ASAP7_75t_SL g276 ( 
.A(n_257),
.B(n_238),
.C(n_237),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_226),
.B(n_225),
.C(n_216),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_238),
.A2(n_191),
.B(n_204),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_259),
.A2(n_228),
.B(n_234),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_226),
.B(n_196),
.C(n_209),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_261),
.B(n_232),
.C(n_231),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_234),
.B(n_227),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_262),
.B(n_263),
.Y(n_279)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_230),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_265),
.B(n_277),
.Y(n_286)
);

INVxp67_ASAP7_75t_SL g266 ( 
.A(n_262),
.Y(n_266)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_266),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_271),
.A2(n_248),
.B(n_241),
.Y(n_293)
);

INVxp33_ASAP7_75t_L g272 ( 
.A(n_255),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_272),
.A2(n_259),
.B(n_254),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_275),
.B(n_273),
.C(n_277),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_276),
.B(n_278),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_244),
.B(n_240),
.Y(n_277)
);

NOR3xp33_ASAP7_75t_SL g278 ( 
.A(n_257),
.B(n_199),
.C(n_235),
.Y(n_278)
);

MAJx2_ASAP7_75t_L g280 ( 
.A(n_258),
.B(n_237),
.C(n_218),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_280),
.B(n_249),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_280),
.B(n_247),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_282),
.B(n_283),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_264),
.A2(n_242),
.B1(n_229),
.B2(n_248),
.Y(n_283)
);

MAJx2_ASAP7_75t_L g284 ( 
.A(n_273),
.B(n_260),
.C(n_261),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_284),
.B(n_287),
.Y(n_303)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_285),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_278),
.A2(n_252),
.B(n_246),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_288),
.B(n_289),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_267),
.A2(n_260),
.B(n_242),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_269),
.A2(n_252),
.B(n_243),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_290),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_291),
.B(n_292),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_268),
.B(n_229),
.Y(n_292)
);

A2O1A1Ixp33_ASAP7_75t_SL g297 ( 
.A1(n_293),
.A2(n_276),
.B(n_272),
.C(n_221),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_291),
.B(n_275),
.C(n_267),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_295),
.B(n_301),
.Y(n_307)
);

OAI21x1_ASAP7_75t_L g306 ( 
.A1(n_297),
.A2(n_289),
.B(n_283),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_282),
.B(n_284),
.C(n_287),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_286),
.B(n_265),
.C(n_274),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_304),
.B(n_286),
.C(n_239),
.Y(n_311)
);

AO22x1_ASAP7_75t_L g305 ( 
.A1(n_293),
.A2(n_279),
.B1(n_233),
.B2(n_274),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_305),
.A2(n_223),
.B(n_205),
.Y(n_313)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_306),
.Y(n_316)
);

AOI322xp5_ASAP7_75t_L g308 ( 
.A1(n_302),
.A2(n_281),
.A3(n_294),
.B1(n_270),
.B2(n_253),
.C1(n_263),
.C2(n_251),
.Y(n_308)
);

XOR2x2_ASAP7_75t_L g314 ( 
.A(n_308),
.B(n_310),
.Y(n_314)
);

BUFx24_ASAP7_75t_SL g309 ( 
.A(n_299),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_309),
.Y(n_317)
);

AOI322xp5_ASAP7_75t_L g310 ( 
.A1(n_300),
.A2(n_305),
.A3(n_298),
.B1(n_297),
.B2(n_250),
.C1(n_296),
.C2(n_223),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_311),
.B(n_296),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_303),
.A2(n_222),
.B(n_219),
.Y(n_312)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_312),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_313),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_315),
.B(n_297),
.Y(n_322)
);

HB1xp67_ASAP7_75t_L g318 ( 
.A(n_307),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_316),
.A2(n_297),
.B1(n_303),
.B2(n_219),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_321),
.A2(n_324),
.B1(n_214),
.B2(n_215),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_322),
.B(n_323),
.C(n_203),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_314),
.B(n_214),
.C(n_215),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_L g324 ( 
.A1(n_320),
.A2(n_319),
.B1(n_318),
.B2(n_317),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_325),
.B(n_326),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_323),
.Y(n_328)
);


endmodule