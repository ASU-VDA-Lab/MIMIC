module fake_jpeg_27664_n_295 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_295);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_295;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

INVx3_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx2_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_17),
.B(n_21),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_36),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_18),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx2_ASAP7_75t_SL g39 ( 
.A(n_27),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g46 ( 
.A(n_39),
.Y(n_46)
);

INVx6_ASAP7_75t_SL g40 ( 
.A(n_17),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_26),
.B(n_8),
.Y(n_42)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_42),
.B(n_26),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_61),
.Y(n_69)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_39),
.A2(n_26),
.B1(n_16),
.B2(n_30),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_47),
.A2(n_48),
.B1(n_54),
.B2(n_59),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_39),
.A2(n_16),
.B1(n_26),
.B2(n_30),
.Y(n_48)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_52),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_39),
.A2(n_16),
.B1(n_32),
.B2(n_28),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_39),
.A2(n_18),
.B1(n_32),
.B2(n_28),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_19),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_36),
.B(n_19),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_62),
.B(n_36),
.Y(n_71)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_65),
.A2(n_31),
.B1(n_24),
.B2(n_29),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_67),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_71),
.B(n_83),
.Y(n_107)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_43),
.A2(n_35),
.B1(n_39),
.B2(n_38),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_73),
.A2(n_80),
.B1(n_46),
.B2(n_77),
.Y(n_95)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_74),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_35),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_77),
.B(n_70),
.C(n_68),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_58),
.A2(n_39),
.B1(n_35),
.B2(n_34),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_78),
.A2(n_52),
.B1(n_57),
.B2(n_45),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_50),
.A2(n_34),
.B1(n_37),
.B2(n_25),
.Y(n_80)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_56),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_50),
.B(n_42),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_41),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_51),
.B(n_21),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_85),
.B(n_89),
.Y(n_91)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_86),
.Y(n_101)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_63),
.B(n_60),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_72),
.B(n_60),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_92),
.B(n_115),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_95),
.A2(n_111),
.B1(n_90),
.B2(n_40),
.Y(n_136)
);

AOI21xp33_ASAP7_75t_L g96 ( 
.A1(n_69),
.A2(n_24),
.B(n_31),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_96),
.A2(n_20),
.B(n_25),
.Y(n_142)
);

OAI32xp33_ASAP7_75t_L g97 ( 
.A1(n_76),
.A2(n_34),
.A3(n_33),
.B1(n_29),
.B2(n_58),
.Y(n_97)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_97),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_86),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_109),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_99),
.B(n_114),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_89),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_100),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_67),
.B(n_21),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_105),
.B(n_33),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_73),
.A2(n_46),
.B1(n_49),
.B2(n_34),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_106),
.A2(n_79),
.B1(n_90),
.B2(n_75),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_85),
.A2(n_46),
.B1(n_37),
.B2(n_55),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_108),
.A2(n_68),
.B1(n_70),
.B2(n_79),
.Y(n_129)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_81),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_66),
.Y(n_110)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_110),
.Y(n_122)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_66),
.Y(n_112)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_112),
.Y(n_128)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_81),
.Y(n_113)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_113),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_80),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_77),
.B(n_60),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_116),
.B(n_21),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_117),
.B(n_127),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_120),
.A2(n_125),
.B(n_139),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_121),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g124 ( 
.A(n_116),
.B(n_60),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_124),
.B(n_138),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_104),
.A2(n_87),
.B(n_82),
.Y(n_125)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_109),
.Y(n_126)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_126),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_107),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_129),
.A2(n_106),
.B1(n_95),
.B2(n_93),
.Y(n_146)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_108),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_132),
.B(n_135),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_133),
.A2(n_136),
.B1(n_141),
.B2(n_103),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_100),
.B(n_81),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_91),
.B(n_81),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_137),
.B(n_140),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_115),
.B(n_92),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_104),
.A2(n_33),
.B(n_29),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_91),
.B(n_74),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_114),
.A2(n_88),
.B1(n_75),
.B2(n_40),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_142),
.B(n_139),
.Y(n_145)
);

O2A1O1Ixp33_ASAP7_75t_L g143 ( 
.A1(n_97),
.A2(n_20),
.B(n_40),
.C(n_25),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_143),
.A2(n_23),
.B(n_27),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_144),
.B(n_145),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_146),
.A2(n_165),
.B1(n_170),
.B2(n_120),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_125),
.A2(n_118),
.B(n_134),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_148),
.Y(n_173)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_135),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_150),
.B(n_153),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_124),
.B(n_93),
.C(n_94),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_151),
.B(n_157),
.Y(n_197)
);

A2O1A1Ixp33_ASAP7_75t_SL g152 ( 
.A1(n_131),
.A2(n_102),
.B(n_94),
.C(n_103),
.Y(n_152)
);

AO21x2_ASAP7_75t_L g179 ( 
.A1(n_152),
.A2(n_168),
.B(n_128),
.Y(n_179)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_119),
.Y(n_153)
);

OA21x2_ASAP7_75t_L g155 ( 
.A1(n_118),
.A2(n_102),
.B(n_101),
.Y(n_155)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_155),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_131),
.A2(n_101),
.B(n_113),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_156),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_138),
.B(n_112),
.C(n_110),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_126),
.A2(n_88),
.B1(n_23),
.B2(n_2),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_158),
.B(n_159),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_132),
.A2(n_0),
.B(n_1),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_140),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_160),
.B(n_161),
.Y(n_186)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_137),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_162),
.B(n_167),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_143),
.A2(n_23),
.B(n_22),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_163),
.B(n_122),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_133),
.A2(n_27),
.B1(n_22),
.B2(n_10),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_129),
.B(n_22),
.Y(n_166)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_166),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_141),
.Y(n_167)
);

AOI22x1_ASAP7_75t_L g168 ( 
.A1(n_123),
.A2(n_27),
.B1(n_1),
.B2(n_2),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_127),
.A2(n_123),
.B1(n_142),
.B2(n_120),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_175),
.A2(n_179),
.B1(n_167),
.B2(n_144),
.Y(n_206)
);

FAx1_ASAP7_75t_SL g178 ( 
.A(n_151),
.B(n_130),
.CI(n_128),
.CON(n_178),
.SN(n_178)
);

FAx1_ASAP7_75t_SL g202 ( 
.A(n_178),
.B(n_154),
.CI(n_155),
.CON(n_202),
.SN(n_202)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_164),
.B(n_130),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_180),
.B(n_184),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_183),
.A2(n_166),
.B(n_163),
.Y(n_209)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_169),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_156),
.Y(n_185)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_185),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_172),
.B(n_169),
.Y(n_188)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_188),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_147),
.Y(n_189)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_189),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_159),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_R g200 ( 
.A(n_190),
.B(n_168),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_147),
.B(n_122),
.Y(n_191)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_191),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_149),
.B(n_7),
.Y(n_193)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_193),
.Y(n_217)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_155),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_194),
.A2(n_195),
.B1(n_196),
.B2(n_165),
.Y(n_212)
);

INVx8_ASAP7_75t_L g195 ( 
.A(n_168),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_148),
.B(n_0),
.Y(n_196)
);

XOR2x2_ASAP7_75t_L g198 ( 
.A(n_171),
.B(n_7),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_198),
.B(n_5),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_200),
.A2(n_209),
.B(n_219),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_197),
.B(n_157),
.C(n_171),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_201),
.B(n_203),
.C(n_204),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_202),
.B(n_220),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_197),
.B(n_178),
.C(n_184),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_178),
.B(n_154),
.C(n_166),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_206),
.A2(n_179),
.B1(n_194),
.B2(n_192),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_175),
.B(n_198),
.C(n_181),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_207),
.B(n_214),
.C(n_215),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_177),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_210),
.B(n_186),
.Y(n_223)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_212),
.Y(n_226)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_179),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_213),
.B(n_192),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_181),
.B(n_152),
.C(n_162),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_188),
.B(n_152),
.C(n_8),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_176),
.A2(n_152),
.B1(n_8),
.B2(n_11),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_216),
.A2(n_195),
.B1(n_179),
.B2(n_176),
.Y(n_225)
);

AOI21xp33_ASAP7_75t_L g219 ( 
.A1(n_173),
.A2(n_196),
.B(n_187),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_174),
.B(n_5),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_221),
.B(n_183),
.Y(n_231)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_223),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_225),
.B(n_227),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_218),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_202),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_228),
.B(n_229),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_199),
.A2(n_182),
.B(n_173),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_230),
.B(n_233),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_231),
.B(n_204),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_213),
.A2(n_190),
.B1(n_182),
.B2(n_179),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_232),
.A2(n_225),
.B1(n_226),
.B2(n_200),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_205),
.B(n_192),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_234),
.B(n_236),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_210),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_217),
.B(n_11),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_237),
.B(n_239),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_215),
.B(n_15),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_214),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_240),
.B(n_201),
.Y(n_252)
);

BUFx2_ASAP7_75t_L g241 ( 
.A(n_227),
.Y(n_241)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_241),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_243),
.A2(n_251),
.B1(n_235),
.B2(n_12),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_244),
.B(n_224),
.Y(n_255)
);

NAND3xp33_ASAP7_75t_L g250 ( 
.A(n_223),
.B(n_221),
.C(n_203),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_250),
.B(n_252),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_232),
.A2(n_211),
.B1(n_207),
.B2(n_208),
.Y(n_251)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_229),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_253),
.B(n_233),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_224),
.B(n_209),
.C(n_220),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_254),
.B(n_222),
.C(n_231),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_255),
.B(n_261),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_251),
.B(n_222),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_257),
.B(n_263),
.Y(n_270)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_259),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_246),
.A2(n_238),
.B1(n_242),
.B2(n_243),
.Y(n_260)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_260),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_253),
.A2(n_238),
.B(n_230),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_262),
.B(n_241),
.C(n_4),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_247),
.A2(n_235),
.B(n_12),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_264),
.B(n_265),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_249),
.A2(n_245),
.B(n_248),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_254),
.B(n_4),
.C(n_14),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_266),
.B(n_4),
.C(n_13),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_256),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_267),
.B(n_258),
.Y(n_280)
);

NOR2xp67_ASAP7_75t_SL g269 ( 
.A(n_257),
.B(n_244),
.Y(n_269)
);

OAI21x1_ASAP7_75t_SL g278 ( 
.A1(n_269),
.A2(n_274),
.B(n_263),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_271),
.B(n_266),
.Y(n_277)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_272),
.Y(n_283)
);

NOR2xp67_ASAP7_75t_L g274 ( 
.A(n_262),
.B(n_3),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_277),
.B(n_279),
.Y(n_285)
);

AOI21x1_ASAP7_75t_L g287 ( 
.A1(n_278),
.A2(n_273),
.B(n_275),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_272),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_280),
.B(n_281),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_270),
.A2(n_261),
.B1(n_255),
.B2(n_13),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_268),
.B(n_12),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_282),
.B(n_13),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_283),
.A2(n_267),
.B(n_276),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_284),
.Y(n_289)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g290 ( 
.A1(n_287),
.A2(n_288),
.B(n_279),
.C(n_275),
.D(n_15),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_290),
.B(n_286),
.Y(n_291)
);

AOI21x1_ASAP7_75t_SL g292 ( 
.A1(n_291),
.A2(n_289),
.B(n_285),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_292),
.A2(n_15),
.B(n_1),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_293),
.B(n_0),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_294),
.B(n_2),
.Y(n_295)
);


endmodule