module fake_netlist_1_9044_n_48 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_14, n_7, n_15, n_10, n_8, n_0, n_48);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_14;
input n_7;
input n_15;
input n_10;
input n_8;
input n_0;
output n_48;
wire n_45;
wire n_20;
wire n_38;
wire n_44;
wire n_36;
wire n_47;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_46;
wire n_25;
wire n_30;
wire n_26;
wire n_16;
wire n_33;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_17;
wire n_42;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_43;
wire n_40;
wire n_27;
wire n_39;
BUFx6f_ASAP7_75t_L g16 ( .A(n_5), .Y(n_16) );
AND2x2_ASAP7_75t_SL g17 ( .A(n_5), .B(n_7), .Y(n_17) );
INVx2_ASAP7_75t_SL g18 ( .A(n_13), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_9), .Y(n_19) );
NAND2xp5_ASAP7_75t_L g20 ( .A(n_2), .B(n_14), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_1), .Y(n_21) );
INVx2_ASAP7_75t_L g22 ( .A(n_2), .Y(n_22) );
NAND2x1_ASAP7_75t_L g23 ( .A(n_11), .B(n_15), .Y(n_23) );
INVx2_ASAP7_75t_SL g24 ( .A(n_18), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_19), .Y(n_25) );
NAND2xp5_ASAP7_75t_SL g26 ( .A(n_18), .B(n_0), .Y(n_26) );
NAND2xp5_ASAP7_75t_L g27 ( .A(n_21), .B(n_0), .Y(n_27) );
OAI21xp5_ASAP7_75t_L g28 ( .A1(n_25), .A2(n_19), .B(n_23), .Y(n_28) );
AO31x2_ASAP7_75t_L g29 ( .A1(n_25), .A2(n_22), .A3(n_20), .B(n_17), .Y(n_29) );
INVx1_ASAP7_75t_L g30 ( .A(n_27), .Y(n_30) );
AOI221xp5_ASAP7_75t_L g31 ( .A1(n_30), .A2(n_27), .B1(n_26), .B2(n_24), .C(n_22), .Y(n_31) );
AND2x2_ASAP7_75t_L g32 ( .A(n_30), .B(n_17), .Y(n_32) );
INVx4_ASAP7_75t_L g33 ( .A(n_32), .Y(n_33) );
AND2x2_ASAP7_75t_L g34 ( .A(n_31), .B(n_29), .Y(n_34) );
AOI221xp5_ASAP7_75t_L g35 ( .A1(n_34), .A2(n_28), .B1(n_24), .B2(n_16), .C(n_29), .Y(n_35) );
HB1xp67_ASAP7_75t_L g36 ( .A(n_33), .Y(n_36) );
A2O1A1Ixp33_ASAP7_75t_L g37 ( .A1(n_34), .A2(n_23), .B(n_16), .C(n_29), .Y(n_37) );
AOI21xp5_ASAP7_75t_L g38 ( .A1(n_37), .A2(n_33), .B(n_16), .Y(n_38) );
AOI221xp5_ASAP7_75t_L g39 ( .A1(n_35), .A2(n_33), .B1(n_16), .B2(n_29), .C(n_6), .Y(n_39) );
AOI321xp33_ASAP7_75t_L g40 ( .A1(n_36), .A2(n_29), .A3(n_3), .B1(n_4), .B2(n_6), .C(n_7), .Y(n_40) );
OR5x1_ASAP7_75t_L g41 ( .A(n_40), .B(n_1), .C(n_3), .D(n_4), .E(n_8), .Y(n_41) );
NAND4xp25_ASAP7_75t_L g42 ( .A(n_39), .B(n_29), .C(n_8), .D(n_16), .Y(n_42) );
AND2x2_ASAP7_75t_L g43 ( .A(n_38), .B(n_10), .Y(n_43) );
INVx1_ASAP7_75t_L g44 ( .A(n_43), .Y(n_44) );
INVx1_ASAP7_75t_L g45 ( .A(n_42), .Y(n_45) );
OAI21x1_ASAP7_75t_L g46 ( .A1(n_41), .A2(n_12), .B(n_38), .Y(n_46) );
OAI21x1_ASAP7_75t_L g47 ( .A1(n_46), .A2(n_44), .B(n_45), .Y(n_47) );
OAI21xp5_ASAP7_75t_L g48 ( .A1(n_47), .A2(n_46), .B(n_44), .Y(n_48) );
endmodule