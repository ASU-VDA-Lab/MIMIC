module fake_netlist_1_5562_n_491 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_491);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_491;
wire n_117;
wire n_361;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_73;
wire n_119;
wire n_141;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_312;
wire n_455;
wire n_137;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_390;
wire n_120;
wire n_486;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_283;
wire n_76;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_458;
wire n_418;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g73 ( .A(n_70), .Y(n_73) );
CKINVDCx20_ASAP7_75t_R g74 ( .A(n_65), .Y(n_74) );
CKINVDCx16_ASAP7_75t_R g75 ( .A(n_46), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_59), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_43), .Y(n_77) );
INVxp33_ASAP7_75t_L g78 ( .A(n_67), .Y(n_78) );
INVx1_ASAP7_75t_SL g79 ( .A(n_12), .Y(n_79) );
CKINVDCx5p33_ASAP7_75t_R g80 ( .A(n_26), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_31), .Y(n_81) );
INVxp33_ASAP7_75t_L g82 ( .A(n_4), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_21), .Y(n_83) );
CKINVDCx20_ASAP7_75t_R g84 ( .A(n_27), .Y(n_84) );
INVx2_ASAP7_75t_L g85 ( .A(n_37), .Y(n_85) );
INVxp67_ASAP7_75t_SL g86 ( .A(n_19), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_63), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_62), .Y(n_88) );
BUFx6f_ASAP7_75t_L g89 ( .A(n_21), .Y(n_89) );
BUFx3_ASAP7_75t_L g90 ( .A(n_15), .Y(n_90) );
CKINVDCx14_ASAP7_75t_R g91 ( .A(n_35), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_45), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_52), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_44), .Y(n_94) );
CKINVDCx20_ASAP7_75t_R g95 ( .A(n_68), .Y(n_95) );
CKINVDCx20_ASAP7_75t_R g96 ( .A(n_5), .Y(n_96) );
INVxp33_ASAP7_75t_L g97 ( .A(n_16), .Y(n_97) );
INVxp33_ASAP7_75t_SL g98 ( .A(n_55), .Y(n_98) );
INVxp33_ASAP7_75t_L g99 ( .A(n_17), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_47), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_49), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_3), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_15), .Y(n_103) );
INVx2_ASAP7_75t_L g104 ( .A(n_14), .Y(n_104) );
BUFx5_ASAP7_75t_L g105 ( .A(n_39), .Y(n_105) );
BUFx2_ASAP7_75t_L g106 ( .A(n_90), .Y(n_106) );
INVx2_ASAP7_75t_L g107 ( .A(n_105), .Y(n_107) );
AND2x4_ASAP7_75t_L g108 ( .A(n_104), .B(n_0), .Y(n_108) );
INVx3_ASAP7_75t_L g109 ( .A(n_85), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_75), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g111 ( .A(n_96), .Y(n_111) );
AND2x2_ASAP7_75t_L g112 ( .A(n_82), .B(n_0), .Y(n_112) );
INVx3_ASAP7_75t_L g113 ( .A(n_85), .Y(n_113) );
BUFx3_ASAP7_75t_L g114 ( .A(n_105), .Y(n_114) );
AND2x4_ASAP7_75t_L g115 ( .A(n_104), .B(n_1), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_76), .Y(n_116) );
BUFx6f_ASAP7_75t_L g117 ( .A(n_89), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_75), .Y(n_118) );
BUFx2_ASAP7_75t_L g119 ( .A(n_90), .Y(n_119) );
NAND2xp33_ASAP7_75t_L g120 ( .A(n_105), .B(n_30), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_76), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_77), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_74), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_84), .Y(n_124) );
HB1xp67_ASAP7_75t_L g125 ( .A(n_83), .Y(n_125) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_89), .Y(n_126) );
HB1xp67_ASAP7_75t_L g127 ( .A(n_83), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_102), .B(n_1), .Y(n_128) );
BUFx3_ASAP7_75t_L g129 ( .A(n_106), .Y(n_129) );
NAND2xp5_ASAP7_75t_SL g130 ( .A(n_118), .B(n_78), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_106), .B(n_77), .Y(n_131) );
INVx4_ASAP7_75t_L g132 ( .A(n_114), .Y(n_132) );
NOR3xp33_ASAP7_75t_L g133 ( .A(n_128), .B(n_86), .C(n_102), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_107), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_117), .Y(n_135) );
INVx3_ASAP7_75t_L g136 ( .A(n_108), .Y(n_136) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_117), .Y(n_137) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_117), .Y(n_138) );
NOR2xp33_ASAP7_75t_L g139 ( .A(n_106), .B(n_81), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_107), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_117), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_107), .Y(n_142) );
NAND2xp5_ASAP7_75t_SL g143 ( .A(n_118), .B(n_73), .Y(n_143) );
INVx2_ASAP7_75t_SL g144 ( .A(n_114), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_119), .B(n_81), .Y(n_145) );
BUFx2_ASAP7_75t_L g146 ( .A(n_110), .Y(n_146) );
NAND3x1_ASAP7_75t_L g147 ( .A(n_128), .B(n_112), .C(n_116), .Y(n_147) );
NOR2xp33_ASAP7_75t_L g148 ( .A(n_119), .B(n_87), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_107), .Y(n_149) );
INVx4_ASAP7_75t_L g150 ( .A(n_114), .Y(n_150) );
INVx1_ASAP7_75t_SL g151 ( .A(n_119), .Y(n_151) );
OR2x6_ASAP7_75t_L g152 ( .A(n_108), .B(n_103), .Y(n_152) );
INVx2_ASAP7_75t_SL g153 ( .A(n_114), .Y(n_153) );
BUFx8_ASAP7_75t_L g154 ( .A(n_146), .Y(n_154) );
NAND2x1p5_ASAP7_75t_L g155 ( .A(n_136), .B(n_108), .Y(n_155) );
NAND2xp33_ASAP7_75t_SL g156 ( .A(n_146), .B(n_95), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_136), .Y(n_157) );
NOR3xp33_ASAP7_75t_SL g158 ( .A(n_130), .B(n_124), .C(n_80), .Y(n_158) );
CKINVDCx5p33_ASAP7_75t_R g159 ( .A(n_151), .Y(n_159) );
BUFx2_ASAP7_75t_L g160 ( .A(n_129), .Y(n_160) );
CKINVDCx5p33_ASAP7_75t_R g161 ( .A(n_151), .Y(n_161) );
CKINVDCx20_ASAP7_75t_R g162 ( .A(n_129), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_129), .B(n_116), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_143), .B(n_125), .Y(n_164) );
BUFx3_ASAP7_75t_L g165 ( .A(n_152), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_139), .B(n_121), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_136), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_139), .B(n_121), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_134), .Y(n_169) );
CKINVDCx5p33_ASAP7_75t_R g170 ( .A(n_152), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_148), .B(n_121), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_134), .Y(n_172) );
NOR2xp67_ASAP7_75t_L g173 ( .A(n_136), .B(n_122), .Y(n_173) );
CKINVDCx5p33_ASAP7_75t_R g174 ( .A(n_152), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_140), .Y(n_175) );
NOR3xp33_ASAP7_75t_SL g176 ( .A(n_148), .B(n_103), .C(n_100), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_140), .Y(n_177) );
BUFx2_ASAP7_75t_L g178 ( .A(n_152), .Y(n_178) );
BUFx3_ASAP7_75t_L g179 ( .A(n_152), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_152), .Y(n_180) );
CKINVDCx5p33_ASAP7_75t_R g181 ( .A(n_131), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_147), .B(n_122), .Y(n_182) );
BUFx4f_ASAP7_75t_L g183 ( .A(n_142), .Y(n_183) );
HB1xp67_ASAP7_75t_L g184 ( .A(n_147), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_142), .Y(n_185) );
AND2x4_ASAP7_75t_L g186 ( .A(n_133), .B(n_108), .Y(n_186) );
AND2x4_ASAP7_75t_L g187 ( .A(n_133), .B(n_108), .Y(n_187) );
AND2x4_ASAP7_75t_L g188 ( .A(n_165), .B(n_108), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_166), .A2(n_153), .B(n_144), .Y(n_189) );
HB1xp67_ASAP7_75t_L g190 ( .A(n_159), .Y(n_190) );
HB1xp67_ASAP7_75t_L g191 ( .A(n_161), .Y(n_191) );
AND2x4_ASAP7_75t_L g192 ( .A(n_165), .B(n_115), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_169), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_166), .A2(n_153), .B(n_144), .Y(n_194) );
AND2x2_ASAP7_75t_L g195 ( .A(n_181), .B(n_112), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_186), .B(n_147), .Y(n_196) );
BUFx4f_ASAP7_75t_SL g197 ( .A(n_154), .Y(n_197) );
HB1xp67_ASAP7_75t_L g198 ( .A(n_162), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_169), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_164), .B(n_131), .Y(n_200) );
AND2x2_ASAP7_75t_L g201 ( .A(n_165), .B(n_112), .Y(n_201) );
INVx1_ASAP7_75t_SL g202 ( .A(n_179), .Y(n_202) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_168), .A2(n_153), .B(n_144), .Y(n_203) );
AOI22xp33_ASAP7_75t_L g204 ( .A1(n_187), .A2(n_145), .B1(n_115), .B2(n_125), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_169), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_172), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_172), .Y(n_207) );
A2O1A1Ixp33_ASAP7_75t_L g208 ( .A1(n_173), .A2(n_145), .B(n_115), .C(n_122), .Y(n_208) );
INVx5_ASAP7_75t_L g209 ( .A(n_179), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_172), .Y(n_210) );
OAI22xp5_ASAP7_75t_L g211 ( .A1(n_179), .A2(n_123), .B1(n_115), .B2(n_127), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_175), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_168), .A2(n_132), .B(n_150), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_175), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_175), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_177), .Y(n_216) );
OAI22x1_ASAP7_75t_L g217 ( .A1(n_184), .A2(n_115), .B1(n_127), .B2(n_79), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_186), .B(n_115), .Y(n_218) );
BUFx6f_ASAP7_75t_L g219 ( .A(n_183), .Y(n_219) );
CKINVDCx8_ASAP7_75t_R g220 ( .A(n_170), .Y(n_220) );
AND2x6_ASAP7_75t_L g221 ( .A(n_202), .B(n_180), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_193), .B(n_186), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_193), .Y(n_223) );
AND2x2_ASAP7_75t_L g224 ( .A(n_199), .B(n_178), .Y(n_224) );
INVx4_ASAP7_75t_L g225 ( .A(n_209), .Y(n_225) );
INVxp67_ASAP7_75t_SL g226 ( .A(n_205), .Y(n_226) );
OR2x2_ASAP7_75t_L g227 ( .A(n_211), .B(n_163), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_199), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_207), .B(n_186), .Y(n_229) );
AOI22xp33_ASAP7_75t_L g230 ( .A1(n_200), .A2(n_187), .B1(n_184), .B2(n_182), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_205), .B(n_183), .Y(n_231) );
AOI22xp33_ASAP7_75t_L g232 ( .A1(n_196), .A2(n_187), .B1(n_182), .B2(n_160), .Y(n_232) );
AND2x4_ASAP7_75t_L g233 ( .A(n_209), .B(n_178), .Y(n_233) );
HB1xp67_ASAP7_75t_L g234 ( .A(n_209), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_207), .Y(n_235) );
INVx3_ASAP7_75t_L g236 ( .A(n_209), .Y(n_236) );
OAI211xp5_ASAP7_75t_SL g237 ( .A1(n_204), .A2(n_176), .B(n_158), .C(n_171), .Y(n_237) );
BUFx3_ASAP7_75t_L g238 ( .A(n_209), .Y(n_238) );
OAI21x1_ASAP7_75t_L g239 ( .A1(n_189), .A2(n_163), .B(n_155), .Y(n_239) );
CKINVDCx5p33_ASAP7_75t_R g240 ( .A(n_197), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_210), .Y(n_241) );
BUFx3_ASAP7_75t_L g242 ( .A(n_209), .Y(n_242) );
AOI22xp33_ASAP7_75t_L g243 ( .A1(n_195), .A2(n_187), .B1(n_160), .B2(n_155), .Y(n_243) );
OAI22xp33_ASAP7_75t_L g244 ( .A1(n_210), .A2(n_174), .B1(n_171), .B2(n_123), .Y(n_244) );
AOI22xp33_ASAP7_75t_L g245 ( .A1(n_195), .A2(n_155), .B1(n_157), .B2(n_167), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_212), .Y(n_246) );
OAI22xp5_ASAP7_75t_L g247 ( .A1(n_227), .A2(n_216), .B1(n_215), .B2(n_214), .Y(n_247) );
INVx2_ASAP7_75t_L g248 ( .A(n_226), .Y(n_248) );
AOI22xp33_ASAP7_75t_L g249 ( .A1(n_237), .A2(n_154), .B1(n_156), .B2(n_191), .Y(n_249) );
AND2x2_ASAP7_75t_L g250 ( .A(n_224), .B(n_212), .Y(n_250) );
BUFx3_ASAP7_75t_L g251 ( .A(n_238), .Y(n_251) );
AOI22xp33_ASAP7_75t_L g252 ( .A1(n_237), .A2(n_154), .B1(n_190), .B2(n_198), .Y(n_252) );
AOI211xp5_ASAP7_75t_L g253 ( .A1(n_244), .A2(n_97), .B(n_99), .C(n_201), .Y(n_253) );
AOI221xp5_ASAP7_75t_L g254 ( .A1(n_244), .A2(n_217), .B1(n_176), .B2(n_218), .C(n_208), .Y(n_254) );
AO31x2_ASAP7_75t_L g255 ( .A1(n_223), .A2(n_217), .A3(n_205), .B(n_206), .Y(n_255) );
AOI222xp33_ASAP7_75t_L g256 ( .A1(n_243), .A2(n_154), .B1(n_201), .B2(n_111), .C1(n_215), .C2(n_214), .Y(n_256) );
OAI211xp5_ASAP7_75t_SL g257 ( .A1(n_243), .A2(n_158), .B(n_220), .C(n_120), .Y(n_257) );
AOI22xp33_ASAP7_75t_L g258 ( .A1(n_227), .A2(n_192), .B1(n_188), .B2(n_111), .Y(n_258) );
AOI22xp5_ASAP7_75t_L g259 ( .A1(n_227), .A2(n_216), .B1(n_206), .B2(n_188), .Y(n_259) );
AOI21xp5_ASAP7_75t_SL g260 ( .A1(n_226), .A2(n_206), .B(n_219), .Y(n_260) );
AOI21xp33_ASAP7_75t_L g261 ( .A1(n_231), .A2(n_120), .B(n_202), .Y(n_261) );
OA21x2_ASAP7_75t_L g262 ( .A1(n_239), .A2(n_194), .B(n_203), .Y(n_262) );
OAI21x1_ASAP7_75t_L g263 ( .A1(n_239), .A2(n_213), .B(n_155), .Y(n_263) );
AO21x2_ASAP7_75t_L g264 ( .A1(n_239), .A2(n_173), .B(n_88), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_223), .Y(n_265) );
AOI221xp5_ASAP7_75t_L g266 ( .A1(n_230), .A2(n_222), .B1(n_229), .B2(n_245), .C(n_232), .Y(n_266) );
OAI21x1_ASAP7_75t_L g267 ( .A1(n_263), .A2(n_231), .B(n_236), .Y(n_267) );
INVx3_ASAP7_75t_L g268 ( .A(n_248), .Y(n_268) );
AOI22xp33_ASAP7_75t_L g269 ( .A1(n_256), .A2(n_245), .B1(n_232), .B2(n_224), .Y(n_269) );
NOR2xp33_ASAP7_75t_L g270 ( .A(n_249), .B(n_220), .Y(n_270) );
AOI21xp5_ASAP7_75t_L g271 ( .A1(n_248), .A2(n_260), .B(n_247), .Y(n_271) );
NOR4xp25_ASAP7_75t_SL g272 ( .A(n_257), .B(n_240), .C(n_228), .D(n_241), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_265), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_265), .Y(n_274) );
OAI211xp5_ASAP7_75t_L g275 ( .A1(n_253), .A2(n_91), .B(n_234), .C(n_94), .Y(n_275) );
OAI321xp33_ASAP7_75t_L g276 ( .A1(n_254), .A2(n_252), .A3(n_258), .B1(n_247), .B2(n_259), .C(n_266), .Y(n_276) );
OAI221xp5_ASAP7_75t_L g277 ( .A1(n_256), .A2(n_246), .B1(n_228), .B2(n_235), .C(n_183), .Y(n_277) );
AOI21xp5_ASAP7_75t_L g278 ( .A1(n_248), .A2(n_235), .B(n_183), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_250), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_250), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_255), .Y(n_281) );
OAI211xp5_ASAP7_75t_L g282 ( .A1(n_254), .A2(n_234), .B(n_101), .C(n_88), .Y(n_282) );
AOI22xp33_ASAP7_75t_L g283 ( .A1(n_266), .A2(n_224), .B1(n_233), .B2(n_221), .Y(n_283) );
NOR4xp25_ASAP7_75t_SL g284 ( .A(n_261), .B(n_100), .C(n_87), .D(n_92), .Y(n_284) );
OA21x2_ASAP7_75t_L g285 ( .A1(n_263), .A2(n_261), .B(n_259), .Y(n_285) );
OR2x2_ASAP7_75t_L g286 ( .A(n_255), .B(n_233), .Y(n_286) );
AND2x2_ASAP7_75t_L g287 ( .A(n_255), .B(n_236), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_273), .Y(n_288) );
AND2x2_ASAP7_75t_L g289 ( .A(n_268), .B(n_264), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_268), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_268), .Y(n_291) );
INVx2_ASAP7_75t_SL g292 ( .A(n_268), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_273), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_274), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_274), .Y(n_295) );
HB1xp67_ASAP7_75t_L g296 ( .A(n_286), .Y(n_296) );
AND2x2_ASAP7_75t_L g297 ( .A(n_287), .B(n_264), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_281), .Y(n_298) );
INVx6_ASAP7_75t_L g299 ( .A(n_286), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_281), .Y(n_300) );
AND2x2_ASAP7_75t_L g301 ( .A(n_287), .B(n_264), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_279), .B(n_255), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_279), .Y(n_303) );
OR2x2_ASAP7_75t_L g304 ( .A(n_280), .B(n_255), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_280), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_271), .Y(n_306) );
BUFx2_ASAP7_75t_L g307 ( .A(n_267), .Y(n_307) );
AND2x2_ASAP7_75t_L g308 ( .A(n_285), .B(n_264), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_267), .Y(n_309) );
OAI211xp5_ASAP7_75t_SL g310 ( .A1(n_275), .A2(n_93), .B(n_113), .C(n_109), .Y(n_310) );
OR2x2_ASAP7_75t_L g311 ( .A(n_283), .B(n_255), .Y(n_311) );
AOI22xp33_ASAP7_75t_L g312 ( .A1(n_277), .A2(n_233), .B1(n_221), .B2(n_251), .Y(n_312) );
NAND3xp33_ASAP7_75t_L g313 ( .A(n_284), .B(n_93), .C(n_89), .Y(n_313) );
OAI21xp5_ASAP7_75t_SL g314 ( .A1(n_269), .A2(n_233), .B(n_236), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_285), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_285), .Y(n_316) );
AND2x2_ASAP7_75t_L g317 ( .A(n_285), .B(n_251), .Y(n_317) );
CKINVDCx5p33_ASAP7_75t_R g318 ( .A(n_299), .Y(n_318) );
BUFx2_ASAP7_75t_L g319 ( .A(n_299), .Y(n_319) );
OR2x2_ASAP7_75t_L g320 ( .A(n_296), .B(n_251), .Y(n_320) );
OR2x2_ASAP7_75t_L g321 ( .A(n_304), .B(n_278), .Y(n_321) );
INVx3_ASAP7_75t_L g322 ( .A(n_292), .Y(n_322) );
OR2x2_ASAP7_75t_L g323 ( .A(n_304), .B(n_89), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_303), .B(n_282), .Y(n_324) );
NAND4xp25_ASAP7_75t_L g325 ( .A(n_312), .B(n_270), .C(n_109), .D(n_113), .Y(n_325) );
NOR2xp33_ASAP7_75t_L g326 ( .A(n_303), .B(n_276), .Y(n_326) );
NAND4xp25_ASAP7_75t_L g327 ( .A(n_314), .B(n_109), .C(n_113), .D(n_98), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_288), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_305), .B(n_89), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_293), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_293), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_294), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_297), .B(n_105), .Y(n_333) );
CKINVDCx20_ASAP7_75t_R g334 ( .A(n_299), .Y(n_334) );
AOI22xp33_ASAP7_75t_L g335 ( .A1(n_299), .A2(n_89), .B1(n_221), .B2(n_238), .Y(n_335) );
NAND2xp5_ASAP7_75t_SL g336 ( .A(n_292), .B(n_276), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_295), .Y(n_337) );
NOR2xp33_ASAP7_75t_L g338 ( .A(n_305), .B(n_2), .Y(n_338) );
NOR2xp67_ASAP7_75t_SL g339 ( .A(n_313), .B(n_260), .Y(n_339) );
AOI22x1_ASAP7_75t_L g340 ( .A1(n_289), .A2(n_225), .B1(n_109), .B2(n_113), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_298), .B(n_272), .Y(n_341) );
OR2x2_ASAP7_75t_L g342 ( .A(n_302), .B(n_262), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_298), .B(n_272), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_297), .B(n_105), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_300), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_300), .Y(n_346) );
NOR3xp33_ASAP7_75t_SL g347 ( .A(n_310), .B(n_2), .C(n_3), .Y(n_347) );
OR2x2_ASAP7_75t_L g348 ( .A(n_301), .B(n_262), .Y(n_348) );
OAI33xp33_ASAP7_75t_L g349 ( .A1(n_311), .A2(n_4), .A3(n_5), .B1(n_6), .B2(n_7), .B3(n_8), .Y(n_349) );
INVx3_ASAP7_75t_L g350 ( .A(n_290), .Y(n_350) );
AND2x4_ASAP7_75t_L g351 ( .A(n_317), .B(n_238), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_301), .B(n_105), .Y(n_352) );
NOR4xp25_ASAP7_75t_SL g353 ( .A(n_307), .B(n_284), .C(n_7), .D(n_8), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_311), .B(n_109), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_290), .Y(n_355) );
OAI21xp5_ASAP7_75t_L g356 ( .A1(n_313), .A2(n_109), .B(n_113), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_291), .Y(n_357) );
OAI31xp33_ASAP7_75t_SL g358 ( .A1(n_317), .A2(n_233), .A3(n_192), .B(n_10), .Y(n_358) );
AND2x4_ASAP7_75t_L g359 ( .A(n_334), .B(n_319), .Y(n_359) );
NOR2xp33_ASAP7_75t_SL g360 ( .A(n_318), .B(n_225), .Y(n_360) );
OR2x2_ASAP7_75t_L g361 ( .A(n_323), .B(n_291), .Y(n_361) );
AOI21xp5_ASAP7_75t_L g362 ( .A1(n_340), .A2(n_306), .B(n_308), .Y(n_362) );
OAI22xp5_ASAP7_75t_L g363 ( .A1(n_334), .A2(n_308), .B1(n_306), .B2(n_307), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_333), .B(n_315), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_318), .B(n_315), .Y(n_365) );
AOI221xp5_ASAP7_75t_L g366 ( .A1(n_326), .A2(n_113), .B1(n_316), .B2(n_309), .C(n_117), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_333), .B(n_316), .Y(n_367) );
OAI321xp33_ASAP7_75t_L g368 ( .A1(n_336), .A2(n_309), .A3(n_126), .B1(n_117), .B2(n_105), .C(n_12), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_332), .Y(n_369) );
OAI21xp33_ASAP7_75t_L g370 ( .A1(n_358), .A2(n_117), .B(n_126), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_337), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_319), .B(n_105), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_344), .B(n_6), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_344), .B(n_9), .Y(n_374) );
OAI322xp33_ASAP7_75t_L g375 ( .A1(n_323), .A2(n_117), .A3(n_126), .B1(n_11), .B2(n_13), .C1(n_14), .C2(n_16), .Y(n_375) );
INVxp67_ASAP7_75t_SL g376 ( .A(n_320), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_328), .Y(n_377) );
OAI222xp33_ASAP7_75t_L g378 ( .A1(n_336), .A2(n_225), .B1(n_236), .B2(n_238), .C1(n_242), .C2(n_192), .Y(n_378) );
AOI22xp5_ASAP7_75t_L g379 ( .A1(n_327), .A2(n_221), .B1(n_225), .B2(n_236), .Y(n_379) );
AOI322xp5_ASAP7_75t_L g380 ( .A1(n_352), .A2(n_117), .A3(n_126), .B1(n_11), .B2(n_13), .C1(n_17), .C2(n_18), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_328), .Y(n_381) );
AOI221xp5_ASAP7_75t_L g382 ( .A1(n_349), .A2(n_126), .B1(n_225), .B2(n_185), .C(n_22), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_330), .Y(n_383) );
XOR2x2_ASAP7_75t_L g384 ( .A(n_338), .B(n_9), .Y(n_384) );
NOR2x1p5_ASAP7_75t_SL g385 ( .A(n_342), .B(n_135), .Y(n_385) );
A2O1A1Ixp33_ASAP7_75t_L g386 ( .A1(n_347), .A2(n_242), .B(n_219), .C(n_126), .Y(n_386) );
OAI22xp5_ASAP7_75t_L g387 ( .A1(n_324), .A2(n_242), .B1(n_262), .B2(n_219), .Y(n_387) );
AOI211xp5_ASAP7_75t_L g388 ( .A1(n_325), .A2(n_126), .B(n_242), .C(n_219), .Y(n_388) );
OAI21xp5_ASAP7_75t_L g389 ( .A1(n_356), .A2(n_221), .B(n_262), .Y(n_389) );
NAND2xp33_ASAP7_75t_SL g390 ( .A(n_339), .B(n_219), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_330), .Y(n_391) );
NOR2xp33_ASAP7_75t_L g392 ( .A(n_354), .B(n_19), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_346), .B(n_20), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_331), .B(n_126), .Y(n_394) );
OAI21xp5_ASAP7_75t_SL g395 ( .A1(n_335), .A2(n_126), .B(n_22), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_331), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_345), .B(n_20), .Y(n_397) );
NAND4xp25_ASAP7_75t_L g398 ( .A(n_341), .B(n_23), .C(n_24), .D(n_185), .Y(n_398) );
INVx2_ASAP7_75t_SL g399 ( .A(n_351), .Y(n_399) );
AOI32xp33_ASAP7_75t_L g400 ( .A1(n_351), .A2(n_23), .A3(n_24), .B1(n_177), .B2(n_221), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_348), .B(n_25), .Y(n_401) );
OAI221xp5_ASAP7_75t_SL g402 ( .A1(n_321), .A2(n_167), .B1(n_157), .B2(n_221), .C(n_141), .Y(n_402) );
NOR3xp33_ASAP7_75t_SL g403 ( .A(n_398), .B(n_343), .C(n_329), .Y(n_403) );
AOI21xp5_ASAP7_75t_L g404 ( .A1(n_390), .A2(n_321), .B(n_342), .Y(n_404) );
XNOR2xp5_ASAP7_75t_L g405 ( .A(n_384), .B(n_345), .Y(n_405) );
AOI22xp33_ASAP7_75t_L g406 ( .A1(n_370), .A2(n_322), .B1(n_350), .B2(n_357), .Y(n_406) );
OAI33xp33_ASAP7_75t_L g407 ( .A1(n_363), .A2(n_355), .A3(n_353), .B1(n_322), .B2(n_350), .B3(n_141), .Y(n_407) );
AOI322xp5_ASAP7_75t_L g408 ( .A1(n_376), .A2(n_350), .A3(n_221), .B1(n_141), .B2(n_135), .C1(n_34), .C2(n_36), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_369), .Y(n_409) );
CKINVDCx5p33_ASAP7_75t_R g410 ( .A(n_359), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_371), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_372), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_377), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_381), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_383), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_391), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_396), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_365), .B(n_28), .Y(n_418) );
OAI211xp5_ASAP7_75t_SL g419 ( .A1(n_400), .A2(n_135), .B(n_149), .C(n_33), .Y(n_419) );
AOI21xp33_ASAP7_75t_L g420 ( .A1(n_373), .A2(n_29), .B(n_32), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_394), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_364), .B(n_38), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_397), .Y(n_423) );
OR2x2_ASAP7_75t_L g424 ( .A(n_364), .B(n_40), .Y(n_424) );
AND2x4_ASAP7_75t_L g425 ( .A(n_399), .B(n_41), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_397), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_367), .B(n_42), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_367), .Y(n_428) );
INVxp67_ASAP7_75t_SL g429 ( .A(n_363), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_394), .Y(n_430) );
OR2x2_ASAP7_75t_L g431 ( .A(n_361), .B(n_48), .Y(n_431) );
XNOR2x1_ASAP7_75t_L g432 ( .A(n_374), .B(n_50), .Y(n_432) );
OR2x2_ASAP7_75t_L g433 ( .A(n_387), .B(n_51), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_393), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_385), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_387), .B(n_53), .Y(n_436) );
INVx4_ASAP7_75t_L g437 ( .A(n_401), .Y(n_437) );
NAND2xp5_ASAP7_75t_SL g438 ( .A(n_360), .B(n_362), .Y(n_438) );
INVx2_ASAP7_75t_SL g439 ( .A(n_410), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_429), .B(n_382), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_428), .B(n_366), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_423), .B(n_380), .Y(n_442) );
AOI22xp5_ASAP7_75t_L g443 ( .A1(n_432), .A2(n_392), .B1(n_395), .B2(n_379), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_426), .B(n_389), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_409), .Y(n_445) );
OAI22xp5_ASAP7_75t_L g446 ( .A1(n_437), .A2(n_388), .B1(n_402), .B2(n_386), .Y(n_446) );
AOI22xp33_ASAP7_75t_SL g447 ( .A1(n_437), .A2(n_378), .B1(n_375), .B2(n_368), .Y(n_447) );
INVx2_ASAP7_75t_SL g448 ( .A(n_410), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_434), .B(n_54), .Y(n_449) );
INVx1_ASAP7_75t_SL g450 ( .A(n_425), .Y(n_450) );
AOI21xp5_ASAP7_75t_L g451 ( .A1(n_438), .A2(n_149), .B(n_138), .Y(n_451) );
NOR2x1_ASAP7_75t_L g452 ( .A(n_438), .B(n_56), .Y(n_452) );
OR2x2_ASAP7_75t_L g453 ( .A(n_413), .B(n_57), .Y(n_453) );
AOI32xp33_ASAP7_75t_L g454 ( .A1(n_437), .A2(n_58), .A3(n_60), .B1(n_61), .B2(n_64), .Y(n_454) );
OAI221xp5_ASAP7_75t_L g455 ( .A1(n_403), .A2(n_138), .B1(n_137), .B2(n_71), .C(n_72), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_430), .B(n_66), .Y(n_456) );
XOR2x2_ASAP7_75t_L g457 ( .A(n_405), .B(n_69), .Y(n_457) );
NOR3xp33_ASAP7_75t_L g458 ( .A(n_407), .B(n_150), .C(n_132), .Y(n_458) );
NAND3xp33_ASAP7_75t_L g459 ( .A(n_403), .B(n_137), .C(n_138), .Y(n_459) );
OAI22xp5_ASAP7_75t_L g460 ( .A1(n_439), .A2(n_406), .B1(n_404), .B2(n_435), .Y(n_460) );
OAI21xp5_ASAP7_75t_SL g461 ( .A1(n_447), .A2(n_406), .B(n_419), .Y(n_461) );
NAND4xp25_ASAP7_75t_SL g462 ( .A(n_443), .B(n_408), .C(n_418), .D(n_436), .Y(n_462) );
AOI221xp5_ASAP7_75t_L g463 ( .A1(n_440), .A2(n_411), .B1(n_412), .B2(n_415), .C(n_417), .Y(n_463) );
BUFx2_ASAP7_75t_L g464 ( .A(n_448), .Y(n_464) );
NAND2x1p5_ASAP7_75t_L g465 ( .A(n_452), .B(n_425), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_440), .B(n_416), .Y(n_466) );
NAND2xp33_ASAP7_75t_L g467 ( .A(n_454), .B(n_418), .Y(n_467) );
AOI22xp5_ASAP7_75t_L g468 ( .A1(n_446), .A2(n_442), .B1(n_450), .B2(n_457), .Y(n_468) );
AOI332xp33_ASAP7_75t_L g469 ( .A1(n_445), .A2(n_414), .A3(n_421), .B1(n_422), .B2(n_427), .B3(n_424), .C1(n_433), .C2(n_431), .Y(n_469) );
OAI21xp33_ASAP7_75t_L g470 ( .A1(n_444), .A2(n_422), .B(n_420), .Y(n_470) );
AND2x4_ASAP7_75t_L g471 ( .A(n_450), .B(n_137), .Y(n_471) );
NAND3xp33_ASAP7_75t_SL g472 ( .A(n_446), .B(n_150), .C(n_132), .Y(n_472) );
OAI211xp5_ASAP7_75t_SL g473 ( .A1(n_441), .A2(n_137), .B(n_138), .C(n_150), .Y(n_473) );
NAND4xp25_ASAP7_75t_L g474 ( .A(n_459), .B(n_137), .C(n_138), .D(n_455), .Y(n_474) );
OAI211xp5_ASAP7_75t_L g475 ( .A1(n_441), .A2(n_138), .B(n_451), .C(n_449), .Y(n_475) );
OAI22xp5_ASAP7_75t_SL g476 ( .A1(n_453), .A2(n_405), .B1(n_448), .B2(n_439), .Y(n_476) );
NOR3xp33_ASAP7_75t_L g477 ( .A(n_456), .B(n_440), .C(n_459), .Y(n_477) );
OAI221xp5_ASAP7_75t_L g478 ( .A1(n_458), .A2(n_429), .B1(n_440), .B2(n_447), .C(n_442), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_477), .B(n_463), .Y(n_479) );
NAND3xp33_ASAP7_75t_SL g480 ( .A(n_468), .B(n_461), .C(n_478), .Y(n_480) );
XOR2xp5_ASAP7_75t_L g481 ( .A(n_468), .B(n_476), .Y(n_481) );
INVx1_ASAP7_75t_SL g482 ( .A(n_464), .Y(n_482) );
NAND3xp33_ASAP7_75t_SL g483 ( .A(n_475), .B(n_469), .C(n_465), .Y(n_483) );
NAND4xp75_ASAP7_75t_L g484 ( .A(n_479), .B(n_466), .C(n_462), .D(n_472), .Y(n_484) );
XNOR2xp5_ASAP7_75t_L g485 ( .A(n_481), .B(n_460), .Y(n_485) );
AND2x2_ASAP7_75t_SL g486 ( .A(n_480), .B(n_467), .Y(n_486) );
INVxp67_ASAP7_75t_SL g487 ( .A(n_485), .Y(n_487) );
CKINVDCx20_ASAP7_75t_R g488 ( .A(n_486), .Y(n_488) );
INVxp67_ASAP7_75t_L g489 ( .A(n_487), .Y(n_489) );
AOI322xp5_ASAP7_75t_L g490 ( .A1(n_489), .A2(n_488), .A3(n_486), .B1(n_482), .B2(n_483), .C1(n_484), .C2(n_470), .Y(n_490) );
O2A1O1Ixp33_ASAP7_75t_L g491 ( .A1(n_490), .A2(n_474), .B(n_473), .C(n_471), .Y(n_491) );
endmodule