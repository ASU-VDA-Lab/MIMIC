module fake_jpeg_12676_n_559 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_559);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_559;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_479;
wire n_415;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_18),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_8),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

INVx8_ASAP7_75t_SL g41 ( 
.A(n_7),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_3),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_4),
.Y(n_46)
);

BUFx4f_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

CKINVDCx14_ASAP7_75t_R g48 ( 
.A(n_6),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_18),
.Y(n_50)
);

BUFx16f_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_16),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_53),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_42),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_54),
.B(n_66),
.Y(n_142)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_55),
.Y(n_136)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_56),
.Y(n_148)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g143 ( 
.A(n_57),
.Y(n_143)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_58),
.Y(n_109)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx13_ASAP7_75t_L g113 ( 
.A(n_59),
.Y(n_113)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_60),
.Y(n_120)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_61),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_41),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_62),
.B(n_72),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_63),
.Y(n_119)
);

AND2x2_ASAP7_75t_SL g64 ( 
.A(n_30),
.B(n_0),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_64),
.B(n_44),
.C(n_32),
.Y(n_175)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g125 ( 
.A(n_65),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_9),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_67),
.Y(n_153)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_68),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g111 ( 
.A(n_69),
.Y(n_111)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_70),
.Y(n_122)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_71),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_30),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_22),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_73),
.Y(n_146)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_74),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_24),
.B(n_9),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_75),
.B(n_85),
.Y(n_139)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_76),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_9),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_77),
.B(n_80),
.Y(n_134)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_30),
.Y(n_78)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_78),
.Y(n_171)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_79),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_8),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_81),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_23),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_82),
.Y(n_145)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_21),
.Y(n_83)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_83),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_30),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g170 ( 
.A(n_84),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_24),
.B(n_18),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_21),
.Y(n_86)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_86),
.Y(n_138)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_22),
.Y(n_87)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_87),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_23),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_88),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_22),
.Y(n_89)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_89),
.Y(n_110)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_31),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_90),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_33),
.B(n_18),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_91),
.B(n_102),
.Y(n_140)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_31),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_92),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_25),
.Y(n_93)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_93),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_31),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_94),
.Y(n_173)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_25),
.Y(n_95)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_95),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_51),
.B(n_33),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_96),
.B(n_100),
.Y(n_151)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_97),
.Y(n_172)
);

INVx3_ASAP7_75t_SL g98 ( 
.A(n_30),
.Y(n_98)
);

INVx2_ASAP7_75t_SL g162 ( 
.A(n_98),
.Y(n_162)
);

INVx2_ASAP7_75t_SL g99 ( 
.A(n_30),
.Y(n_99)
);

BUFx2_ASAP7_75t_R g166 ( 
.A(n_99),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_25),
.B(n_8),
.Y(n_100)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_30),
.Y(n_101)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_101),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_19),
.B(n_26),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_31),
.Y(n_103)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_103),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_36),
.Y(n_104)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_104),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_19),
.B(n_8),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_105),
.B(n_49),
.Y(n_147)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_21),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_106),
.B(n_107),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_32),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_21),
.Y(n_108)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_108),
.Y(n_144)
);

BUFx10_ASAP7_75t_L g115 ( 
.A(n_59),
.Y(n_115)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_115),
.Y(n_240)
);

INVx11_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

INVx5_ASAP7_75t_SL g228 ( 
.A(n_117),
.Y(n_228)
);

OAI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_108),
.A2(n_36),
.B1(n_37),
.B2(n_25),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_127),
.A2(n_55),
.B1(n_67),
.B2(n_71),
.Y(n_192)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_84),
.Y(n_128)
);

INVx5_ASAP7_75t_L g226 ( 
.A(n_128),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_59),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_132),
.B(n_133),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_79),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_58),
.A2(n_37),
.B1(n_36),
.B2(n_40),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_135),
.A2(n_152),
.B1(n_161),
.B2(n_98),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_147),
.B(n_156),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_97),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_149),
.B(n_176),
.Y(n_197)
);

OAI22xp33_ASAP7_75t_L g152 ( 
.A1(n_90),
.A2(n_37),
.B1(n_36),
.B2(n_28),
.Y(n_152)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_63),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_155),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_73),
.B(n_26),
.Y(n_156)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_68),
.Y(n_157)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_157),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_64),
.A2(n_44),
.B(n_32),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_159),
.A2(n_78),
.B(n_93),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_73),
.B(n_26),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_160),
.B(n_164),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_92),
.A2(n_104),
.B1(n_103),
.B2(n_94),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_68),
.B(n_20),
.Y(n_164)
);

BUFx10_ASAP7_75t_L g168 ( 
.A(n_65),
.Y(n_168)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_168),
.Y(n_187)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_69),
.Y(n_174)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_174),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_175),
.B(n_101),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_53),
.Y(n_176)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_124),
.Y(n_178)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_178),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_166),
.Y(n_179)
);

INVx4_ASAP7_75t_SL g289 ( 
.A(n_179),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_152),
.A2(n_88),
.B1(n_82),
.B2(n_52),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_180),
.A2(n_192),
.B1(n_212),
.B2(n_45),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_139),
.B(n_64),
.C(n_81),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_181),
.B(n_239),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_115),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_182),
.B(n_216),
.Y(n_254)
);

BUFx12f_ASAP7_75t_L g184 ( 
.A(n_146),
.Y(n_184)
);

INVx4_ASAP7_75t_L g252 ( 
.A(n_184),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_185),
.A2(n_207),
.B1(n_213),
.B2(n_215),
.Y(n_244)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_136),
.Y(n_186)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_186),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_188),
.B(n_112),
.Y(n_241)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_116),
.Y(n_189)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_189),
.Y(n_248)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_153),
.Y(n_190)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_190),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_147),
.B(n_140),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_191),
.B(n_201),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_141),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_193),
.B(n_196),
.Y(n_253)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_131),
.Y(n_195)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_195),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_143),
.Y(n_196)
);

BUFx12f_ASAP7_75t_L g198 ( 
.A(n_146),
.Y(n_198)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_198),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_111),
.Y(n_199)
);

INVx5_ASAP7_75t_L g284 ( 
.A(n_199),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_119),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_200),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_165),
.B(n_138),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_154),
.Y(n_202)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_202),
.Y(n_260)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_122),
.Y(n_203)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_203),
.Y(n_249)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_137),
.Y(n_205)
);

BUFx2_ASAP7_75t_L g256 ( 
.A(n_205),
.Y(n_256)
);

CKINVDCx12_ASAP7_75t_R g206 ( 
.A(n_115),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_206),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_135),
.A2(n_76),
.B1(n_89),
.B2(n_95),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_119),
.Y(n_208)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_208),
.Y(n_259)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_137),
.Y(n_209)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_209),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_151),
.A2(n_44),
.B1(n_49),
.B2(n_43),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_210),
.A2(n_211),
.B1(n_34),
.B2(n_20),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_134),
.A2(n_49),
.B1(n_43),
.B2(n_40),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_127),
.A2(n_20),
.B1(n_38),
.B2(n_34),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_161),
.A2(n_19),
.B1(n_46),
.B2(n_45),
.Y(n_213)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_110),
.Y(n_214)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_214),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_142),
.A2(n_37),
.B1(n_28),
.B2(n_50),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_123),
.B(n_50),
.Y(n_216)
);

OR2x2_ASAP7_75t_L g217 ( 
.A(n_120),
.B(n_40),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_217),
.B(n_227),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_167),
.B(n_28),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_218),
.B(n_222),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_219),
.A2(n_129),
.B(n_112),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_148),
.A2(n_52),
.B1(n_50),
.B2(n_46),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_220),
.A2(n_45),
.B1(n_34),
.B2(n_38),
.Y(n_277)
);

CKINVDCx9p33_ASAP7_75t_R g221 ( 
.A(n_117),
.Y(n_221)
);

OR2x2_ASAP7_75t_L g266 ( 
.A(n_221),
.B(n_231),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_172),
.B(n_28),
.Y(n_222)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_126),
.Y(n_224)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_224),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_145),
.Y(n_225)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_225),
.Y(n_251)
);

CKINVDCx12_ASAP7_75t_R g227 ( 
.A(n_113),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_150),
.B(n_27),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_229),
.B(n_237),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_145),
.Y(n_230)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_230),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_144),
.B(n_52),
.Y(n_231)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_110),
.Y(n_232)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_232),
.Y(n_267)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_111),
.Y(n_233)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_233),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_111),
.Y(n_234)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_234),
.Y(n_280)
);

INVx5_ASAP7_75t_L g236 ( 
.A(n_129),
.Y(n_236)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_236),
.Y(n_282)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_171),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_144),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_238),
.B(n_162),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_118),
.B(n_46),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_241),
.B(n_243),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_179),
.A2(n_168),
.B(n_166),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_192),
.A2(n_109),
.B1(n_169),
.B2(n_163),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_245),
.A2(n_290),
.B1(n_291),
.B2(n_228),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_247),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_188),
.B(n_162),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g296 ( 
.A(n_263),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_215),
.A2(n_168),
.B1(n_174),
.B2(n_157),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_268),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_272),
.B(n_276),
.Y(n_311)
);

CKINVDCx14_ASAP7_75t_R g314 ( 
.A(n_274),
.Y(n_314)
);

O2A1O1Ixp33_ASAP7_75t_SL g276 ( 
.A1(n_219),
.A2(n_113),
.B(n_128),
.C(n_170),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_277),
.A2(n_278),
.B1(n_286),
.B2(n_228),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_207),
.A2(n_118),
.B1(n_155),
.B2(n_121),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_281),
.B(n_288),
.Y(n_326)
);

OA22x2_ASAP7_75t_L g283 ( 
.A1(n_221),
.A2(n_114),
.B1(n_169),
.B2(n_163),
.Y(n_283)
);

OA22x2_ASAP7_75t_L g324 ( 
.A1(n_283),
.A2(n_204),
.B1(n_223),
.B2(n_205),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_L g286 ( 
.A1(n_217),
.A2(n_121),
.B1(n_158),
.B2(n_173),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_183),
.B(n_130),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_287),
.B(n_187),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_235),
.A2(n_38),
.B(n_27),
.Y(n_288)
);

OAI22xp33_ASAP7_75t_L g290 ( 
.A1(n_239),
.A2(n_158),
.B1(n_173),
.B2(n_109),
.Y(n_290)
);

OAI22xp33_ASAP7_75t_L g291 ( 
.A1(n_201),
.A2(n_130),
.B1(n_43),
.B2(n_27),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_249),
.Y(n_292)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_292),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_253),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_293),
.B(n_295),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_254),
.B(n_177),
.Y(n_294)
);

CKINVDCx14_ASAP7_75t_R g344 ( 
.A(n_294),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_271),
.Y(n_295)
);

BUFx12f_ASAP7_75t_L g297 ( 
.A(n_258),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_297),
.B(n_300),
.Y(n_359)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_261),
.Y(n_298)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_298),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_299),
.A2(n_323),
.B1(n_332),
.B2(n_336),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_285),
.B(n_181),
.C(n_219),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_301),
.B(n_331),
.C(n_243),
.Y(n_337)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_249),
.Y(n_302)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_302),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g340 ( 
.A(n_303),
.B(n_324),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_248),
.B(n_246),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_304),
.B(n_305),
.Y(n_363)
);

AND2x6_ASAP7_75t_L g305 ( 
.A(n_285),
.B(n_191),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_269),
.B(n_197),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_306),
.B(n_307),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_269),
.B(n_186),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_267),
.Y(n_308)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_308),
.Y(n_356)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_242),
.Y(n_309)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_309),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_255),
.B(n_224),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_312),
.Y(n_350)
);

INVx6_ASAP7_75t_L g315 ( 
.A(n_273),
.Y(n_315)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_315),
.Y(n_367)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_242),
.Y(n_316)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_316),
.Y(n_371)
);

AND2x6_ASAP7_75t_L g317 ( 
.A(n_276),
.B(n_226),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_317),
.B(n_319),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_262),
.B(n_178),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_273),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_320),
.Y(n_362)
);

AND2x6_ASAP7_75t_L g321 ( 
.A(n_241),
.B(n_226),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_321),
.B(n_329),
.Y(n_366)
);

CKINVDCx9p33_ASAP7_75t_R g322 ( 
.A(n_289),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g341 ( 
.A(n_322),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_290),
.A2(n_194),
.B1(n_190),
.B2(n_202),
.Y(n_323)
);

INVx4_ASAP7_75t_L g325 ( 
.A(n_261),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_325),
.B(n_328),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_244),
.A2(n_194),
.B1(n_200),
.B2(n_208),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_327),
.A2(n_330),
.B1(n_251),
.B2(n_265),
.Y(n_338)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_250),
.Y(n_328)
);

INVx1_ASAP7_75t_SL g329 ( 
.A(n_263),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_244),
.A2(n_230),
.B1(n_225),
.B2(n_209),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_263),
.B(n_240),
.C(n_214),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_245),
.A2(n_232),
.B1(n_236),
.B2(n_223),
.Y(n_332)
);

INVx1_ASAP7_75t_SL g333 ( 
.A(n_241),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_333),
.B(n_334),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_266),
.B(n_240),
.Y(n_334)
);

INVx5_ASAP7_75t_L g335 ( 
.A(n_259),
.Y(n_335)
);

CKINVDCx16_ASAP7_75t_R g343 ( 
.A(n_335),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_266),
.B(n_204),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_337),
.B(n_339),
.Y(n_387)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_338),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_301),
.B(n_281),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_311),
.A2(n_291),
.B1(n_268),
.B2(n_288),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_345),
.A2(n_346),
.B1(n_357),
.B2(n_358),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_311),
.A2(n_283),
.B1(n_278),
.B2(n_267),
.Y(n_346)
);

AOI22xp33_ASAP7_75t_L g347 ( 
.A1(n_327),
.A2(n_283),
.B1(n_289),
.B2(n_265),
.Y(n_347)
);

AOI22xp33_ASAP7_75t_SL g379 ( 
.A1(n_347),
.A2(n_351),
.B1(n_324),
.B2(n_325),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_296),
.B(n_329),
.C(n_305),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_348),
.Y(n_377)
);

OAI22x1_ASAP7_75t_L g351 ( 
.A1(n_317),
.A2(n_283),
.B1(n_277),
.B2(n_252),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_322),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_353),
.B(n_297),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_311),
.A2(n_251),
.B1(n_282),
.B2(n_259),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_313),
.A2(n_318),
.B1(n_296),
.B2(n_333),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_313),
.A2(n_318),
.B1(n_310),
.B2(n_326),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_SL g376 ( 
.A1(n_361),
.A2(n_326),
.B(n_331),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_299),
.A2(n_282),
.B1(n_264),
.B2(n_275),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_365),
.A2(n_309),
.B1(n_298),
.B2(n_335),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_310),
.A2(n_264),
.B1(n_256),
.B2(n_275),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_368),
.A2(n_373),
.B1(n_332),
.B2(n_323),
.Y(n_388)
);

XNOR2x1_ASAP7_75t_L g372 ( 
.A(n_310),
.B(n_256),
.Y(n_372)
);

XOR2x2_ASAP7_75t_L g393 ( 
.A(n_372),
.B(n_374),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_326),
.A2(n_250),
.B1(n_260),
.B2(n_257),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_307),
.B(n_280),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g431 ( 
.A1(n_376),
.A2(n_390),
.B(n_398),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_352),
.B(n_314),
.Y(n_378)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_378),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g432 ( 
.A1(n_379),
.A2(n_383),
.B1(n_392),
.B2(n_397),
.Y(n_432)
);

BUFx12f_ASAP7_75t_L g380 ( 
.A(n_341),
.Y(n_380)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_380),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g381 ( 
.A1(n_361),
.A2(n_321),
.B(n_324),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_381),
.Y(n_418)
);

NOR3xp33_ASAP7_75t_L g429 ( 
.A(n_382),
.B(n_384),
.C(n_391),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_344),
.B(n_297),
.Y(n_384)
);

AND2x2_ASAP7_75t_SL g386 ( 
.A(n_370),
.B(n_324),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g425 ( 
.A1(n_386),
.A2(n_395),
.B(n_364),
.Y(n_425)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_388),
.Y(n_414)
);

OR2x2_ASAP7_75t_L g389 ( 
.A(n_370),
.B(n_252),
.Y(n_389)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_389),
.Y(n_416)
);

AOI21xp5_ASAP7_75t_L g390 ( 
.A1(n_366),
.A2(n_279),
.B(n_280),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_342),
.B(n_260),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_340),
.A2(n_315),
.B1(n_320),
.B2(n_279),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_358),
.B(n_257),
.Y(n_394)
);

NAND2x1p5_ASAP7_75t_L g438 ( 
.A(n_394),
.B(n_375),
.Y(n_438)
);

A2O1A1O1Ixp25_ASAP7_75t_L g395 ( 
.A1(n_348),
.A2(n_125),
.B(n_170),
.C(n_284),
.D(n_270),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_352),
.B(n_284),
.Y(n_396)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_396),
.Y(n_422)
);

AOI22xp33_ASAP7_75t_SL g397 ( 
.A1(n_365),
.A2(n_270),
.B1(n_234),
.B2(n_233),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_SL g398 ( 
.A1(n_366),
.A2(n_199),
.B(n_170),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_374),
.B(n_350),
.Y(n_399)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_399),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_350),
.B(n_0),
.Y(n_400)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_400),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_349),
.B(n_198),
.Y(n_401)
);

NOR3xp33_ASAP7_75t_L g430 ( 
.A(n_401),
.B(n_404),
.C(n_405),
.Y(n_430)
);

BUFx12f_ASAP7_75t_L g402 ( 
.A(n_343),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_402),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_340),
.A2(n_198),
.B1(n_184),
.B2(n_0),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_403),
.A2(n_338),
.B1(n_373),
.B2(n_371),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_349),
.B(n_184),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_355),
.B(n_359),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_355),
.B(n_7),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_406),
.B(n_407),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_356),
.B(n_7),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_357),
.B(n_0),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_408),
.B(n_368),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_346),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_409),
.A2(n_369),
.B1(n_340),
.B2(n_354),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_387),
.B(n_393),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_413),
.B(n_420),
.Y(n_458)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_417),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_378),
.B(n_356),
.Y(n_419)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_419),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_387),
.B(n_339),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_396),
.B(n_364),
.Y(n_421)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_421),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_L g452 ( 
.A1(n_423),
.A2(n_389),
.B1(n_408),
.B2(n_383),
.Y(n_452)
);

CKINVDCx16_ASAP7_75t_R g424 ( 
.A(n_382),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_424),
.B(n_440),
.Y(n_451)
);

AOI21xp5_ASAP7_75t_L g455 ( 
.A1(n_425),
.A2(n_398),
.B(n_394),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_399),
.B(n_337),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_426),
.B(n_435),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_377),
.B(n_372),
.C(n_363),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_427),
.B(n_384),
.C(n_391),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_410),
.B(n_371),
.Y(n_428)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_428),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_434),
.A2(n_388),
.B1(n_394),
.B2(n_386),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_393),
.B(n_345),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_385),
.A2(n_351),
.B1(n_367),
.B2(n_354),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_436),
.A2(n_389),
.B1(n_392),
.B2(n_403),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_L g463 ( 
.A1(n_438),
.A2(n_406),
.B(n_407),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_SL g439 ( 
.A(n_393),
.B(n_375),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_439),
.B(n_386),
.Y(n_448)
);

HAxp5_ASAP7_75t_SL g440 ( 
.A(n_376),
.B(n_375),
.CON(n_440),
.SN(n_440)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_410),
.B(n_360),
.Y(n_442)
);

CKINVDCx16_ASAP7_75t_R g457 ( 
.A(n_442),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_SL g443 ( 
.A(n_413),
.B(n_385),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_SL g473 ( 
.A(n_443),
.B(n_446),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_SL g446 ( 
.A(n_420),
.B(n_405),
.Y(n_446)
);

OAI31xp33_ASAP7_75t_L g447 ( 
.A1(n_416),
.A2(n_386),
.A3(n_381),
.B(n_390),
.Y(n_447)
);

AOI21xp5_ASAP7_75t_L g475 ( 
.A1(n_447),
.A2(n_463),
.B(n_431),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_448),
.B(n_459),
.Y(n_489)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_441),
.Y(n_449)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_449),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_450),
.A2(n_452),
.B1(n_434),
.B2(n_414),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_453),
.B(n_468),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_L g477 ( 
.A1(n_454),
.A2(n_460),
.B1(n_423),
.B2(n_436),
.Y(n_477)
);

INVxp67_ASAP7_75t_L g479 ( 
.A(n_455),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g456 ( 
.A(n_433),
.Y(n_456)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_456),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_SL g459 ( 
.A(n_426),
.B(n_435),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_414),
.A2(n_409),
.B1(n_395),
.B2(n_400),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_427),
.B(n_395),
.C(n_404),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_461),
.B(n_462),
.C(n_465),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_439),
.B(n_401),
.C(n_360),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_433),
.B(n_367),
.C(n_362),
.Y(n_465)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_422),
.Y(n_467)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_467),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_421),
.B(n_425),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_L g493 ( 
.A1(n_471),
.A2(n_482),
.B1(n_491),
.B2(n_454),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_445),
.B(n_429),
.Y(n_474)
);

CKINVDCx14_ASAP7_75t_R g497 ( 
.A(n_474),
.Y(n_497)
);

OAI21xp5_ASAP7_75t_L g507 ( 
.A1(n_475),
.A2(n_455),
.B(n_448),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_458),
.B(n_418),
.C(n_431),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_476),
.B(n_478),
.Y(n_506)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_477),
.B(n_460),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_458),
.B(n_418),
.C(n_442),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_446),
.B(n_419),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_481),
.B(n_490),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_450),
.A2(n_432),
.B1(n_416),
.B2(n_412),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_466),
.B(n_428),
.C(n_438),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_483),
.B(n_453),
.C(n_462),
.Y(n_503)
);

OAI21xp5_ASAP7_75t_SL g486 ( 
.A1(n_451),
.A2(n_430),
.B(n_412),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_486),
.B(n_487),
.Y(n_501)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_469),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_444),
.Y(n_488)
);

BUFx2_ASAP7_75t_L g494 ( 
.A(n_488),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_466),
.B(n_422),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_457),
.A2(n_437),
.B1(n_417),
.B2(n_438),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_464),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_492),
.B(n_437),
.Y(n_495)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_493),
.Y(n_517)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_495),
.Y(n_523)
);

AOI21xp33_ASAP7_75t_L g496 ( 
.A1(n_479),
.A2(n_463),
.B(n_461),
.Y(n_496)
);

OAI21xp33_ASAP7_75t_SL g520 ( 
.A1(n_496),
.A2(n_504),
.B(n_505),
.Y(n_520)
);

NOR3xp33_ASAP7_75t_SL g498 ( 
.A(n_484),
.B(n_411),
.C(n_447),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_498),
.B(n_500),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g515 ( 
.A(n_499),
.B(n_473),
.Y(n_515)
);

CKINVDCx16_ASAP7_75t_R g500 ( 
.A(n_491),
.Y(n_500)
);

BUFx12_ASAP7_75t_L g502 ( 
.A(n_478),
.Y(n_502)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_502),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_503),
.B(n_459),
.Y(n_518)
);

BUFx12f_ASAP7_75t_SL g504 ( 
.A(n_476),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_485),
.B(n_465),
.Y(n_505)
);

OAI21xp5_ASAP7_75t_L g512 ( 
.A1(n_507),
.A2(n_475),
.B(n_470),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_L g508 ( 
.A1(n_482),
.A2(n_443),
.B1(n_468),
.B2(n_415),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_508),
.A2(n_479),
.B1(n_493),
.B2(n_483),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_503),
.B(n_470),
.C(n_480),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g526 ( 
.A(n_510),
.B(n_513),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_SL g530 ( 
.A1(n_511),
.A2(n_508),
.B1(n_504),
.B2(n_499),
.Y(n_530)
);

OAI21xp5_ASAP7_75t_L g529 ( 
.A1(n_512),
.A2(n_507),
.B(n_514),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_506),
.B(n_480),
.C(n_490),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_SL g514 ( 
.A1(n_501),
.A2(n_471),
.B1(n_472),
.B2(n_481),
.Y(n_514)
);

AOI22xp33_ASAP7_75t_SL g528 ( 
.A1(n_514),
.A2(n_523),
.B1(n_511),
.B2(n_517),
.Y(n_528)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_515),
.Y(n_533)
);

OAI21x1_ASAP7_75t_L g525 ( 
.A1(n_518),
.A2(n_519),
.B(n_516),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g519 ( 
.A(n_509),
.B(n_473),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_505),
.B(n_489),
.C(n_362),
.Y(n_522)
);

CKINVDCx16_ASAP7_75t_R g527 ( 
.A(n_522),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_509),
.B(n_489),
.C(n_411),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_524),
.Y(n_534)
);

AOI21xp5_ASAP7_75t_L g541 ( 
.A1(n_525),
.A2(n_529),
.B(n_532),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_SL g540 ( 
.A1(n_528),
.A2(n_522),
.B1(n_524),
.B2(n_515),
.Y(n_540)
);

XOR2xp5_ASAP7_75t_L g542 ( 
.A(n_530),
.B(n_519),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_SL g531 ( 
.A1(n_521),
.A2(n_498),
.B1(n_495),
.B2(n_497),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_531),
.B(n_536),
.Y(n_537)
);

OAI21x1_ASAP7_75t_L g532 ( 
.A1(n_520),
.A2(n_502),
.B(n_494),
.Y(n_532)
);

OAI21xp5_ASAP7_75t_SL g535 ( 
.A1(n_512),
.A2(n_502),
.B(n_494),
.Y(n_535)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_535),
.Y(n_539)
);

FAx1_ASAP7_75t_SL g536 ( 
.A(n_510),
.B(n_380),
.CI(n_402),
.CON(n_536),
.SN(n_536)
);

AOI31xp67_ASAP7_75t_L g543 ( 
.A1(n_536),
.A2(n_380),
.A3(n_402),
.B(n_5),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_537),
.B(n_538),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_526),
.B(n_513),
.Y(n_538)
);

AOI322xp5_ASAP7_75t_L g547 ( 
.A1(n_540),
.A2(n_542),
.A3(n_543),
.B1(n_544),
.B2(n_535),
.C1(n_530),
.C2(n_531),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_SL g544 ( 
.A(n_526),
.B(n_402),
.Y(n_544)
);

OAI21xp5_ASAP7_75t_SL g545 ( 
.A1(n_541),
.A2(n_534),
.B(n_527),
.Y(n_545)
);

AOI21xp5_ASAP7_75t_L g550 ( 
.A1(n_545),
.A2(n_17),
.B(n_2),
.Y(n_550)
);

XNOR2x1_ASAP7_75t_L g552 ( 
.A(n_547),
.B(n_5),
.Y(n_552)
);

AOI322xp5_ASAP7_75t_L g548 ( 
.A1(n_539),
.A2(n_543),
.A3(n_536),
.B1(n_529),
.B2(n_533),
.C1(n_542),
.C2(n_402),
.Y(n_548)
);

AO21x1_ASAP7_75t_L g551 ( 
.A1(n_548),
.A2(n_549),
.B(n_1),
.Y(n_551)
);

AOI322xp5_ASAP7_75t_L g549 ( 
.A1(n_539),
.A2(n_380),
.A3(n_2),
.B1(n_5),
.B2(n_6),
.C1(n_10),
.C2(n_1),
.Y(n_549)
);

OAI21xp5_ASAP7_75t_SL g554 ( 
.A1(n_550),
.A2(n_546),
.B(n_14),
.Y(n_554)
);

AOI322xp5_ASAP7_75t_L g553 ( 
.A1(n_551),
.A2(n_552),
.A3(n_5),
.B1(n_10),
.B2(n_12),
.C1(n_14),
.C2(n_15),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_553),
.B(n_554),
.C(n_12),
.Y(n_555)
);

OAI21xp5_ASAP7_75t_L g556 ( 
.A1(n_555),
.A2(n_12),
.B(n_15),
.Y(n_556)
);

NAND3xp33_ASAP7_75t_L g557 ( 
.A(n_556),
.B(n_15),
.C(n_16),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_557),
.B(n_17),
.C(n_15),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_558),
.B(n_16),
.C(n_17),
.Y(n_559)
);


endmodule