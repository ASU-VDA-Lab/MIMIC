module fake_jpeg_30807_n_157 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_157);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_157;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_138;
wire n_101;
wire n_149;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_17),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_37),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_45),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_1),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_26),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

BUFx6f_ASAP7_75t_SL g61 ( 
.A(n_13),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_7),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_3),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_49),
.B(n_21),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

BUFx12_ASAP7_75t_L g67 ( 
.A(n_11),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_38),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_6),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_22),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_48),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_2),
.B(n_7),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_55),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_76),
.Y(n_87)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_73),
.B(n_0),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_70),
.Y(n_77)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_4),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_81),
.Y(n_89)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_79),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_65),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_52),
.B(n_4),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_82),
.B(n_51),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_82),
.B(n_63),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_88),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_77),
.B(n_50),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_93),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_83),
.B(n_56),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_91),
.B(n_94),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_80),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_75),
.B(n_59),
.Y(n_94)
);

INVx13_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_95),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_76),
.B(n_56),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_97),
.B(n_5),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_87),
.A2(n_72),
.B1(n_50),
.B2(n_59),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_98),
.A2(n_100),
.B1(n_15),
.B2(n_16),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_95),
.A2(n_62),
.B1(n_51),
.B2(n_72),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_92),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_114),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_97),
.B(n_60),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_102),
.B(n_108),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_87),
.A2(n_68),
.B(n_58),
.Y(n_105)
);

AND2x2_ASAP7_75t_SL g123 ( 
.A(n_105),
.B(n_8),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_91),
.A2(n_62),
.B(n_54),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_106),
.A2(n_110),
.B(n_116),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_53),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_107),
.B(n_109),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_71),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_96),
.A2(n_27),
.B(n_44),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_96),
.B(n_5),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_111),
.B(n_115),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_84),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_113),
.B(n_28),
.Y(n_120)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_86),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_97),
.B(n_6),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_87),
.A2(n_67),
.B(n_8),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_120),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_103),
.B(n_99),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_121),
.B(n_126),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_123),
.B(n_128),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_101),
.Y(n_124)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_124),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_104),
.B(n_67),
.Y(n_126)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_110),
.Y(n_127)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_127),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_105),
.B(n_9),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_112),
.A2(n_10),
.B1(n_12),
.B2(n_14),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_129),
.A2(n_127),
.B1(n_131),
.B2(n_123),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_130),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_100),
.A2(n_18),
.B1(n_20),
.B2(n_25),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_131),
.A2(n_31),
.B(n_32),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_43),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_132),
.B(n_30),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_116),
.B(n_29),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_SL g136 ( 
.A(n_133),
.B(n_125),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_136),
.B(n_140),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_142),
.A2(n_118),
.B(n_122),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_143),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_119),
.B(n_33),
.C(n_34),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_144),
.B(n_118),
.Y(n_147)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_134),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_145),
.B(n_146),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_147),
.B(n_137),
.C(n_135),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_150),
.B(n_152),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_147),
.B(n_139),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_153),
.B(n_141),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_154),
.A2(n_148),
.B(n_151),
.Y(n_155)
);

OAI321xp33_ASAP7_75t_L g156 ( 
.A1(n_155),
.A2(n_149),
.A3(n_138),
.B1(n_141),
.B2(n_117),
.C(n_39),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_156),
.B(n_41),
.Y(n_157)
);


endmodule