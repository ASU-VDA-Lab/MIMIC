module fake_jpeg_19833_n_101 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_101);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_101;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx8_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

INVx2_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

HB1xp67_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_18),
.B(n_0),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_24),
.B(n_26),
.Y(n_36)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_18),
.B(n_0),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_18),
.B(n_0),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_32),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_12),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_29)
);

A2O1A1Ixp33_ASAP7_75t_SL g51 ( 
.A1(n_29),
.A2(n_2),
.B(n_21),
.C(n_22),
.Y(n_51)
);

AND2x2_ASAP7_75t_SL g30 ( 
.A(n_22),
.B(n_1),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_30),
.B(n_14),
.C(n_19),
.Y(n_49)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_13),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_13),
.B(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_14),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_20),
.Y(n_40)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_32),
.Y(n_34)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_27),
.A2(n_12),
.B1(n_17),
.B2(n_16),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_38),
.A2(n_51),
.B1(n_20),
.B2(n_8),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_41),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g41 ( 
.A(n_24),
.Y(n_41)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_26),
.B(n_16),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_28),
.B(n_23),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_46),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_23),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_47),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_31),
.B(n_17),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_48),
.A2(n_50),
.B1(n_4),
.B2(n_10),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_4),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_29),
.B(n_15),
.Y(n_50)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_43),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_34),
.A2(n_30),
.B1(n_19),
.B2(n_15),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_55),
.A2(n_56),
.B1(n_58),
.B2(n_63),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_45),
.A2(n_30),
.B1(n_25),
.B2(n_21),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_51),
.A2(n_30),
.B1(n_20),
.B2(n_10),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_64),
.B(n_11),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_66),
.B(n_36),
.C(n_49),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_69),
.Y(n_82)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_37),
.Y(n_69)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_72),
.A2(n_73),
.B(n_74),
.Y(n_85)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_36),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_53),
.B(n_42),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_75),
.B(n_60),
.C(n_52),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_61),
.B(n_11),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_76),
.A2(n_77),
.B1(n_62),
.B2(n_42),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_57),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_81),
.C(n_39),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_79),
.B(n_39),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_69),
.A2(n_53),
.B1(n_51),
.B2(n_52),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_80),
.B(n_75),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_66),
.C(n_35),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_86),
.B(n_87),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_83),
.B(n_68),
.Y(n_87)
);

AOI221xp5_ASAP7_75t_L g88 ( 
.A1(n_82),
.A2(n_71),
.B1(n_75),
.B2(n_51),
.C(n_62),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_88),
.A2(n_82),
.B(n_85),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_89),
.B(n_90),
.C(n_81),
.Y(n_92)
);

MAJx2_ASAP7_75t_L g95 ( 
.A(n_91),
.B(n_51),
.C(n_54),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_92),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_88),
.B(n_78),
.C(n_84),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_94),
.B(n_35),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_95),
.A2(n_93),
.B(n_96),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_97),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_35),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_100),
.B(n_98),
.Y(n_101)
);


endmodule