module fake_jpeg_8424_n_39 (n_3, n_2, n_1, n_0, n_4, n_5, n_39);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_39;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g6 ( 
.A(n_2),
.Y(n_6)
);

INVx1_ASAP7_75t_L g7 ( 
.A(n_4),
.Y(n_7)
);

INVx3_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_L g9 ( 
.A(n_1),
.B(n_4),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

INVx6_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

INVx8_ASAP7_75t_L g12 ( 
.A(n_10),
.Y(n_12)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx6_ASAP7_75t_SL g13 ( 
.A(n_8),
.Y(n_13)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_9),
.B(n_0),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_14),
.B(n_15),
.Y(n_19)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_6),
.B(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_6),
.B(n_0),
.Y(n_17)
);

NOR2x1_ASAP7_75t_L g22 ( 
.A(n_17),
.B(n_7),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_22),
.B(n_7),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_19),
.B(n_15),
.C(n_14),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_25),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_18),
.B(n_16),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_24),
.B(n_26),
.Y(n_27)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_23),
.A2(n_21),
.B1(n_12),
.B2(n_11),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_SL g31 ( 
.A(n_28),
.B(n_11),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_29),
.B(n_20),
.C(n_13),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_30),
.B(n_32),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_31),
.A2(n_8),
.B1(n_12),
.B2(n_21),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_28),
.B(n_27),
.C(n_18),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_34),
.Y(n_35)
);

OR2x2_ASAP7_75t_L g36 ( 
.A(n_35),
.B(n_33),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_36),
.Y(n_37)
);

O2A1O1Ixp33_ASAP7_75t_SL g38 ( 
.A1(n_37),
.A2(n_10),
.B(n_1),
.C(n_5),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_38),
.B(n_5),
.Y(n_39)
);


endmodule