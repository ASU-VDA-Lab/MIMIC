module real_jpeg_18882_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_83;
wire n_78;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_292;
wire n_221;
wire n_249;
wire n_288;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_184;
wire n_56;
wire n_48;
wire n_164;
wire n_200;
wire n_293;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_188;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_298;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_205;
wire n_195;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_259;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_240;
wire n_297;
wire n_55;
wire n_185;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_209;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_216;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_244;
wire n_295;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_283;
wire n_85;
wire n_102;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;
wire n_16;

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_0),
.A2(n_165),
.B1(n_166),
.B2(n_168),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_0),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_0),
.A2(n_165),
.B1(n_240),
.B2(n_242),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_1),
.A2(n_62),
.B1(n_66),
.B2(n_67),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_1),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_1),
.A2(n_66),
.B1(n_184),
.B2(n_188),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_1),
.A2(n_66),
.B1(n_259),
.B2(n_261),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_3),
.Y(n_145)
);

BUFx5_ASAP7_75t_L g151 ( 
.A(n_3),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_3),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_3),
.Y(n_161)
);

OAI22x1_ASAP7_75t_SL g91 ( 
.A1(n_4),
.A2(n_92),
.B1(n_94),
.B2(n_95),
.Y(n_91)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_4),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_5),
.A2(n_129),
.B1(n_134),
.B2(n_135),
.Y(n_128)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_5),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_5),
.A2(n_117),
.B1(n_134),
.B2(n_175),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_6),
.A2(n_50),
.B1(n_55),
.B2(n_59),
.Y(n_49)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_6),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_6),
.A2(n_59),
.B1(n_231),
.B2(n_235),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_6),
.A2(n_59),
.B1(n_282),
.B2(n_283),
.Y(n_281)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_7),
.Y(n_88)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_7),
.Y(n_104)
);

BUFx5_ASAP7_75t_L g288 ( 
.A(n_7),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_8),
.B(n_71),
.Y(n_70)
);

OAI32xp33_ASAP7_75t_L g113 ( 
.A1(n_8),
.A2(n_24),
.A3(n_114),
.B1(n_117),
.B2(n_120),
.Y(n_113)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_8),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_8),
.A2(n_121),
.B1(n_196),
.B2(n_199),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_8),
.B(n_60),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_8),
.A2(n_85),
.B1(n_265),
.B2(n_281),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_9),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_9),
.Y(n_156)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_9),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_9),
.Y(n_191)
);

OAI22xp33_ASAP7_75t_L g105 ( 
.A1(n_10),
.A2(n_106),
.B1(n_107),
.B2(n_108),
.Y(n_105)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_10),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_11),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_11),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_12),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_13),
.Y(n_90)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_13),
.Y(n_100)
);

BUFx4f_ASAP7_75t_L g137 ( 
.A(n_13),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_13),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_206),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_205),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

NOR2xp67_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_179),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_18),
.B(n_179),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_20),
.B1(n_110),
.B2(n_111),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_69),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_48),
.B1(n_60),
.B2(n_61),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_23),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_23),
.A2(n_49),
.B1(n_195),
.B2(n_204),
.Y(n_194)
);

AO21x2_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_33),
.B(n_41),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_28),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_38),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_43),
.B1(n_45),
.B2(n_46),
.Y(n_41)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_42),
.Y(n_167)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_46),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVxp67_ASAP7_75t_SL g119 ( 
.A(n_47),
.Y(n_119)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx2_ASAP7_75t_SL g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_53),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_54),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_58),
.Y(n_198)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_60),
.Y(n_204)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_65),
.Y(n_68)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_65),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_83),
.Y(n_69)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

AOI22x1_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_76),
.B1(n_78),
.B2(n_81),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

AOI22x1_ASAP7_75t_SL g83 ( 
.A1(n_84),
.A2(n_91),
.B1(n_101),
.B2(n_105),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_84),
.A2(n_91),
.B1(n_128),
.B2(n_138),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_84),
.A2(n_257),
.B1(n_264),
.B2(n_266),
.Y(n_256)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_85),
.A2(n_239),
.B1(n_247),
.B2(n_248),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_85),
.A2(n_258),
.B1(n_281),
.B2(n_286),
.Y(n_285)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_89),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_88),
.Y(n_247)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_89),
.Y(n_106)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_89),
.Y(n_213)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_90),
.Y(n_93)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_90),
.Y(n_133)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_90),
.Y(n_146)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_90),
.Y(n_282)
);

BUFx2_ASAP7_75t_L g283 ( 
.A(n_92),
.Y(n_283)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_98),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_99),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_102),
.B(n_121),
.Y(n_279)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_103),
.Y(n_138)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_112),
.A2(n_139),
.B1(n_177),
.B2(n_178),
.Y(n_111)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_112),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_126),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_113),
.A2(n_126),
.B1(n_127),
.B2(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_113),
.Y(n_181)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_122),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_121),
.B(n_216),
.Y(n_215)
);

OAI21xp33_ASAP7_75t_SL g226 ( 
.A1(n_121),
.A2(n_215),
.B(n_227),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_121),
.B(n_172),
.Y(n_289)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_122),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_123),
.Y(n_176)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_128),
.Y(n_248)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_137),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_137),
.Y(n_241)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_138),
.Y(n_265)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_139),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_163),
.B1(n_172),
.B2(n_173),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_141),
.A2(n_164),
.B1(n_183),
.B2(n_192),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_141),
.A2(n_192),
.B1(n_226),
.B2(n_230),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_141),
.A2(n_183),
.B1(n_192),
.B2(n_230),
.Y(n_252)
);

AND2x2_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_152),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_142),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_146),
.B1(n_147),
.B2(n_150),
.Y(n_142)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_149),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g260 ( 
.A(n_149),
.Y(n_260)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_149),
.Y(n_278)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_151),
.Y(n_220)
);

OAI22xp33_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_157),
.B1(n_160),
.B2(n_162),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_155),
.Y(n_162)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_156),
.Y(n_171)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_160),
.Y(n_214)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_167),
.Y(n_229)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_172),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_182),
.C(n_193),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_180),
.B(n_296),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_182),
.A2(n_193),
.B1(n_194),
.B2(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_182),
.Y(n_297)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_187),
.Y(n_234)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_187),
.Y(n_236)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

BUFx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

BUFx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

AOI21x1_ASAP7_75t_SL g206 ( 
.A1(n_207),
.A2(n_293),
.B(n_298),
.Y(n_206)
);

OAI21x1_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_254),
.B(n_292),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_237),
.Y(n_208)
);

OR2x2_ASAP7_75t_L g292 ( 
.A(n_209),
.B(n_237),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_224),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_210),
.A2(n_224),
.B1(n_225),
.B2(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_210),
.Y(n_268)
);

OAI32xp33_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_213),
.A3(n_214),
.B1(n_215),
.B2(n_217),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_221),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_249),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_238),
.B(n_251),
.C(n_253),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_239),
.Y(n_266)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

BUFx2_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_252),
.B2(n_253),
.Y(n_249)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_250),
.Y(n_253)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_255),
.A2(n_269),
.B(n_291),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_267),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_256),
.B(n_267),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx2_ASAP7_75t_SL g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_284),
.B(n_290),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_280),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_279),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_289),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_285),
.B(n_289),
.Y(n_290)
);

INVx6_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

BUFx12f_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_294),
.B(n_295),
.Y(n_298)
);


endmodule