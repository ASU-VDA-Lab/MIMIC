module fake_jpeg_27492_n_270 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_270);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_270;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx11_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_17),
.B(n_8),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_40),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_25),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_32),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_30),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_30),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_42),
.B(n_22),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_43),
.B(n_46),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_41),
.A2(n_25),
.B1(n_23),
.B2(n_26),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_44),
.A2(n_19),
.B1(n_22),
.B2(n_24),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_40),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_34),
.A2(n_23),
.B1(n_16),
.B2(n_33),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_49),
.A2(n_60),
.B1(n_28),
.B2(n_27),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_20),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_50),
.B(n_56),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_34),
.A2(n_23),
.B1(n_16),
.B2(n_33),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_51),
.A2(n_18),
.B1(n_31),
.B2(n_20),
.Y(n_68)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_59),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_42),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_55),
.B(n_58),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_20),
.Y(n_56)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_37),
.A2(n_23),
.B1(n_31),
.B2(n_18),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

HAxp5_ASAP7_75t_SL g62 ( 
.A(n_39),
.B(n_17),
.CON(n_62),
.SN(n_62)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_62),
.B(n_29),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_37),
.A2(n_24),
.B1(n_22),
.B2(n_19),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_63),
.A2(n_27),
.B1(n_19),
.B2(n_28),
.Y(n_76)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_37),
.Y(n_73)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_65),
.B(n_69),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_46),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_67),
.B(n_81),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_68),
.B(n_77),
.Y(n_110)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_43),
.A2(n_50),
.B(n_60),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_70),
.A2(n_87),
.B(n_32),
.Y(n_108)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_49),
.A2(n_18),
.B1(n_31),
.B2(n_24),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_74),
.A2(n_75),
.B1(n_76),
.B2(n_78),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_53),
.A2(n_28),
.B1(n_27),
.B2(n_39),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_79),
.B(n_82),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_55),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_53),
.A2(n_39),
.B1(n_37),
.B2(n_29),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_88),
.Y(n_101)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_48),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_52),
.B(n_32),
.Y(n_88)
);

AOI32xp33_ASAP7_75t_L g90 ( 
.A1(n_87),
.A2(n_52),
.A3(n_39),
.B1(n_63),
.B2(n_26),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_90),
.A2(n_94),
.B(n_108),
.Y(n_131)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_91),
.B(n_95),
.Y(n_138)
);

AND2x6_ASAP7_75t_L g92 ( 
.A(n_87),
.B(n_15),
.Y(n_92)
);

AND2x6_ASAP7_75t_L g133 ( 
.A(n_92),
.B(n_10),
.Y(n_133)
);

OA21x2_ASAP7_75t_L g94 ( 
.A1(n_71),
.A2(n_59),
.B(n_56),
.Y(n_94)
);

INVx13_ASAP7_75t_L g95 ( 
.A(n_65),
.Y(n_95)
);

BUFx24_ASAP7_75t_SL g97 ( 
.A(n_85),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_97),
.Y(n_117)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_69),
.Y(n_98)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_71),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_99),
.B(n_100),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_80),
.B(n_26),
.Y(n_100)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_65),
.Y(n_102)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_102),
.Y(n_116)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

INVx13_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_105),
.Y(n_125)
);

AO22x1_ASAP7_75t_SL g107 ( 
.A1(n_70),
.A2(n_57),
.B1(n_64),
.B2(n_54),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_107),
.A2(n_76),
.B1(n_57),
.B2(n_79),
.Y(n_120)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_73),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_112),
.Y(n_132)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_78),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_80),
.B(n_32),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_94),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_112),
.A2(n_88),
.B1(n_86),
.B2(n_81),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_114),
.A2(n_120),
.B1(n_121),
.B2(n_124),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_110),
.A2(n_77),
.B1(n_74),
.B2(n_68),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_115),
.A2(n_118),
.B1(n_136),
.B2(n_91),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_110),
.A2(n_83),
.B1(n_67),
.B2(n_86),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_108),
.B(n_113),
.C(n_96),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_119),
.B(n_130),
.C(n_98),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_101),
.A2(n_61),
.B1(n_72),
.B2(n_45),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_101),
.A2(n_61),
.B1(n_72),
.B2(n_48),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_110),
.A2(n_72),
.B1(n_84),
.B2(n_85),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_127),
.A2(n_134),
.B1(n_120),
.B2(n_121),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_106),
.B(n_107),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_128),
.A2(n_129),
.B(n_135),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_96),
.A2(n_17),
.B1(n_29),
.B2(n_21),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_109),
.Y(n_130)
);

NAND3xp33_ASAP7_75t_L g156 ( 
.A(n_133),
.B(n_3),
.C(n_4),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_107),
.A2(n_29),
.B1(n_21),
.B2(n_32),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_94),
.A2(n_1),
.B(n_2),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_107),
.A2(n_32),
.B1(n_4),
.B2(n_5),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_137),
.B(n_94),
.Y(n_145)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_89),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_139),
.B(n_99),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_127),
.B(n_111),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_140),
.B(n_151),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_142),
.A2(n_148),
.B(n_149),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_126),
.B(n_111),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_143),
.B(n_144),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_145),
.B(n_146),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_132),
.B(n_100),
.Y(n_146)
);

A2O1A1O1Ixp25_ASAP7_75t_L g148 ( 
.A1(n_131),
.A2(n_90),
.B(n_92),
.C(n_103),
.D(n_93),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_131),
.A2(n_93),
.B(n_105),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_150),
.A2(n_128),
.B1(n_134),
.B2(n_136),
.Y(n_170)
);

INVx2_ASAP7_75t_SL g151 ( 
.A(n_123),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_132),
.B(n_91),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_152),
.A2(n_154),
.B(n_3),
.Y(n_181)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_138),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_153),
.B(n_158),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_135),
.A2(n_105),
.B(n_102),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_123),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_155),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_156),
.A2(n_165),
.B(n_133),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_157),
.B(n_115),
.C(n_125),
.Y(n_179)
);

OR2x2_ASAP7_75t_L g158 ( 
.A(n_126),
.B(n_32),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_139),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_159),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_137),
.B(n_102),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_160),
.B(n_161),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_130),
.B(n_95),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_124),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_162),
.B(n_163),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_129),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_122),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_164),
.Y(n_189)
);

AOI32xp33_ASAP7_75t_L g165 ( 
.A1(n_119),
.A2(n_95),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_165)
);

BUFx12f_ASAP7_75t_L g166 ( 
.A(n_116),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_166),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_168),
.A2(n_170),
.B1(n_166),
.B2(n_9),
.Y(n_207)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_152),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_171),
.B(n_175),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_157),
.B(n_161),
.C(n_149),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_172),
.B(n_179),
.C(n_147),
.Y(n_198)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_152),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_141),
.A2(n_128),
.B(n_118),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_176),
.A2(n_186),
.B(n_154),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_142),
.A2(n_125),
.B1(n_117),
.B2(n_7),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_180),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_R g201 ( 
.A(n_181),
.Y(n_201)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_160),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_182),
.B(n_185),
.Y(n_204)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_151),
.Y(n_185)
);

XOR2x2_ASAP7_75t_L g186 ( 
.A(n_145),
.B(n_6),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_190),
.A2(n_197),
.B(n_199),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_172),
.B(n_141),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_191),
.B(n_192),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_172),
.B(n_150),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_179),
.B(n_146),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_193),
.B(n_196),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_188),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_194),
.B(n_203),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_177),
.B(n_148),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_180),
.A2(n_163),
.B1(n_162),
.B2(n_147),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_198),
.B(n_185),
.C(n_167),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_170),
.A2(n_159),
.B1(n_158),
.B2(n_151),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_176),
.B(n_166),
.Y(n_200)
);

FAx1_ASAP7_75t_SL g214 ( 
.A(n_200),
.B(n_187),
.CI(n_181),
.CON(n_214),
.SN(n_214)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_202),
.A2(n_178),
.B1(n_169),
.B2(n_182),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_183),
.A2(n_168),
.B1(n_186),
.B2(n_184),
.Y(n_203)
);

BUFx4f_ASAP7_75t_SL g205 ( 
.A(n_173),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_205),
.Y(n_217)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_183),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_206),
.B(n_208),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_207),
.A2(n_186),
.B1(n_178),
.B2(n_189),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_184),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_187),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_209),
.B(n_175),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_194),
.A2(n_177),
.B(n_188),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_210),
.B(n_212),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_211),
.A2(n_174),
.B1(n_205),
.B2(n_155),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_214),
.B(n_191),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_196),
.B(n_169),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_215),
.B(n_216),
.Y(n_235)
);

AND2x4_ASAP7_75t_L g218 ( 
.A(n_200),
.B(n_171),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_218),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_220),
.B(n_204),
.C(n_201),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_202),
.B(n_166),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_224),
.B(n_225),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_193),
.B(n_167),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_226),
.B(n_227),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_213),
.B(n_198),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_213),
.B(n_192),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_228),
.B(n_230),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_220),
.B(n_195),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_231),
.B(n_234),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_223),
.B(n_197),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_233),
.B(n_218),
.Y(n_247)
);

FAx1_ASAP7_75t_SL g236 ( 
.A(n_212),
.B(n_205),
.CI(n_9),
.CON(n_236),
.SN(n_236)
);

FAx1_ASAP7_75t_SL g240 ( 
.A(n_236),
.B(n_211),
.CI(n_219),
.CON(n_240),
.SN(n_240)
);

OR2x2_ASAP7_75t_L g249 ( 
.A(n_240),
.B(n_241),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_229),
.A2(n_217),
.B1(n_210),
.B2(n_218),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_237),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_242),
.B(n_244),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_230),
.B(n_222),
.Y(n_243)
);

OR2x2_ASAP7_75t_L g252 ( 
.A(n_243),
.B(n_247),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_235),
.A2(n_218),
.B(n_214),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_236),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_245),
.B(n_242),
.Y(n_254)
);

CKINVDCx14_ASAP7_75t_R g248 ( 
.A(n_238),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_248),
.B(n_250),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_246),
.B(n_227),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_246),
.B(n_231),
.C(n_228),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_251),
.B(n_255),
.C(n_221),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_254),
.A2(n_240),
.B(n_214),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_239),
.B(n_226),
.C(n_221),
.Y(n_255)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_256),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_248),
.B(n_245),
.C(n_232),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_SL g263 ( 
.A(n_257),
.B(n_249),
.C(n_10),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_252),
.B(n_232),
.Y(n_258)
);

AOI31xp67_ASAP7_75t_SL g262 ( 
.A1(n_258),
.A2(n_259),
.A3(n_261),
.B(n_254),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_253),
.Y(n_261)
);

AOI322xp5_ASAP7_75t_L g267 ( 
.A1(n_262),
.A2(n_263),
.A3(n_11),
.B1(n_12),
.B2(n_13),
.C1(n_14),
.C2(n_15),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_260),
.A2(n_8),
.B1(n_11),
.B2(n_12),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_265),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_267),
.B(n_264),
.C(n_12),
.Y(n_268)
);

NOR2x1_ASAP7_75t_L g269 ( 
.A(n_268),
.B(n_266),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_269),
.B(n_15),
.Y(n_270)
);


endmodule