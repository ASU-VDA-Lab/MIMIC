module fake_jpeg_26352_n_396 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_396);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_396;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_12),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_40),
.Y(n_91)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_41),
.Y(n_84)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_43),
.Y(n_115)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_23),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_45),
.A2(n_34),
.B1(n_32),
.B2(n_28),
.Y(n_90)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_46),
.Y(n_95)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_49),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_51),
.B(n_54),
.Y(n_76)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_52),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_24),
.B(n_11),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_53),
.B(n_55),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_30),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_24),
.B(n_14),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_57),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_58),
.B(n_61),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_19),
.B(n_0),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_59),
.B(n_28),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_62),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_63),
.B(n_67),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g113 ( 
.A(n_64),
.Y(n_113)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_65),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_66),
.Y(n_114)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_68),
.Y(n_104)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_69),
.B(n_71),
.Y(n_97)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_22),
.Y(n_70)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_70),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_18),
.Y(n_71)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_73),
.B(n_37),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_56),
.A2(n_32),
.B1(n_34),
.B2(n_19),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_74),
.A2(n_42),
.B1(n_75),
.B2(n_40),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_59),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_79),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_61),
.A2(n_31),
.B1(n_33),
.B2(n_16),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_85),
.A2(n_86),
.B1(n_90),
.B2(n_17),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_52),
.A2(n_33),
.B1(n_17),
.B2(n_16),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_87),
.B(n_92),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_45),
.B(n_36),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_88),
.B(n_93),
.Y(n_128)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_43),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_54),
.A2(n_46),
.B1(n_49),
.B2(n_48),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_94),
.B(n_107),
.Y(n_133)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_68),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_101),
.B(n_109),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_106),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_70),
.B(n_36),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_57),
.B(n_29),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_111),
.B(n_112),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_72),
.B(n_29),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_116),
.A2(n_98),
.B1(n_82),
.B2(n_110),
.Y(n_168)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_117),
.B(n_120),
.Y(n_183)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_118),
.B(n_122),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_77),
.Y(n_119)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_119),
.Y(n_171)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_95),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_86),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_123),
.B(n_124),
.Y(n_193)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_91),
.Y(n_125)
);

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_125),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_107),
.B(n_25),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_126),
.B(n_136),
.Y(n_162)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_91),
.Y(n_129)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_129),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_100),
.B(n_50),
.C(n_66),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_130),
.B(n_3),
.C(n_5),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_103),
.A2(n_41),
.B1(n_104),
.B2(n_80),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_132),
.Y(n_160)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_89),
.Y(n_135)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_135),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_90),
.B(n_18),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_76),
.Y(n_137)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_137),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_75),
.A2(n_47),
.B1(n_25),
.B2(n_64),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_138),
.A2(n_1),
.B1(n_3),
.B2(n_5),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_103),
.A2(n_37),
.B1(n_26),
.B2(n_25),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_139),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_74),
.B(n_0),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_140),
.B(n_149),
.Y(n_186)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_115),
.Y(n_141)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_141),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_104),
.A2(n_26),
.B1(n_10),
.B2(n_11),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_142),
.Y(n_176)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_84),
.Y(n_144)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_144),
.Y(n_173)
);

A2O1A1Ixp33_ASAP7_75t_L g145 ( 
.A1(n_81),
.A2(n_73),
.B(n_60),
.C(n_58),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_145),
.B(n_151),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_78),
.A2(n_51),
.B(n_2),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_146),
.A2(n_8),
.B(n_133),
.Y(n_192)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_97),
.Y(n_147)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_147),
.Y(n_180)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_96),
.Y(n_148)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_148),
.Y(n_181)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_85),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g150 ( 
.A(n_98),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_150),
.B(n_144),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_84),
.B(n_71),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_99),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_152),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_99),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_153),
.Y(n_185)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_108),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_154),
.B(n_155),
.Y(n_188)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_108),
.Y(n_155)
);

AOI32xp33_ASAP7_75t_L g156 ( 
.A1(n_105),
.A2(n_71),
.A3(n_65),
.B1(n_63),
.B2(n_4),
.Y(n_156)
);

AOI32xp33_ASAP7_75t_L g169 ( 
.A1(n_156),
.A2(n_114),
.A3(n_113),
.B1(n_82),
.B2(n_4),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_77),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_157),
.Y(n_194)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_115),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_158),
.B(n_9),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_117),
.A2(n_80),
.B1(n_105),
.B2(n_83),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_159),
.Y(n_213)
);

OAI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_149),
.A2(n_83),
.B1(n_110),
.B2(n_102),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_163),
.A2(n_175),
.B1(n_184),
.B2(n_155),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_168),
.A2(n_189),
.B(n_192),
.Y(n_218)
);

OAI21xp33_ASAP7_75t_L g223 ( 
.A1(n_169),
.A2(n_178),
.B(n_190),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_143),
.A2(n_77),
.B1(n_113),
.B2(n_114),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_172),
.A2(n_174),
.B1(n_118),
.B2(n_124),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_135),
.A2(n_114),
.B1(n_113),
.B2(n_102),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_123),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_179),
.A2(n_152),
.B1(n_153),
.B2(n_150),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_182),
.B(n_184),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_136),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_133),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_187),
.A2(n_191),
.B1(n_196),
.B2(n_189),
.Y(n_201)
);

O2A1O1Ixp33_ASAP7_75t_L g189 ( 
.A1(n_140),
.A2(n_6),
.B(n_8),
.C(n_9),
.Y(n_189)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_190),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_133),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_195),
.A2(n_197),
.B(n_185),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_128),
.A2(n_121),
.B1(n_126),
.B2(n_154),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_198),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_180),
.B(n_127),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_199),
.B(n_200),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_180),
.B(n_148),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_201),
.B(n_205),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_181),
.B(n_137),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_203),
.B(n_206),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_162),
.B(n_134),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_204),
.B(n_212),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_181),
.B(n_166),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_188),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_207),
.B(n_219),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_186),
.A2(n_130),
.B1(n_146),
.B2(n_121),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_208),
.A2(n_209),
.B1(n_217),
.B2(n_220),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_186),
.A2(n_158),
.B1(n_122),
.B2(n_141),
.Y(n_209)
);

BUFx8_ASAP7_75t_L g210 ( 
.A(n_165),
.Y(n_210)
);

INVx6_ASAP7_75t_L g242 ( 
.A(n_210),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_166),
.B(n_147),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_211),
.B(n_214),
.Y(n_246)
);

OR2x2_ASAP7_75t_L g212 ( 
.A(n_178),
.B(n_145),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_164),
.B(n_131),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_162),
.B(n_125),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_215),
.B(n_231),
.Y(n_247)
);

INVx8_ASAP7_75t_L g216 ( 
.A(n_171),
.Y(n_216)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_216),
.Y(n_243)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_188),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_183),
.A2(n_129),
.B1(n_119),
.B2(n_157),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_192),
.B(n_196),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_221),
.B(n_224),
.Y(n_255)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_171),
.Y(n_222)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_222),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_223),
.A2(n_195),
.B(n_175),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_183),
.B(n_187),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_164),
.B(n_177),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_225),
.B(n_161),
.Y(n_253)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_165),
.Y(n_226)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_226),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_193),
.A2(n_160),
.B1(n_168),
.B2(n_170),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_227),
.A2(n_229),
.B1(n_232),
.B2(n_235),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_177),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_228),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_193),
.A2(n_179),
.B1(n_169),
.B2(n_176),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_230),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_191),
.B(n_189),
.Y(n_231)
);

BUFx2_ASAP7_75t_L g233 ( 
.A(n_173),
.Y(n_233)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_233),
.Y(n_251)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_197),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_234),
.B(n_209),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_163),
.A2(n_182),
.B1(n_185),
.B2(n_167),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_228),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_240),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_230),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_249),
.B(n_252),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_250),
.A2(n_231),
.B1(n_218),
.B2(n_212),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_233),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_253),
.B(n_262),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_221),
.B(n_195),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_254),
.B(n_232),
.C(n_224),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_212),
.A2(n_195),
.B(n_194),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_258),
.Y(n_271)
);

O2A1O1Ixp33_ASAP7_75t_L g259 ( 
.A1(n_213),
.A2(n_161),
.B(n_173),
.C(n_167),
.Y(n_259)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_259),
.Y(n_269)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_233),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_260),
.B(n_261),
.Y(n_270)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_216),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_222),
.B(n_216),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_263),
.B(n_247),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_215),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_266),
.B(n_267),
.Y(n_277)
);

BUFx24_ASAP7_75t_SL g267 ( 
.A(n_204),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_213),
.A2(n_218),
.B(n_227),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_268),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_236),
.A2(n_205),
.B1(n_219),
.B2(n_207),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_273),
.A2(n_288),
.B1(n_291),
.B2(n_293),
.Y(n_316)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_263),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_275),
.B(n_276),
.Y(n_305)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_259),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_278),
.B(n_280),
.Y(n_307)
);

INVx1_ASAP7_75t_SL g279 ( 
.A(n_247),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_279),
.B(n_282),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_268),
.Y(n_280)
);

XNOR2x1_ASAP7_75t_L g299 ( 
.A(n_281),
.B(n_250),
.Y(n_299)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_259),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_266),
.B(n_202),
.Y(n_284)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_284),
.Y(n_301)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_257),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_286),
.B(n_287),
.Y(n_302)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_257),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_236),
.A2(n_229),
.B1(n_235),
.B2(n_208),
.Y(n_288)
);

OA22x2_ASAP7_75t_L g289 ( 
.A1(n_237),
.A2(n_240),
.B1(n_238),
.B2(n_217),
.Y(n_289)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_289),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_290),
.B(n_295),
.C(n_255),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_238),
.A2(n_220),
.B1(n_234),
.B2(n_202),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_237),
.B(n_201),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_292),
.A2(n_256),
.B(n_258),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_249),
.A2(n_232),
.B1(n_226),
.B2(n_210),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_241),
.B(n_210),
.Y(n_294)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_294),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_255),
.B(n_210),
.C(n_254),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_270),
.Y(n_296)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_296),
.Y(n_331)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_297),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_285),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_298),
.B(n_265),
.Y(n_328)
);

XNOR2x2_ASAP7_75t_L g338 ( 
.A(n_299),
.B(n_289),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_300),
.B(n_304),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_290),
.B(n_239),
.C(n_241),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_304),
.B(n_309),
.C(n_314),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_270),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_306),
.B(n_308),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_277),
.B(n_264),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_295),
.B(n_239),
.C(n_251),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_272),
.A2(n_245),
.B(n_244),
.Y(n_310)
);

CKINVDCx14_ASAP7_75t_R g332 ( 
.A(n_310),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_274),
.B(n_246),
.Y(n_311)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_311),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_272),
.A2(n_280),
.B1(n_271),
.B2(n_292),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_313),
.B(n_317),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_288),
.B(n_251),
.C(n_260),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_271),
.A2(n_242),
.B1(n_252),
.B2(n_243),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_294),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_318),
.B(n_279),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_293),
.B(n_264),
.C(n_243),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_319),
.B(n_292),
.C(n_283),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_320),
.B(n_326),
.Y(n_354)
);

FAx1_ASAP7_75t_SL g324 ( 
.A(n_299),
.B(n_276),
.CI(n_284),
.CON(n_324),
.SN(n_324)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_324),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_325),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_326),
.B(n_329),
.C(n_314),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_298),
.B(n_273),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_327),
.B(n_334),
.Y(n_353)
);

INVxp33_ASAP7_75t_L g344 ( 
.A(n_328),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_309),
.B(n_287),
.C(n_286),
.Y(n_329)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_305),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_302),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_335),
.B(n_336),
.Y(n_346)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_305),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_319),
.B(n_248),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_SL g349 ( 
.A(n_337),
.B(n_301),
.Y(n_349)
);

XNOR2x1_ASAP7_75t_L g352 ( 
.A(n_338),
.B(n_313),
.Y(n_352)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_303),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_339),
.A2(n_275),
.B1(n_301),
.B2(n_312),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_341),
.B(n_351),
.C(n_320),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_323),
.B(n_300),
.C(n_315),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_342),
.B(n_343),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_323),
.B(n_315),
.C(n_317),
.Y(n_343)
);

INVxp33_ASAP7_75t_L g360 ( 
.A(n_345),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_L g348 ( 
.A1(n_338),
.A2(n_307),
.B(n_297),
.Y(n_348)
);

AOI211xp5_ASAP7_75t_L g355 ( 
.A1(n_348),
.A2(n_332),
.B(n_321),
.C(n_322),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_349),
.B(n_324),
.Y(n_365)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_322),
.A2(n_307),
.B(n_310),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_350),
.B(n_324),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_329),
.B(n_316),
.C(n_312),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_352),
.A2(n_339),
.B1(n_331),
.B2(n_334),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_354),
.B(n_316),
.Y(n_359)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_355),
.Y(n_374)
);

A2O1A1Ixp33_ASAP7_75t_SL g356 ( 
.A1(n_352),
.A2(n_289),
.B(n_321),
.C(n_269),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_356),
.A2(n_361),
.B1(n_364),
.B2(n_282),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_358),
.B(n_354),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_359),
.B(n_348),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_362),
.B(n_344),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_342),
.B(n_333),
.C(n_328),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_363),
.B(n_365),
.Y(n_371)
);

A2O1A1Ixp33_ASAP7_75t_SL g364 ( 
.A1(n_343),
.A2(n_289),
.B(n_278),
.C(n_269),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_341),
.B(n_330),
.C(n_336),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_366),
.B(n_353),
.Y(n_373)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_367),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_368),
.B(n_369),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_357),
.B(n_351),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_364),
.B(n_346),
.C(n_340),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_370),
.B(n_375),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_SL g372 ( 
.A1(n_365),
.A2(n_347),
.B(n_350),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_372),
.A2(n_373),
.B(n_364),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_376),
.B(n_370),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_377),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_371),
.B(n_360),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_378),
.B(n_380),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_374),
.B(n_248),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_SL g389 ( 
.A(n_382),
.B(n_344),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_368),
.B(n_356),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_383),
.B(n_367),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_379),
.B(n_369),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_386),
.B(n_389),
.Y(n_391)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_387),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_SL g390 ( 
.A1(n_385),
.A2(n_378),
.B(n_381),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_390),
.B(n_388),
.Y(n_393)
);

AOI322xp5_ASAP7_75t_L g394 ( 
.A1(n_393),
.A2(n_385),
.A3(n_392),
.B1(n_391),
.B2(n_384),
.C1(n_242),
.C2(n_261),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_L g395 ( 
.A1(n_394),
.A2(n_265),
.B(n_356),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_395),
.B(n_242),
.Y(n_396)
);


endmodule