module real_aes_9784_n_6 (n_4, n_0, n_3, n_5, n_2, n_1, n_6);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_1;
output n_6;
wire n_17;
wire n_22;
wire n_13;
wire n_24;
wire n_12;
wire n_19;
wire n_25;
wire n_14;
wire n_11;
wire n_16;
wire n_15;
wire n_9;
wire n_23;
wire n_20;
wire n_26;
wire n_18;
wire n_21;
wire n_7;
wire n_8;
wire n_10;
AOI21xp33_ASAP7_75t_L g16 ( .A1(n_0), .A2(n_1), .B(n_2), .Y(n_16) );
INVx1_ASAP7_75t_L g23 ( .A(n_0), .Y(n_23) );
INVx1_ASAP7_75t_L g12 ( .A(n_1), .Y(n_12) );
AOI21xp5_ASAP7_75t_L g13 ( .A1(n_1), .A2(n_14), .B(n_15), .Y(n_13) );
AND2x2_ASAP7_75t_L g25 ( .A(n_2), .B(n_26), .Y(n_25) );
INVx1_ASAP7_75t_L g14 ( .A(n_3), .Y(n_14) );
AND2x2_ASAP7_75t_L g15 ( .A(n_3), .B(n_12), .Y(n_15) );
BUFx2_ASAP7_75t_L g11 ( .A(n_4), .Y(n_11) );
INVx1_ASAP7_75t_L g24 ( .A(n_4), .Y(n_24) );
O2A1O1Ixp33_ASAP7_75t_R g6 ( .A1(n_5), .A2(n_7), .B(n_16), .C(n_17), .Y(n_6) );
INVx1_ASAP7_75t_L g26 ( .A(n_5), .Y(n_26) );
CKINVDCx20_ASAP7_75t_R g7 ( .A(n_8), .Y(n_7) );
AOI21xp5_ASAP7_75t_L g8 ( .A1(n_9), .A2(n_12), .B(n_13), .Y(n_8) );
INVx1_ASAP7_75t_L g9 ( .A(n_10), .Y(n_9) );
BUFx8_ASAP7_75t_SL g10 ( .A(n_11), .Y(n_10) );
INVx4_ASAP7_75t_L g22 ( .A(n_15), .Y(n_22) );
INVx2_ASAP7_75t_L g17 ( .A(n_18), .Y(n_17) );
BUFx12f_ASAP7_75t_L g18 ( .A(n_19), .Y(n_18) );
INVx4_ASAP7_75t_L g19 ( .A(n_20), .Y(n_19) );
AND2x2_ASAP7_75t_SL g20 ( .A(n_21), .B(n_25), .Y(n_20) );
NOR3xp33_ASAP7_75t_L g21 ( .A(n_22), .B(n_23), .C(n_24), .Y(n_21) );
endmodule