module fake_jpeg_11061_n_525 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_525);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_525;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_387;
wire n_270;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_393;
wire n_288;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_2),
.B(n_17),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_15),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_7),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_17),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_16),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_12),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_0),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_5),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_9),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_9),
.Y(n_55)
);

BUFx24_ASAP7_75t_L g56 ( 
.A(n_8),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_57),
.Y(n_126)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_58),
.Y(n_130)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_59),
.Y(n_140)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_60),
.Y(n_124)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_56),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_61),
.Y(n_148)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_22),
.B(n_0),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_62),
.B(n_63),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_35),
.B(n_2),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_64),
.Y(n_143)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_65),
.Y(n_179)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_56),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_66),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_67),
.Y(n_150)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g139 ( 
.A(n_68),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_69),
.Y(n_134)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_28),
.Y(n_70)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_70),
.Y(n_147)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_71),
.Y(n_132)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_25),
.Y(n_72)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_72),
.Y(n_133)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_25),
.Y(n_73)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_73),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_74),
.Y(n_142)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_75),
.Y(n_145)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_19),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_76),
.Y(n_153)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_28),
.Y(n_77)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_77),
.Y(n_164)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_28),
.Y(n_78)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_78),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_35),
.B(n_3),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_79),
.B(n_91),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_45),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_80),
.A2(n_50),
.B1(n_52),
.B2(n_32),
.Y(n_131)
);

INVx4_ASAP7_75t_SL g81 ( 
.A(n_56),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_81),
.Y(n_163)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_22),
.Y(n_82)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_82),
.Y(n_123)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_83),
.Y(n_183)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_30),
.Y(n_84)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_84),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_85),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_19),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_86),
.Y(n_167)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_36),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_87),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_36),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_88),
.Y(n_192)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_20),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_89),
.Y(n_171)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_30),
.Y(n_90)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_90),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_45),
.B(n_16),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_23),
.Y(n_92)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_92),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_36),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_93),
.Y(n_201)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_30),
.Y(n_94)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_94),
.Y(n_157)
);

INVx3_ASAP7_75t_SL g95 ( 
.A(n_20),
.Y(n_95)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_95),
.Y(n_186)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_41),
.Y(n_96)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_96),
.Y(n_188)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_97),
.Y(n_169)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_20),
.Y(n_98)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_98),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_34),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_99),
.B(n_111),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_36),
.Y(n_100)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_100),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_43),
.Y(n_101)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_101),
.Y(n_136)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_20),
.Y(n_102)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_102),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_55),
.Y(n_103)
);

INVx5_ASAP7_75t_L g177 ( 
.A(n_103),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_43),
.Y(n_104)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_104),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_55),
.Y(n_105)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_105),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_43),
.Y(n_106)
);

INVx6_ASAP7_75t_L g187 ( 
.A(n_106),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_43),
.Y(n_107)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_107),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_53),
.Y(n_108)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_108),
.Y(n_129)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_20),
.Y(n_109)
);

BUFx2_ASAP7_75t_L g175 ( 
.A(n_109),
.Y(n_175)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_41),
.Y(n_110)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_110),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_50),
.B(n_4),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_55),
.Y(n_112)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_112),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_50),
.B(n_5),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_113),
.B(n_119),
.Y(n_158)
);

BUFx5_ASAP7_75t_L g114 ( 
.A(n_20),
.Y(n_114)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_114),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_53),
.Y(n_115)
);

INVx8_ASAP7_75t_L g162 ( 
.A(n_115),
.Y(n_162)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_53),
.Y(n_116)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_116),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_53),
.Y(n_117)
);

INVx8_ASAP7_75t_L g173 ( 
.A(n_117),
.Y(n_173)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_18),
.Y(n_118)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_118),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_21),
.B(n_6),
.Y(n_119)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_18),
.Y(n_120)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_120),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_18),
.Y(n_121)
);

INVx3_ASAP7_75t_SL g160 ( 
.A(n_121),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_62),
.A2(n_42),
.B1(n_52),
.B2(n_38),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_122),
.A2(n_154),
.B1(n_200),
.B2(n_44),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_111),
.B(n_32),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_125),
.B(n_155),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_113),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_128),
.B(n_135),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_131),
.A2(n_37),
.B1(n_54),
.B2(n_24),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_69),
.B(n_26),
.Y(n_135)
);

INVxp67_ASAP7_75t_SL g138 ( 
.A(n_81),
.Y(n_138)
);

INVx11_ASAP7_75t_L g246 ( 
.A(n_138),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_76),
.A2(n_26),
.B1(n_48),
.B2(n_21),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_61),
.B(n_31),
.Y(n_155)
);

INVx2_ASAP7_75t_SL g161 ( 
.A(n_69),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_161),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_66),
.B(n_31),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_168),
.B(n_172),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_85),
.B(n_33),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_68),
.A2(n_29),
.B1(n_49),
.B2(n_47),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_180),
.A2(n_199),
.B(n_49),
.Y(n_242)
);

INVx2_ASAP7_75t_SL g185 ( 
.A(n_105),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_185),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_89),
.B(n_33),
.Y(n_190)
);

A2O1A1Ixp33_ASAP7_75t_L g225 ( 
.A1(n_190),
.A2(n_37),
.B(n_54),
.C(n_23),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_116),
.B(n_38),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_193),
.B(n_46),
.Y(n_244)
);

INVx2_ASAP7_75t_SL g196 ( 
.A(n_95),
.Y(n_196)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_196),
.Y(n_204)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_87),
.Y(n_197)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_197),
.Y(n_206)
);

INVx2_ASAP7_75t_SL g198 ( 
.A(n_109),
.Y(n_198)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_198),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_121),
.A2(n_29),
.B1(n_49),
.B2(n_47),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_64),
.A2(n_44),
.B1(n_48),
.B2(n_46),
.Y(n_200)
);

BUFx2_ASAP7_75t_L g202 ( 
.A(n_152),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_202),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_203),
.B(n_235),
.Y(n_296)
);

INVx5_ASAP7_75t_L g205 ( 
.A(n_134),
.Y(n_205)
);

INVx4_ASAP7_75t_L g312 ( 
.A(n_205),
.Y(n_312)
);

BUFx3_ASAP7_75t_L g207 ( 
.A(n_161),
.Y(n_207)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_207),
.Y(n_269)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_123),
.Y(n_210)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_210),
.Y(n_281)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_159),
.Y(n_211)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_211),
.Y(n_284)
);

INVx6_ASAP7_75t_L g213 ( 
.A(n_127),
.Y(n_213)
);

INVx8_ASAP7_75t_L g279 ( 
.A(n_213),
.Y(n_279)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_181),
.Y(n_214)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_214),
.Y(n_286)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_165),
.Y(n_215)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_215),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_152),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_218),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_158),
.A2(n_117),
.B1(n_115),
.B2(n_108),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_219),
.A2(n_227),
.B1(n_163),
.B2(n_160),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_136),
.A2(n_107),
.B1(n_106),
.B2(n_104),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_220),
.A2(n_232),
.B1(n_239),
.B2(n_258),
.Y(n_302)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_138),
.Y(n_221)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_221),
.Y(n_299)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_186),
.Y(n_222)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_222),
.Y(n_301)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_182),
.Y(n_223)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_223),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_225),
.B(n_228),
.Y(n_285)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_156),
.Y(n_226)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_226),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_190),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_126),
.Y(n_229)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_229),
.Y(n_277)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_178),
.Y(n_230)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_230),
.Y(n_282)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_130),
.Y(n_231)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_231),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_L g232 ( 
.A1(n_174),
.A2(n_101),
.B1(n_100),
.B2(n_93),
.Y(n_232)
);

INVx6_ASAP7_75t_L g233 ( 
.A(n_187),
.Y(n_233)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_233),
.Y(n_319)
);

XNOR2x1_ASAP7_75t_L g234 ( 
.A(n_146),
.B(n_158),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_234),
.B(n_264),
.Y(n_298)
);

INVx2_ASAP7_75t_SL g235 ( 
.A(n_148),
.Y(n_235)
);

INVx6_ASAP7_75t_L g236 ( 
.A(n_195),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_236),
.B(n_237),
.Y(n_311)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_140),
.Y(n_237)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_124),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_238),
.B(n_243),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_147),
.A2(n_88),
.B1(n_86),
.B2(n_67),
.Y(n_239)
);

INVx2_ASAP7_75t_SL g240 ( 
.A(n_177),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_240),
.Y(n_314)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_132),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_241),
.Y(n_287)
);

O2A1O1Ixp33_ASAP7_75t_L g275 ( 
.A1(n_242),
.A2(n_253),
.B(n_139),
.C(n_160),
.Y(n_275)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_133),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_244),
.B(n_248),
.Y(n_310)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_137),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_245),
.Y(n_291)
);

INVx6_ASAP7_75t_L g247 ( 
.A(n_143),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g305 ( 
.A1(n_247),
.A2(n_252),
.B1(n_254),
.B2(n_255),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_146),
.B(n_39),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_149),
.B(n_39),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_249),
.B(n_259),
.Y(n_315)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_164),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_250),
.Y(n_272)
);

INVx4_ASAP7_75t_L g251 ( 
.A(n_145),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_251),
.Y(n_280)
);

INVx5_ASAP7_75t_L g252 ( 
.A(n_142),
.Y(n_252)
);

OA22x2_ASAP7_75t_L g253 ( 
.A1(n_149),
.A2(n_47),
.B1(n_29),
.B2(n_24),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_143),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_179),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_166),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_256),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_150),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_257),
.A2(n_260),
.B1(n_265),
.B2(n_266),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_169),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_144),
.B(n_7),
.Y(n_259)
);

INVx5_ASAP7_75t_L g260 ( 
.A(n_170),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_144),
.B(n_8),
.Y(n_261)
);

BUFx24_ASAP7_75t_SL g297 ( 
.A(n_261),
.Y(n_297)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_183),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_262),
.B(n_10),
.Y(n_317)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_176),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_263),
.B(n_267),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_188),
.B(n_9),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_150),
.Y(n_265)
);

BUFx12f_ASAP7_75t_L g266 ( 
.A(n_163),
.Y(n_266)
);

INVx4_ASAP7_75t_L g267 ( 
.A(n_129),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_196),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_268),
.B(n_185),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_216),
.A2(n_199),
.B1(n_180),
.B2(n_184),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_271),
.A2(n_290),
.B1(n_293),
.B2(n_294),
.Y(n_349)
);

NAND2xp33_ASAP7_75t_SL g348 ( 
.A(n_273),
.B(n_275),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_264),
.A2(n_184),
.B1(n_153),
.B2(n_173),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_274),
.A2(n_313),
.B1(n_246),
.B2(n_247),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_217),
.A2(n_139),
.B(n_151),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_289),
.A2(n_308),
.B(n_207),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_232),
.A2(n_153),
.B1(n_192),
.B2(n_167),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_209),
.A2(n_167),
.B1(n_192),
.B2(n_201),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_253),
.A2(n_201),
.B1(n_162),
.B2(n_191),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g322 ( 
.A(n_304),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_253),
.B(n_189),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_306),
.B(n_309),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_258),
.A2(n_157),
.B1(n_141),
.B2(n_198),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_307),
.A2(n_316),
.B1(n_40),
.B2(n_12),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_246),
.A2(n_175),
.B(n_171),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_206),
.B(n_10),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_213),
.A2(n_175),
.B1(n_171),
.B2(n_194),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_255),
.A2(n_233),
.B1(n_236),
.B2(n_208),
.Y(n_316)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_317),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_299),
.Y(n_321)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_321),
.Y(n_359)
);

INVxp67_ASAP7_75t_SL g386 ( 
.A(n_323),
.Y(n_386)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_299),
.Y(n_324)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_324),
.Y(n_360)
);

AO22x1_ASAP7_75t_SL g325 ( 
.A1(n_275),
.A2(n_204),
.B1(n_202),
.B2(n_267),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_325),
.B(n_351),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_295),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_326),
.B(n_338),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_298),
.B(n_218),
.C(n_224),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_327),
.B(n_330),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_306),
.A2(n_265),
.B1(n_257),
.B2(n_254),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_328),
.A2(n_336),
.B1(n_347),
.B2(n_354),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_279),
.Y(n_329)
);

INVx3_ASAP7_75t_L g375 ( 
.A(n_329),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_298),
.B(n_224),
.C(n_212),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_285),
.B(n_315),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_331),
.Y(n_378)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_276),
.Y(n_332)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_332),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_296),
.B(n_212),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_333),
.B(n_342),
.Y(n_380)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_278),
.Y(n_334)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_334),
.Y(n_384)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_276),
.Y(n_335)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_335),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_273),
.A2(n_251),
.B1(n_241),
.B2(n_240),
.Y(n_336)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_301),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_304),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_339),
.B(n_345),
.Y(n_368)
);

AOI22xp33_ASAP7_75t_L g340 ( 
.A1(n_294),
.A2(n_230),
.B1(n_226),
.B2(n_235),
.Y(n_340)
);

AOI22xp33_ASAP7_75t_SL g365 ( 
.A1(n_340),
.A2(n_344),
.B1(n_307),
.B2(n_316),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_310),
.B(n_266),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_341),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_296),
.B(n_266),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g372 ( 
.A1(n_343),
.A2(n_300),
.B(n_287),
.Y(n_372)
);

AOI22xp33_ASAP7_75t_SL g344 ( 
.A1(n_271),
.A2(n_34),
.B1(n_40),
.B2(n_13),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_301),
.Y(n_345)
);

NAND2x1_ASAP7_75t_SL g346 ( 
.A(n_289),
.B(n_34),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_L g361 ( 
.A1(n_346),
.A2(n_343),
.B(n_348),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_274),
.A2(n_34),
.B1(n_40),
.B2(n_13),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_281),
.B(n_10),
.Y(n_350)
);

CKINVDCx14_ASAP7_75t_R g373 ( 
.A(n_350),
.Y(n_373)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_281),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_278),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_352),
.B(n_353),
.Y(n_383)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_284),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_296),
.A2(n_34),
.B1(n_40),
.B2(n_14),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_355),
.A2(n_300),
.B1(n_313),
.B2(n_309),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_305),
.A2(n_40),
.B1(n_12),
.B2(n_14),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_356),
.A2(n_314),
.B1(n_312),
.B2(n_280),
.Y(n_382)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_284),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_357),
.B(n_358),
.Y(n_385)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_286),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_L g396 ( 
.A1(n_361),
.A2(n_367),
.B(n_370),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_336),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_362),
.B(n_354),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_364),
.A2(n_386),
.B1(n_362),
.B2(n_328),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_365),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_L g367 ( 
.A1(n_346),
.A2(n_308),
.B(n_318),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_332),
.A2(n_302),
.B1(n_293),
.B2(n_290),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_372),
.B(n_387),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_L g376 ( 
.A1(n_346),
.A2(n_317),
.B(n_286),
.Y(n_376)
);

CKINVDCx16_ASAP7_75t_R g400 ( 
.A(n_376),
.Y(n_400)
);

MAJx2_ASAP7_75t_L g377 ( 
.A(n_330),
.B(n_297),
.C(n_311),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_377),
.B(n_327),
.C(n_320),
.Y(n_399)
);

O2A1O1Ixp33_ASAP7_75t_L g381 ( 
.A1(n_325),
.A2(n_287),
.B(n_291),
.C(n_280),
.Y(n_381)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_381),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_382),
.A2(n_390),
.B1(n_355),
.B2(n_352),
.Y(n_398)
);

AO22x1_ASAP7_75t_SL g387 ( 
.A1(n_322),
.A2(n_319),
.B1(n_303),
.B2(n_277),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_339),
.B(n_283),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_388),
.B(n_345),
.Y(n_412)
);

AOI22xp33_ASAP7_75t_SL g390 ( 
.A1(n_334),
.A2(n_292),
.B1(n_312),
.B2(n_282),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_SL g391 ( 
.A(n_378),
.B(n_320),
.Y(n_391)
);

NAND3xp33_ASAP7_75t_L g434 ( 
.A(n_391),
.B(n_373),
.C(n_360),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_393),
.A2(n_410),
.B1(n_414),
.B2(n_416),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_370),
.A2(n_349),
.B1(n_335),
.B2(n_337),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_397),
.A2(n_398),
.B1(n_403),
.B2(n_406),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_399),
.B(n_270),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_369),
.B(n_380),
.C(n_377),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_401),
.B(n_404),
.C(n_377),
.Y(n_418)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_375),
.Y(n_402)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_402),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_386),
.A2(n_349),
.B1(n_337),
.B2(n_322),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_369),
.B(n_333),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_385),
.Y(n_405)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_405),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_374),
.A2(n_325),
.B1(n_342),
.B2(n_324),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_374),
.A2(n_321),
.B1(n_323),
.B2(n_358),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_407),
.A2(n_415),
.B1(n_403),
.B2(n_359),
.Y(n_430)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_385),
.Y(n_408)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_408),
.Y(n_431)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_409),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_364),
.A2(n_347),
.B1(n_356),
.B2(n_353),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_366),
.Y(n_411)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_411),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_412),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_SL g413 ( 
.A(n_380),
.B(n_357),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_SL g421 ( 
.A(n_413),
.B(n_368),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_381),
.A2(n_351),
.B1(n_338),
.B2(n_326),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_371),
.A2(n_319),
.B1(n_329),
.B2(n_279),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_381),
.A2(n_329),
.B1(n_283),
.B2(n_272),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_366),
.Y(n_417)
);

AOI22xp33_ASAP7_75t_SL g437 ( 
.A1(n_417),
.A2(n_384),
.B1(n_387),
.B2(n_292),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_418),
.B(n_401),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_L g419 ( 
.A1(n_396),
.A2(n_361),
.B(n_367),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_419),
.B(n_422),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_393),
.A2(n_363),
.B1(n_389),
.B2(n_371),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_420),
.A2(n_423),
.B1(n_432),
.B2(n_406),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_SL g449 ( 
.A(n_421),
.B(n_427),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_SL g422 ( 
.A1(n_395),
.A2(n_368),
.B(n_388),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_410),
.A2(n_389),
.B1(n_363),
.B2(n_376),
.Y(n_423)
);

OA22x2_ASAP7_75t_L g424 ( 
.A1(n_392),
.A2(n_382),
.B1(n_372),
.B2(n_387),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_424),
.B(n_434),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_SL g427 ( 
.A(n_404),
.B(n_379),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_391),
.B(n_373),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_SL g452 ( 
.A(n_429),
.B(n_411),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_L g455 ( 
.A1(n_430),
.A2(n_437),
.B1(n_439),
.B2(n_409),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_392),
.A2(n_359),
.B1(n_360),
.B2(n_383),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_397),
.A2(n_383),
.B1(n_375),
.B2(n_387),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_436),
.A2(n_440),
.B1(n_416),
.B2(n_414),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_L g439 ( 
.A1(n_394),
.A2(n_384),
.B1(n_272),
.B2(n_303),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_407),
.A2(n_282),
.B1(n_269),
.B2(n_277),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_442),
.B(n_413),
.C(n_399),
.Y(n_448)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_443),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_444),
.B(n_447),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_446),
.B(n_448),
.C(n_454),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_428),
.A2(n_408),
.B1(n_405),
.B2(n_396),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_427),
.B(n_417),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_450),
.B(n_460),
.Y(n_465)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_438),
.Y(n_451)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_451),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_452),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_418),
.B(n_400),
.C(n_412),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_455),
.B(n_459),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_426),
.A2(n_395),
.B1(n_400),
.B2(n_398),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_456),
.B(n_457),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_L g457 ( 
.A1(n_426),
.A2(n_415),
.B1(n_402),
.B2(n_291),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_442),
.B(n_269),
.C(n_270),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_458),
.B(n_440),
.C(n_425),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_L g459 ( 
.A1(n_433),
.A2(n_288),
.B1(n_10),
.B2(n_16),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_421),
.B(n_288),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_420),
.A2(n_16),
.B1(n_433),
.B2(n_423),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_461),
.B(n_462),
.Y(n_469)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_438),
.Y(n_462)
);

AOI21xp5_ASAP7_75t_L g466 ( 
.A1(n_453),
.A2(n_422),
.B(n_419),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_SL g482 ( 
.A1(n_466),
.A2(n_445),
.B(n_443),
.Y(n_482)
);

XOR2x1_ASAP7_75t_L g467 ( 
.A(n_447),
.B(n_436),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_467),
.B(n_472),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_454),
.B(n_425),
.C(n_431),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_475),
.B(n_476),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_446),
.B(n_431),
.C(n_430),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_SL g477 ( 
.A(n_452),
.B(n_441),
.Y(n_477)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_477),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_470),
.A2(n_444),
.B1(n_456),
.B2(n_457),
.Y(n_479)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_479),
.Y(n_490)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_463),
.Y(n_480)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_480),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_469),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_481),
.B(n_482),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_473),
.A2(n_461),
.B1(n_441),
.B2(n_451),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_483),
.B(n_487),
.Y(n_494)
);

BUFx24_ASAP7_75t_SL g485 ( 
.A(n_464),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_SL g492 ( 
.A(n_485),
.B(n_488),
.Y(n_492)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_475),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_474),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_470),
.A2(n_462),
.B1(n_424),
.B2(n_432),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_489),
.B(n_467),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_SL g493 ( 
.A(n_478),
.B(n_465),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_493),
.B(n_499),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_484),
.B(n_478),
.C(n_471),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_496),
.B(n_498),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_SL g497 ( 
.A(n_486),
.B(n_466),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_497),
.B(n_465),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_484),
.B(n_471),
.C(n_476),
.Y(n_498)
);

NAND4xp25_ASAP7_75t_L g500 ( 
.A(n_495),
.B(n_494),
.C(n_490),
.D(n_491),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_500),
.B(n_501),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_496),
.B(n_482),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_SL g509 ( 
.A(n_503),
.B(n_506),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_498),
.B(n_483),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_504),
.B(n_505),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_493),
.B(n_479),
.C(n_474),
.Y(n_505)
);

OAI21xp5_ASAP7_75t_L g506 ( 
.A1(n_492),
.A2(n_489),
.B(n_448),
.Y(n_506)
);

OAI21x1_ASAP7_75t_L g508 ( 
.A1(n_502),
.A2(n_468),
.B(n_424),
.Y(n_508)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_508),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_507),
.B(n_472),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_510),
.B(n_511),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_505),
.B(n_499),
.C(n_458),
.Y(n_511)
);

AOI21xp5_ASAP7_75t_SL g514 ( 
.A1(n_513),
.A2(n_507),
.B(n_480),
.Y(n_514)
);

AOI31xp33_ASAP7_75t_L g518 ( 
.A1(n_514),
.A2(n_512),
.A3(n_509),
.B(n_450),
.Y(n_518)
);

OAI21xp5_ASAP7_75t_SL g517 ( 
.A1(n_512),
.A2(n_435),
.B(n_424),
.Y(n_517)
);

INVxp67_ASAP7_75t_L g519 ( 
.A(n_517),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_L g520 ( 
.A1(n_518),
.A2(n_516),
.B(n_515),
.Y(n_520)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_520),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_519),
.B(n_435),
.Y(n_521)
);

AOI21xp5_ASAP7_75t_L g523 ( 
.A1(n_522),
.A2(n_521),
.B(n_460),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_523),
.B(n_449),
.Y(n_524)
);

XOR2xp5_ASAP7_75t_L g525 ( 
.A(n_524),
.B(n_449),
.Y(n_525)
);


endmodule