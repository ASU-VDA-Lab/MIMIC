module fake_netlist_1_7633_n_33 (n_1, n_2, n_6, n_4, n_3, n_5, n_7, n_0, n_33);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_7;
input n_0;
output n_33;
wire n_20;
wire n_23;
wire n_28;
wire n_8;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_18;
wire n_32;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
NAND2xp33_ASAP7_75t_R g8 ( .A(n_7), .B(n_6), .Y(n_8) );
CKINVDCx5p33_ASAP7_75t_R g9 ( .A(n_0), .Y(n_9) );
CKINVDCx5p33_ASAP7_75t_R g10 ( .A(n_2), .Y(n_10) );
INVx1_ASAP7_75t_L g11 ( .A(n_0), .Y(n_11) );
CKINVDCx16_ASAP7_75t_R g12 ( .A(n_5), .Y(n_12) );
INVx3_ASAP7_75t_L g13 ( .A(n_4), .Y(n_13) );
NOR2xp33_ASAP7_75t_L g14 ( .A(n_13), .B(n_1), .Y(n_14) );
NAND2xp5_ASAP7_75t_SL g15 ( .A(n_13), .B(n_12), .Y(n_15) );
BUFx3_ASAP7_75t_L g16 ( .A(n_13), .Y(n_16) );
NAND2xp5_ASAP7_75t_SL g17 ( .A(n_12), .B(n_1), .Y(n_17) );
BUFx2_ASAP7_75t_L g18 ( .A(n_9), .Y(n_18) );
INVxp67_ASAP7_75t_L g19 ( .A(n_18), .Y(n_19) );
HB1xp67_ASAP7_75t_L g20 ( .A(n_16), .Y(n_20) );
INVx2_ASAP7_75t_L g21 ( .A(n_14), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_14), .Y(n_22) );
NAND2xp5_ASAP7_75t_L g23 ( .A(n_20), .B(n_15), .Y(n_23) );
OR2x2_ASAP7_75t_L g24 ( .A(n_19), .B(n_17), .Y(n_24) );
HB1xp67_ASAP7_75t_L g25 ( .A(n_19), .Y(n_25) );
NAND3xp33_ASAP7_75t_L g26 ( .A(n_25), .B(n_22), .C(n_21), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_23), .Y(n_27) );
INVx1_ASAP7_75t_L g28 ( .A(n_27), .Y(n_28) );
INVx1_ASAP7_75t_L g29 ( .A(n_26), .Y(n_29) );
HB1xp67_ASAP7_75t_L g30 ( .A(n_28), .Y(n_30) );
NOR3xp33_ASAP7_75t_L g31 ( .A(n_29), .B(n_24), .C(n_11), .Y(n_31) );
NAND2xp5_ASAP7_75t_SL g32 ( .A(n_30), .B(n_31), .Y(n_32) );
AOI22xp5_ASAP7_75t_L g33 ( .A1(n_32), .A2(n_8), .B1(n_10), .B2(n_3), .Y(n_33) );
endmodule