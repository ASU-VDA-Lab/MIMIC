module fake_jpeg_16602_n_149 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_149);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_149;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx3_ASAP7_75t_SL g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_17),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_38),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_39),
.B(n_40),
.Y(n_42)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_21),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_47),
.B(n_49),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_30),
.B(n_28),
.Y(n_48)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_16),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_32),
.B(n_28),
.Y(n_52)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_25),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_54),
.B(n_57),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_14),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_56),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_31),
.B(n_14),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_34),
.B(n_29),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_58),
.Y(n_81)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

A2O1A1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_55),
.A2(n_15),
.B(n_26),
.C(n_16),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_61),
.B(n_75),
.Y(n_79)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_62),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_47),
.A2(n_40),
.B1(n_19),
.B2(n_23),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_64),
.A2(n_71),
.B1(n_73),
.B2(n_75),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_23),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_24),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_50),
.A2(n_15),
.B1(n_26),
.B2(n_25),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_67),
.A2(n_72),
.B1(n_43),
.B2(n_24),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_44),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_68),
.B(n_70),
.Y(n_86)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_74),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_41),
.B(n_18),
.Y(n_70)
);

AND2x6_ASAP7_75t_L g71 ( 
.A(n_49),
.B(n_0),
.Y(n_71)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_49),
.A2(n_38),
.B1(n_35),
.B2(n_17),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_42),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_50),
.A2(n_29),
.B1(n_20),
.B2(n_18),
.Y(n_75)
);

AND2x6_ASAP7_75t_L g78 ( 
.A(n_51),
.B(n_0),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_78),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_79),
.A2(n_94),
.B1(n_80),
.B2(n_86),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_63),
.B(n_20),
.Y(n_80)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_83),
.B(n_61),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_46),
.Y(n_84)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_89),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_65),
.B(n_46),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_87),
.A2(n_77),
.B1(n_64),
.B2(n_68),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_59),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_58),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_46),
.Y(n_95)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_95),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_90),
.A2(n_71),
.B1(n_73),
.B2(n_77),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_97),
.B(n_107),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_SL g114 ( 
.A(n_98),
.B(n_101),
.Y(n_114)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_93),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_100),
.B(n_105),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_95),
.B(n_66),
.C(n_34),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_86),
.Y(n_112)
);

OA21x2_ASAP7_75t_L g105 ( 
.A1(n_79),
.A2(n_84),
.B(n_91),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_87),
.A2(n_90),
.B1(n_91),
.B2(n_83),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_106),
.A2(n_109),
.B(n_98),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_108),
.A2(n_10),
.B(n_11),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_87),
.A2(n_78),
.B1(n_69),
.B2(n_44),
.Y(n_109)
);

INVxp67_ASAP7_75t_SL g110 ( 
.A(n_100),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_110),
.B(n_72),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_111),
.A2(n_113),
.B(n_118),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_112),
.B(n_106),
.C(n_99),
.Y(n_125)
);

A2O1A1O1Ixp25_ASAP7_75t_L g113 ( 
.A1(n_105),
.A2(n_88),
.B(n_92),
.C(n_82),
.D(n_81),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_81),
.Y(n_116)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_116),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_103),
.B(n_104),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_119),
.B(n_97),
.Y(n_128)
);

A2O1A1O1Ixp25_ASAP7_75t_L g120 ( 
.A1(n_105),
.A2(n_82),
.B(n_93),
.C(n_60),
.D(n_34),
.Y(n_120)
);

NOR3xp33_ASAP7_75t_SL g124 ( 
.A(n_120),
.B(n_109),
.C(n_101),
.Y(n_124)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_122),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_124),
.A2(n_114),
.B(n_96),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_125),
.B(n_126),
.C(n_114),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_115),
.B(n_99),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_113),
.Y(n_127)
);

OAI221xp5_ASAP7_75t_L g132 ( 
.A1(n_127),
.A2(n_128),
.B1(n_110),
.B2(n_22),
.C(n_9),
.Y(n_132)
);

OAI321xp33_ASAP7_75t_L g129 ( 
.A1(n_124),
.A2(n_117),
.A3(n_120),
.B1(n_121),
.B2(n_96),
.C(n_125),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_129),
.B(n_130),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_131),
.B(n_1),
.Y(n_138)
);

AOI31xp67_ASAP7_75t_L g136 ( 
.A1(n_132),
.A2(n_8),
.A3(n_2),
.B(n_3),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g133 ( 
.A(n_121),
.B(n_22),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_133),
.A2(n_1),
.B(n_2),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_136),
.B(n_138),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_134),
.A2(n_123),
.B1(n_53),
.B2(n_3),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_137),
.A2(n_4),
.B(n_5),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_139),
.B(n_133),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_135),
.B(n_4),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_141),
.B(n_143),
.Y(n_144)
);

AOI322xp5_ASAP7_75t_L g145 ( 
.A1(n_142),
.A2(n_5),
.A3(n_6),
.B1(n_7),
.B2(n_53),
.C1(n_137),
.C2(n_140),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_143),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_146),
.A2(n_147),
.B(n_5),
.Y(n_148)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_144),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_7),
.Y(n_149)
);


endmodule