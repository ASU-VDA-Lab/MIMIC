module fake_aes_2253_n_1572 (n_117, n_44, n_185, n_22, n_57, n_26, n_284, n_278, n_60, n_114, n_41, n_94, n_125, n_9, n_161, n_177, n_130, n_189, n_311, n_19, n_292, n_309, n_160, n_154, n_7, n_29, n_229, n_252, n_152, n_113, n_206, n_17, n_288, n_6, n_296, n_157, n_79, n_202, n_38, n_142, n_232, n_316, n_31, n_211, n_275, n_0, n_131, n_112, n_205, n_162, n_163, n_105, n_227, n_231, n_298, n_144, n_27, n_53, n_183, n_199, n_83, n_28, n_48, n_100, n_305, n_228, n_236, n_150, n_3, n_18, n_301, n_66, n_222, n_234, n_286, n_15, n_190, n_246, n_39, n_279, n_303, n_289, n_249, n_244, n_50, n_73, n_49, n_119, n_141, n_97, n_167, n_171, n_65, n_196, n_192, n_312, n_137, n_277, n_45, n_85, n_250, n_314, n_237, n_181, n_101, n_62, n_255, n_36, n_37, n_91, n_108, n_116, n_230, n_209, n_274, n_16, n_282, n_319, n_241, n_95, n_238, n_318, n_293, n_135, n_42, n_24, n_247, n_304, n_294, n_313, n_210, n_184, n_310, n_191, n_307, n_46, n_32, n_235, n_243, n_268, n_174, n_248, n_72, n_299, n_43, n_89, n_256, n_67, n_77, n_20, n_54, n_172, n_251, n_59, n_218, n_1, n_271, n_302, n_270, n_153, n_61, n_259, n_308, n_93, n_140, n_207, n_224, n_96, n_219, n_133, n_149, n_81, n_69, n_214, n_204, n_88, n_33, n_107, n_254, n_262, n_10, n_239, n_87, n_98, n_276, n_320, n_285, n_195, n_165, n_34, n_5, n_23, n_8, n_217, n_139, n_193, n_273, n_120, n_70, n_245, n_90, n_260, n_78, n_197, n_201, n_317, n_4, n_40, n_111, n_64, n_265, n_264, n_200, n_208, n_126, n_178, n_118, n_179, n_315, n_86, n_143, n_295, n_263, n_166, n_186, n_75, n_136, n_283, n_76, n_216, n_147, n_148, n_212, n_92, n_11, n_168, n_134, n_233, n_82, n_106, n_173, n_51, n_225, n_220, n_267, n_221, n_203, n_52, n_102, n_115, n_80, n_300, n_158, n_121, n_35, n_240, n_103, n_180, n_104, n_74, n_272, n_146, n_306, n_47, n_215, n_242, n_155, n_13, n_198, n_169, n_156, n_124, n_297, n_128, n_129, n_63, n_14, n_71, n_56, n_188, n_127, n_291, n_170, n_281, n_58, n_122, n_187, n_138, n_258, n_253, n_84, n_266, n_55, n_12, n_213, n_182, n_226, n_159, n_176, n_68, n_2, n_123, n_223, n_25, n_30, n_194, n_287, n_110, n_261, n_164, n_175, n_145, n_290, n_280, n_21, n_99, n_109, n_132, n_151, n_257, n_269, n_1572);
input n_117;
input n_44;
input n_185;
input n_22;
input n_57;
input n_26;
input n_284;
input n_278;
input n_60;
input n_114;
input n_41;
input n_94;
input n_125;
input n_9;
input n_161;
input n_177;
input n_130;
input n_189;
input n_311;
input n_19;
input n_292;
input n_309;
input n_160;
input n_154;
input n_7;
input n_29;
input n_229;
input n_252;
input n_152;
input n_113;
input n_206;
input n_17;
input n_288;
input n_6;
input n_296;
input n_157;
input n_79;
input n_202;
input n_38;
input n_142;
input n_232;
input n_316;
input n_31;
input n_211;
input n_275;
input n_0;
input n_131;
input n_112;
input n_205;
input n_162;
input n_163;
input n_105;
input n_227;
input n_231;
input n_298;
input n_144;
input n_27;
input n_53;
input n_183;
input n_199;
input n_83;
input n_28;
input n_48;
input n_100;
input n_305;
input n_228;
input n_236;
input n_150;
input n_3;
input n_18;
input n_301;
input n_66;
input n_222;
input n_234;
input n_286;
input n_15;
input n_190;
input n_246;
input n_39;
input n_279;
input n_303;
input n_289;
input n_249;
input n_244;
input n_50;
input n_73;
input n_49;
input n_119;
input n_141;
input n_97;
input n_167;
input n_171;
input n_65;
input n_196;
input n_192;
input n_312;
input n_137;
input n_277;
input n_45;
input n_85;
input n_250;
input n_314;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_37;
input n_91;
input n_108;
input n_116;
input n_230;
input n_209;
input n_274;
input n_16;
input n_282;
input n_319;
input n_241;
input n_95;
input n_238;
input n_318;
input n_293;
input n_135;
input n_42;
input n_24;
input n_247;
input n_304;
input n_294;
input n_313;
input n_210;
input n_184;
input n_310;
input n_191;
input n_307;
input n_46;
input n_32;
input n_235;
input n_243;
input n_268;
input n_174;
input n_248;
input n_72;
input n_299;
input n_43;
input n_89;
input n_256;
input n_67;
input n_77;
input n_20;
input n_54;
input n_172;
input n_251;
input n_59;
input n_218;
input n_1;
input n_271;
input n_302;
input n_270;
input n_153;
input n_61;
input n_259;
input n_308;
input n_93;
input n_140;
input n_207;
input n_224;
input n_96;
input n_219;
input n_133;
input n_149;
input n_81;
input n_69;
input n_214;
input n_204;
input n_88;
input n_33;
input n_107;
input n_254;
input n_262;
input n_10;
input n_239;
input n_87;
input n_98;
input n_276;
input n_320;
input n_285;
input n_195;
input n_165;
input n_34;
input n_5;
input n_23;
input n_8;
input n_217;
input n_139;
input n_193;
input n_273;
input n_120;
input n_70;
input n_245;
input n_90;
input n_260;
input n_78;
input n_197;
input n_201;
input n_317;
input n_4;
input n_40;
input n_111;
input n_64;
input n_265;
input n_264;
input n_200;
input n_208;
input n_126;
input n_178;
input n_118;
input n_179;
input n_315;
input n_86;
input n_143;
input n_295;
input n_263;
input n_166;
input n_186;
input n_75;
input n_136;
input n_283;
input n_76;
input n_216;
input n_147;
input n_148;
input n_212;
input n_92;
input n_11;
input n_168;
input n_134;
input n_233;
input n_82;
input n_106;
input n_173;
input n_51;
input n_225;
input n_220;
input n_267;
input n_221;
input n_203;
input n_52;
input n_102;
input n_115;
input n_80;
input n_300;
input n_158;
input n_121;
input n_35;
input n_240;
input n_103;
input n_180;
input n_104;
input n_74;
input n_272;
input n_146;
input n_306;
input n_47;
input n_215;
input n_242;
input n_155;
input n_13;
input n_198;
input n_169;
input n_156;
input n_124;
input n_297;
input n_128;
input n_129;
input n_63;
input n_14;
input n_71;
input n_56;
input n_188;
input n_127;
input n_291;
input n_170;
input n_281;
input n_58;
input n_122;
input n_187;
input n_138;
input n_258;
input n_253;
input n_84;
input n_266;
input n_55;
input n_12;
input n_213;
input n_182;
input n_226;
input n_159;
input n_176;
input n_68;
input n_2;
input n_123;
input n_223;
input n_25;
input n_30;
input n_194;
input n_287;
input n_110;
input n_261;
input n_164;
input n_175;
input n_145;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_132;
input n_151;
input n_257;
input n_269;
output n_1572;
wire n_1309;
wire n_1497;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_646;
wire n_1334;
wire n_829;
wire n_1198;
wire n_1571;
wire n_1382;
wire n_667;
wire n_988;
wire n_1477;
wire n_1363;
wire n_655;
wire n_1298;
wire n_1391;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1527;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_1445;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_1528;
wire n_789;
wire n_1197;
wire n_1163;
wire n_1404;
wire n_387;
wire n_452;
wire n_518;
wire n_1336;
wire n_411;
wire n_1341;
wire n_1381;
wire n_860;
wire n_1208;
wire n_1201;
wire n_1342;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1352;
wire n_1503;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_1355;
wire n_915;
wire n_1536;
wire n_367;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1407;
wire n_1475;
wire n_1505;
wire n_1018;
wire n_979;
wire n_499;
wire n_1349;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_1561;
wire n_1337;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1525;
wire n_1448;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1414;
wire n_1500;
wire n_1209;
wire n_1399;
wire n_1441;
wire n_926;
wire n_1274;
wire n_1569;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1406;
wire n_1099;
wire n_1328;
wire n_1369;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1443;
wire n_1313;
wire n_954;
wire n_574;
wire n_822;
wire n_706;
wire n_823;
wire n_1181;
wire n_1438;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1547;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1377;
wire n_1079;
wire n_409;
wire n_1321;
wire n_677;
wire n_1354;
wire n_1242;
wire n_756;
wire n_1385;
wire n_1240;
wire n_1139;
wire n_577;
wire n_1394;
wire n_870;
wire n_1324;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_1551;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_1388;
wire n_327;
wire n_1102;
wire n_723;
wire n_972;
wire n_1522;
wire n_1499;
wire n_1437;
wire n_997;
wire n_1387;
wire n_1244;
wire n_1464;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_1452;
wire n_359;
wire n_1402;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1447;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_1510;
wire n_1467;
wire n_994;
wire n_930;
wire n_1413;
wire n_410;
wire n_774;
wire n_1207;
wire n_1463;
wire n_377;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1365;
wire n_1164;
wire n_1533;
wire n_451;
wire n_487;
wire n_748;
wire n_1373;
wire n_1563;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1461;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_1542;
wire n_1311;
wire n_1558;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_1412;
wire n_1502;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_1306;
wire n_958;
wire n_468;
wire n_1453;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_1333;
wire n_1361;
wire n_1557;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_1345;
wire n_661;
wire n_890;
wire n_787;
wire n_1488;
wire n_1015;
wire n_548;
wire n_1048;
wire n_1564;
wire n_1521;
wire n_973;
wire n_587;
wire n_1468;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_1435;
wire n_1539;
wire n_796;
wire n_1216;
wire n_927;
wire n_1405;
wire n_1433;
wire n_840;
wire n_846;
wire n_968;
wire n_1543;
wire n_512;
wire n_1330;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_1515;
wire n_897;
wire n_1188;
wire n_1496;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_1415;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_1062;
wire n_708;
wire n_1271;
wire n_634;
wire n_1537;
wire n_1520;
wire n_696;
wire n_1203;
wire n_1546;
wire n_1524;
wire n_1013;
wire n_1000;
wire n_1370;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_1465;
wire n_329;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_1540;
wire n_952;
wire n_685;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_1472;
wire n_943;
wire n_1326;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1346;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1427;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1153;
wire n_816;
wire n_522;
wire n_898;
wire n_1562;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_1514;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_1060;
wire n_721;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_1440;
wire n_1541;
wire n_1397;
wire n_1356;
wire n_836;
wire n_561;
wire n_1096;
wire n_1553;
wire n_594;
wire n_531;
wire n_1136;
wire n_1007;
wire n_1117;
wire n_1408;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1339;
wire n_1432;
wire n_1315;
wire n_1490;
wire n_867;
wire n_1070;
wire n_1529;
wire n_1270;
wire n_1474;
wire n_1512;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1507;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_323;
wire n_347;
wire n_515;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1449;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_1495;
wire n_606;
wire n_332;
wire n_1292;
wire n_1425;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1416;
wire n_1566;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_1559;
wire n_1483;
wire n_496;
wire n_1362;
wire n_801;
wire n_1059;
wire n_701;
wire n_1530;
wire n_612;
wire n_1513;
wire n_1418;
wire n_1032;
wire n_1284;
wire n_1358;
wire n_336;
wire n_464;
wire n_1243;
wire n_1196;
wire n_1338;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_1554;
wire n_400;
wire n_1455;
wire n_386;
wire n_432;
wire n_659;
wire n_1329;
wire n_1509;
wire n_1185;
wire n_1511;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_330;
wire n_1087;
wire n_662;
wire n_1372;
wire n_1460;
wire n_1451;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_1459;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_1319;
wire n_596;
wire n_1215;
wire n_951;
wire n_321;
wire n_1024;
wire n_1016;
wire n_652;
wire n_333;
wire n_1417;
wire n_1357;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1380;
wire n_1254;
wire n_764;
wire n_426;
wire n_1508;
wire n_1375;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_1458;
wire n_381;
wire n_1255;
wire n_322;
wire n_1299;
wire n_1450;
wire n_1332;
wire n_1480;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_1429;
wire n_805;
wire n_729;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_1470;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_1526;
wire n_788;
wire n_1454;
wire n_1471;
wire n_1383;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_420;
wire n_1089;
wire n_1434;
wire n_1058;
wire n_388;
wire n_1396;
wire n_1400;
wire n_1517;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_1473;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1351;
wire n_1318;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1478;
wire n_1068;
wire n_1565;
wire n_1149;
wire n_1430;
wire n_615;
wire n_1386;
wire n_1552;
wire n_1170;
wire n_1523;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_1492;
wire n_440;
wire n_1550;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_1395;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_1340;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1325;
wire n_1043;
wire n_1283;
wire n_346;
wire n_1489;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1516;
wire n_1027;
wire n_1040;
wire n_1367;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1538;
wire n_1073;
wire n_868;
wire n_1466;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_1393;
wire n_538;
wire n_492;
wire n_1426;
wire n_1555;
wire n_1150;
wire n_1462;
wire n_1327;
wire n_368;
wire n_1444;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1436;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_1378;
wire n_1570;
wire n_385;
wire n_1127;
wire n_1348;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_1409;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_1158;
wire n_1493;
wire n_1544;
wire n_328;
wire n_743;
wire n_757;
wire n_1568;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1498;
wire n_1224;
wire n_383;
wire n_762;
wire n_1422;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_1376;
wire n_765;
wire n_1177;
wire n_1545;
wire n_1310;
wire n_462;
wire n_1347;
wire n_1384;
wire n_783;
wire n_1074;
wire n_1374;
wire n_463;
wire n_1379;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_1534;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_1501;
wire n_777;
wire n_1504;
wire n_351;
wire n_401;
wire n_345;
wire n_360;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1479;
wire n_1360;
wire n_1486;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_326;
wire n_1081;
wire n_1457;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_1518;
wire n_945;
wire n_554;
wire n_726;
wire n_1519;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_1389;
wire n_630;
wire n_1180;
wire n_647;
wire n_1364;
wire n_1350;
wire n_844;
wire n_1403;
wire n_1160;
wire n_1420;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_895;
wire n_1481;
wire n_798;
wire n_887;
wire n_471;
wire n_1476;
wire n_1014;
wire n_1410;
wire n_1442;
wire n_665;
wire n_1154;
wire n_1560;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_1491;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_935;
wire n_910;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1485;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_1532;
wire n_889;
wire n_689;
wire n_902;
wire n_1423;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_1368;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1482;
wire n_1343;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_1494;
wire n_622;
wire n_601;
wire n_1331;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_1506;
wire n_1469;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_1535;
wire n_1439;
wire n_374;
wire n_718;
wire n_1484;
wire n_1567;
wire n_1238;
wire n_1411;
wire n_1114;
wire n_1304;
wire n_948;
wire n_1286;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1359;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_398;
wire n_445;
wire n_656;
wire n_1230;
wire n_553;
wire n_1431;
wire n_325;
wire n_349;
wire n_1021;
wire n_1456;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1353;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_1424;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1239;
wire n_1335;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_1344;
wire n_335;
wire n_700;
wire n_534;
wire n_1401;
wire n_1296;
wire n_1428;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_1549;
wire n_1053;
wire n_1223;
wire n_1421;
wire n_1390;
wire n_967;
wire n_1419;
wire n_1258;
wire n_1487;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_1531;
wire n_371;
wire n_1548;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_1371;
wire n_929;
wire n_1111;
wire n_976;
wire n_1446;
wire n_695;
wire n_1104;
wire n_1392;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_1366;
wire n_480;
wire n_453;
wire n_833;
wire n_1556;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_1398;
wire n_491;
wire n_1291;
INVx1_ASAP7_75t_L g321 ( .A(n_30), .Y(n_321) );
CKINVDCx5p33_ASAP7_75t_R g322 ( .A(n_273), .Y(n_322) );
CKINVDCx16_ASAP7_75t_R g323 ( .A(n_315), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_91), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_30), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_0), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_150), .Y(n_327) );
CKINVDCx16_ASAP7_75t_R g328 ( .A(n_0), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_124), .Y(n_329) );
CKINVDCx5p33_ASAP7_75t_R g330 ( .A(n_157), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_231), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_226), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_134), .Y(n_333) );
CKINVDCx5p33_ASAP7_75t_R g334 ( .A(n_71), .Y(n_334) );
CKINVDCx20_ASAP7_75t_R g335 ( .A(n_286), .Y(n_335) );
BUFx2_ASAP7_75t_L g336 ( .A(n_242), .Y(n_336) );
CKINVDCx5p33_ASAP7_75t_R g337 ( .A(n_317), .Y(n_337) );
CKINVDCx5p33_ASAP7_75t_R g338 ( .A(n_101), .Y(n_338) );
NOR2xp67_ASAP7_75t_L g339 ( .A(n_292), .B(n_303), .Y(n_339) );
BUFx3_ASAP7_75t_L g340 ( .A(n_196), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_237), .Y(n_341) );
CKINVDCx20_ASAP7_75t_R g342 ( .A(n_227), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_122), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_176), .Y(n_344) );
CKINVDCx5p33_ASAP7_75t_R g345 ( .A(n_264), .Y(n_345) );
INVxp67_ASAP7_75t_SL g346 ( .A(n_295), .Y(n_346) );
CKINVDCx5p33_ASAP7_75t_R g347 ( .A(n_266), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_130), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_249), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_210), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_288), .Y(n_351) );
CKINVDCx16_ASAP7_75t_R g352 ( .A(n_174), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_205), .Y(n_353) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_140), .Y(n_354) );
CKINVDCx20_ASAP7_75t_R g355 ( .A(n_189), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_99), .Y(n_356) );
CKINVDCx16_ASAP7_75t_R g357 ( .A(n_47), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_225), .Y(n_358) );
CKINVDCx16_ASAP7_75t_R g359 ( .A(n_39), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_256), .Y(n_360) );
CKINVDCx5p33_ASAP7_75t_R g361 ( .A(n_138), .Y(n_361) );
CKINVDCx20_ASAP7_75t_R g362 ( .A(n_27), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_98), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_143), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_298), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_240), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_147), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_52), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_170), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_181), .Y(n_370) );
INVxp67_ASAP7_75t_SL g371 ( .A(n_310), .Y(n_371) );
INVxp67_ASAP7_75t_SL g372 ( .A(n_123), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_86), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_97), .Y(n_374) );
CKINVDCx5p33_ASAP7_75t_R g375 ( .A(n_262), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_164), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_207), .Y(n_377) );
BUFx6f_ASAP7_75t_L g378 ( .A(n_57), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_224), .Y(n_379) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_291), .Y(n_380) );
CKINVDCx14_ASAP7_75t_R g381 ( .A(n_239), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_47), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_203), .Y(n_383) );
INVxp67_ASAP7_75t_SL g384 ( .A(n_14), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_129), .Y(n_385) );
CKINVDCx5p33_ASAP7_75t_R g386 ( .A(n_8), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_36), .Y(n_387) );
INVxp67_ASAP7_75t_L g388 ( .A(n_32), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_105), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_20), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_13), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_282), .Y(n_392) );
CKINVDCx5p33_ASAP7_75t_R g393 ( .A(n_192), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_222), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_162), .Y(n_395) );
INVx2_ASAP7_75t_SL g396 ( .A(n_259), .Y(n_396) );
INVxp33_ASAP7_75t_L g397 ( .A(n_121), .Y(n_397) );
BUFx3_ASAP7_75t_L g398 ( .A(n_109), .Y(n_398) );
CKINVDCx16_ASAP7_75t_R g399 ( .A(n_248), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_250), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_61), .Y(n_401) );
BUFx3_ASAP7_75t_L g402 ( .A(n_220), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_145), .Y(n_403) );
CKINVDCx20_ASAP7_75t_R g404 ( .A(n_19), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_101), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_33), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_20), .Y(n_407) );
INVxp33_ASAP7_75t_SL g408 ( .A(n_319), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_75), .Y(n_409) );
CKINVDCx20_ASAP7_75t_R g410 ( .A(n_7), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_93), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_309), .Y(n_412) );
CKINVDCx20_ASAP7_75t_R g413 ( .A(n_301), .Y(n_413) );
BUFx6f_ASAP7_75t_L g414 ( .A(n_221), .Y(n_414) );
INVxp67_ASAP7_75t_SL g415 ( .A(n_34), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_253), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_275), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_57), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_269), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_230), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_17), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_184), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_116), .Y(n_423) );
BUFx3_ASAP7_75t_L g424 ( .A(n_190), .Y(n_424) );
INVxp33_ASAP7_75t_SL g425 ( .A(n_168), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_154), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_38), .Y(n_427) );
NOR2xp67_ASAP7_75t_L g428 ( .A(n_149), .B(n_63), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_22), .Y(n_429) );
BUFx6f_ASAP7_75t_L g430 ( .A(n_215), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_320), .Y(n_431) );
HB1xp67_ASAP7_75t_L g432 ( .A(n_179), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_12), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_6), .Y(n_434) );
INVxp33_ASAP7_75t_SL g435 ( .A(n_24), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_204), .Y(n_436) );
INVx1_ASAP7_75t_SL g437 ( .A(n_297), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_62), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_17), .Y(n_439) );
CKINVDCx20_ASAP7_75t_R g440 ( .A(n_188), .Y(n_440) );
CKINVDCx5p33_ASAP7_75t_R g441 ( .A(n_28), .Y(n_441) );
CKINVDCx5p33_ASAP7_75t_R g442 ( .A(n_167), .Y(n_442) );
CKINVDCx14_ASAP7_75t_R g443 ( .A(n_61), .Y(n_443) );
CKINVDCx16_ASAP7_75t_R g444 ( .A(n_132), .Y(n_444) );
CKINVDCx5p33_ASAP7_75t_R g445 ( .A(n_314), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_48), .Y(n_446) );
BUFx3_ASAP7_75t_L g447 ( .A(n_213), .Y(n_447) );
CKINVDCx5p33_ASAP7_75t_R g448 ( .A(n_308), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_232), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_283), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_263), .Y(n_451) );
CKINVDCx5p33_ASAP7_75t_R g452 ( .A(n_276), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_307), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_209), .Y(n_454) );
BUFx2_ASAP7_75t_L g455 ( .A(n_281), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_7), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_50), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_180), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_77), .Y(n_459) );
CKINVDCx5p33_ASAP7_75t_R g460 ( .A(n_208), .Y(n_460) );
INVxp67_ASAP7_75t_L g461 ( .A(n_41), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_78), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_69), .Y(n_463) );
CKINVDCx5p33_ASAP7_75t_R g464 ( .A(n_217), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_115), .Y(n_465) );
INVx1_ASAP7_75t_SL g466 ( .A(n_223), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_153), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_219), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_142), .Y(n_469) );
INVx1_ASAP7_75t_SL g470 ( .A(n_98), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_268), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_218), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_304), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_169), .B(n_247), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_278), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_177), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_117), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_23), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_272), .Y(n_479) );
CKINVDCx5p33_ASAP7_75t_R g480 ( .A(n_93), .Y(n_480) );
INVx2_ASAP7_75t_SL g481 ( .A(n_299), .Y(n_481) );
BUFx2_ASAP7_75t_L g482 ( .A(n_78), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_214), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_110), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_148), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_48), .Y(n_486) );
BUFx3_ASAP7_75t_L g487 ( .A(n_313), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_271), .Y(n_488) );
CKINVDCx20_ASAP7_75t_R g489 ( .A(n_71), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_10), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_171), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_119), .Y(n_492) );
BUFx6f_ASAP7_75t_L g493 ( .A(n_414), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_364), .Y(n_494) );
BUFx6f_ASAP7_75t_L g495 ( .A(n_414), .Y(n_495) );
INVx3_ASAP7_75t_L g496 ( .A(n_378), .Y(n_496) );
INVx2_ASAP7_75t_L g497 ( .A(n_414), .Y(n_497) );
HB1xp67_ASAP7_75t_L g498 ( .A(n_443), .Y(n_498) );
BUFx3_ASAP7_75t_L g499 ( .A(n_336), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_414), .Y(n_500) );
INVx3_ASAP7_75t_L g501 ( .A(n_378), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_364), .Y(n_502) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_336), .B(n_1), .Y(n_503) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_455), .B(n_1), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_365), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_455), .B(n_2), .Y(n_506) );
CKINVDCx5p33_ASAP7_75t_R g507 ( .A(n_443), .Y(n_507) );
AND3x1_ASAP7_75t_L g508 ( .A(n_373), .B(n_2), .C(n_3), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_365), .Y(n_509) );
AND2x4_ASAP7_75t_L g510 ( .A(n_396), .B(n_3), .Y(n_510) );
OA21x2_ASAP7_75t_L g511 ( .A1(n_366), .A2(n_4), .B(n_5), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_482), .B(n_4), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_366), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_414), .Y(n_514) );
CKINVDCx5p33_ASAP7_75t_R g515 ( .A(n_323), .Y(n_515) );
CKINVDCx5p33_ASAP7_75t_R g516 ( .A(n_352), .Y(n_516) );
INVx2_ASAP7_75t_L g517 ( .A(n_430), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_482), .B(n_5), .Y(n_518) );
CKINVDCx20_ASAP7_75t_R g519 ( .A(n_328), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_397), .B(n_6), .Y(n_520) );
BUFx6f_ASAP7_75t_L g521 ( .A(n_430), .Y(n_521) );
CKINVDCx5p33_ASAP7_75t_R g522 ( .A(n_399), .Y(n_522) );
INVx1_ASAP7_75t_SL g523 ( .A(n_335), .Y(n_523) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_397), .B(n_8), .Y(n_524) );
BUFx3_ASAP7_75t_L g525 ( .A(n_340), .Y(n_525) );
AND2x4_ASAP7_75t_L g526 ( .A(n_396), .B(n_481), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_367), .Y(n_527) );
INVx6_ASAP7_75t_L g528 ( .A(n_340), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_430), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_381), .B(n_9), .Y(n_530) );
INVx2_ASAP7_75t_L g531 ( .A(n_430), .Y(n_531) );
AOI22xp5_ASAP7_75t_L g532 ( .A1(n_435), .A2(n_11), .B1(n_9), .B2(n_10), .Y(n_532) );
INVx2_ASAP7_75t_L g533 ( .A(n_493), .Y(n_533) );
OAI22xp33_ASAP7_75t_SL g534 ( .A1(n_532), .A2(n_359), .B1(n_357), .B2(n_435), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_511), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_511), .Y(n_536) );
INVx3_ASAP7_75t_L g537 ( .A(n_510), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_511), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_511), .Y(n_539) );
INVx1_ASAP7_75t_SL g540 ( .A(n_498), .Y(n_540) );
INVx2_ASAP7_75t_L g541 ( .A(n_493), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_499), .B(n_498), .Y(n_542) );
AND2x6_ASAP7_75t_L g543 ( .A(n_510), .B(n_474), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_499), .B(n_444), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_493), .Y(n_545) );
INVx5_ASAP7_75t_L g546 ( .A(n_528), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_511), .Y(n_547) );
INVx5_ASAP7_75t_R g548 ( .A(n_515), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_499), .B(n_354), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_511), .Y(n_550) );
INVx2_ASAP7_75t_L g551 ( .A(n_493), .Y(n_551) );
NOR2xp33_ASAP7_75t_L g552 ( .A(n_499), .B(n_380), .Y(n_552) );
INVx2_ASAP7_75t_L g553 ( .A(n_493), .Y(n_553) );
BUFx3_ASAP7_75t_L g554 ( .A(n_510), .Y(n_554) );
AO22x2_ASAP7_75t_L g555 ( .A1(n_510), .A2(n_367), .B1(n_415), .B2(n_384), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_526), .B(n_432), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_512), .B(n_381), .Y(n_557) );
INVx2_ASAP7_75t_SL g558 ( .A(n_530), .Y(n_558) );
NOR2xp33_ASAP7_75t_L g559 ( .A(n_526), .B(n_481), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_496), .Y(n_560) );
NOR2xp33_ASAP7_75t_L g561 ( .A(n_526), .B(n_408), .Y(n_561) );
NOR2xp33_ASAP7_75t_L g562 ( .A(n_526), .B(n_408), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_496), .Y(n_563) );
NAND2xp5_ASAP7_75t_SL g564 ( .A(n_507), .B(n_322), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_526), .B(n_334), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_496), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_496), .Y(n_567) );
CKINVDCx20_ASAP7_75t_R g568 ( .A(n_519), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_496), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_501), .Y(n_570) );
INVxp33_ASAP7_75t_SL g571 ( .A(n_515), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_512), .A2(n_324), .B1(n_325), .B2(n_321), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_501), .Y(n_573) );
AND2x6_ASAP7_75t_L g574 ( .A(n_510), .B(n_474), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_512), .B(n_373), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_501), .Y(n_576) );
AND2x6_ASAP7_75t_L g577 ( .A(n_510), .B(n_398), .Y(n_577) );
INVx4_ASAP7_75t_L g578 ( .A(n_528), .Y(n_578) );
BUFx6f_ASAP7_75t_L g579 ( .A(n_493), .Y(n_579) );
INVx2_ASAP7_75t_L g580 ( .A(n_493), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_520), .B(n_387), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_501), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_542), .Y(n_583) );
INVx4_ASAP7_75t_L g584 ( .A(n_543), .Y(n_584) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_543), .A2(n_502), .B1(n_505), .B2(n_494), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_542), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_540), .B(n_516), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_557), .B(n_520), .Y(n_588) );
OAI22xp5_ASAP7_75t_L g589 ( .A1(n_555), .A2(n_523), .B1(n_335), .B2(n_355), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_557), .B(n_520), .Y(n_590) );
INVx5_ASAP7_75t_L g591 ( .A(n_577), .Y(n_591) );
OAI22xp33_ASAP7_75t_L g592 ( .A1(n_558), .A2(n_532), .B1(n_518), .B2(n_506), .Y(n_592) );
OAI22xp5_ASAP7_75t_SL g593 ( .A1(n_568), .A2(n_404), .B1(n_410), .B2(n_362), .Y(n_593) );
BUFx5_ASAP7_75t_L g594 ( .A(n_577), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_558), .Y(n_595) );
INVxp67_ASAP7_75t_L g596 ( .A(n_544), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_555), .Y(n_597) );
NAND2xp5_ASAP7_75t_SL g598 ( .A(n_561), .B(n_530), .Y(n_598) );
NAND2xp5_ASAP7_75t_SL g599 ( .A(n_562), .B(n_565), .Y(n_599) );
NAND2xp5_ASAP7_75t_SL g600 ( .A(n_549), .B(n_530), .Y(n_600) );
BUFx12f_ASAP7_75t_L g601 ( .A(n_548), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_555), .A2(n_504), .B1(n_503), .B2(n_494), .Y(n_602) );
INVx2_ASAP7_75t_SL g603 ( .A(n_581), .Y(n_603) );
NAND2xp5_ASAP7_75t_SL g604 ( .A(n_556), .B(n_507), .Y(n_604) );
O2A1O1Ixp33_ASAP7_75t_L g605 ( .A1(n_534), .A2(n_518), .B(n_505), .C(n_509), .Y(n_605) );
AOI22xp5_ASAP7_75t_L g606 ( .A1(n_555), .A2(n_504), .B1(n_503), .B2(n_524), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_581), .Y(n_607) );
AO22x1_ASAP7_75t_L g608 ( .A1(n_571), .A2(n_523), .B1(n_516), .B2(n_522), .Y(n_608) );
INVx3_ASAP7_75t_L g609 ( .A(n_554), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_575), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_552), .B(n_575), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g612 ( .A1(n_543), .A2(n_509), .B1(n_513), .B2(n_502), .Y(n_612) );
INVx5_ASAP7_75t_L g613 ( .A(n_577), .Y(n_613) );
AO22x1_ASAP7_75t_L g614 ( .A1(n_548), .A2(n_522), .B1(n_425), .B2(n_506), .Y(n_614) );
BUFx6f_ASAP7_75t_L g615 ( .A(n_554), .Y(n_615) );
INVxp67_ASAP7_75t_L g616 ( .A(n_543), .Y(n_616) );
HB1xp67_ASAP7_75t_L g617 ( .A(n_554), .Y(n_617) );
BUFx3_ASAP7_75t_L g618 ( .A(n_577), .Y(n_618) );
AND2x4_ASAP7_75t_L g619 ( .A(n_564), .B(n_508), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g620 ( .A1(n_543), .A2(n_527), .B1(n_513), .B2(n_525), .Y(n_620) );
CKINVDCx5p33_ASAP7_75t_R g621 ( .A(n_572), .Y(n_621) );
NOR2xp33_ASAP7_75t_L g622 ( .A(n_559), .B(n_537), .Y(n_622) );
OAI22xp5_ASAP7_75t_L g623 ( .A1(n_537), .A2(n_355), .B1(n_413), .B2(n_342), .Y(n_623) );
INVx2_ASAP7_75t_L g624 ( .A(n_537), .Y(n_624) );
INVxp33_ASAP7_75t_L g625 ( .A(n_535), .Y(n_625) );
NAND2xp5_ASAP7_75t_SL g626 ( .A(n_535), .B(n_322), .Y(n_626) );
AND2x4_ASAP7_75t_L g627 ( .A(n_543), .B(n_508), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_543), .Y(n_628) );
BUFx6f_ASAP7_75t_SL g629 ( .A(n_577), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_574), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_574), .B(n_527), .Y(n_631) );
NAND2xp5_ASAP7_75t_SL g632 ( .A(n_536), .B(n_330), .Y(n_632) );
AOI22xp5_ASAP7_75t_L g633 ( .A1(n_574), .A2(n_413), .B1(n_440), .B2(n_342), .Y(n_633) );
INVx4_ASAP7_75t_L g634 ( .A(n_574), .Y(n_634) );
AOI22xp33_ASAP7_75t_L g635 ( .A1(n_574), .A2(n_525), .B1(n_356), .B2(n_363), .Y(n_635) );
AOI22xp33_ASAP7_75t_L g636 ( .A1(n_574), .A2(n_525), .B1(n_368), .B2(n_374), .Y(n_636) );
BUFx2_ASAP7_75t_L g637 ( .A(n_574), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_577), .Y(n_638) );
INVx3_ASAP7_75t_L g639 ( .A(n_577), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_578), .B(n_525), .Y(n_640) );
INVx2_ASAP7_75t_L g641 ( .A(n_578), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_578), .B(n_330), .Y(n_642) );
AOI22xp33_ASAP7_75t_L g643 ( .A1(n_536), .A2(n_425), .B1(n_528), .B2(n_382), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_538), .Y(n_644) );
CKINVDCx5p33_ASAP7_75t_R g645 ( .A(n_538), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_578), .B(n_337), .Y(n_646) );
INVx2_ASAP7_75t_L g647 ( .A(n_560), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_539), .B(n_337), .Y(n_648) );
INVxp67_ASAP7_75t_SL g649 ( .A(n_547), .Y(n_649) );
INVx2_ASAP7_75t_SL g650 ( .A(n_547), .Y(n_650) );
AOI22xp5_ASAP7_75t_L g651 ( .A1(n_550), .A2(n_440), .B1(n_334), .B2(n_386), .Y(n_651) );
AOI22xp33_ASAP7_75t_L g652 ( .A1(n_550), .A2(n_528), .B1(n_389), .B2(n_390), .Y(n_652) );
OAI21xp5_ASAP7_75t_L g653 ( .A1(n_560), .A2(n_329), .B(n_327), .Y(n_653) );
NOR2xp33_ASAP7_75t_L g654 ( .A(n_546), .B(n_519), .Y(n_654) );
AND2x2_ASAP7_75t_L g655 ( .A(n_546), .B(n_338), .Y(n_655) );
NOR2xp33_ASAP7_75t_L g656 ( .A(n_546), .B(n_345), .Y(n_656) );
CKINVDCx20_ASAP7_75t_R g657 ( .A(n_546), .Y(n_657) );
INVx2_ASAP7_75t_L g658 ( .A(n_563), .Y(n_658) );
AND2x4_ASAP7_75t_L g659 ( .A(n_546), .B(n_388), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_563), .B(n_347), .Y(n_660) );
AND2x4_ASAP7_75t_L g661 ( .A(n_566), .B(n_461), .Y(n_661) );
INVx2_ASAP7_75t_SL g662 ( .A(n_566), .Y(n_662) );
NOR2x1_ASAP7_75t_L g663 ( .A(n_567), .B(n_331), .Y(n_663) );
AOI22xp33_ASAP7_75t_L g664 ( .A1(n_567), .A2(n_391), .B1(n_401), .B2(n_326), .Y(n_664) );
INVxp67_ASAP7_75t_SL g665 ( .A(n_569), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_569), .B(n_347), .Y(n_666) );
BUFx6f_ASAP7_75t_L g667 ( .A(n_579), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_570), .Y(n_668) );
CKINVDCx5p33_ASAP7_75t_R g669 ( .A(n_570), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_573), .B(n_361), .Y(n_670) );
INVx3_ASAP7_75t_L g671 ( .A(n_573), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_576), .Y(n_672) );
OAI22xp5_ASAP7_75t_SL g673 ( .A1(n_576), .A2(n_404), .B1(n_410), .B2(n_362), .Y(n_673) );
NOR2xp33_ASAP7_75t_L g674 ( .A(n_582), .B(n_361), .Y(n_674) );
INVx2_ASAP7_75t_SL g675 ( .A(n_582), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_533), .Y(n_676) );
INVx2_ASAP7_75t_SL g677 ( .A(n_579), .Y(n_677) );
AOI22xp33_ASAP7_75t_L g678 ( .A1(n_533), .A2(n_406), .B1(n_407), .B2(n_405), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_533), .B(n_375), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_541), .B(n_375), .Y(n_680) );
INVxp67_ASAP7_75t_L g681 ( .A(n_541), .Y(n_681) );
OAI22xp33_ASAP7_75t_L g682 ( .A1(n_541), .A2(n_489), .B1(n_338), .B2(n_441), .Y(n_682) );
NOR2x1p5_ASAP7_75t_L g683 ( .A(n_545), .B(n_386), .Y(n_683) );
AOI22xp5_ASAP7_75t_L g684 ( .A1(n_545), .A2(n_480), .B1(n_441), .B2(n_470), .Y(n_684) );
OAI22xp5_ASAP7_75t_SL g685 ( .A1(n_593), .A2(n_489), .B1(n_480), .B2(n_442), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_596), .B(n_409), .Y(n_686) );
BUFx2_ASAP7_75t_L g687 ( .A(n_587), .Y(n_687) );
BUFx12f_ASAP7_75t_L g688 ( .A(n_601), .Y(n_688) );
AO22x1_ASAP7_75t_L g689 ( .A1(n_623), .A2(n_442), .B1(n_445), .B2(n_393), .Y(n_689) );
BUFx2_ASAP7_75t_L g690 ( .A(n_627), .Y(n_690) );
BUFx6f_ASAP7_75t_L g691 ( .A(n_591), .Y(n_691) );
A2O1A1Ixp33_ASAP7_75t_L g692 ( .A1(n_622), .A2(n_411), .B(n_421), .C(n_418), .Y(n_692) );
INVx2_ASAP7_75t_SL g693 ( .A(n_661), .Y(n_693) );
AOI21x1_ASAP7_75t_L g694 ( .A1(n_648), .A2(n_551), .B(n_545), .Y(n_694) );
AOI21xp5_ASAP7_75t_L g695 ( .A1(n_649), .A2(n_371), .B(n_346), .Y(n_695) );
O2A1O1Ixp33_ASAP7_75t_L g696 ( .A1(n_592), .A2(n_433), .B(n_438), .C(n_429), .Y(n_696) );
OAI22xp5_ASAP7_75t_L g697 ( .A1(n_585), .A2(n_446), .B1(n_456), .B2(n_439), .Y(n_697) );
BUFx2_ASAP7_75t_L g698 ( .A(n_627), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_595), .Y(n_699) );
NAND2xp33_ASAP7_75t_SL g700 ( .A(n_584), .B(n_393), .Y(n_700) );
NOR2xp33_ASAP7_75t_L g701 ( .A(n_596), .B(n_457), .Y(n_701) );
BUFx3_ASAP7_75t_L g702 ( .A(n_610), .Y(n_702) );
AND2x2_ASAP7_75t_L g703 ( .A(n_603), .B(n_459), .Y(n_703) );
INVx5_ASAP7_75t_L g704 ( .A(n_584), .Y(n_704) );
AOI21xp5_ASAP7_75t_L g705 ( .A1(n_649), .A2(n_372), .B(n_343), .Y(n_705) );
CKINVDCx5p33_ASAP7_75t_R g706 ( .A(n_608), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_588), .B(n_590), .Y(n_707) );
NAND2x1_ASAP7_75t_SL g708 ( .A(n_633), .B(n_428), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g709 ( .A1(n_597), .A2(n_528), .B1(n_462), .B2(n_478), .Y(n_709) );
OAI22xp5_ASAP7_75t_L g710 ( .A1(n_585), .A2(n_486), .B1(n_490), .B2(n_463), .Y(n_710) );
BUFx3_ASAP7_75t_L g711 ( .A(n_607), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_583), .Y(n_712) );
A2O1A1Ixp33_ASAP7_75t_L g713 ( .A1(n_605), .A2(n_427), .B(n_434), .C(n_387), .Y(n_713) );
INVx1_ASAP7_75t_L g714 ( .A(n_586), .Y(n_714) );
INVx1_ASAP7_75t_L g715 ( .A(n_665), .Y(n_715) );
BUFx3_ASAP7_75t_L g716 ( .A(n_619), .Y(n_716) );
INVx5_ASAP7_75t_L g717 ( .A(n_634), .Y(n_717) );
AND2x2_ASAP7_75t_L g718 ( .A(n_651), .B(n_427), .Y(n_718) );
OAI22xp5_ASAP7_75t_L g719 ( .A1(n_612), .A2(n_434), .B1(n_528), .B2(n_378), .Y(n_719) );
AOI22xp33_ASAP7_75t_SL g720 ( .A1(n_589), .A2(n_445), .B1(n_452), .B2(n_448), .Y(n_720) );
NAND2xp5_ASAP7_75t_SL g721 ( .A(n_634), .B(n_448), .Y(n_721) );
CKINVDCx5p33_ASAP7_75t_R g722 ( .A(n_673), .Y(n_722) );
BUFx3_ASAP7_75t_L g723 ( .A(n_619), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_612), .B(n_452), .Y(n_724) );
INVxp67_ASAP7_75t_SL g725 ( .A(n_617), .Y(n_725) );
NOR2xp33_ASAP7_75t_L g726 ( .A(n_604), .B(n_460), .Y(n_726) );
BUFx12f_ASAP7_75t_L g727 ( .A(n_621), .Y(n_727) );
HB1xp67_ASAP7_75t_L g728 ( .A(n_682), .Y(n_728) );
BUFx3_ASAP7_75t_L g729 ( .A(n_657), .Y(n_729) );
AOI22xp33_ASAP7_75t_L g730 ( .A1(n_602), .A2(n_378), .B1(n_344), .B2(n_348), .Y(n_730) );
BUFx3_ASAP7_75t_L g731 ( .A(n_661), .Y(n_731) );
OR2x2_ASAP7_75t_L g732 ( .A(n_682), .B(n_460), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_599), .B(n_464), .Y(n_733) );
AOI21xp5_ASAP7_75t_L g734 ( .A1(n_625), .A2(n_349), .B(n_332), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_611), .B(n_464), .Y(n_735) );
INVx1_ASAP7_75t_L g736 ( .A(n_665), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_624), .Y(n_737) );
AND2x4_ASAP7_75t_L g738 ( .A(n_616), .B(n_350), .Y(n_738) );
NOR2xp67_ASAP7_75t_SL g739 ( .A(n_591), .B(n_398), .Y(n_739) );
BUFx6f_ASAP7_75t_L g740 ( .A(n_591), .Y(n_740) );
AOI21xp5_ASAP7_75t_L g741 ( .A1(n_650), .A2(n_353), .B(n_351), .Y(n_741) );
AND2x2_ASAP7_75t_L g742 ( .A(n_600), .B(n_378), .Y(n_742) );
O2A1O1Ixp33_ASAP7_75t_SL g743 ( .A1(n_626), .A2(n_360), .B(n_369), .C(n_358), .Y(n_743) );
INVx3_ASAP7_75t_L g744 ( .A(n_615), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_645), .B(n_376), .Y(n_745) );
AOI22xp5_ASAP7_75t_L g746 ( .A1(n_592), .A2(n_379), .B1(n_383), .B2(n_377), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_644), .B(n_385), .Y(n_747) );
CKINVDCx5p33_ASAP7_75t_R g748 ( .A(n_614), .Y(n_748) );
INVx1_ASAP7_75t_L g749 ( .A(n_631), .Y(n_749) );
BUFx6f_ASAP7_75t_L g750 ( .A(n_591), .Y(n_750) );
CKINVDCx5p33_ASAP7_75t_R g751 ( .A(n_606), .Y(n_751) );
BUFx6f_ASAP7_75t_L g752 ( .A(n_613), .Y(n_752) );
O2A1O1Ixp33_ASAP7_75t_L g753 ( .A1(n_598), .A2(n_395), .B(n_400), .C(n_394), .Y(n_753) );
BUFx6f_ASAP7_75t_L g754 ( .A(n_613), .Y(n_754) );
NAND2xp5_ASAP7_75t_SL g755 ( .A(n_613), .B(n_437), .Y(n_755) );
INVx1_ASAP7_75t_SL g756 ( .A(n_613), .Y(n_756) );
INVx3_ASAP7_75t_L g757 ( .A(n_609), .Y(n_757) );
INVx2_ASAP7_75t_L g758 ( .A(n_609), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_620), .B(n_403), .Y(n_759) );
BUFx3_ASAP7_75t_L g760 ( .A(n_659), .Y(n_760) );
INVx1_ASAP7_75t_L g761 ( .A(n_668), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_620), .B(n_412), .Y(n_762) );
HB1xp67_ASAP7_75t_L g763 ( .A(n_683), .Y(n_763) );
AND2x4_ASAP7_75t_L g764 ( .A(n_616), .B(n_416), .Y(n_764) );
INVx2_ASAP7_75t_L g765 ( .A(n_671), .Y(n_765) );
BUFx2_ASAP7_75t_L g766 ( .A(n_637), .Y(n_766) );
AND2x4_ASAP7_75t_L g767 ( .A(n_628), .B(n_630), .Y(n_767) );
INVx1_ASAP7_75t_L g768 ( .A(n_672), .Y(n_768) );
AND2x2_ASAP7_75t_SL g769 ( .A(n_635), .B(n_417), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_617), .B(n_419), .Y(n_770) );
INVx2_ASAP7_75t_L g771 ( .A(n_671), .Y(n_771) );
BUFx6f_ASAP7_75t_L g772 ( .A(n_618), .Y(n_772) );
OAI22xp5_ASAP7_75t_L g773 ( .A1(n_635), .A2(n_422), .B1(n_423), .B2(n_420), .Y(n_773) );
INVxp67_ASAP7_75t_L g774 ( .A(n_684), .Y(n_774) );
BUFx2_ASAP7_75t_L g775 ( .A(n_655), .Y(n_775) );
INVx1_ASAP7_75t_L g776 ( .A(n_669), .Y(n_776) );
INVx3_ASAP7_75t_L g777 ( .A(n_639), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_636), .B(n_426), .Y(n_778) );
INVx2_ASAP7_75t_L g779 ( .A(n_641), .Y(n_779) );
O2A1O1Ixp33_ASAP7_75t_L g780 ( .A1(n_653), .A2(n_449), .B(n_450), .C(n_431), .Y(n_780) );
INVx1_ASAP7_75t_L g781 ( .A(n_659), .Y(n_781) );
AOI22xp33_ASAP7_75t_SL g782 ( .A1(n_629), .A2(n_424), .B1(n_447), .B2(n_402), .Y(n_782) );
OR2x2_ASAP7_75t_L g783 ( .A(n_664), .B(n_11), .Y(n_783) );
INVx2_ASAP7_75t_L g784 ( .A(n_647), .Y(n_784) );
CKINVDCx6p67_ASAP7_75t_R g785 ( .A(n_629), .Y(n_785) );
BUFx6f_ASAP7_75t_L g786 ( .A(n_639), .Y(n_786) );
AOI221x1_ASAP7_75t_L g787 ( .A1(n_638), .A2(n_476), .B1(n_451), .B2(n_453), .C(n_454), .Y(n_787) );
HB1xp67_ASAP7_75t_L g788 ( .A(n_654), .Y(n_788) );
INVxp67_ASAP7_75t_L g789 ( .A(n_660), .Y(n_789) );
OAI22xp5_ASAP7_75t_L g790 ( .A1(n_636), .A2(n_465), .B1(n_467), .B2(n_458), .Y(n_790) );
INVxp67_ASAP7_75t_SL g791 ( .A(n_594), .Y(n_791) );
AOI21xp5_ASAP7_75t_L g792 ( .A1(n_632), .A2(n_469), .B(n_468), .Y(n_792) );
INVx1_ASAP7_75t_SL g793 ( .A(n_594), .Y(n_793) );
INVx2_ASAP7_75t_L g794 ( .A(n_658), .Y(n_794) );
OR2x6_ASAP7_75t_L g795 ( .A(n_663), .B(n_339), .Y(n_795) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_643), .B(n_471), .Y(n_796) );
O2A1O1Ixp33_ASAP7_75t_L g797 ( .A1(n_664), .A2(n_473), .B(n_475), .C(n_472), .Y(n_797) );
NOR2xp33_ASAP7_75t_L g798 ( .A(n_666), .B(n_466), .Y(n_798) );
OAI22xp5_ASAP7_75t_L g799 ( .A1(n_678), .A2(n_484), .B1(n_485), .B2(n_477), .Y(n_799) );
INVx3_ASAP7_75t_L g800 ( .A(n_594), .Y(n_800) );
INVx3_ASAP7_75t_L g801 ( .A(n_594), .Y(n_801) );
BUFx5_ASAP7_75t_L g802 ( .A(n_676), .Y(n_802) );
HB1xp67_ASAP7_75t_L g803 ( .A(n_670), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g804 ( .A(n_594), .B(n_488), .Y(n_804) );
INVx1_ASAP7_75t_L g805 ( .A(n_678), .Y(n_805) );
NOR2xp33_ASAP7_75t_L g806 ( .A(n_642), .B(n_646), .Y(n_806) );
INVx4_ASAP7_75t_L g807 ( .A(n_594), .Y(n_807) );
AND2x2_ASAP7_75t_L g808 ( .A(n_674), .B(n_12), .Y(n_808) );
BUFx6f_ASAP7_75t_L g809 ( .A(n_667), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_652), .B(n_491), .Y(n_810) );
INVx3_ASAP7_75t_L g811 ( .A(n_662), .Y(n_811) );
AOI21xp5_ASAP7_75t_L g812 ( .A1(n_640), .A2(n_492), .B(n_341), .Y(n_812) );
INVx1_ASAP7_75t_L g813 ( .A(n_679), .Y(n_813) );
BUFx6f_ASAP7_75t_L g814 ( .A(n_667), .Y(n_814) );
INVx3_ASAP7_75t_L g815 ( .A(n_675), .Y(n_815) );
AOI22xp5_ASAP7_75t_L g816 ( .A1(n_656), .A2(n_370), .B1(n_392), .B2(n_333), .Y(n_816) );
AOI22xp33_ASAP7_75t_L g817 ( .A1(n_680), .A2(n_424), .B1(n_447), .B2(n_402), .Y(n_817) );
AND2x6_ASAP7_75t_L g818 ( .A(n_667), .B(n_487), .Y(n_818) );
AOI22xp33_ASAP7_75t_L g819 ( .A1(n_681), .A2(n_487), .B1(n_436), .B2(n_479), .Y(n_819) );
AOI22xp5_ASAP7_75t_L g820 ( .A1(n_677), .A2(n_436), .B1(n_479), .B2(n_392), .Y(n_820) );
INVx4_ASAP7_75t_L g821 ( .A(n_667), .Y(n_821) );
BUFx3_ASAP7_75t_L g822 ( .A(n_601), .Y(n_822) );
INVx3_ASAP7_75t_L g823 ( .A(n_615), .Y(n_823) );
INVx1_ASAP7_75t_L g824 ( .A(n_595), .Y(n_824) );
INVx3_ASAP7_75t_L g825 ( .A(n_615), .Y(n_825) );
INVx2_ASAP7_75t_L g826 ( .A(n_615), .Y(n_826) );
O2A1O1Ixp5_ASAP7_75t_L g827 ( .A1(n_599), .A2(n_483), .B(n_580), .C(n_553), .Y(n_827) );
BUFx2_ASAP7_75t_L g828 ( .A(n_587), .Y(n_828) );
INVx2_ASAP7_75t_L g829 ( .A(n_615), .Y(n_829) );
INVx1_ASAP7_75t_L g830 ( .A(n_595), .Y(n_830) );
OAI22xp5_ASAP7_75t_L g831 ( .A1(n_585), .A2(n_501), .B1(n_497), .B2(n_500), .Y(n_831) );
INVx1_ASAP7_75t_L g832 ( .A(n_595), .Y(n_832) );
NAND2xp5_ASAP7_75t_SL g833 ( .A(n_584), .B(n_430), .Y(n_833) );
INVx1_ASAP7_75t_L g834 ( .A(n_595), .Y(n_834) );
BUFx3_ASAP7_75t_L g835 ( .A(n_601), .Y(n_835) );
AOI21xp5_ASAP7_75t_L g836 ( .A1(n_649), .A2(n_553), .B(n_551), .Y(n_836) );
BUFx2_ASAP7_75t_L g837 ( .A(n_587), .Y(n_837) );
BUFx12f_ASAP7_75t_L g838 ( .A(n_601), .Y(n_838) );
INVx2_ASAP7_75t_SL g839 ( .A(n_587), .Y(n_839) );
AOI21xp5_ASAP7_75t_L g840 ( .A1(n_649), .A2(n_553), .B(n_551), .Y(n_840) );
NAND2xp5_ASAP7_75t_L g841 ( .A(n_596), .B(n_497), .Y(n_841) );
BUFx3_ASAP7_75t_L g842 ( .A(n_601), .Y(n_842) );
O2A1O1Ixp33_ASAP7_75t_L g843 ( .A1(n_611), .A2(n_500), .B(n_514), .C(n_497), .Y(n_843) );
INVx2_ASAP7_75t_L g844 ( .A(n_802), .Y(n_844) );
OAI22xp5_ASAP7_75t_L g845 ( .A1(n_769), .A2(n_514), .B1(n_517), .B2(n_500), .Y(n_845) );
OR2x6_ASAP7_75t_L g846 ( .A(n_688), .B(n_514), .Y(n_846) );
NAND2x1p5_ASAP7_75t_L g847 ( .A(n_704), .B(n_717), .Y(n_847) );
AOI21xp33_ASAP7_75t_L g848 ( .A1(n_732), .A2(n_13), .B(n_14), .Y(n_848) );
OAI21x1_ASAP7_75t_L g849 ( .A1(n_694), .A2(n_840), .B(n_836), .Y(n_849) );
OAI22xp5_ASAP7_75t_L g850 ( .A1(n_728), .A2(n_529), .B1(n_531), .B2(n_517), .Y(n_850) );
OAI22xp5_ASAP7_75t_L g851 ( .A1(n_715), .A2(n_736), .B1(n_745), .B2(n_746), .Y(n_851) );
INVx1_ASAP7_75t_L g852 ( .A(n_702), .Y(n_852) );
O2A1O1Ixp33_ASAP7_75t_L g853 ( .A1(n_713), .A2(n_529), .B(n_531), .C(n_517), .Y(n_853) );
HB1xp67_ASAP7_75t_L g854 ( .A(n_704), .Y(n_854) );
NAND2x1p5_ASAP7_75t_L g855 ( .A(n_704), .B(n_517), .Y(n_855) );
OR2x6_ASAP7_75t_L g856 ( .A(n_838), .B(n_529), .Y(n_856) );
AO21x2_ASAP7_75t_L g857 ( .A1(n_812), .A2(n_531), .B(n_495), .Y(n_857) );
NOR2xp67_ASAP7_75t_L g858 ( .A(n_822), .B(n_15), .Y(n_858) );
AND2x2_ASAP7_75t_L g859 ( .A(n_687), .B(n_15), .Y(n_859) );
INVx8_ASAP7_75t_L g860 ( .A(n_704), .Y(n_860) );
INVx1_ASAP7_75t_L g861 ( .A(n_711), .Y(n_861) );
AOI22xp5_ASAP7_75t_L g862 ( .A1(n_751), .A2(n_495), .B1(n_521), .B2(n_493), .Y(n_862) );
INVx1_ASAP7_75t_L g863 ( .A(n_712), .Y(n_863) );
AND2x2_ASAP7_75t_L g864 ( .A(n_828), .B(n_16), .Y(n_864) );
INVx1_ASAP7_75t_L g865 ( .A(n_714), .Y(n_865) );
OAI22xp5_ASAP7_75t_L g866 ( .A1(n_745), .A2(n_521), .B1(n_495), .B2(n_19), .Y(n_866) );
OAI22xp5_ASAP7_75t_L g867 ( .A1(n_805), .A2(n_521), .B1(n_495), .B2(n_21), .Y(n_867) );
AND2x2_ASAP7_75t_L g868 ( .A(n_837), .B(n_16), .Y(n_868) );
OAI21x1_ASAP7_75t_L g869 ( .A1(n_827), .A2(n_521), .B(n_495), .Y(n_869) );
OA21x2_ASAP7_75t_L g870 ( .A1(n_787), .A2(n_521), .B(n_579), .Y(n_870) );
INVx1_ASAP7_75t_L g871 ( .A(n_699), .Y(n_871) );
AND2x2_ASAP7_75t_L g872 ( .A(n_839), .B(n_18), .Y(n_872) );
AOI222xp33_ASAP7_75t_L g873 ( .A1(n_685), .A2(n_18), .B1(n_21), .B2(n_23), .C1(n_24), .C2(n_25), .Y(n_873) );
AND2x4_ASAP7_75t_L g874 ( .A(n_716), .B(n_25), .Y(n_874) );
CKINVDCx6p67_ASAP7_75t_R g875 ( .A(n_835), .Y(n_875) );
INVx2_ASAP7_75t_L g876 ( .A(n_802), .Y(n_876) );
INVx3_ASAP7_75t_L g877 ( .A(n_717), .Y(n_877) );
OA21x2_ASAP7_75t_L g878 ( .A1(n_812), .A2(n_579), .B(n_107), .Y(n_878) );
NAND2xp5_ASAP7_75t_L g879 ( .A(n_707), .B(n_26), .Y(n_879) );
AND2x2_ASAP7_75t_L g880 ( .A(n_693), .B(n_26), .Y(n_880) );
INVx1_ASAP7_75t_L g881 ( .A(n_824), .Y(n_881) );
BUFx10_ASAP7_75t_L g882 ( .A(n_776), .Y(n_882) );
OA21x2_ASAP7_75t_L g883 ( .A1(n_804), .A2(n_108), .B(n_106), .Y(n_883) );
INVx1_ASAP7_75t_L g884 ( .A(n_830), .Y(n_884) );
INVx2_ASAP7_75t_L g885 ( .A(n_802), .Y(n_885) );
O2A1O1Ixp33_ASAP7_75t_L g886 ( .A1(n_696), .A2(n_27), .B(n_28), .C(n_29), .Y(n_886) );
OAI21x1_ASAP7_75t_L g887 ( .A1(n_800), .A2(n_112), .B(n_111), .Y(n_887) );
OA21x2_ASAP7_75t_L g888 ( .A1(n_804), .A2(n_114), .B(n_113), .Y(n_888) );
INVx1_ASAP7_75t_L g889 ( .A(n_832), .Y(n_889) );
AOI21xp5_ASAP7_75t_L g890 ( .A1(n_707), .A2(n_120), .B(n_118), .Y(n_890) );
NOR2xp67_ASAP7_75t_L g891 ( .A(n_842), .B(n_29), .Y(n_891) );
NOR2x1_ASAP7_75t_SL g892 ( .A(n_717), .B(n_31), .Y(n_892) );
AOI22xp5_ASAP7_75t_L g893 ( .A1(n_774), .A2(n_31), .B1(n_32), .B2(n_33), .Y(n_893) );
BUFx6f_ASAP7_75t_L g894 ( .A(n_809), .Y(n_894) );
NAND2xp5_ASAP7_75t_L g895 ( .A(n_735), .B(n_34), .Y(n_895) );
AOI22x1_ASAP7_75t_L g896 ( .A1(n_741), .A2(n_163), .B1(n_316), .B2(n_312), .Y(n_896) );
NAND2xp5_ASAP7_75t_L g897 ( .A(n_735), .B(n_35), .Y(n_897) );
INVx1_ASAP7_75t_L g898 ( .A(n_834), .Y(n_898) );
INVx2_ASAP7_75t_L g899 ( .A(n_802), .Y(n_899) );
AO21x2_ASAP7_75t_L g900 ( .A1(n_734), .A2(n_126), .B(n_125), .Y(n_900) );
HB1xp67_ASAP7_75t_L g901 ( .A(n_717), .Y(n_901) );
AND2x2_ASAP7_75t_L g902 ( .A(n_731), .B(n_35), .Y(n_902) );
OAI21x1_ASAP7_75t_L g903 ( .A1(n_801), .A2(n_128), .B(n_127), .Y(n_903) );
AOI22xp5_ASAP7_75t_L g904 ( .A1(n_789), .A2(n_36), .B1(n_37), .B2(n_38), .Y(n_904) );
AOI22xp33_ASAP7_75t_L g905 ( .A1(n_783), .A2(n_697), .B1(n_710), .B2(n_718), .Y(n_905) );
NAND2xp5_ASAP7_75t_L g906 ( .A(n_686), .B(n_37), .Y(n_906) );
OA21x2_ASAP7_75t_L g907 ( .A1(n_747), .A2(n_133), .B(n_131), .Y(n_907) );
INVx2_ASAP7_75t_L g908 ( .A(n_802), .Y(n_908) );
OAI21x1_ASAP7_75t_L g909 ( .A1(n_843), .A2(n_136), .B(n_135), .Y(n_909) );
INVx1_ASAP7_75t_L g910 ( .A(n_742), .Y(n_910) );
CKINVDCx5p33_ASAP7_75t_R g911 ( .A(n_706), .Y(n_911) );
OA21x2_ASAP7_75t_L g912 ( .A1(n_747), .A2(n_139), .B(n_137), .Y(n_912) );
OAI22xp5_ASAP7_75t_L g913 ( .A1(n_725), .A2(n_39), .B1(n_40), .B2(n_41), .Y(n_913) );
INVx2_ASAP7_75t_L g914 ( .A(n_784), .Y(n_914) );
OAI21x1_ASAP7_75t_L g915 ( .A1(n_843), .A2(n_144), .B(n_141), .Y(n_915) );
NAND2xp5_ASAP7_75t_SL g916 ( .A(n_793), .B(n_146), .Y(n_916) );
AO21x2_ASAP7_75t_L g917 ( .A1(n_734), .A2(n_152), .B(n_151), .Y(n_917) );
INVx2_ASAP7_75t_L g918 ( .A(n_794), .Y(n_918) );
NAND2xp5_ASAP7_75t_L g919 ( .A(n_686), .B(n_40), .Y(n_919) );
OAI21x1_ASAP7_75t_L g920 ( .A1(n_833), .A2(n_156), .B(n_155), .Y(n_920) );
OAI221xp5_ASAP7_75t_L g921 ( .A1(n_720), .A2(n_42), .B1(n_43), .B2(n_44), .C(n_45), .Y(n_921) );
OAI22xp5_ASAP7_75t_L g922 ( .A1(n_770), .A2(n_42), .B1(n_43), .B2(n_44), .Y(n_922) );
OAI21x1_ASAP7_75t_SL g923 ( .A1(n_719), .A2(n_45), .B(n_46), .Y(n_923) );
INVx2_ASAP7_75t_L g924 ( .A(n_761), .Y(n_924) );
INVx1_ASAP7_75t_L g925 ( .A(n_841), .Y(n_925) );
OAI21x1_ASAP7_75t_L g926 ( .A1(n_741), .A2(n_159), .B(n_158), .Y(n_926) );
INVx3_ASAP7_75t_L g927 ( .A(n_811), .Y(n_927) );
AND2x4_ASAP7_75t_L g928 ( .A(n_723), .B(n_46), .Y(n_928) );
INVx3_ASAP7_75t_L g929 ( .A(n_811), .Y(n_929) );
OAI21xp5_ASAP7_75t_L g930 ( .A1(n_705), .A2(n_161), .B(n_160), .Y(n_930) );
AO32x2_ASAP7_75t_L g931 ( .A1(n_719), .A2(n_49), .A3(n_50), .B1(n_51), .B2(n_52), .Y(n_931) );
A2O1A1Ixp33_ASAP7_75t_L g932 ( .A1(n_780), .A2(n_49), .B(n_51), .C(n_53), .Y(n_932) );
AOI22xp33_ASAP7_75t_L g933 ( .A1(n_697), .A2(n_53), .B1(n_54), .B2(n_55), .Y(n_933) );
NAND2xp5_ASAP7_75t_L g934 ( .A(n_701), .B(n_54), .Y(n_934) );
OAI21xp5_ASAP7_75t_L g935 ( .A1(n_705), .A2(n_695), .B(n_813), .Y(n_935) );
OAI22xp5_ASAP7_75t_L g936 ( .A1(n_770), .A2(n_55), .B1(n_56), .B2(n_58), .Y(n_936) );
AND2x2_ASAP7_75t_SL g937 ( .A(n_690), .B(n_56), .Y(n_937) );
INVx2_ASAP7_75t_SL g938 ( .A(n_729), .Y(n_938) );
INVx1_ASAP7_75t_L g939 ( .A(n_841), .Y(n_939) );
INVx1_ASAP7_75t_L g940 ( .A(n_703), .Y(n_940) );
NAND2xp5_ASAP7_75t_SL g941 ( .A(n_793), .B(n_165), .Y(n_941) );
AND2x4_ASAP7_75t_L g942 ( .A(n_698), .B(n_58), .Y(n_942) );
INVx2_ASAP7_75t_L g943 ( .A(n_768), .Y(n_943) );
NAND2xp5_ASAP7_75t_L g944 ( .A(n_692), .B(n_59), .Y(n_944) );
A2O1A1Ixp33_ASAP7_75t_L g945 ( .A1(n_753), .A2(n_59), .B(n_60), .C(n_62), .Y(n_945) );
CKINVDCx5p33_ASAP7_75t_R g946 ( .A(n_785), .Y(n_946) );
INVx4_ASAP7_75t_L g947 ( .A(n_815), .Y(n_947) );
INVx1_ASAP7_75t_SL g948 ( .A(n_689), .Y(n_948) );
OAI21xp5_ASAP7_75t_L g949 ( .A1(n_695), .A2(n_202), .B(n_311), .Y(n_949) );
AND2x4_ASAP7_75t_L g950 ( .A(n_815), .B(n_60), .Y(n_950) );
A2O1A1Ixp33_ASAP7_75t_L g951 ( .A1(n_797), .A2(n_63), .B(n_64), .C(n_65), .Y(n_951) );
INVx1_ASAP7_75t_L g952 ( .A(n_803), .Y(n_952) );
INVx2_ASAP7_75t_L g953 ( .A(n_765), .Y(n_953) );
INVx1_ASAP7_75t_L g954 ( .A(n_763), .Y(n_954) );
AOI21xp5_ASAP7_75t_L g955 ( .A1(n_792), .A2(n_201), .B(n_306), .Y(n_955) );
OAI22xp5_ASAP7_75t_L g956 ( .A1(n_788), .A2(n_64), .B1(n_65), .B2(n_66), .Y(n_956) );
INVx2_ASAP7_75t_L g957 ( .A(n_771), .Y(n_957) );
INVx1_ASAP7_75t_SL g958 ( .A(n_708), .Y(n_958) );
CKINVDCx5p33_ASAP7_75t_R g959 ( .A(n_727), .Y(n_959) );
BUFx2_ASAP7_75t_SL g960 ( .A(n_818), .Y(n_960) );
AO21x2_ASAP7_75t_L g961 ( .A1(n_792), .A2(n_206), .B(n_305), .Y(n_961) );
OA21x2_ASAP7_75t_L g962 ( .A1(n_817), .A2(n_200), .B(n_302), .Y(n_962) );
CKINVDCx6p67_ASAP7_75t_R g963 ( .A(n_818), .Y(n_963) );
AOI22xp33_ASAP7_75t_L g964 ( .A1(n_710), .A2(n_66), .B1(n_67), .B2(n_68), .Y(n_964) );
OAI21x1_ASAP7_75t_SL g965 ( .A1(n_807), .A2(n_762), .B(n_759), .Y(n_965) );
OAI21x1_ASAP7_75t_L g966 ( .A1(n_744), .A2(n_199), .B(n_300), .Y(n_966) );
BUFx3_ASAP7_75t_L g967 ( .A(n_691), .Y(n_967) );
AND2x4_ASAP7_75t_L g968 ( .A(n_767), .B(n_67), .Y(n_968) );
AND2x2_ASAP7_75t_L g969 ( .A(n_722), .B(n_68), .Y(n_969) );
INVx1_ASAP7_75t_L g970 ( .A(n_737), .Y(n_970) );
BUFx2_ASAP7_75t_L g971 ( .A(n_760), .Y(n_971) );
INVx1_ASAP7_75t_L g972 ( .A(n_796), .Y(n_972) );
OAI21x1_ASAP7_75t_L g973 ( .A1(n_744), .A2(n_198), .B(n_296), .Y(n_973) );
OAI21x1_ASAP7_75t_L g974 ( .A1(n_823), .A2(n_197), .B(n_294), .Y(n_974) );
INVx1_ASAP7_75t_L g975 ( .A(n_796), .Y(n_975) );
OAI21x1_ASAP7_75t_L g976 ( .A1(n_823), .A2(n_195), .B(n_293), .Y(n_976) );
INVx2_ASAP7_75t_L g977 ( .A(n_809), .Y(n_977) );
OAI21x1_ASAP7_75t_L g978 ( .A1(n_825), .A2(n_194), .B(n_290), .Y(n_978) );
INVx3_ASAP7_75t_L g979 ( .A(n_772), .Y(n_979) );
INVx2_ASAP7_75t_L g980 ( .A(n_809), .Y(n_980) );
OAI21x1_ASAP7_75t_L g981 ( .A1(n_825), .A2(n_193), .B(n_289), .Y(n_981) );
BUFx4f_ASAP7_75t_L g982 ( .A(n_818), .Y(n_982) );
BUFx10_ASAP7_75t_L g983 ( .A(n_818), .Y(n_983) );
AOI21x1_ASAP7_75t_L g984 ( .A1(n_739), .A2(n_191), .B(n_287), .Y(n_984) );
AND2x4_ASAP7_75t_L g985 ( .A(n_767), .B(n_69), .Y(n_985) );
INVx2_ASAP7_75t_L g986 ( .A(n_814), .Y(n_986) );
OA21x2_ASAP7_75t_L g987 ( .A1(n_816), .A2(n_211), .B(n_285), .Y(n_987) );
O2A1O1Ixp33_ASAP7_75t_L g988 ( .A1(n_773), .A2(n_70), .B(n_72), .C(n_73), .Y(n_988) );
AO32x2_ASAP7_75t_L g989 ( .A1(n_773), .A2(n_70), .A3(n_72), .B1(n_73), .B2(n_74), .Y(n_989) );
INVx1_ASAP7_75t_SL g990 ( .A(n_775), .Y(n_990) );
OAI21xp5_ASAP7_75t_L g991 ( .A1(n_749), .A2(n_212), .B(n_284), .Y(n_991) );
INVx2_ASAP7_75t_L g992 ( .A(n_814), .Y(n_992) );
INVx2_ASAP7_75t_L g993 ( .A(n_814), .Y(n_993) );
NAND2xp5_ASAP7_75t_L g994 ( .A(n_730), .B(n_74), .Y(n_994) );
HB1xp67_ASAP7_75t_L g995 ( .A(n_766), .Y(n_995) );
NAND2xp5_ASAP7_75t_L g996 ( .A(n_724), .B(n_75), .Y(n_996) );
BUFx3_ASAP7_75t_L g997 ( .A(n_691), .Y(n_997) );
INVx1_ASAP7_75t_L g998 ( .A(n_808), .Y(n_998) );
INVx1_ASAP7_75t_L g999 ( .A(n_738), .Y(n_999) );
AOI22xp33_ASAP7_75t_L g1000 ( .A1(n_790), .A2(n_76), .B1(n_77), .B2(n_79), .Y(n_1000) );
INVx2_ASAP7_75t_L g1001 ( .A(n_779), .Y(n_1001) );
AND2x4_ASAP7_75t_L g1002 ( .A(n_781), .B(n_76), .Y(n_1002) );
AND2x6_ASAP7_75t_L g1003 ( .A(n_772), .B(n_166), .Y(n_1003) );
AND2x4_ASAP7_75t_L g1004 ( .A(n_757), .B(n_79), .Y(n_1004) );
AOI22xp33_ASAP7_75t_L g1005 ( .A1(n_790), .A2(n_80), .B1(n_81), .B2(n_82), .Y(n_1005) );
AND2x2_ASAP7_75t_L g1006 ( .A(n_726), .B(n_80), .Y(n_1006) );
INVx1_ASAP7_75t_L g1007 ( .A(n_738), .Y(n_1007) );
BUFx5_ASAP7_75t_L g1008 ( .A(n_764), .Y(n_1008) );
CKINVDCx5p33_ASAP7_75t_R g1009 ( .A(n_748), .Y(n_1009) );
OR2x2_ASAP7_75t_L g1010 ( .A(n_733), .B(n_81), .Y(n_1010) );
INVx1_ASAP7_75t_L g1011 ( .A(n_764), .Y(n_1011) );
INVx3_ASAP7_75t_L g1012 ( .A(n_772), .Y(n_1012) );
O2A1O1Ixp33_ASAP7_75t_SL g1013 ( .A1(n_755), .A2(n_216), .B(n_280), .C(n_279), .Y(n_1013) );
INVx1_ASAP7_75t_L g1014 ( .A(n_810), .Y(n_1014) );
OA21x2_ASAP7_75t_L g1015 ( .A1(n_820), .A2(n_187), .B(n_277), .Y(n_1015) );
AOI221xp5_ASAP7_75t_L g1016 ( .A1(n_940), .A2(n_799), .B1(n_798), .B2(n_778), .C(n_762), .Y(n_1016) );
AO21x2_ASAP7_75t_L g1017 ( .A1(n_965), .A2(n_759), .B(n_778), .Y(n_1017) );
AOI22xp33_ASAP7_75t_L g1018 ( .A1(n_937), .A2(n_799), .B1(n_795), .B2(n_810), .Y(n_1018) );
NAND2xp5_ASAP7_75t_L g1019 ( .A(n_905), .B(n_733), .Y(n_1019) );
INVx1_ASAP7_75t_L g1020 ( .A(n_871), .Y(n_1020) );
INVx2_ASAP7_75t_L g1021 ( .A(n_924), .Y(n_1021) );
OAI211xp5_ASAP7_75t_L g1022 ( .A1(n_873), .A2(n_782), .B(n_819), .C(n_743), .Y(n_1022) );
INVx3_ASAP7_75t_L g1023 ( .A(n_860), .Y(n_1023) );
OAI22xp5_ASAP7_75t_L g1024 ( .A1(n_905), .A2(n_724), .B1(n_709), .B2(n_795), .Y(n_1024) );
OAI21xp5_ASAP7_75t_L g1025 ( .A1(n_851), .A2(n_721), .B(n_700), .Y(n_1025) );
BUFx3_ASAP7_75t_L g1026 ( .A(n_875), .Y(n_1026) );
AOI221xp5_ASAP7_75t_L g1027 ( .A1(n_998), .A2(n_831), .B1(n_757), .B2(n_758), .C(n_777), .Y(n_1027) );
AOI21xp5_ASAP7_75t_L g1028 ( .A1(n_849), .A2(n_791), .B(n_829), .Y(n_1028) );
OAI22xp5_ASAP7_75t_L g1029 ( .A1(n_925), .A2(n_795), .B1(n_807), .B2(n_756), .Y(n_1029) );
AOI21xp5_ASAP7_75t_L g1030 ( .A1(n_869), .A2(n_826), .B(n_821), .Y(n_1030) );
AND2x2_ASAP7_75t_L g1031 ( .A(n_937), .B(n_82), .Y(n_1031) );
INVx2_ASAP7_75t_L g1032 ( .A(n_924), .Y(n_1032) );
INVx2_ASAP7_75t_L g1033 ( .A(n_943), .Y(n_1033) );
AOI22xp33_ASAP7_75t_L g1034 ( .A1(n_935), .A2(n_831), .B1(n_777), .B2(n_786), .Y(n_1034) );
AOI22xp33_ASAP7_75t_L g1035 ( .A1(n_944), .A2(n_786), .B1(n_756), .B2(n_752), .Y(n_1035) );
NOR3xp33_ASAP7_75t_L g1036 ( .A(n_886), .B(n_821), .C(n_84), .Y(n_1036) );
OAI221xp5_ASAP7_75t_L g1037 ( .A1(n_990), .A2(n_786), .B1(n_754), .B2(n_752), .C(n_750), .Y(n_1037) );
AOI222xp33_ASAP7_75t_L g1038 ( .A1(n_863), .A2(n_754), .B1(n_752), .B2(n_750), .C1(n_740), .C2(n_691), .Y(n_1038) );
AOI22xp33_ASAP7_75t_L g1039 ( .A1(n_972), .A2(n_754), .B1(n_750), .B2(n_740), .Y(n_1039) );
INVx1_ASAP7_75t_L g1040 ( .A(n_881), .Y(n_1040) );
AOI221xp5_ASAP7_75t_L g1041 ( .A1(n_865), .A2(n_740), .B1(n_84), .B2(n_85), .C(n_86), .Y(n_1041) );
INVx2_ASAP7_75t_L g1042 ( .A(n_943), .Y(n_1042) );
INVx2_ASAP7_75t_L g1043 ( .A(n_914), .Y(n_1043) );
HB1xp67_ASAP7_75t_L g1044 ( .A(n_995), .Y(n_1044) );
OAI22xp5_ASAP7_75t_L g1045 ( .A1(n_939), .A2(n_83), .B1(n_85), .B2(n_87), .Y(n_1045) );
INVx1_ASAP7_75t_L g1046 ( .A(n_884), .Y(n_1046) );
NAND3xp33_ASAP7_75t_L g1047 ( .A(n_932), .B(n_83), .C(n_87), .Y(n_1047) );
BUFx2_ASAP7_75t_L g1048 ( .A(n_846), .Y(n_1048) );
AOI22xp33_ASAP7_75t_L g1049 ( .A1(n_942), .A2(n_88), .B1(n_89), .B2(n_90), .Y(n_1049) );
AOI221xp5_ASAP7_75t_L g1050 ( .A1(n_952), .A2(n_88), .B1(n_89), .B2(n_90), .C(n_91), .Y(n_1050) );
OAI22xp5_ASAP7_75t_L g1051 ( .A1(n_942), .A2(n_92), .B1(n_94), .B2(n_95), .Y(n_1051) );
INVx1_ASAP7_75t_L g1052 ( .A(n_889), .Y(n_1052) );
BUFx4f_ASAP7_75t_SL g1053 ( .A(n_963), .Y(n_1053) );
AOI222xp33_ASAP7_75t_L g1054 ( .A1(n_969), .A2(n_92), .B1(n_94), .B2(n_95), .C1(n_96), .C2(n_97), .Y(n_1054) );
INVx1_ASAP7_75t_L g1055 ( .A(n_898), .Y(n_1055) );
BUFx4f_ASAP7_75t_SL g1056 ( .A(n_938), .Y(n_1056) );
OAI22xp5_ASAP7_75t_L g1057 ( .A1(n_942), .A2(n_96), .B1(n_99), .B2(n_100), .Y(n_1057) );
INVx2_ASAP7_75t_L g1058 ( .A(n_914), .Y(n_1058) );
AOI221xp5_ASAP7_75t_L g1059 ( .A1(n_886), .A2(n_100), .B1(n_102), .B2(n_103), .C(n_104), .Y(n_1059) );
A2O1A1Ixp33_ASAP7_75t_L g1060 ( .A1(n_988), .A2(n_102), .B(n_103), .C(n_104), .Y(n_1060) );
AOI21xp5_ASAP7_75t_L g1061 ( .A1(n_895), .A2(n_243), .B(n_172), .Y(n_1061) );
INVx1_ASAP7_75t_L g1062 ( .A(n_970), .Y(n_1062) );
OAI22xp5_ASAP7_75t_L g1063 ( .A1(n_1002), .A2(n_105), .B1(n_173), .B2(n_175), .Y(n_1063) );
OAI22xp5_ASAP7_75t_SL g1064 ( .A1(n_911), .A2(n_178), .B1(n_182), .B2(n_183), .Y(n_1064) );
AOI22xp5_ASAP7_75t_L g1065 ( .A1(n_874), .A2(n_185), .B1(n_186), .B2(n_228), .Y(n_1065) );
OAI22xp5_ASAP7_75t_L g1066 ( .A1(n_1002), .A2(n_229), .B1(n_233), .B2(n_234), .Y(n_1066) );
AND2x2_ASAP7_75t_L g1067 ( .A(n_995), .B(n_235), .Y(n_1067) );
AND2x2_ASAP7_75t_L g1068 ( .A(n_859), .B(n_236), .Y(n_1068) );
AOI221xp5_ASAP7_75t_L g1069 ( .A1(n_975), .A2(n_238), .B1(n_241), .B2(n_244), .C(n_245), .Y(n_1069) );
AOI221xp5_ASAP7_75t_L g1070 ( .A1(n_848), .A2(n_246), .B1(n_251), .B2(n_252), .C(n_254), .Y(n_1070) );
INVx4_ASAP7_75t_L g1071 ( .A(n_860), .Y(n_1071) );
HB1xp67_ASAP7_75t_L g1072 ( .A(n_1004), .Y(n_1072) );
AOI21xp5_ASAP7_75t_L g1073 ( .A1(n_897), .A2(n_255), .B(n_257), .Y(n_1073) );
A2O1A1Ixp33_ASAP7_75t_L g1074 ( .A1(n_988), .A2(n_258), .B(n_260), .C(n_261), .Y(n_1074) );
INVx3_ASAP7_75t_L g1075 ( .A(n_860), .Y(n_1075) );
AND2x2_ASAP7_75t_L g1076 ( .A(n_864), .B(n_265), .Y(n_1076) );
AOI221xp5_ASAP7_75t_L g1077 ( .A1(n_868), .A2(n_267), .B1(n_270), .B2(n_274), .C(n_318), .Y(n_1077) );
AOI21xp33_ASAP7_75t_L g1078 ( .A1(n_996), .A2(n_879), .B(n_934), .Y(n_1078) );
BUFx12f_ASAP7_75t_L g1079 ( .A(n_946), .Y(n_1079) );
OAI22xp5_ASAP7_75t_L g1080 ( .A1(n_1002), .A2(n_968), .B1(n_985), .B2(n_919), .Y(n_1080) );
OAI221xp5_ASAP7_75t_L g1081 ( .A1(n_958), .A2(n_948), .B1(n_906), .B2(n_893), .C(n_945), .Y(n_1081) );
INVxp67_ASAP7_75t_L g1082 ( .A(n_950), .Y(n_1082) );
INVx1_ASAP7_75t_L g1083 ( .A(n_872), .Y(n_1083) );
HB1xp67_ASAP7_75t_L g1084 ( .A(n_1004), .Y(n_1084) );
OAI22xp5_ASAP7_75t_L g1085 ( .A1(n_968), .A2(n_985), .B1(n_928), .B2(n_874), .Y(n_1085) );
AOI221xp5_ASAP7_75t_L g1086 ( .A1(n_1014), .A2(n_956), .B1(n_954), .B2(n_922), .C(n_936), .Y(n_1086) );
INVx3_ASAP7_75t_L g1087 ( .A(n_847), .Y(n_1087) );
INVx1_ASAP7_75t_L g1088 ( .A(n_874), .Y(n_1088) );
OAI22xp5_ASAP7_75t_L g1089 ( .A1(n_968), .A2(n_985), .B1(n_928), .B2(n_964), .Y(n_1089) );
INVx1_ASAP7_75t_L g1090 ( .A(n_928), .Y(n_1090) );
OAI211xp5_ASAP7_75t_L g1091 ( .A1(n_933), .A2(n_964), .B(n_904), .C(n_1000), .Y(n_1091) );
AOI21xp33_ASAP7_75t_L g1092 ( .A1(n_1010), .A2(n_853), .B(n_845), .Y(n_1092) );
AOI22xp5_ASAP7_75t_L g1093 ( .A1(n_950), .A2(n_1006), .B1(n_999), .B2(n_1011), .Y(n_1093) );
AOI22xp33_ASAP7_75t_L g1094 ( .A1(n_921), .A2(n_933), .B1(n_1005), .B2(n_1000), .Y(n_1094) );
NAND2xp5_ASAP7_75t_L g1095 ( .A(n_1007), .B(n_852), .Y(n_1095) );
AOI22xp33_ASAP7_75t_L g1096 ( .A1(n_1005), .A2(n_950), .B1(n_913), .B2(n_910), .Y(n_1096) );
NAND2xp33_ASAP7_75t_SL g1097 ( .A(n_854), .B(n_901), .Y(n_1097) );
AOI22xp33_ASAP7_75t_L g1098 ( .A1(n_923), .A2(n_1004), .B1(n_994), .B2(n_880), .Y(n_1098) );
OAI22xp5_ASAP7_75t_L g1099 ( .A1(n_982), .A2(n_856), .B1(n_846), .B2(n_918), .Y(n_1099) );
AOI21xp5_ASAP7_75t_L g1100 ( .A1(n_857), .A2(n_916), .B(n_941), .Y(n_1100) );
AOI222xp33_ASAP7_75t_L g1101 ( .A1(n_911), .A2(n_861), .B1(n_1009), .B2(n_902), .C1(n_959), .C2(n_891), .Y(n_1101) );
AOI21xp5_ASAP7_75t_L g1102 ( .A1(n_916), .A2(n_941), .B(n_853), .Y(n_1102) );
OAI22xp33_ASAP7_75t_L g1103 ( .A1(n_846), .A2(n_856), .B1(n_982), .B2(n_858), .Y(n_1103) );
NAND2xp5_ASAP7_75t_L g1104 ( .A(n_1008), .B(n_947), .Y(n_1104) );
INVx1_ASAP7_75t_L g1105 ( .A(n_989), .Y(n_1105) );
AOI221xp5_ASAP7_75t_L g1106 ( .A1(n_866), .A2(n_945), .B1(n_951), .B2(n_932), .C(n_971), .Y(n_1106) );
OAI21xp33_ASAP7_75t_L g1107 ( .A1(n_951), .A2(n_862), .B(n_930), .Y(n_1107) );
AND2x4_ASAP7_75t_L g1108 ( .A(n_947), .B(n_927), .Y(n_1108) );
AOI22xp33_ASAP7_75t_L g1109 ( .A1(n_1008), .A2(n_856), .B1(n_1001), .B2(n_867), .Y(n_1109) );
BUFx3_ASAP7_75t_L g1110 ( .A(n_946), .Y(n_1110) );
AOI22xp33_ASAP7_75t_L g1111 ( .A1(n_1008), .A2(n_957), .B1(n_953), .B2(n_949), .Y(n_1111) );
OAI22xp5_ASAP7_75t_L g1112 ( .A1(n_960), .A2(n_901), .B1(n_854), .B2(n_908), .Y(n_1112) );
AOI221xp5_ASAP7_75t_L g1113 ( .A1(n_1009), .A2(n_850), .B1(n_959), .B2(n_927), .C(n_929), .Y(n_1113) );
INVx1_ASAP7_75t_L g1114 ( .A(n_989), .Y(n_1114) );
INVx2_ASAP7_75t_L g1115 ( .A(n_953), .Y(n_1115) );
OA21x2_ASAP7_75t_L g1116 ( .A1(n_909), .A2(n_915), .B(n_991), .Y(n_1116) );
AOI22xp33_ASAP7_75t_L g1117 ( .A1(n_1008), .A2(n_957), .B1(n_882), .B2(n_1003), .Y(n_1117) );
INVx2_ASAP7_75t_L g1118 ( .A(n_967), .Y(n_1118) );
AOI22xp33_ASAP7_75t_L g1119 ( .A1(n_1008), .A2(n_882), .B1(n_929), .B2(n_877), .Y(n_1119) );
NAND2xp5_ASAP7_75t_L g1120 ( .A(n_1008), .B(n_979), .Y(n_1120) );
AOI22xp33_ASAP7_75t_L g1121 ( .A1(n_1003), .A2(n_900), .B1(n_917), .B2(n_961), .Y(n_1121) );
INVx4_ASAP7_75t_SL g1122 ( .A(n_1003), .Y(n_1122) );
OAI22xp5_ASAP7_75t_L g1123 ( .A1(n_844), .A2(n_885), .B1(n_908), .B2(n_899), .Y(n_1123) );
INVx2_ASAP7_75t_L g1124 ( .A(n_967), .Y(n_1124) );
OAI221xp5_ASAP7_75t_L g1125 ( .A1(n_955), .A2(n_890), .B1(n_896), .B2(n_962), .C(n_987), .Y(n_1125) );
NAND2xp5_ASAP7_75t_L g1126 ( .A(n_979), .B(n_1012), .Y(n_1126) );
AOI22xp33_ASAP7_75t_L g1127 ( .A1(n_877), .A2(n_844), .B1(n_885), .B2(n_899), .Y(n_1127) );
NAND2xp5_ASAP7_75t_L g1128 ( .A(n_1012), .B(n_997), .Y(n_1128) );
AOI22xp33_ASAP7_75t_L g1129 ( .A1(n_1003), .A2(n_917), .B1(n_900), .B2(n_961), .Y(n_1129) );
INVx2_ASAP7_75t_L g1130 ( .A(n_997), .Y(n_1130) );
OAI221xp5_ASAP7_75t_L g1131 ( .A1(n_955), .A2(n_962), .B1(n_987), .B2(n_1015), .C(n_847), .Y(n_1131) );
AOI21xp5_ASAP7_75t_L g1132 ( .A1(n_878), .A2(n_977), .B(n_992), .Y(n_1132) );
INVx3_ASAP7_75t_L g1133 ( .A(n_983), .Y(n_1133) );
OAI221xp5_ASAP7_75t_L g1134 ( .A1(n_1015), .A2(n_870), .B1(n_855), .B2(n_876), .C(n_883), .Y(n_1134) );
INVx2_ASAP7_75t_L g1135 ( .A(n_966), .Y(n_1135) );
NAND2xp5_ASAP7_75t_L g1136 ( .A(n_876), .B(n_892), .Y(n_1136) );
OAI22xp5_ASAP7_75t_L g1137 ( .A1(n_855), .A2(n_870), .B1(n_894), .B2(n_1015), .Y(n_1137) );
AOI21xp5_ASAP7_75t_L g1138 ( .A1(n_878), .A2(n_977), .B(n_993), .Y(n_1138) );
AOI31xp33_ASAP7_75t_L g1139 ( .A1(n_1013), .A2(n_983), .A3(n_931), .B(n_1003), .Y(n_1139) );
OAI21xp5_ASAP7_75t_L g1140 ( .A1(n_926), .A2(n_920), .B(n_992), .Y(n_1140) );
OAI221xp5_ASAP7_75t_L g1141 ( .A1(n_883), .A2(n_888), .B1(n_912), .B2(n_907), .C(n_1013), .Y(n_1141) );
NAND2xp5_ASAP7_75t_L g1142 ( .A(n_980), .B(n_986), .Y(n_1142) );
BUFx6f_ASAP7_75t_L g1143 ( .A(n_894), .Y(n_1143) );
NAND2xp5_ASAP7_75t_L g1144 ( .A(n_980), .B(n_986), .Y(n_1144) );
AOI22xp33_ASAP7_75t_L g1145 ( .A1(n_907), .A2(n_912), .B1(n_888), .B2(n_887), .Y(n_1145) );
OAI221xp5_ASAP7_75t_SL g1146 ( .A1(n_989), .A2(n_931), .B1(n_903), .B2(n_974), .C(n_973), .Y(n_1146) );
OAI21xp33_ASAP7_75t_L g1147 ( .A1(n_976), .A2(n_978), .B(n_981), .Y(n_1147) );
AND2x4_ASAP7_75t_L g1148 ( .A(n_894), .B(n_984), .Y(n_1148) );
A2O1A1Ixp33_ASAP7_75t_L g1149 ( .A1(n_894), .A2(n_935), .B(n_886), .C(n_806), .Y(n_1149) );
AOI22xp33_ASAP7_75t_L g1150 ( .A1(n_931), .A2(n_937), .B1(n_751), .B2(n_905), .Y(n_1150) );
NAND2xp5_ASAP7_75t_L g1151 ( .A(n_989), .B(n_931), .Y(n_1151) );
OAI221xp5_ASAP7_75t_L g1152 ( .A1(n_905), .A2(n_605), .B1(n_839), .B2(n_828), .C(n_837), .Y(n_1152) );
AOI22xp33_ASAP7_75t_SL g1153 ( .A1(n_937), .A2(n_623), .B1(n_589), .B2(n_593), .Y(n_1153) );
OR2x2_ASAP7_75t_L g1154 ( .A(n_990), .B(n_523), .Y(n_1154) );
NAND2xp5_ASAP7_75t_L g1155 ( .A(n_905), .B(n_592), .Y(n_1155) );
INVx1_ASAP7_75t_L g1156 ( .A(n_871), .Y(n_1156) );
OAI22xp5_ASAP7_75t_L g1157 ( .A1(n_905), .A2(n_769), .B1(n_633), .B2(n_851), .Y(n_1157) );
INVx1_ASAP7_75t_L g1158 ( .A(n_871), .Y(n_1158) );
INVx1_ASAP7_75t_L g1159 ( .A(n_871), .Y(n_1159) );
AOI22xp33_ASAP7_75t_L g1160 ( .A1(n_937), .A2(n_751), .B1(n_905), .B2(n_851), .Y(n_1160) );
BUFx2_ASAP7_75t_L g1161 ( .A(n_846), .Y(n_1161) );
OAI211xp5_ASAP7_75t_L g1162 ( .A1(n_873), .A2(n_708), .B(n_746), .C(n_602), .Y(n_1162) );
AOI22xp33_ASAP7_75t_L g1163 ( .A1(n_937), .A2(n_751), .B1(n_905), .B2(n_851), .Y(n_1163) );
BUFx2_ASAP7_75t_L g1164 ( .A(n_846), .Y(n_1164) );
OAI22xp33_ASAP7_75t_L g1165 ( .A1(n_851), .A2(n_633), .B1(n_623), .B2(n_589), .Y(n_1165) );
OR2x2_ASAP7_75t_L g1166 ( .A(n_990), .B(n_523), .Y(n_1166) );
INVx1_ASAP7_75t_L g1167 ( .A(n_871), .Y(n_1167) );
BUFx3_ASAP7_75t_L g1168 ( .A(n_1071), .Y(n_1168) );
OR2x2_ASAP7_75t_L g1169 ( .A(n_1085), .B(n_1155), .Y(n_1169) );
AND2x2_ASAP7_75t_L g1170 ( .A(n_1021), .B(n_1032), .Y(n_1170) );
INVx2_ASAP7_75t_L g1171 ( .A(n_1033), .Y(n_1171) );
AND2x2_ASAP7_75t_L g1172 ( .A(n_1042), .B(n_1043), .Y(n_1172) );
HB1xp67_ASAP7_75t_L g1173 ( .A(n_1044), .Y(n_1173) );
INVxp67_ASAP7_75t_L g1174 ( .A(n_1154), .Y(n_1174) );
INVx1_ASAP7_75t_L g1175 ( .A(n_1058), .Y(n_1175) );
INVx1_ASAP7_75t_L g1176 ( .A(n_1115), .Y(n_1176) );
OR2x2_ASAP7_75t_L g1177 ( .A(n_1089), .B(n_1044), .Y(n_1177) );
BUFx6f_ASAP7_75t_L g1178 ( .A(n_1143), .Y(n_1178) );
NOR2xp33_ASAP7_75t_L g1179 ( .A(n_1153), .B(n_1152), .Y(n_1179) );
HB1xp67_ASAP7_75t_L g1180 ( .A(n_1087), .Y(n_1180) );
AND2x2_ASAP7_75t_L g1181 ( .A(n_1020), .B(n_1040), .Y(n_1181) );
INVx1_ASAP7_75t_L g1182 ( .A(n_1105), .Y(n_1182) );
OAI31xp33_ASAP7_75t_SL g1183 ( .A1(n_1153), .A2(n_1157), .A3(n_1103), .B(n_1165), .Y(n_1183) );
INVx1_ASAP7_75t_L g1184 ( .A(n_1114), .Y(n_1184) );
AND2x2_ASAP7_75t_L g1185 ( .A(n_1046), .B(n_1052), .Y(n_1185) );
AND2x2_ASAP7_75t_L g1186 ( .A(n_1055), .B(n_1156), .Y(n_1186) );
INVx1_ASAP7_75t_L g1187 ( .A(n_1151), .Y(n_1187) );
NAND2xp5_ASAP7_75t_L g1188 ( .A(n_1160), .B(n_1163), .Y(n_1188) );
INVx1_ASAP7_75t_L g1189 ( .A(n_1158), .Y(n_1189) );
NOR2xp33_ASAP7_75t_L g1190 ( .A(n_1166), .B(n_1162), .Y(n_1190) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1159), .Y(n_1191) );
INVx1_ASAP7_75t_L g1192 ( .A(n_1167), .Y(n_1192) );
AND2x2_ASAP7_75t_L g1193 ( .A(n_1062), .B(n_1160), .Y(n_1193) );
OR2x2_ASAP7_75t_L g1194 ( .A(n_1019), .B(n_1072), .Y(n_1194) );
INVxp67_ASAP7_75t_SL g1195 ( .A(n_1072), .Y(n_1195) );
HB1xp67_ASAP7_75t_L g1196 ( .A(n_1087), .Y(n_1196) );
AND2x2_ASAP7_75t_L g1197 ( .A(n_1163), .B(n_1084), .Y(n_1197) );
OR2x2_ASAP7_75t_L g1198 ( .A(n_1084), .B(n_1080), .Y(n_1198) );
INVxp67_ASAP7_75t_SL g1199 ( .A(n_1082), .Y(n_1199) );
AND2x2_ASAP7_75t_L g1200 ( .A(n_1150), .B(n_1031), .Y(n_1200) );
AND2x2_ASAP7_75t_L g1201 ( .A(n_1150), .B(n_1082), .Y(n_1201) );
INVx1_ASAP7_75t_L g1202 ( .A(n_1142), .Y(n_1202) );
INVx2_ASAP7_75t_L g1203 ( .A(n_1148), .Y(n_1203) );
INVx2_ASAP7_75t_SL g1204 ( .A(n_1071), .Y(n_1204) );
OR2x2_ASAP7_75t_L g1205 ( .A(n_1088), .B(n_1090), .Y(n_1205) );
AND2x4_ASAP7_75t_L g1206 ( .A(n_1122), .B(n_1117), .Y(n_1206) );
AND2x2_ASAP7_75t_L g1207 ( .A(n_1096), .B(n_1018), .Y(n_1207) );
INVx1_ASAP7_75t_L g1208 ( .A(n_1144), .Y(n_1208) );
INVx1_ASAP7_75t_L g1209 ( .A(n_1017), .Y(n_1209) );
AND2x2_ASAP7_75t_L g1210 ( .A(n_1096), .B(n_1018), .Y(n_1210) );
AND2x2_ASAP7_75t_L g1211 ( .A(n_1067), .B(n_1036), .Y(n_1211) );
NAND2xp5_ASAP7_75t_L g1212 ( .A(n_1165), .B(n_1016), .Y(n_1212) );
AND2x2_ASAP7_75t_L g1213 ( .A(n_1036), .B(n_1083), .Y(n_1213) );
INVx3_ASAP7_75t_SL g1214 ( .A(n_1122), .Y(n_1214) );
NAND2xp5_ASAP7_75t_L g1215 ( .A(n_1086), .B(n_1093), .Y(n_1215) );
INVx2_ASAP7_75t_SL g1216 ( .A(n_1023), .Y(n_1216) );
INVx1_ASAP7_75t_L g1217 ( .A(n_1017), .Y(n_1217) );
OR2x2_ASAP7_75t_L g1218 ( .A(n_1048), .B(n_1161), .Y(n_1218) );
NAND2xp5_ASAP7_75t_L g1219 ( .A(n_1101), .B(n_1054), .Y(n_1219) );
INVx1_ASAP7_75t_L g1220 ( .A(n_1136), .Y(n_1220) );
INVx1_ASAP7_75t_L g1221 ( .A(n_1123), .Y(n_1221) );
INVx1_ASAP7_75t_L g1222 ( .A(n_1122), .Y(n_1222) );
AND2x2_ASAP7_75t_L g1223 ( .A(n_1024), .B(n_1060), .Y(n_1223) );
INVx1_ASAP7_75t_SL g1224 ( .A(n_1056), .Y(n_1224) );
AND2x4_ASAP7_75t_L g1225 ( .A(n_1117), .B(n_1118), .Y(n_1225) );
AND2x2_ASAP7_75t_L g1226 ( .A(n_1068), .B(n_1076), .Y(n_1226) );
HB1xp67_ASAP7_75t_L g1227 ( .A(n_1023), .Y(n_1227) );
AND2x2_ASAP7_75t_L g1228 ( .A(n_1124), .B(n_1130), .Y(n_1228) );
INVx1_ASAP7_75t_L g1229 ( .A(n_1097), .Y(n_1229) );
BUFx3_ASAP7_75t_L g1230 ( .A(n_1075), .Y(n_1230) );
NAND2xp5_ASAP7_75t_L g1231 ( .A(n_1095), .B(n_1094), .Y(n_1231) );
AND2x2_ASAP7_75t_L g1232 ( .A(n_1049), .B(n_1094), .Y(n_1232) );
INVxp67_ASAP7_75t_SL g1233 ( .A(n_1099), .Y(n_1233) );
INVx1_ASAP7_75t_L g1234 ( .A(n_1135), .Y(n_1234) );
AND2x2_ASAP7_75t_L g1235 ( .A(n_1075), .B(n_1108), .Y(n_1235) );
AND2x2_ASAP7_75t_L g1236 ( .A(n_1108), .B(n_1164), .Y(n_1236) );
OAI211xp5_ASAP7_75t_SL g1237 ( .A1(n_1113), .A2(n_1081), .B(n_1050), .C(n_1059), .Y(n_1237) );
AND2x2_ASAP7_75t_L g1238 ( .A(n_1149), .B(n_1078), .Y(n_1238) );
INVx3_ASAP7_75t_L g1239 ( .A(n_1148), .Y(n_1239) );
HB1xp67_ASAP7_75t_L g1240 ( .A(n_1056), .Y(n_1240) );
INVx3_ASAP7_75t_L g1241 ( .A(n_1133), .Y(n_1241) );
NOR2x1_ASAP7_75t_SL g1242 ( .A(n_1112), .B(n_1137), .Y(n_1242) );
INVx1_ASAP7_75t_L g1243 ( .A(n_1139), .Y(n_1243) );
CKINVDCx20_ASAP7_75t_R g1244 ( .A(n_1026), .Y(n_1244) );
AND2x2_ASAP7_75t_L g1245 ( .A(n_1098), .B(n_1104), .Y(n_1245) );
AND2x2_ASAP7_75t_L g1246 ( .A(n_1098), .B(n_1120), .Y(n_1246) );
AND2x2_ASAP7_75t_L g1247 ( .A(n_1106), .B(n_1057), .Y(n_1247) );
AND2x2_ASAP7_75t_L g1248 ( .A(n_1051), .B(n_1038), .Y(n_1248) );
OR2x2_ASAP7_75t_L g1249 ( .A(n_1128), .B(n_1091), .Y(n_1249) );
NOR2x1_ASAP7_75t_SL g1250 ( .A(n_1029), .B(n_1066), .Y(n_1250) );
HB1xp67_ASAP7_75t_L g1251 ( .A(n_1053), .Y(n_1251) );
HB1xp67_ASAP7_75t_L g1252 ( .A(n_1053), .Y(n_1252) );
INVx2_ASAP7_75t_SL g1253 ( .A(n_1133), .Y(n_1253) );
BUFx2_ASAP7_75t_L g1254 ( .A(n_1140), .Y(n_1254) );
OR2x2_ASAP7_75t_L g1255 ( .A(n_1126), .B(n_1103), .Y(n_1255) );
INVx1_ASAP7_75t_L g1256 ( .A(n_1146), .Y(n_1256) );
NOR2x1p5_ASAP7_75t_L g1257 ( .A(n_1047), .B(n_1110), .Y(n_1257) );
INVx1_ASAP7_75t_L g1258 ( .A(n_1146), .Y(n_1258) );
AND2x2_ASAP7_75t_L g1259 ( .A(n_1039), .B(n_1127), .Y(n_1259) );
BUFx3_ASAP7_75t_L g1260 ( .A(n_1037), .Y(n_1260) );
INVx1_ASAP7_75t_L g1261 ( .A(n_1134), .Y(n_1261) );
HB1xp67_ASAP7_75t_L g1262 ( .A(n_1045), .Y(n_1262) );
AND2x4_ASAP7_75t_L g1263 ( .A(n_1039), .B(n_1028), .Y(n_1263) );
AND2x2_ASAP7_75t_L g1264 ( .A(n_1119), .B(n_1034), .Y(n_1264) );
BUFx2_ASAP7_75t_L g1265 ( .A(n_1025), .Y(n_1265) );
OR2x2_ASAP7_75t_L g1266 ( .A(n_1111), .B(n_1107), .Y(n_1266) );
NAND2xp5_ASAP7_75t_L g1267 ( .A(n_1022), .B(n_1041), .Y(n_1267) );
INVx2_ASAP7_75t_L g1268 ( .A(n_1141), .Y(n_1268) );
INVx2_ASAP7_75t_L g1269 ( .A(n_1116), .Y(n_1269) );
NAND4xp25_ASAP7_75t_L g1270 ( .A(n_1121), .B(n_1129), .C(n_1074), .D(n_1109), .Y(n_1270) );
HB1xp67_ASAP7_75t_L g1271 ( .A(n_1063), .Y(n_1271) );
AND2x2_ASAP7_75t_L g1272 ( .A(n_1034), .B(n_1027), .Y(n_1272) );
INVx2_ASAP7_75t_L g1273 ( .A(n_1131), .Y(n_1273) );
AND2x2_ASAP7_75t_L g1274 ( .A(n_1111), .B(n_1065), .Y(n_1274) );
NAND2xp5_ASAP7_75t_L g1275 ( .A(n_1212), .B(n_1121), .Y(n_1275) );
BUFx2_ASAP7_75t_L g1276 ( .A(n_1206), .Y(n_1276) );
NAND2xp5_ASAP7_75t_L g1277 ( .A(n_1207), .B(n_1129), .Y(n_1277) );
AND2x2_ASAP7_75t_L g1278 ( .A(n_1246), .B(n_1145), .Y(n_1278) );
AOI22xp33_ASAP7_75t_L g1279 ( .A1(n_1179), .A2(n_1109), .B1(n_1092), .B2(n_1064), .Y(n_1279) );
INVx1_ASAP7_75t_L g1280 ( .A(n_1182), .Y(n_1280) );
AND2x2_ASAP7_75t_L g1281 ( .A(n_1246), .B(n_1145), .Y(n_1281) );
INVx1_ASAP7_75t_L g1282 ( .A(n_1182), .Y(n_1282) );
INVx3_ASAP7_75t_L g1283 ( .A(n_1206), .Y(n_1283) );
AND2x4_ASAP7_75t_L g1284 ( .A(n_1206), .B(n_1132), .Y(n_1284) );
INVx1_ASAP7_75t_L g1285 ( .A(n_1184), .Y(n_1285) );
HB1xp67_ASAP7_75t_L g1286 ( .A(n_1173), .Y(n_1286) );
INVx1_ASAP7_75t_L g1287 ( .A(n_1184), .Y(n_1287) );
OAI33xp33_ASAP7_75t_L g1288 ( .A1(n_1256), .A2(n_1147), .A3(n_1079), .B1(n_1070), .B2(n_1125), .B3(n_1077), .Y(n_1288) );
INVx1_ASAP7_75t_L g1289 ( .A(n_1187), .Y(n_1289) );
AND2x2_ASAP7_75t_L g1290 ( .A(n_1256), .B(n_1138), .Y(n_1290) );
INVxp67_ASAP7_75t_L g1291 ( .A(n_1204), .Y(n_1291) );
NAND2xp5_ASAP7_75t_L g1292 ( .A(n_1207), .B(n_1035), .Y(n_1292) );
OAI221xp5_ASAP7_75t_L g1293 ( .A1(n_1183), .A2(n_1035), .B1(n_1069), .B2(n_1102), .C(n_1100), .Y(n_1293) );
AND2x2_ASAP7_75t_L g1294 ( .A(n_1258), .B(n_1030), .Y(n_1294) );
AND2x2_ASAP7_75t_L g1295 ( .A(n_1258), .B(n_1061), .Y(n_1295) );
AND2x2_ASAP7_75t_L g1296 ( .A(n_1245), .B(n_1073), .Y(n_1296) );
INVx1_ASAP7_75t_L g1297 ( .A(n_1187), .Y(n_1297) );
INVx1_ASAP7_75t_L g1298 ( .A(n_1234), .Y(n_1298) );
OAI321xp33_ASAP7_75t_L g1299 ( .A1(n_1219), .A2(n_1237), .A3(n_1188), .B1(n_1270), .B2(n_1265), .C(n_1190), .Y(n_1299) );
AND2x2_ASAP7_75t_L g1300 ( .A(n_1245), .B(n_1238), .Y(n_1300) );
NAND2x1_ASAP7_75t_L g1301 ( .A(n_1206), .B(n_1239), .Y(n_1301) );
NAND2xp5_ASAP7_75t_L g1302 ( .A(n_1210), .B(n_1238), .Y(n_1302) );
NOR2x1_ASAP7_75t_SL g1303 ( .A(n_1222), .B(n_1168), .Y(n_1303) );
OR2x2_ASAP7_75t_L g1304 ( .A(n_1177), .B(n_1194), .Y(n_1304) );
HB1xp67_ASAP7_75t_L g1305 ( .A(n_1170), .Y(n_1305) );
AND2x2_ASAP7_75t_L g1306 ( .A(n_1201), .B(n_1210), .Y(n_1306) );
INVxp67_ASAP7_75t_L g1307 ( .A(n_1204), .Y(n_1307) );
AND2x2_ASAP7_75t_L g1308 ( .A(n_1201), .B(n_1193), .Y(n_1308) );
INVx2_ASAP7_75t_SL g1309 ( .A(n_1168), .Y(n_1309) );
INVx1_ASAP7_75t_L g1310 ( .A(n_1221), .Y(n_1310) );
AND2x2_ASAP7_75t_L g1311 ( .A(n_1193), .B(n_1170), .Y(n_1311) );
CKINVDCx20_ASAP7_75t_R g1312 ( .A(n_1244), .Y(n_1312) );
AOI221xp5_ASAP7_75t_L g1313 ( .A1(n_1215), .A2(n_1213), .B1(n_1174), .B2(n_1247), .C(n_1231), .Y(n_1313) );
AND2x2_ASAP7_75t_L g1314 ( .A(n_1172), .B(n_1197), .Y(n_1314) );
INVx1_ASAP7_75t_L g1315 ( .A(n_1221), .Y(n_1315) );
AND2x2_ASAP7_75t_L g1316 ( .A(n_1172), .B(n_1197), .Y(n_1316) );
HB1xp67_ASAP7_75t_L g1317 ( .A(n_1180), .Y(n_1317) );
AND2x2_ASAP7_75t_L g1318 ( .A(n_1200), .B(n_1181), .Y(n_1318) );
INVx1_ASAP7_75t_L g1319 ( .A(n_1209), .Y(n_1319) );
AND2x2_ASAP7_75t_L g1320 ( .A(n_1200), .B(n_1181), .Y(n_1320) );
AND2x2_ASAP7_75t_L g1321 ( .A(n_1185), .B(n_1186), .Y(n_1321) );
INVx1_ASAP7_75t_L g1322 ( .A(n_1217), .Y(n_1322) );
OAI33xp33_ASAP7_75t_L g1323 ( .A1(n_1189), .A2(n_1191), .A3(n_1192), .B1(n_1249), .B2(n_1267), .B3(n_1220), .Y(n_1323) );
INVx1_ASAP7_75t_L g1324 ( .A(n_1217), .Y(n_1324) );
INVx1_ASAP7_75t_L g1325 ( .A(n_1189), .Y(n_1325) );
AND2x2_ASAP7_75t_L g1326 ( .A(n_1185), .B(n_1186), .Y(n_1326) );
AND2x2_ASAP7_75t_L g1327 ( .A(n_1171), .B(n_1191), .Y(n_1327) );
INVx2_ASAP7_75t_SL g1328 ( .A(n_1168), .Y(n_1328) );
INVx1_ASAP7_75t_L g1329 ( .A(n_1192), .Y(n_1329) );
INVx1_ASAP7_75t_L g1330 ( .A(n_1175), .Y(n_1330) );
INVx2_ASAP7_75t_SL g1331 ( .A(n_1230), .Y(n_1331) );
HB1xp67_ASAP7_75t_L g1332 ( .A(n_1196), .Y(n_1332) );
INVx2_ASAP7_75t_L g1333 ( .A(n_1269), .Y(n_1333) );
AND2x2_ASAP7_75t_L g1334 ( .A(n_1171), .B(n_1175), .Y(n_1334) );
NAND2xp67_ASAP7_75t_L g1335 ( .A(n_1213), .B(n_1248), .Y(n_1335) );
NAND2xp5_ASAP7_75t_L g1336 ( .A(n_1169), .B(n_1265), .Y(n_1336) );
BUFx2_ASAP7_75t_L g1337 ( .A(n_1239), .Y(n_1337) );
INVx1_ASAP7_75t_L g1338 ( .A(n_1176), .Y(n_1338) );
AND2x2_ASAP7_75t_L g1339 ( .A(n_1176), .B(n_1169), .Y(n_1339) );
HB1xp67_ASAP7_75t_L g1340 ( .A(n_1227), .Y(n_1340) );
AND2x2_ASAP7_75t_L g1341 ( .A(n_1243), .B(n_1261), .Y(n_1341) );
OAI21xp5_ASAP7_75t_L g1342 ( .A1(n_1232), .A2(n_1247), .B(n_1262), .Y(n_1342) );
NAND2xp5_ASAP7_75t_L g1343 ( .A(n_1194), .B(n_1202), .Y(n_1343) );
NAND2xp5_ASAP7_75t_L g1344 ( .A(n_1202), .B(n_1208), .Y(n_1344) );
NAND2xp5_ASAP7_75t_L g1345 ( .A(n_1208), .B(n_1220), .Y(n_1345) );
INVxp67_ASAP7_75t_L g1346 ( .A(n_1240), .Y(n_1346) );
AND2x2_ASAP7_75t_L g1347 ( .A(n_1243), .B(n_1261), .Y(n_1347) );
INVx1_ASAP7_75t_L g1348 ( .A(n_1325), .Y(n_1348) );
OR2x2_ASAP7_75t_L g1349 ( .A(n_1304), .B(n_1177), .Y(n_1349) );
OR2x2_ASAP7_75t_L g1350 ( .A(n_1304), .B(n_1249), .Y(n_1350) );
NAND2xp5_ASAP7_75t_L g1351 ( .A(n_1321), .B(n_1232), .Y(n_1351) );
NAND2xp5_ASAP7_75t_L g1352 ( .A(n_1321), .B(n_1211), .Y(n_1352) );
INVx1_ASAP7_75t_L g1353 ( .A(n_1325), .Y(n_1353) );
NAND2xp5_ASAP7_75t_L g1354 ( .A(n_1326), .B(n_1211), .Y(n_1354) );
INVx1_ASAP7_75t_L g1355 ( .A(n_1329), .Y(n_1355) );
INVx2_ASAP7_75t_L g1356 ( .A(n_1333), .Y(n_1356) );
AND2x2_ASAP7_75t_L g1357 ( .A(n_1300), .B(n_1273), .Y(n_1357) );
NAND2xp5_ASAP7_75t_L g1358 ( .A(n_1326), .B(n_1223), .Y(n_1358) );
INVx6_ASAP7_75t_L g1359 ( .A(n_1334), .Y(n_1359) );
INVx1_ASAP7_75t_L g1360 ( .A(n_1329), .Y(n_1360) );
INVx1_ASAP7_75t_SL g1361 ( .A(n_1312), .Y(n_1361) );
INVxp67_ASAP7_75t_L g1362 ( .A(n_1340), .Y(n_1362) );
OR2x2_ASAP7_75t_L g1363 ( .A(n_1302), .B(n_1198), .Y(n_1363) );
NOR2xp33_ASAP7_75t_L g1364 ( .A(n_1346), .B(n_1224), .Y(n_1364) );
INVx1_ASAP7_75t_L g1365 ( .A(n_1286), .Y(n_1365) );
NAND2xp5_ASAP7_75t_L g1366 ( .A(n_1318), .B(n_1223), .Y(n_1366) );
NAND2xp5_ASAP7_75t_L g1367 ( .A(n_1318), .B(n_1272), .Y(n_1367) );
INVx1_ASAP7_75t_L g1368 ( .A(n_1330), .Y(n_1368) );
INVx1_ASAP7_75t_L g1369 ( .A(n_1330), .Y(n_1369) );
NAND2xp5_ASAP7_75t_L g1370 ( .A(n_1320), .B(n_1272), .Y(n_1370) );
NAND2xp5_ASAP7_75t_L g1371 ( .A(n_1320), .B(n_1228), .Y(n_1371) );
HB1xp67_ASAP7_75t_L g1372 ( .A(n_1317), .Y(n_1372) );
NOR3xp33_ASAP7_75t_L g1373 ( .A(n_1299), .B(n_1241), .C(n_1253), .Y(n_1373) );
INVx1_ASAP7_75t_L g1374 ( .A(n_1338), .Y(n_1374) );
OAI21xp33_ASAP7_75t_L g1375 ( .A1(n_1335), .A2(n_1270), .B(n_1248), .Y(n_1375) );
OR2x2_ASAP7_75t_L g1376 ( .A(n_1302), .B(n_1198), .Y(n_1376) );
AND2x2_ASAP7_75t_L g1377 ( .A(n_1300), .B(n_1273), .Y(n_1377) );
NAND2x1p5_ASAP7_75t_L g1378 ( .A(n_1309), .B(n_1260), .Y(n_1378) );
AND2x2_ASAP7_75t_L g1379 ( .A(n_1278), .B(n_1281), .Y(n_1379) );
INVx1_ASAP7_75t_L g1380 ( .A(n_1338), .Y(n_1380) );
AND2x2_ASAP7_75t_L g1381 ( .A(n_1278), .B(n_1203), .Y(n_1381) );
INVx1_ASAP7_75t_L g1382 ( .A(n_1280), .Y(n_1382) );
NAND2xp33_ASAP7_75t_SL g1383 ( .A(n_1301), .B(n_1214), .Y(n_1383) );
NOR2x1_ASAP7_75t_L g1384 ( .A(n_1344), .B(n_1257), .Y(n_1384) );
INVx1_ASAP7_75t_L g1385 ( .A(n_1280), .Y(n_1385) );
NOR2xp67_ASAP7_75t_L g1386 ( .A(n_1309), .B(n_1251), .Y(n_1386) );
INVx1_ASAP7_75t_SL g1387 ( .A(n_1328), .Y(n_1387) );
NOR3xp33_ASAP7_75t_SL g1388 ( .A(n_1299), .B(n_1222), .C(n_1229), .Y(n_1388) );
NAND2x1p5_ASAP7_75t_L g1389 ( .A(n_1328), .B(n_1260), .Y(n_1389) );
NAND2xp5_ASAP7_75t_L g1390 ( .A(n_1305), .B(n_1228), .Y(n_1390) );
NAND2xp5_ASAP7_75t_L g1391 ( .A(n_1313), .B(n_1271), .Y(n_1391) );
OAI211xp5_ASAP7_75t_L g1392 ( .A1(n_1342), .A2(n_1233), .B(n_1252), .C(n_1226), .Y(n_1392) );
AND2x2_ASAP7_75t_L g1393 ( .A(n_1281), .B(n_1203), .Y(n_1393) );
HB1xp67_ASAP7_75t_L g1394 ( .A(n_1332), .Y(n_1394) );
NAND2xp5_ASAP7_75t_L g1395 ( .A(n_1306), .B(n_1218), .Y(n_1395) );
INVx1_ASAP7_75t_L g1396 ( .A(n_1282), .Y(n_1396) );
INVx1_ASAP7_75t_L g1397 ( .A(n_1282), .Y(n_1397) );
AND2x2_ASAP7_75t_L g1398 ( .A(n_1314), .B(n_1316), .Y(n_1398) );
NOR2xp33_ASAP7_75t_L g1399 ( .A(n_1291), .B(n_1235), .Y(n_1399) );
NAND2xp5_ASAP7_75t_L g1400 ( .A(n_1306), .B(n_1218), .Y(n_1400) );
BUFx2_ASAP7_75t_L g1401 ( .A(n_1337), .Y(n_1401) );
INVx1_ASAP7_75t_L g1402 ( .A(n_1285), .Y(n_1402) );
AND2x2_ASAP7_75t_L g1403 ( .A(n_1314), .B(n_1203), .Y(n_1403) );
BUFx2_ASAP7_75t_L g1404 ( .A(n_1337), .Y(n_1404) );
AND2x2_ASAP7_75t_L g1405 ( .A(n_1316), .B(n_1268), .Y(n_1405) );
OR2x2_ASAP7_75t_L g1406 ( .A(n_1336), .B(n_1268), .Y(n_1406) );
INVx1_ASAP7_75t_L g1407 ( .A(n_1285), .Y(n_1407) );
AND2x2_ASAP7_75t_L g1408 ( .A(n_1311), .B(n_1239), .Y(n_1408) );
INVx1_ASAP7_75t_L g1409 ( .A(n_1287), .Y(n_1409) );
NAND2xp5_ASAP7_75t_L g1410 ( .A(n_1379), .B(n_1351), .Y(n_1410) );
NAND2xp33_ASAP7_75t_SL g1411 ( .A(n_1388), .B(n_1276), .Y(n_1411) );
NAND2xp5_ASAP7_75t_L g1412 ( .A(n_1379), .B(n_1341), .Y(n_1412) );
OR2x2_ASAP7_75t_L g1413 ( .A(n_1398), .B(n_1350), .Y(n_1413) );
NOR3xp33_ASAP7_75t_L g1414 ( .A(n_1375), .B(n_1288), .C(n_1307), .Y(n_1414) );
INVx1_ASAP7_75t_L g1415 ( .A(n_1372), .Y(n_1415) );
INVx1_ASAP7_75t_SL g1416 ( .A(n_1361), .Y(n_1416) );
NAND2xp5_ASAP7_75t_L g1417 ( .A(n_1367), .B(n_1341), .Y(n_1417) );
OR2x2_ASAP7_75t_L g1418 ( .A(n_1398), .B(n_1350), .Y(n_1418) );
NAND2xp5_ASAP7_75t_L g1419 ( .A(n_1370), .B(n_1347), .Y(n_1419) );
INVx3_ASAP7_75t_SL g1420 ( .A(n_1387), .Y(n_1420) );
INVx1_ASAP7_75t_L g1421 ( .A(n_1394), .Y(n_1421) );
INVx1_ASAP7_75t_L g1422 ( .A(n_1365), .Y(n_1422) );
OR2x2_ASAP7_75t_L g1423 ( .A(n_1371), .B(n_1336), .Y(n_1423) );
OR2x2_ASAP7_75t_L g1424 ( .A(n_1352), .B(n_1311), .Y(n_1424) );
INVx1_ASAP7_75t_L g1425 ( .A(n_1348), .Y(n_1425) );
OR2x2_ASAP7_75t_L g1426 ( .A(n_1354), .B(n_1308), .Y(n_1426) );
AND2x4_ASAP7_75t_L g1427 ( .A(n_1408), .B(n_1276), .Y(n_1427) );
NAND2xp5_ASAP7_75t_L g1428 ( .A(n_1357), .B(n_1347), .Y(n_1428) );
AND2x2_ASAP7_75t_L g1429 ( .A(n_1408), .B(n_1308), .Y(n_1429) );
INVx1_ASAP7_75t_L g1430 ( .A(n_1353), .Y(n_1430) );
NAND2xp5_ASAP7_75t_L g1431 ( .A(n_1357), .B(n_1342), .Y(n_1431) );
INVx1_ASAP7_75t_L g1432 ( .A(n_1355), .Y(n_1432) );
INVx2_ASAP7_75t_SL g1433 ( .A(n_1359), .Y(n_1433) );
INVx2_ASAP7_75t_L g1434 ( .A(n_1356), .Y(n_1434) );
AND2x2_ASAP7_75t_L g1435 ( .A(n_1403), .B(n_1290), .Y(n_1435) );
NOR2xp33_ASAP7_75t_L g1436 ( .A(n_1391), .B(n_1335), .Y(n_1436) );
OR2x2_ASAP7_75t_L g1437 ( .A(n_1349), .B(n_1292), .Y(n_1437) );
OR2x2_ASAP7_75t_L g1438 ( .A(n_1349), .B(n_1292), .Y(n_1438) );
NAND2xp5_ASAP7_75t_L g1439 ( .A(n_1377), .B(n_1339), .Y(n_1439) );
AND2x2_ASAP7_75t_L g1440 ( .A(n_1403), .B(n_1290), .Y(n_1440) );
AND2x2_ASAP7_75t_L g1441 ( .A(n_1381), .B(n_1283), .Y(n_1441) );
OR2x2_ASAP7_75t_L g1442 ( .A(n_1363), .B(n_1277), .Y(n_1442) );
OAI31xp33_ASAP7_75t_L g1443 ( .A1(n_1392), .A2(n_1257), .A3(n_1293), .B(n_1226), .Y(n_1443) );
AND2x2_ASAP7_75t_L g1444 ( .A(n_1381), .B(n_1283), .Y(n_1444) );
NAND2xp5_ASAP7_75t_L g1445 ( .A(n_1377), .B(n_1339), .Y(n_1445) );
NAND2xp5_ASAP7_75t_L g1446 ( .A(n_1366), .B(n_1343), .Y(n_1446) );
OR2x2_ASAP7_75t_L g1447 ( .A(n_1363), .B(n_1277), .Y(n_1447) );
NAND2xp5_ASAP7_75t_L g1448 ( .A(n_1358), .B(n_1343), .Y(n_1448) );
NAND2xp5_ASAP7_75t_L g1449 ( .A(n_1376), .B(n_1327), .Y(n_1449) );
INVx1_ASAP7_75t_L g1450 ( .A(n_1360), .Y(n_1450) );
INVx2_ASAP7_75t_L g1451 ( .A(n_1356), .Y(n_1451) );
NOR3xp33_ASAP7_75t_L g1452 ( .A(n_1373), .B(n_1323), .C(n_1293), .Y(n_1452) );
INVx1_ASAP7_75t_L g1453 ( .A(n_1382), .Y(n_1453) );
OR2x2_ASAP7_75t_L g1454 ( .A(n_1376), .B(n_1283), .Y(n_1454) );
NAND3xp33_ASAP7_75t_L g1455 ( .A(n_1362), .B(n_1279), .C(n_1294), .Y(n_1455) );
INVx1_ASAP7_75t_L g1456 ( .A(n_1385), .Y(n_1456) );
INVx1_ASAP7_75t_SL g1457 ( .A(n_1359), .Y(n_1457) );
AND2x2_ASAP7_75t_L g1458 ( .A(n_1429), .B(n_1393), .Y(n_1458) );
AOI22xp5_ASAP7_75t_L g1459 ( .A1(n_1414), .A2(n_1384), .B1(n_1386), .B2(n_1399), .Y(n_1459) );
NOR2xp67_ASAP7_75t_L g1460 ( .A(n_1433), .B(n_1364), .Y(n_1460) );
OR2x2_ASAP7_75t_L g1461 ( .A(n_1413), .B(n_1406), .Y(n_1461) );
OAI21xp5_ASAP7_75t_SL g1462 ( .A1(n_1443), .A2(n_1389), .B(n_1378), .Y(n_1462) );
INVx1_ASAP7_75t_L g1463 ( .A(n_1422), .Y(n_1463) );
INVx1_ASAP7_75t_L g1464 ( .A(n_1425), .Y(n_1464) );
AND2x2_ASAP7_75t_L g1465 ( .A(n_1435), .B(n_1393), .Y(n_1465) );
OAI22xp5_ASAP7_75t_L g1466 ( .A1(n_1420), .A2(n_1389), .B1(n_1378), .B2(n_1359), .Y(n_1466) );
INVx1_ASAP7_75t_L g1467 ( .A(n_1430), .Y(n_1467) );
INVxp67_ASAP7_75t_SL g1468 ( .A(n_1434), .Y(n_1468) );
AOI22xp5_ASAP7_75t_L g1469 ( .A1(n_1414), .A2(n_1405), .B1(n_1359), .B2(n_1283), .Y(n_1469) );
NOR2xp33_ASAP7_75t_L g1470 ( .A(n_1436), .B(n_1395), .Y(n_1470) );
OAI221xp5_ASAP7_75t_L g1471 ( .A1(n_1452), .A2(n_1389), .B1(n_1378), .B2(n_1383), .C(n_1406), .Y(n_1471) );
INVx1_ASAP7_75t_L g1472 ( .A(n_1432), .Y(n_1472) );
OAI21xp33_ASAP7_75t_L g1473 ( .A1(n_1452), .A2(n_1405), .B(n_1400), .Y(n_1473) );
NOR2xp33_ASAP7_75t_SL g1474 ( .A(n_1420), .B(n_1214), .Y(n_1474) );
A2O1A1Ixp33_ASAP7_75t_L g1475 ( .A1(n_1411), .A2(n_1383), .B(n_1301), .C(n_1331), .Y(n_1475) );
INVx1_ASAP7_75t_L g1476 ( .A(n_1450), .Y(n_1476) );
NAND2xp5_ASAP7_75t_L g1477 ( .A(n_1435), .B(n_1294), .Y(n_1477) );
INVx1_ASAP7_75t_L g1478 ( .A(n_1453), .Y(n_1478) );
INVx1_ASAP7_75t_L g1479 ( .A(n_1456), .Y(n_1479) );
OAI22xp5_ASAP7_75t_L g1480 ( .A1(n_1418), .A2(n_1390), .B1(n_1331), .B2(n_1404), .Y(n_1480) );
OAI32xp33_ASAP7_75t_L g1481 ( .A1(n_1411), .A2(n_1260), .A3(n_1229), .B1(n_1255), .B2(n_1275), .Y(n_1481) );
OAI311xp33_ASAP7_75t_L g1482 ( .A1(n_1455), .A2(n_1255), .A3(n_1345), .B1(n_1275), .C1(n_1344), .Y(n_1482) );
AND2x2_ASAP7_75t_L g1483 ( .A(n_1440), .B(n_1284), .Y(n_1483) );
AND2x2_ASAP7_75t_L g1484 ( .A(n_1440), .B(n_1401), .Y(n_1484) );
NOR2xp33_ASAP7_75t_L g1485 ( .A(n_1436), .B(n_1396), .Y(n_1485) );
INVx2_ASAP7_75t_SL g1486 ( .A(n_1433), .Y(n_1486) );
AO22x1_ASAP7_75t_L g1487 ( .A1(n_1457), .A2(n_1214), .B1(n_1404), .B2(n_1401), .Y(n_1487) );
AOI22xp33_ASAP7_75t_L g1488 ( .A1(n_1415), .A2(n_1295), .B1(n_1296), .B2(n_1284), .Y(n_1488) );
INVx1_ASAP7_75t_L g1489 ( .A(n_1421), .Y(n_1489) );
NOR2x1_ASAP7_75t_L g1490 ( .A(n_1416), .B(n_1241), .Y(n_1490) );
AOI222xp33_ASAP7_75t_L g1491 ( .A1(n_1473), .A2(n_1431), .B1(n_1419), .B2(n_1417), .C1(n_1448), .C2(n_1446), .Y(n_1491) );
O2A1O1Ixp33_ASAP7_75t_L g1492 ( .A1(n_1482), .A2(n_1345), .B(n_1412), .C(n_1410), .Y(n_1492) );
INVx1_ASAP7_75t_L g1493 ( .A(n_1464), .Y(n_1493) );
INVx1_ASAP7_75t_L g1494 ( .A(n_1467), .Y(n_1494) );
NAND2xp5_ASAP7_75t_L g1495 ( .A(n_1485), .B(n_1428), .Y(n_1495) );
NAND2xp5_ASAP7_75t_L g1496 ( .A(n_1485), .B(n_1437), .Y(n_1496) );
INVx1_ASAP7_75t_L g1497 ( .A(n_1472), .Y(n_1497) );
NOR2xp33_ASAP7_75t_L g1498 ( .A(n_1470), .B(n_1426), .Y(n_1498) );
INVx1_ASAP7_75t_L g1499 ( .A(n_1476), .Y(n_1499) );
OAI21xp5_ASAP7_75t_L g1500 ( .A1(n_1459), .A2(n_1295), .B(n_1427), .Y(n_1500) );
NAND2xp5_ASAP7_75t_L g1501 ( .A(n_1465), .B(n_1438), .Y(n_1501) );
AOI22xp5_ASAP7_75t_L g1502 ( .A1(n_1469), .A2(n_1427), .B1(n_1442), .B2(n_1447), .Y(n_1502) );
NAND2xp5_ASAP7_75t_L g1503 ( .A(n_1465), .B(n_1439), .Y(n_1503) );
INVx1_ASAP7_75t_L g1504 ( .A(n_1478), .Y(n_1504) );
BUFx2_ASAP7_75t_L g1505 ( .A(n_1486), .Y(n_1505) );
OR2x2_ASAP7_75t_L g1506 ( .A(n_1461), .B(n_1423), .Y(n_1506) );
INVx1_ASAP7_75t_L g1507 ( .A(n_1479), .Y(n_1507) );
INVx1_ASAP7_75t_L g1508 ( .A(n_1463), .Y(n_1508) );
XNOR2x2_ASAP7_75t_SL g1509 ( .A(n_1460), .B(n_1424), .Y(n_1509) );
INVx1_ASAP7_75t_L g1510 ( .A(n_1489), .Y(n_1510) );
INVx2_ASAP7_75t_L g1511 ( .A(n_1468), .Y(n_1511) );
NAND2xp33_ASAP7_75t_R g1512 ( .A(n_1474), .B(n_1427), .Y(n_1512) );
A2O1A1Ixp33_ASAP7_75t_L g1513 ( .A1(n_1462), .A2(n_1445), .B(n_1454), .C(n_1230), .Y(n_1513) );
OAI221xp5_ASAP7_75t_L g1514 ( .A1(n_1513), .A2(n_1475), .B1(n_1471), .B2(n_1480), .C(n_1486), .Y(n_1514) );
OAI211xp5_ASAP7_75t_SL g1515 ( .A1(n_1491), .A2(n_1475), .B(n_1488), .C(n_1490), .Y(n_1515) );
OAI322xp33_ASAP7_75t_L g1516 ( .A1(n_1498), .A2(n_1470), .A3(n_1477), .B1(n_1449), .B2(n_1484), .C1(n_1483), .C2(n_1466), .Y(n_1516) );
AOI22xp5_ASAP7_75t_L g1517 ( .A1(n_1512), .A2(n_1483), .B1(n_1488), .B2(n_1458), .Y(n_1517) );
INVx1_ASAP7_75t_L g1518 ( .A(n_1493), .Y(n_1518) );
INVx1_ASAP7_75t_L g1519 ( .A(n_1494), .Y(n_1519) );
BUFx2_ASAP7_75t_L g1520 ( .A(n_1505), .Y(n_1520) );
OAI31xp33_ASAP7_75t_L g1521 ( .A1(n_1513), .A2(n_1458), .A3(n_1481), .B(n_1444), .Y(n_1521) );
AOI21xp33_ASAP7_75t_SL g1522 ( .A1(n_1512), .A2(n_1487), .B(n_1253), .Y(n_1522) );
AOI221xp5_ASAP7_75t_L g1523 ( .A1(n_1492), .A2(n_1444), .B1(n_1441), .B2(n_1402), .C(n_1409), .Y(n_1523) );
OAI22xp5_ASAP7_75t_L g1524 ( .A1(n_1498), .A2(n_1441), .B1(n_1380), .B2(n_1374), .Y(n_1524) );
AOI21xp5_ASAP7_75t_L g1525 ( .A1(n_1509), .A2(n_1500), .B(n_1511), .Y(n_1525) );
AOI21xp5_ASAP7_75t_L g1526 ( .A1(n_1511), .A2(n_1303), .B(n_1250), .Y(n_1526) );
AOI21xp33_ASAP7_75t_L g1527 ( .A1(n_1510), .A2(n_1216), .B(n_1368), .Y(n_1527) );
NAND3x2_ASAP7_75t_L g1528 ( .A(n_1506), .B(n_1284), .C(n_1254), .Y(n_1528) );
INVx1_ASAP7_75t_L g1529 ( .A(n_1497), .Y(n_1529) );
AOI21xp33_ASAP7_75t_L g1530 ( .A1(n_1528), .A2(n_1508), .B(n_1507), .Y(n_1530) );
AOI22xp33_ASAP7_75t_L g1531 ( .A1(n_1515), .A2(n_1496), .B1(n_1502), .B2(n_1495), .Y(n_1531) );
NOR3xp33_ASAP7_75t_L g1532 ( .A(n_1514), .B(n_1241), .C(n_1504), .Y(n_1532) );
AOI211xp5_ASAP7_75t_SL g1533 ( .A1(n_1525), .A2(n_1516), .B(n_1517), .C(n_1523), .Y(n_1533) );
AOI221xp5_ASAP7_75t_L g1534 ( .A1(n_1524), .A2(n_1499), .B1(n_1501), .B2(n_1503), .C(n_1397), .Y(n_1534) );
XOR2xp5_ASAP7_75t_L g1535 ( .A(n_1520), .B(n_1303), .Y(n_1535) );
AOI22xp5_ASAP7_75t_L g1536 ( .A1(n_1524), .A2(n_1284), .B1(n_1296), .B2(n_1407), .Y(n_1536) );
OAI211xp5_ASAP7_75t_SL g1537 ( .A1(n_1521), .A2(n_1266), .B(n_1241), .C(n_1369), .Y(n_1537) );
AOI221xp5_ASAP7_75t_L g1538 ( .A1(n_1522), .A2(n_1297), .B1(n_1289), .B2(n_1310), .C(n_1315), .Y(n_1538) );
AOI22xp33_ASAP7_75t_L g1539 ( .A1(n_1527), .A2(n_1315), .B1(n_1310), .B2(n_1236), .Y(n_1539) );
NOR4xp25_ASAP7_75t_L g1540 ( .A(n_1518), .B(n_1236), .C(n_1216), .D(n_1235), .Y(n_1540) );
O2A1O1Ixp33_ASAP7_75t_L g1541 ( .A1(n_1533), .A2(n_1529), .B(n_1519), .C(n_1526), .Y(n_1541) );
OR2x2_ASAP7_75t_L g1542 ( .A(n_1540), .B(n_1451), .Y(n_1542) );
AND2x2_ASAP7_75t_L g1543 ( .A(n_1532), .B(n_1451), .Y(n_1543) );
INVx1_ASAP7_75t_L g1544 ( .A(n_1535), .Y(n_1544) );
NOR2xp67_ASAP7_75t_L g1545 ( .A(n_1531), .B(n_1434), .Y(n_1545) );
AND2x2_ASAP7_75t_L g1546 ( .A(n_1534), .B(n_1242), .Y(n_1546) );
NAND3xp33_ASAP7_75t_SL g1547 ( .A(n_1538), .B(n_1274), .C(n_1266), .Y(n_1547) );
AOI211xp5_ASAP7_75t_L g1548 ( .A1(n_1537), .A2(n_1230), .B(n_1274), .C(n_1264), .Y(n_1548) );
NOR3xp33_ASAP7_75t_L g1549 ( .A(n_1541), .B(n_1530), .C(n_1536), .Y(n_1549) );
NAND4xp25_ASAP7_75t_L g1550 ( .A(n_1544), .B(n_1539), .C(n_1264), .D(n_1259), .Y(n_1550) );
INVx2_ASAP7_75t_SL g1551 ( .A(n_1546), .Y(n_1551) );
AO22x1_ASAP7_75t_L g1552 ( .A1(n_1543), .A2(n_1199), .B1(n_1195), .B2(n_1225), .Y(n_1552) );
INVx1_ASAP7_75t_L g1553 ( .A(n_1542), .Y(n_1553) );
INVx1_ASAP7_75t_L g1554 ( .A(n_1547), .Y(n_1554) );
NAND4xp25_ASAP7_75t_L g1555 ( .A(n_1549), .B(n_1548), .C(n_1545), .D(n_1259), .Y(n_1555) );
INVx1_ASAP7_75t_L g1556 ( .A(n_1553), .Y(n_1556) );
INVx1_ASAP7_75t_L g1557 ( .A(n_1554), .Y(n_1557) );
NAND2xp5_ASAP7_75t_L g1558 ( .A(n_1551), .B(n_1548), .Y(n_1558) );
INVx3_ASAP7_75t_L g1559 ( .A(n_1556), .Y(n_1559) );
XNOR2xp5_ASAP7_75t_L g1560 ( .A(n_1557), .B(n_1550), .Y(n_1560) );
OAI22xp5_ASAP7_75t_SL g1561 ( .A1(n_1558), .A2(n_1552), .B1(n_1225), .B2(n_1289), .Y(n_1561) );
OAI22xp5_ASAP7_75t_L g1562 ( .A1(n_1555), .A2(n_1297), .B1(n_1287), .B2(n_1324), .Y(n_1562) );
NAND2xp5_ASAP7_75t_L g1563 ( .A(n_1560), .B(n_1327), .Y(n_1563) );
NAND4xp25_ASAP7_75t_SL g1564 ( .A(n_1561), .B(n_1205), .C(n_1319), .D(n_1322), .Y(n_1564) );
HB1xp67_ASAP7_75t_L g1565 ( .A(n_1559), .Y(n_1565) );
AOI21xp5_ASAP7_75t_L g1566 ( .A1(n_1565), .A2(n_1562), .B(n_1250), .Y(n_1566) );
AOI22xp33_ASAP7_75t_L g1567 ( .A1(n_1564), .A2(n_1225), .B1(n_1254), .B2(n_1263), .Y(n_1567) );
AOI22xp33_ASAP7_75t_SL g1568 ( .A1(n_1563), .A2(n_1242), .B1(n_1225), .B2(n_1263), .Y(n_1568) );
NAND2xp5_ASAP7_75t_L g1569 ( .A(n_1566), .B(n_1319), .Y(n_1569) );
NAND3xp33_ASAP7_75t_R g1570 ( .A(n_1568), .B(n_1205), .C(n_1178), .Y(n_1570) );
OAI22xp5_ASAP7_75t_L g1571 ( .A1(n_1567), .A2(n_1322), .B1(n_1324), .B2(n_1298), .Y(n_1571) );
AOI22xp33_ASAP7_75t_L g1572 ( .A1(n_1571), .A2(n_1569), .B1(n_1570), .B2(n_1239), .Y(n_1572) );
endmodule