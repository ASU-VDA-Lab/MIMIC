module real_jpeg_10991_n_18 (n_17, n_8, n_319, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_3, n_320, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_319;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_320;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_1),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_1),
.A2(n_24),
.B1(n_32),
.B2(n_33),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_1),
.A2(n_24),
.B1(n_61),
.B2(n_62),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_1),
.A2(n_24),
.B1(n_46),
.B2(n_47),
.Y(n_254)
);

INVx2_ASAP7_75t_SL g29 ( 
.A(n_2),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_2),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

AOI21xp33_ASAP7_75t_L g172 ( 
.A1(n_2),
.A2(n_11),
.B(n_33),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_3),
.A2(n_61),
.B1(n_62),
.B2(n_142),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_3),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_3),
.A2(n_46),
.B1(n_47),
.B2(n_142),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_3),
.A2(n_32),
.B1(n_33),
.B2(n_142),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_3),
.A2(n_25),
.B1(n_26),
.B2(n_142),
.Y(n_269)
);

BUFx10_ASAP7_75t_L g85 ( 
.A(n_4),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_5),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_6),
.A2(n_25),
.B1(n_26),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_6),
.A2(n_32),
.B1(n_33),
.B2(n_35),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_6),
.A2(n_35),
.B1(n_46),
.B2(n_47),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g220 ( 
.A1(n_6),
.A2(n_35),
.B1(n_61),
.B2(n_62),
.Y(n_220)
);

BUFx6f_ASAP7_75t_SL g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

A2O1A1Ixp33_ASAP7_75t_SL g58 ( 
.A1(n_9),
.A2(n_46),
.B(n_59),
.C(n_60),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_9),
.B(n_46),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_9),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_60)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_9),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_10),
.A2(n_25),
.B1(n_26),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_10),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_10),
.A2(n_54),
.B1(n_61),
.B2(n_62),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_10),
.A2(n_46),
.B1(n_47),
.B2(n_54),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_10),
.A2(n_32),
.B1(n_33),
.B2(n_54),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_11),
.A2(n_46),
.B(n_93),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_11),
.B(n_46),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_11),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_11),
.A2(n_104),
.B1(n_105),
.B2(n_106),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_11),
.A2(n_32),
.B(n_132),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_11),
.B(n_32),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_11),
.B(n_36),
.Y(n_153)
);

OAI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_11),
.A2(n_25),
.B1(n_26),
.B2(n_108),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_12),
.A2(n_46),
.B1(n_47),
.B2(n_95),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_12),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_12),
.A2(n_61),
.B1(n_62),
.B2(n_95),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_12),
.A2(n_32),
.B1(n_33),
.B2(n_95),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_12),
.A2(n_25),
.B1(n_26),
.B2(n_95),
.Y(n_193)
);

BUFx2_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_14),
.A2(n_25),
.B1(n_26),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_14),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_14),
.A2(n_56),
.B1(n_61),
.B2(n_62),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g222 ( 
.A1(n_14),
.A2(n_46),
.B1(n_47),
.B2(n_56),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_14),
.A2(n_32),
.B1(n_33),
.B2(n_56),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_15),
.A2(n_61),
.B1(n_62),
.B2(n_88),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_15),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_15),
.A2(n_46),
.B1(n_47),
.B2(n_88),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_15),
.A2(n_32),
.B1(n_33),
.B2(n_88),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_15),
.A2(n_25),
.B1(n_26),
.B2(n_88),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_16),
.A2(n_61),
.B1(n_62),
.B2(n_124),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_16),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_16),
.A2(n_46),
.B1(n_47),
.B2(n_124),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_16),
.A2(n_32),
.B1(n_33),
.B2(n_124),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_16),
.A2(n_25),
.B1(n_26),
.B2(n_124),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_17),
.A2(n_61),
.B1(n_62),
.B2(n_83),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_17),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_17),
.A2(n_46),
.B1(n_47),
.B2(n_83),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_17),
.A2(n_32),
.B1(n_33),
.B2(n_83),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_17),
.A2(n_25),
.B1(n_26),
.B2(n_83),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_70),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_69),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_37),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_22),
.B(n_37),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_27),
.B1(n_34),
.B2(n_36),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_23),
.A2(n_27),
.B1(n_36),
.B2(n_66),
.Y(n_65)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_25),
.Y(n_26)
);

A2O1A1Ixp33_ASAP7_75t_L g28 ( 
.A1(n_25),
.A2(n_29),
.B(n_30),
.C(n_31),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_29),
.Y(n_30)
);

A2O1A1Ixp33_ASAP7_75t_L g171 ( 
.A1(n_25),
.A2(n_29),
.B(n_108),
.C(n_172),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_27),
.A2(n_36),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_28),
.A2(n_31),
.B1(n_53),
.B2(n_55),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_28),
.A2(n_31),
.B1(n_204),
.B2(n_205),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_28),
.A2(n_31),
.B1(n_205),
.B2(n_230),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_28),
.A2(n_31),
.B1(n_230),
.B2(n_248),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_28),
.A2(n_31),
.B1(n_248),
.B2(n_269),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_28),
.A2(n_31),
.B1(n_53),
.B2(n_269),
.Y(n_291)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

A2O1A1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_32),
.A2(n_43),
.B(n_44),
.C(n_45),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_43),
.Y(n_44)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_65),
.C(n_67),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_38),
.A2(n_39),
.B1(n_312),
.B2(n_314),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_51),
.C(n_57),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_40),
.A2(n_41),
.B1(n_57),
.B2(n_295),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_45),
.B1(n_49),
.B2(n_50),
.Y(n_41)
);

AO21x1_ASAP7_75t_L g68 ( 
.A1(n_42),
.A2(n_45),
.B(n_50),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_42),
.A2(n_45),
.B1(n_131),
.B2(n_133),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_42),
.A2(n_45),
.B1(n_133),
.B2(n_150),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_42),
.A2(n_45),
.B1(n_150),
.B2(n_190),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_42),
.A2(n_45),
.B1(n_190),
.B2(n_201),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_42),
.A2(n_45),
.B1(n_201),
.B2(n_227),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_42),
.A2(n_45),
.B1(n_227),
.B2(n_245),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_42),
.A2(n_45),
.B1(n_245),
.B2(n_262),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_42),
.A2(n_45),
.B1(n_49),
.B2(n_262),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_43),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_43),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_44),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_45),
.B(n_108),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_46),
.B(n_48),
.Y(n_137)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_47),
.A2(n_136),
.B1(n_137),
.B2(n_138),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_51),
.A2(n_52),
.B1(n_302),
.B2(n_303),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_55),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_57),
.A2(n_294),
.B1(n_295),
.B2(n_296),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_57),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_60),
.B(n_64),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_58),
.A2(n_60),
.B1(n_92),
.B2(n_94),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_58),
.A2(n_60),
.B1(n_94),
.B2(n_121),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_58),
.A2(n_60),
.B1(n_121),
.B2(n_129),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_58),
.A2(n_60),
.B1(n_129),
.B2(n_161),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_58),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_58),
.A2(n_60),
.B1(n_212),
.B2(n_213),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_58),
.A2(n_60),
.B1(n_213),
.B2(n_222),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_58),
.A2(n_60),
.B1(n_222),
.B2(n_254),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_58),
.A2(n_60),
.B1(n_64),
.B2(n_254),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_59),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_60),
.B(n_108),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_60),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_61),
.B(n_85),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_61),
.B(n_63),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_61),
.B(n_112),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_62),
.A2(n_97),
.B1(n_98),
.B2(n_99),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_65),
.A2(n_67),
.B1(n_68),
.B2(n_313),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_65),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_71),
.A2(n_310),
.B(n_316),
.Y(n_70)
);

OAI321xp33_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_287),
.A3(n_305),
.B1(n_308),
.B2(n_309),
.C(n_319),
.Y(n_71)
);

AOI321xp33_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_238),
.A3(n_275),
.B1(n_281),
.B2(n_286),
.C(n_320),
.Y(n_72)
);

NOR3xp33_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_195),
.C(n_234),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_165),
.B(n_194),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_76),
.A2(n_144),
.B(n_164),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_126),
.B(n_143),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_78),
.A2(n_115),
.B(n_125),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_101),
.B(n_114),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_89),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_80),
.B(n_89),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_84),
.B1(n_85),
.B2(n_86),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_82),
.A2(n_104),
.B1(n_105),
.B2(n_106),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_84),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_84),
.A2(n_85),
.B1(n_141),
.B2(n_155),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_85),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_87),
.A2(n_105),
.B1(n_106),
.B2(n_123),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_90),
.A2(n_91),
.B1(n_96),
.B2(n_100),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_90),
.B(n_100),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_93),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_96),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_102),
.A2(n_109),
.B(n_113),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_107),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_103),
.B(n_107),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_105),
.A2(n_106),
.B1(n_123),
.B2(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_105),
.A2(n_106),
.B1(n_175),
.B2(n_176),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_105),
.A2(n_106),
.B1(n_176),
.B2(n_210),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_105),
.A2(n_106),
.B1(n_210),
.B2(n_220),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_105),
.A2(n_106),
.B(n_220),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_106),
.B(n_108),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_110),
.B(n_111),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_117),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_116),
.B(n_117),
.Y(n_125)
);

CKINVDCx5p33_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_118),
.B(n_127),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_118),
.B(n_127),
.Y(n_143)
);

FAx1_ASAP7_75t_SL g118 ( 
.A(n_119),
.B(n_120),
.CI(n_122),
.CON(n_118),
.SN(n_118)
);

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_127),
.Y(n_145)
);

FAx1_ASAP7_75t_SL g127 ( 
.A(n_128),
.B(n_130),
.CI(n_134),
.CON(n_127),
.SN(n_127)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_132),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_139),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_135),
.B(n_139),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_145),
.B(n_146),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_147),
.A2(n_148),
.B1(n_157),
.B2(n_158),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_147),
.B(n_160),
.C(n_162),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_151),
.B1(n_152),
.B2(n_156),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_149),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_154),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_153),
.B(n_154),
.C(n_156),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_155),
.Y(n_175)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_159),
.A2(n_160),
.B1(n_162),
.B2(n_163),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_159),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_160),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_161),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_166),
.B(n_167),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_180),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_177),
.B1(n_178),
.B2(n_179),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_169),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_169),
.B(n_179),
.C(n_180),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_171),
.B1(n_173),
.B2(n_174),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_170),
.B(n_174),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_177),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_191),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_183),
.B1(n_188),
.B2(n_189),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_183),
.B(n_188),
.C(n_191),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_185),
.B1(n_186),
.B2(n_187),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_186),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_193),
.Y(n_204)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

AOI21xp33_ASAP7_75t_L g282 ( 
.A1(n_196),
.A2(n_283),
.B(n_284),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_215),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_197),
.B(n_215),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_208),
.C(n_214),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_198),
.B(n_237),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_199),
.B(n_207),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_202),
.B1(n_203),
.B2(n_206),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_200),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_SL g232 ( 
.A(n_202),
.B(n_206),
.C(n_207),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_203),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_208),
.B(n_214),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_211),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_209),
.B(n_211),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_216),
.A2(n_217),
.B1(n_232),
.B2(n_233),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_223),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_218),
.B(n_223),
.C(n_233),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_221),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_219),
.B(n_221),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_224),
.B(n_228),
.C(n_231),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_226),
.A2(n_228),
.B1(n_229),
.B2(n_231),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_226),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_229),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_232),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_235),
.B(n_236),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_257),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_239),
.B(n_257),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_250),
.C(n_256),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_240),
.A2(n_241),
.B1(n_250),
.B2(n_280),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_241),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_242),
.B(n_246),
.C(n_249),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_244),
.A2(n_246),
.B1(n_247),
.B2(n_249),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_244),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_247),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_250),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_253),
.B2(n_255),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_251),
.A2(n_252),
.B1(n_268),
.B2(n_270),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_251),
.A2(n_268),
.B(n_271),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_252),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_252),
.B(n_253),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_253),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_256),
.B(n_279),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_258),
.A2(n_259),
.B1(n_273),
.B2(n_274),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_265),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_260),
.B(n_265),
.C(n_274),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_263),
.B(n_264),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_261),
.B(n_263),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_264),
.B(n_289),
.C(n_297),
.Y(n_288)
);

FAx1_ASAP7_75t_SL g307 ( 
.A(n_264),
.B(n_289),
.CI(n_297),
.CON(n_307),
.SN(n_307)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_267),
.B1(n_271),
.B2(n_272),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_267),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_268),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_272),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_273),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_276),
.A2(n_282),
.B(n_285),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_277),
.B(n_278),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_298),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_288),
.B(n_298),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_291),
.B1(n_292),
.B2(n_293),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_290),
.A2(n_291),
.B1(n_300),
.B2(n_301),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_291),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_291),
.B(n_295),
.C(n_296),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_291),
.B(n_300),
.C(n_304),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_293),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_294),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_304),
.Y(n_298)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_303),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_306),
.B(n_307),
.Y(n_308)
);

BUFx24_ASAP7_75t_SL g318 ( 
.A(n_307),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_315),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_311),
.B(n_315),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_312),
.Y(n_314)
);


endmodule