module fake_netlist_6_670_n_1730 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1730);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1730;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g156 ( 
.A(n_76),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_92),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_145),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_134),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_84),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_91),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_122),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_117),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_143),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_72),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_7),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_138),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_60),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_125),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_14),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_105),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_70),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_112),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_139),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_10),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_114),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_78),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_126),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_102),
.Y(n_179)
);

BUFx2_ASAP7_75t_SL g180 ( 
.A(n_26),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_93),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_121),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_77),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_37),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_50),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_7),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_32),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_57),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_144),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_39),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_32),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_151),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_30),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_115),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_48),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_1),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_47),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_141),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_111),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_90),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_40),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_31),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_43),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_95),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_113),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_47),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_51),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_124),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_128),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_154),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_20),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_106),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_118),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_132),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_33),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_119),
.Y(n_216)
);

INVx2_ASAP7_75t_SL g217 ( 
.A(n_83),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g218 ( 
.A(n_13),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_27),
.Y(n_219)
);

INVx2_ASAP7_75t_SL g220 ( 
.A(n_2),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_136),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_56),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_0),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_39),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_94),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_96),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_142),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_42),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_38),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_103),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_88),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_23),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_99),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_68),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_120),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_109),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_12),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_153),
.Y(n_238)
);

BUFx2_ASAP7_75t_L g239 ( 
.A(n_123),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_69),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_13),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_25),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_58),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_133),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_97),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_87),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_35),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_0),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_40),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_82),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_10),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_9),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_41),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_110),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_21),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_23),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_9),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_50),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_131),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_48),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_52),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_127),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_41),
.Y(n_263)
);

BUFx2_ASAP7_75t_L g264 ( 
.A(n_18),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_14),
.Y(n_265)
);

BUFx8_ASAP7_75t_SL g266 ( 
.A(n_26),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_89),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_55),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_63),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_1),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_66),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_116),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_135),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_85),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_19),
.Y(n_275)
);

BUFx10_ASAP7_75t_L g276 ( 
.A(n_64),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_107),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_18),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_30),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_34),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_29),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_31),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_42),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_8),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_73),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_33),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_152),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_15),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_130),
.Y(n_289)
);

BUFx5_ASAP7_75t_L g290 ( 
.A(n_74),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_19),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_49),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_3),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_29),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_43),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_101),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_6),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_155),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_35),
.Y(n_299)
);

INVx2_ASAP7_75t_SL g300 ( 
.A(n_2),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_59),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_146),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_53),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_21),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_16),
.Y(n_305)
);

BUFx8_ASAP7_75t_SL g306 ( 
.A(n_28),
.Y(n_306)
);

CKINVDCx14_ASAP7_75t_R g307 ( 
.A(n_148),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_86),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_38),
.Y(n_309)
);

INVx1_ASAP7_75t_SL g310 ( 
.A(n_37),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_264),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_160),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_266),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_282),
.Y(n_314)
);

INVxp67_ASAP7_75t_SL g315 ( 
.A(n_243),
.Y(n_315)
);

BUFx10_ASAP7_75t_L g316 ( 
.A(n_287),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_164),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_282),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_282),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_282),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_282),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_165),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_292),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_292),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_204),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_306),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g327 ( 
.A(n_170),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_214),
.Y(n_328)
);

CKINVDCx14_ASAP7_75t_R g329 ( 
.A(n_187),
.Y(n_329)
);

HB1xp67_ASAP7_75t_L g330 ( 
.A(n_170),
.Y(n_330)
);

BUFx2_ASAP7_75t_L g331 ( 
.A(n_190),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_189),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_234),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_292),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_268),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_272),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_194),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_274),
.Y(n_338)
);

INVxp33_ASAP7_75t_L g339 ( 
.A(n_166),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_292),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_285),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_198),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_292),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_180),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_288),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_277),
.Y(n_346)
);

CKINVDCx14_ASAP7_75t_R g347 ( 
.A(n_307),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_288),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_190),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_199),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_200),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_218),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g353 ( 
.A(n_184),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_218),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_208),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_175),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_209),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_210),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_185),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_193),
.Y(n_360)
);

INVxp67_ASAP7_75t_SL g361 ( 
.A(n_239),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_196),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_213),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_221),
.Y(n_364)
);

INVxp33_ASAP7_75t_SL g365 ( 
.A(n_184),
.Y(n_365)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_186),
.Y(n_366)
);

BUFx3_ASAP7_75t_L g367 ( 
.A(n_171),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_222),
.Y(n_368)
);

CKINVDCx14_ASAP7_75t_R g369 ( 
.A(n_276),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_201),
.Y(n_370)
);

INVxp33_ASAP7_75t_SL g371 ( 
.A(n_186),
.Y(n_371)
);

BUFx2_ASAP7_75t_L g372 ( 
.A(n_252),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_225),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_202),
.Y(n_374)
);

INVxp67_ASAP7_75t_SL g375 ( 
.A(n_171),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_206),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_207),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_215),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_219),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_231),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_229),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_236),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_311),
.A2(n_263),
.B1(n_270),
.B2(n_253),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_323),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_375),
.B(n_240),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_315),
.A2(n_256),
.B1(n_309),
.B2(n_305),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_323),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_314),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_314),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_332),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_318),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_318),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_367),
.B(n_220),
.Y(n_393)
);

BUFx8_ASAP7_75t_L g394 ( 
.A(n_372),
.Y(n_394)
);

AND2x4_ASAP7_75t_L g395 ( 
.A(n_319),
.B(n_240),
.Y(n_395)
);

NAND2x1p5_ASAP7_75t_L g396 ( 
.A(n_319),
.B(n_217),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_320),
.B(n_217),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_316),
.B(n_276),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_320),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_321),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_312),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_321),
.Y(n_402)
);

INVxp67_ASAP7_75t_SL g403 ( 
.A(n_379),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_324),
.Y(n_404)
);

OR2x2_ASAP7_75t_L g405 ( 
.A(n_372),
.B(n_220),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_R g406 ( 
.A(n_347),
.B(n_244),
.Y(n_406)
);

OA21x2_ASAP7_75t_L g407 ( 
.A1(n_324),
.A2(n_241),
.B(n_237),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_334),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_337),
.Y(n_409)
);

AND3x2_ASAP7_75t_L g410 ( 
.A(n_361),
.B(n_269),
.C(n_178),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_334),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_340),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_340),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_342),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_343),
.Y(n_415)
);

BUFx3_ASAP7_75t_L g416 ( 
.A(n_367),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_343),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_345),
.Y(n_418)
);

BUFx3_ASAP7_75t_L g419 ( 
.A(n_367),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_356),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_345),
.Y(n_421)
);

INVx3_ASAP7_75t_L g422 ( 
.A(n_348),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_356),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_359),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_346),
.A2(n_281),
.B1(n_309),
.B2(n_305),
.Y(n_425)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_348),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_359),
.Y(n_427)
);

BUFx8_ASAP7_75t_L g428 ( 
.A(n_331),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_349),
.B(n_300),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_360),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_360),
.Y(n_431)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_362),
.Y(n_432)
);

BUFx3_ASAP7_75t_L g433 ( 
.A(n_349),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_362),
.Y(n_434)
);

AND2x6_ASAP7_75t_L g435 ( 
.A(n_352),
.B(n_233),
.Y(n_435)
);

AND2x4_ASAP7_75t_L g436 ( 
.A(n_352),
.B(n_178),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_370),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_350),
.Y(n_438)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_370),
.Y(n_439)
);

HB1xp67_ASAP7_75t_L g440 ( 
.A(n_327),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_374),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_317),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_374),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_376),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_376),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_377),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_339),
.A2(n_310),
.B1(n_255),
.B2(n_279),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_431),
.Y(n_448)
);

INVxp67_ASAP7_75t_SL g449 ( 
.A(n_416),
.Y(n_449)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_384),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_385),
.B(n_393),
.Y(n_451)
);

INVx2_ASAP7_75t_SL g452 ( 
.A(n_416),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_391),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_416),
.B(n_351),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_390),
.B(n_357),
.Y(n_455)
);

INVx2_ASAP7_75t_SL g456 ( 
.A(n_419),
.Y(n_456)
);

INVx3_ASAP7_75t_L g457 ( 
.A(n_384),
.Y(n_457)
);

AND2x4_ASAP7_75t_L g458 ( 
.A(n_419),
.B(n_269),
.Y(n_458)
);

BUFx3_ASAP7_75t_L g459 ( 
.A(n_419),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_391),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_387),
.Y(n_461)
);

NAND3xp33_ASAP7_75t_L g462 ( 
.A(n_407),
.B(n_344),
.C(n_262),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_387),
.Y(n_463)
);

BUFx4f_ASAP7_75t_L g464 ( 
.A(n_407),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_392),
.Y(n_465)
);

AOI22xp33_ASAP7_75t_L g466 ( 
.A1(n_385),
.A2(n_407),
.B1(n_436),
.B2(n_393),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_409),
.Y(n_467)
);

CKINVDCx6p67_ASAP7_75t_R g468 ( 
.A(n_401),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_388),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_414),
.B(n_358),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_385),
.B(n_368),
.Y(n_471)
);

INVxp33_ASAP7_75t_L g472 ( 
.A(n_440),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_388),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_438),
.B(n_373),
.Y(n_474)
);

OR2x6_ASAP7_75t_L g475 ( 
.A(n_396),
.B(n_302),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_398),
.B(n_380),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_388),
.Y(n_477)
);

INVx2_ASAP7_75t_SL g478 ( 
.A(n_405),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_405),
.B(n_365),
.Y(n_479)
);

INVx4_ASAP7_75t_L g480 ( 
.A(n_389),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_399),
.Y(n_481)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_384),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_406),
.B(n_371),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_403),
.B(n_316),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_392),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_399),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_399),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_400),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_408),
.Y(n_489)
);

NAND3xp33_ASAP7_75t_L g490 ( 
.A(n_407),
.B(n_302),
.C(n_377),
.Y(n_490)
);

INVx3_ASAP7_75t_L g491 ( 
.A(n_384),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_431),
.Y(n_492)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_384),
.Y(n_493)
);

BUFx10_ASAP7_75t_L g494 ( 
.A(n_440),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_408),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_433),
.B(n_354),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_408),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_389),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_400),
.Y(n_499)
);

INVx4_ASAP7_75t_L g500 ( 
.A(n_389),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_442),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_389),
.Y(n_502)
);

BUFx4f_ASAP7_75t_L g503 ( 
.A(n_407),
.Y(n_503)
);

NAND2xp33_ASAP7_75t_L g504 ( 
.A(n_396),
.B(n_233),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_402),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_431),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_428),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_R g508 ( 
.A(n_428),
.B(n_355),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_403),
.B(n_316),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_433),
.B(n_329),
.Y(n_510)
);

OR2x2_ASAP7_75t_L g511 ( 
.A(n_425),
.B(n_330),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_425),
.B(n_316),
.Y(n_512)
);

AND2x6_ASAP7_75t_L g513 ( 
.A(n_395),
.B(n_233),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_386),
.B(n_382),
.Y(n_514)
);

BUFx6f_ASAP7_75t_L g515 ( 
.A(n_431),
.Y(n_515)
);

BUFx3_ASAP7_75t_L g516 ( 
.A(n_395),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_402),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_411),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_386),
.B(n_363),
.Y(n_519)
);

OR2x2_ASAP7_75t_L g520 ( 
.A(n_447),
.B(n_353),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_428),
.B(n_364),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_411),
.Y(n_522)
);

INVxp33_ASAP7_75t_L g523 ( 
.A(n_383),
.Y(n_523)
);

INVx5_ASAP7_75t_L g524 ( 
.A(n_435),
.Y(n_524)
);

INVx1_ASAP7_75t_SL g525 ( 
.A(n_429),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_412),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_415),
.Y(n_527)
);

BUFx3_ASAP7_75t_L g528 ( 
.A(n_395),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_415),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_431),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_417),
.Y(n_531)
);

NAND3xp33_ASAP7_75t_L g532 ( 
.A(n_436),
.B(n_378),
.C(n_381),
.Y(n_532)
);

INVx2_ASAP7_75t_SL g533 ( 
.A(n_410),
.Y(n_533)
);

OR2x2_ASAP7_75t_L g534 ( 
.A(n_447),
.B(n_366),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_417),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_432),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_432),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_384),
.Y(n_538)
);

INVx4_ASAP7_75t_L g539 ( 
.A(n_389),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_395),
.B(n_369),
.Y(n_540)
);

AOI22xp33_ASAP7_75t_L g541 ( 
.A1(n_436),
.A2(n_300),
.B1(n_295),
.B2(n_248),
.Y(n_541)
);

AND3x2_ASAP7_75t_L g542 ( 
.A(n_429),
.B(n_331),
.C(n_157),
.Y(n_542)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_384),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_432),
.Y(n_544)
);

INVx2_ASAP7_75t_SL g545 ( 
.A(n_410),
.Y(n_545)
);

CKINVDCx6p67_ASAP7_75t_R g546 ( 
.A(n_433),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_389),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_422),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_422),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_432),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_431),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_422),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_439),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_396),
.B(n_245),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_439),
.Y(n_555)
);

INVx5_ASAP7_75t_L g556 ( 
.A(n_435),
.Y(n_556)
);

AND2x2_ASAP7_75t_SL g557 ( 
.A(n_436),
.B(n_233),
.Y(n_557)
);

INVx4_ASAP7_75t_L g558 ( 
.A(n_389),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_396),
.B(n_246),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_404),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_404),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_404),
.Y(n_562)
);

HB1xp67_ASAP7_75t_L g563 ( 
.A(n_428),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_439),
.B(n_354),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_422),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_439),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_431),
.Y(n_567)
);

AOI22xp33_ASAP7_75t_L g568 ( 
.A1(n_420),
.A2(n_437),
.B1(n_445),
.B2(n_444),
.Y(n_568)
);

AOI22xp33_ASAP7_75t_SL g569 ( 
.A1(n_394),
.A2(n_322),
.B1(n_341),
.B2(n_338),
.Y(n_569)
);

INVx1_ASAP7_75t_SL g570 ( 
.A(n_383),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_426),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_404),
.Y(n_572)
);

BUFx3_ASAP7_75t_L g573 ( 
.A(n_404),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_420),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_423),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_423),
.B(n_378),
.Y(n_576)
);

INVx4_ASAP7_75t_L g577 ( 
.A(n_404),
.Y(n_577)
);

INVx3_ASAP7_75t_L g578 ( 
.A(n_404),
.Y(n_578)
);

CKINVDCx6p67_ASAP7_75t_R g579 ( 
.A(n_394),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_424),
.B(n_313),
.Y(n_580)
);

INVx2_ASAP7_75t_SL g581 ( 
.A(n_397),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_413),
.B(n_250),
.Y(n_582)
);

NAND2xp33_ASAP7_75t_SL g583 ( 
.A(n_397),
.B(n_252),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_413),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_424),
.B(n_326),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_413),
.B(n_296),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_426),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_413),
.B(n_298),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_427),
.B(n_325),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_394),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_394),
.B(n_276),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_426),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_427),
.Y(n_593)
);

NAND3xp33_ASAP7_75t_L g594 ( 
.A(n_479),
.B(n_195),
.C(n_191),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_581),
.B(n_426),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_581),
.B(n_413),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_451),
.B(n_413),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_451),
.B(n_413),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_466),
.B(n_156),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_525),
.B(n_328),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_517),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_557),
.B(n_176),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_517),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_516),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_557),
.B(n_179),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_471),
.B(n_158),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_518),
.Y(n_607)
);

NOR2xp67_ASAP7_75t_L g608 ( 
.A(n_476),
.B(n_430),
.Y(n_608)
);

INVx2_ASAP7_75t_SL g609 ( 
.A(n_494),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_557),
.B(n_181),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_574),
.B(n_183),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_478),
.B(n_158),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_574),
.B(n_575),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_516),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_575),
.B(n_192),
.Y(n_615)
);

NAND2xp33_ASAP7_75t_L g616 ( 
.A(n_554),
.B(n_559),
.Y(n_616)
);

NAND2xp33_ASAP7_75t_L g617 ( 
.A(n_452),
.B(n_456),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_516),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_464),
.B(n_233),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_528),
.Y(n_620)
);

OAI22xp33_ASAP7_75t_L g621 ( 
.A1(n_523),
.A2(n_284),
.B1(n_249),
.B2(n_251),
.Y(n_621)
);

AOI22xp5_ASAP7_75t_L g622 ( 
.A1(n_589),
.A2(n_333),
.B1(n_336),
.B2(n_335),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_518),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_593),
.B(n_205),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_593),
.B(n_452),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_527),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_456),
.B(n_212),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_464),
.B(n_235),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_527),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_564),
.B(n_226),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_478),
.B(n_159),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_564),
.B(n_227),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_464),
.B(n_235),
.Y(n_633)
);

NOR2xp67_ASAP7_75t_L g634 ( 
.A(n_467),
.B(n_446),
.Y(n_634)
);

INVx2_ASAP7_75t_SL g635 ( 
.A(n_494),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_529),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_458),
.B(n_230),
.Y(n_637)
);

AND2x2_ASAP7_75t_SL g638 ( 
.A(n_503),
.B(n_235),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_484),
.B(n_159),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_509),
.B(n_161),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_458),
.B(n_449),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_458),
.B(n_238),
.Y(n_642)
);

INVx3_ASAP7_75t_L g643 ( 
.A(n_528),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_533),
.B(n_161),
.Y(n_644)
);

INVx2_ASAP7_75t_SL g645 ( 
.A(n_494),
.Y(n_645)
);

INVx2_ASAP7_75t_SL g646 ( 
.A(n_494),
.Y(n_646)
);

INVx2_ASAP7_75t_SL g647 ( 
.A(n_496),
.Y(n_647)
);

INVx2_ASAP7_75t_SL g648 ( 
.A(n_496),
.Y(n_648)
);

OAI221xp5_ASAP7_75t_L g649 ( 
.A1(n_541),
.A2(n_280),
.B1(n_247),
.B2(n_258),
.C(n_260),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_576),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_458),
.B(n_259),
.Y(n_651)
);

AOI22xp5_ASAP7_75t_L g652 ( 
.A1(n_533),
.A2(n_174),
.B1(n_308),
.B2(n_303),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_453),
.B(n_267),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_453),
.B(n_271),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_460),
.B(n_273),
.Y(n_655)
);

OR2x2_ASAP7_75t_L g656 ( 
.A(n_511),
.B(n_446),
.Y(n_656)
);

HB1xp67_ASAP7_75t_L g657 ( 
.A(n_545),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_472),
.B(n_430),
.Y(n_658)
);

BUFx6f_ASAP7_75t_L g659 ( 
.A(n_459),
.Y(n_659)
);

BUFx10_ASAP7_75t_L g660 ( 
.A(n_580),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_545),
.B(n_162),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_576),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_460),
.Y(n_663)
);

AOI22xp33_ASAP7_75t_SL g664 ( 
.A1(n_570),
.A2(n_265),
.B1(n_278),
.B2(n_279),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_465),
.B(n_289),
.Y(n_665)
);

NOR2x1p5_ASAP7_75t_L g666 ( 
.A(n_579),
.B(n_590),
.Y(n_666)
);

AOI22xp5_ASAP7_75t_L g667 ( 
.A1(n_462),
.A2(n_168),
.B1(n_308),
.B2(n_303),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_465),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_485),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_585),
.B(n_445),
.Y(n_670)
);

INVxp67_ASAP7_75t_L g671 ( 
.A(n_583),
.Y(n_671)
);

AO22x2_ASAP7_75t_L g672 ( 
.A1(n_511),
.A2(n_283),
.B1(n_299),
.B2(n_301),
.Y(n_672)
);

INVx4_ASAP7_75t_L g673 ( 
.A(n_459),
.Y(n_673)
);

AOI22xp33_ASAP7_75t_L g674 ( 
.A1(n_490),
.A2(n_235),
.B1(n_290),
.B2(n_441),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_503),
.B(n_235),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_485),
.B(n_418),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_454),
.B(n_162),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_488),
.B(n_418),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_488),
.B(n_418),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_499),
.B(n_421),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_499),
.B(n_421),
.Y(n_681)
);

AOI222xp33_ASAP7_75t_L g682 ( 
.A1(n_514),
.A2(n_291),
.B1(n_257),
.B2(n_265),
.C1(n_278),
.C2(n_281),
.Y(n_682)
);

NOR2xp67_ASAP7_75t_L g683 ( 
.A(n_462),
.B(n_444),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_505),
.B(n_421),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_505),
.B(n_434),
.Y(n_685)
);

O2A1O1Ixp33_ASAP7_75t_L g686 ( 
.A1(n_490),
.A2(n_443),
.B(n_441),
.C(n_437),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_522),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_522),
.Y(n_688)
);

INVx3_ASAP7_75t_L g689 ( 
.A(n_459),
.Y(n_689)
);

AND2x6_ASAP7_75t_L g690 ( 
.A(n_536),
.B(n_434),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_529),
.Y(n_691)
);

BUFx6f_ASAP7_75t_L g692 ( 
.A(n_448),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_461),
.Y(n_693)
);

INVxp67_ASAP7_75t_L g694 ( 
.A(n_519),
.Y(n_694)
);

INVx2_ASAP7_75t_SL g695 ( 
.A(n_542),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_531),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_526),
.Y(n_697)
);

BUFx6f_ASAP7_75t_SL g698 ( 
.A(n_579),
.Y(n_698)
);

INVx2_ASAP7_75t_SL g699 ( 
.A(n_520),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_526),
.B(n_443),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_535),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_501),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_503),
.B(n_290),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_535),
.B(n_435),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_536),
.B(n_435),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_537),
.B(n_435),
.Y(n_706)
);

AOI22xp33_ASAP7_75t_L g707 ( 
.A1(n_475),
.A2(n_290),
.B1(n_304),
.B2(n_257),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_537),
.Y(n_708)
);

INVx2_ASAP7_75t_SL g709 ( 
.A(n_520),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_544),
.B(n_435),
.Y(n_710)
);

NAND3xp33_ASAP7_75t_L g711 ( 
.A(n_512),
.B(n_294),
.C(n_197),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_455),
.B(n_163),
.Y(n_712)
);

INVx2_ASAP7_75t_SL g713 ( 
.A(n_534),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_531),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_470),
.B(n_163),
.Y(n_715)
);

AOI22xp5_ASAP7_75t_L g716 ( 
.A1(n_546),
.A2(n_167),
.B1(n_168),
.B2(n_169),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_544),
.B(n_435),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_550),
.B(n_290),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_550),
.B(n_290),
.Y(n_719)
);

NOR3xp33_ASAP7_75t_L g720 ( 
.A(n_591),
.B(n_381),
.C(n_203),
.Y(n_720)
);

AOI22xp5_ASAP7_75t_L g721 ( 
.A1(n_546),
.A2(n_540),
.B1(n_510),
.B2(n_474),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_553),
.B(n_290),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_553),
.Y(n_723)
);

NAND2xp33_ASAP7_75t_L g724 ( 
.A(n_513),
.B(n_290),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_555),
.B(n_435),
.Y(n_725)
);

AOI22xp5_ASAP7_75t_L g726 ( 
.A1(n_475),
.A2(n_167),
.B1(n_169),
.B2(n_172),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_555),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_566),
.B(n_435),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_548),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_566),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_548),
.B(n_172),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_549),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_549),
.B(n_290),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_552),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_552),
.B(n_173),
.Y(n_735)
);

INVxp33_ASAP7_75t_L g736 ( 
.A(n_534),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_565),
.B(n_173),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_565),
.B(n_174),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_571),
.B(n_177),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_571),
.B(n_177),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_587),
.B(n_182),
.Y(n_741)
);

OR2x2_ASAP7_75t_L g742 ( 
.A(n_483),
.B(n_304),
.Y(n_742)
);

INVx3_ASAP7_75t_L g743 ( 
.A(n_587),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_592),
.B(n_182),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_461),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_592),
.B(n_188),
.Y(n_746)
);

OAI221xp5_ASAP7_75t_L g747 ( 
.A1(n_568),
.A2(n_297),
.B1(n_293),
.B2(n_211),
.C(n_223),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_524),
.B(n_188),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_463),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_524),
.B(n_216),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_524),
.B(n_216),
.Y(n_751)
);

INVx2_ASAP7_75t_SL g752 ( 
.A(n_508),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_582),
.B(n_254),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_586),
.B(n_254),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_524),
.B(n_261),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_588),
.B(n_567),
.Y(n_756)
);

OR2x6_ASAP7_75t_L g757 ( 
.A(n_563),
.B(n_3),
.Y(n_757)
);

NOR2x1p5_ASAP7_75t_L g758 ( 
.A(n_468),
.B(n_291),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_463),
.Y(n_759)
);

BUFx3_ASAP7_75t_L g760 ( 
.A(n_702),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_736),
.B(n_521),
.Y(n_761)
);

AND2x6_ASAP7_75t_L g762 ( 
.A(n_643),
.B(n_567),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_658),
.B(n_569),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_698),
.Y(n_764)
);

INVx3_ASAP7_75t_L g765 ( 
.A(n_659),
.Y(n_765)
);

AOI22xp5_ASAP7_75t_L g766 ( 
.A1(n_694),
.A2(n_475),
.B1(n_504),
.B2(n_513),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_708),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_670),
.B(n_475),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_723),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_638),
.B(n_524),
.Y(n_770)
);

AOI22xp33_ASAP7_75t_SL g771 ( 
.A1(n_638),
.A2(n_507),
.B1(n_286),
.B2(n_224),
.Y(n_771)
);

AOI22xp5_ASAP7_75t_L g772 ( 
.A1(n_608),
.A2(n_606),
.B1(n_677),
.B2(n_599),
.Y(n_772)
);

BUFx8_ASAP7_75t_L g773 ( 
.A(n_698),
.Y(n_773)
);

AOI22xp5_ASAP7_75t_L g774 ( 
.A1(n_606),
.A2(n_475),
.B1(n_513),
.B2(n_532),
.Y(n_774)
);

AOI22xp33_ASAP7_75t_L g775 ( 
.A1(n_707),
.A2(n_532),
.B1(n_513),
.B2(n_469),
.Y(n_775)
);

HB1xp67_ASAP7_75t_L g776 ( 
.A(n_657),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_729),
.Y(n_777)
);

NOR2x1p5_ASAP7_75t_L g778 ( 
.A(n_742),
.B(n_468),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_677),
.B(n_573),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_729),
.Y(n_780)
);

INVx1_ASAP7_75t_SL g781 ( 
.A(n_600),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_595),
.B(n_573),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_727),
.Y(n_783)
);

NAND3xp33_ASAP7_75t_SL g784 ( 
.A(n_682),
.B(n_286),
.C(n_228),
.Y(n_784)
);

AOI22xp33_ASAP7_75t_SL g785 ( 
.A1(n_672),
.A2(n_242),
.B1(n_275),
.B2(n_232),
.Y(n_785)
);

OR2x2_ASAP7_75t_L g786 ( 
.A(n_699),
.B(n_261),
.Y(n_786)
);

AND2x4_ASAP7_75t_L g787 ( 
.A(n_647),
.B(n_573),
.Y(n_787)
);

NOR2x2_ASAP7_75t_L g788 ( 
.A(n_757),
.B(n_538),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_663),
.B(n_450),
.Y(n_789)
);

A2O1A1Ixp33_ASAP7_75t_L g790 ( 
.A1(n_683),
.A2(n_538),
.B(n_502),
.C(n_498),
.Y(n_790)
);

AOI22xp33_ASAP7_75t_SL g791 ( 
.A1(n_672),
.A2(n_513),
.B1(n_5),
.B2(n_6),
.Y(n_791)
);

AOI22xp33_ASAP7_75t_L g792 ( 
.A1(n_707),
.A2(n_513),
.B1(n_481),
.B2(n_469),
.Y(n_792)
);

BUFx2_ASAP7_75t_L g793 ( 
.A(n_657),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_668),
.B(n_450),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_730),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_732),
.Y(n_796)
);

AND2x2_ASAP7_75t_L g797 ( 
.A(n_650),
.B(n_473),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_669),
.B(n_450),
.Y(n_798)
);

AOI21x1_ASAP7_75t_L g799 ( 
.A1(n_619),
.A2(n_502),
.B(n_498),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_687),
.B(n_450),
.Y(n_800)
);

BUFx3_ASAP7_75t_L g801 ( 
.A(n_752),
.Y(n_801)
);

INVx4_ASAP7_75t_SL g802 ( 
.A(n_690),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_643),
.B(n_524),
.Y(n_803)
);

AOI22xp5_ASAP7_75t_L g804 ( 
.A1(n_604),
.A2(n_513),
.B1(n_578),
.B2(n_547),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_709),
.B(n_713),
.Y(n_805)
);

OR2x2_ASAP7_75t_SL g806 ( 
.A(n_711),
.B(n_4),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_601),
.Y(n_807)
);

AOI22xp33_ASAP7_75t_L g808 ( 
.A1(n_662),
.A2(n_486),
.B1(n_481),
.B2(n_477),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_601),
.Y(n_809)
);

HB1xp67_ASAP7_75t_L g810 ( 
.A(n_648),
.Y(n_810)
);

OAI22xp5_ASAP7_75t_L g811 ( 
.A1(n_625),
.A2(n_502),
.B1(n_498),
.B2(n_560),
.Y(n_811)
);

AOI22xp33_ASAP7_75t_L g812 ( 
.A1(n_619),
.A2(n_486),
.B1(n_477),
.B2(n_473),
.Y(n_812)
);

BUFx6f_ASAP7_75t_L g813 ( 
.A(n_659),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_732),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_688),
.B(n_457),
.Y(n_815)
);

AND2x4_ASAP7_75t_L g816 ( 
.A(n_634),
.B(n_614),
.Y(n_816)
);

AND2x4_ASAP7_75t_L g817 ( 
.A(n_618),
.B(n_560),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_597),
.B(n_598),
.Y(n_818)
);

AND2x4_ASAP7_75t_L g819 ( 
.A(n_620),
.B(n_560),
.Y(n_819)
);

BUFx3_ASAP7_75t_L g820 ( 
.A(n_695),
.Y(n_820)
);

BUFx6f_ASAP7_75t_L g821 ( 
.A(n_659),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_734),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_603),
.Y(n_823)
);

INVx3_ASAP7_75t_L g824 ( 
.A(n_659),
.Y(n_824)
);

A2O1A1Ixp33_ASAP7_75t_L g825 ( 
.A1(n_639),
.A2(n_562),
.B(n_561),
.C(n_491),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_603),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_656),
.B(n_487),
.Y(n_827)
);

BUFx2_ASAP7_75t_L g828 ( 
.A(n_671),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_607),
.Y(n_829)
);

INVx1_ASAP7_75t_SL g830 ( 
.A(n_622),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_721),
.B(n_556),
.Y(n_831)
);

AOI22xp5_ASAP7_75t_L g832 ( 
.A1(n_616),
.A2(n_547),
.B1(n_578),
.B2(n_572),
.Y(n_832)
);

INVxp67_ASAP7_75t_SL g833 ( 
.A(n_689),
.Y(n_833)
);

AND2x4_ASAP7_75t_L g834 ( 
.A(n_697),
.B(n_701),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_613),
.B(n_457),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_734),
.Y(n_836)
);

AND2x6_ASAP7_75t_L g837 ( 
.A(n_641),
.B(n_561),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_607),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_623),
.B(n_556),
.Y(n_839)
);

INVx3_ASAP7_75t_L g840 ( 
.A(n_689),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_596),
.B(n_482),
.Y(n_841)
);

AND2x4_ASAP7_75t_L g842 ( 
.A(n_673),
.B(n_561),
.Y(n_842)
);

AND2x6_ASAP7_75t_L g843 ( 
.A(n_756),
.B(n_562),
.Y(n_843)
);

AND2x4_ASAP7_75t_L g844 ( 
.A(n_673),
.B(n_562),
.Y(n_844)
);

INVx4_ASAP7_75t_L g845 ( 
.A(n_692),
.Y(n_845)
);

AOI22xp5_ASAP7_75t_L g846 ( 
.A1(n_712),
.A2(n_578),
.B1(n_572),
.B2(n_547),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_623),
.Y(n_847)
);

AND2x4_ASAP7_75t_L g848 ( 
.A(n_720),
.B(n_543),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_612),
.B(n_495),
.Y(n_849)
);

AND3x1_ASAP7_75t_L g850 ( 
.A(n_652),
.B(n_497),
.C(n_487),
.Y(n_850)
);

AND2x4_ASAP7_75t_L g851 ( 
.A(n_666),
.B(n_543),
.Y(n_851)
);

HB1xp67_ASAP7_75t_L g852 ( 
.A(n_757),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_685),
.B(n_491),
.Y(n_853)
);

HB1xp67_ASAP7_75t_L g854 ( 
.A(n_757),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_644),
.B(n_572),
.Y(n_855)
);

INVxp67_ASAP7_75t_L g856 ( 
.A(n_612),
.Y(n_856)
);

AOI22xp33_ASAP7_75t_L g857 ( 
.A1(n_628),
.A2(n_495),
.B1(n_497),
.B2(n_487),
.Y(n_857)
);

AND2x2_ASAP7_75t_L g858 ( 
.A(n_631),
.B(n_495),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_626),
.Y(n_859)
);

INVx3_ASAP7_75t_L g860 ( 
.A(n_743),
.Y(n_860)
);

CKINVDCx8_ASAP7_75t_R g861 ( 
.A(n_712),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_644),
.B(n_500),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_700),
.B(n_482),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_629),
.B(n_556),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_631),
.B(n_482),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_661),
.B(n_482),
.Y(n_866)
);

OAI22xp5_ASAP7_75t_SL g867 ( 
.A1(n_664),
.A2(n_4),
.B1(n_5),
.B2(n_8),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_661),
.B(n_491),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_629),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_660),
.B(n_497),
.Y(n_870)
);

NOR2x2_ASAP7_75t_L g871 ( 
.A(n_672),
.B(n_11),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_636),
.B(n_556),
.Y(n_872)
);

NOR3xp33_ASAP7_75t_SL g873 ( 
.A(n_621),
.B(n_747),
.C(n_649),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_617),
.A2(n_480),
.B(n_577),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_636),
.B(n_556),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_691),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_696),
.B(n_491),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_714),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_714),
.B(n_493),
.Y(n_879)
);

AOI22xp5_ASAP7_75t_L g880 ( 
.A1(n_715),
.A2(n_493),
.B1(n_543),
.B2(n_448),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_743),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_749),
.Y(n_882)
);

NOR2x1_ASAP7_75t_L g883 ( 
.A(n_594),
.B(n_493),
.Y(n_883)
);

OR2x6_ASAP7_75t_L g884 ( 
.A(n_609),
.B(n_515),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_753),
.B(n_493),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_749),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_759),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_692),
.B(n_556),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_639),
.B(n_480),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_759),
.Y(n_890)
);

BUFx3_ASAP7_75t_L g891 ( 
.A(n_635),
.Y(n_891)
);

AO22x1_ASAP7_75t_L g892 ( 
.A1(n_715),
.A2(n_543),
.B1(n_489),
.B2(n_492),
.Y(n_892)
);

AOI22xp33_ASAP7_75t_L g893 ( 
.A1(n_628),
.A2(n_489),
.B1(n_448),
.B2(n_506),
.Y(n_893)
);

AO22x1_ASAP7_75t_L g894 ( 
.A1(n_640),
.A2(n_489),
.B1(n_448),
.B2(n_492),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_676),
.Y(n_895)
);

HB1xp67_ASAP7_75t_L g896 ( 
.A(n_637),
.Y(n_896)
);

AND2x6_ASAP7_75t_SL g897 ( 
.A(n_640),
.B(n_11),
.Y(n_897)
);

OAI22xp5_ASAP7_75t_L g898 ( 
.A1(n_633),
.A2(n_515),
.B1(n_492),
.B2(n_506),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_754),
.B(n_515),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_602),
.B(n_515),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_678),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_605),
.B(n_515),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_693),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_692),
.B(n_703),
.Y(n_904)
);

AOI22xp33_ASAP7_75t_L g905 ( 
.A1(n_633),
.A2(n_530),
.B1(n_492),
.B2(n_506),
.Y(n_905)
);

NAND2xp33_ASAP7_75t_SL g906 ( 
.A(n_645),
.B(n_530),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_646),
.Y(n_907)
);

INVx5_ASAP7_75t_L g908 ( 
.A(n_690),
.Y(n_908)
);

CKINVDCx20_ASAP7_75t_R g909 ( 
.A(n_716),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_610),
.B(n_530),
.Y(n_910)
);

BUFx12f_ASAP7_75t_L g911 ( 
.A(n_758),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_679),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_692),
.B(n_703),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_745),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_667),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_740),
.B(n_448),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_SL g917 ( 
.A(n_704),
.B(n_530),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_611),
.B(n_530),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_615),
.B(n_492),
.Y(n_919)
);

OR2x2_ASAP7_75t_SL g920 ( 
.A(n_621),
.B(n_12),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_SL g921 ( 
.A(n_630),
.B(n_632),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_680),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_675),
.A2(n_539),
.B(n_577),
.Y(n_923)
);

AOI22xp33_ASAP7_75t_L g924 ( 
.A1(n_675),
.A2(n_506),
.B1(n_551),
.B2(n_584),
.Y(n_924)
);

AND2x4_ASAP7_75t_L g925 ( 
.A(n_740),
.B(n_539),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_624),
.B(n_506),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_642),
.A2(n_577),
.B(n_558),
.Y(n_927)
);

HB1xp67_ASAP7_75t_L g928 ( 
.A(n_651),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_726),
.Y(n_929)
);

HB1xp67_ASAP7_75t_L g930 ( 
.A(n_731),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_653),
.B(n_551),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_L g932 ( 
.A(n_744),
.B(n_746),
.Y(n_932)
);

AOI22xp5_ASAP7_75t_L g933 ( 
.A1(n_744),
.A2(n_551),
.B1(n_577),
.B2(n_558),
.Y(n_933)
);

INVx2_ASAP7_75t_SL g934 ( 
.A(n_746),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_SL g935 ( 
.A(n_686),
.B(n_551),
.Y(n_935)
);

INVx2_ASAP7_75t_SL g936 ( 
.A(n_735),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_737),
.B(n_551),
.Y(n_937)
);

NOR3xp33_ASAP7_75t_SL g938 ( 
.A(n_738),
.B(n_15),
.C(n_16),
.Y(n_938)
);

BUFx12f_ASAP7_75t_L g939 ( 
.A(n_690),
.Y(n_939)
);

OR2x6_ASAP7_75t_L g940 ( 
.A(n_760),
.B(n_718),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_921),
.A2(n_684),
.B(n_681),
.Y(n_941)
);

OR2x2_ASAP7_75t_L g942 ( 
.A(n_830),
.B(n_741),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_777),
.Y(n_943)
);

AND2x4_ASAP7_75t_L g944 ( 
.A(n_851),
.B(n_690),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_780),
.Y(n_945)
);

INVx3_ASAP7_75t_L g946 ( 
.A(n_813),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_L g947 ( 
.A(n_856),
.B(n_739),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_796),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_SL g949 ( 
.A(n_856),
.B(n_861),
.Y(n_949)
);

BUFx12f_ASAP7_75t_L g950 ( 
.A(n_773),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_797),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_921),
.A2(n_627),
.B(n_718),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_772),
.B(n_915),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_814),
.Y(n_954)
);

BUFx4f_ASAP7_75t_L g955 ( 
.A(n_911),
.Y(n_955)
);

OR2x2_ASAP7_75t_L g956 ( 
.A(n_781),
.B(n_763),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_900),
.A2(n_719),
.B(n_722),
.Y(n_957)
);

NAND2xp33_ASAP7_75t_L g958 ( 
.A(n_873),
.B(n_690),
.Y(n_958)
);

BUFx2_ASAP7_75t_L g959 ( 
.A(n_828),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_902),
.A2(n_719),
.B(n_722),
.Y(n_960)
);

HB1xp67_ASAP7_75t_L g961 ( 
.A(n_776),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_773),
.Y(n_962)
);

OAI21x1_ASAP7_75t_L g963 ( 
.A1(n_799),
.A2(n_706),
.B(n_705),
.Y(n_963)
);

BUFx2_ASAP7_75t_L g964 ( 
.A(n_793),
.Y(n_964)
);

INVx3_ASAP7_75t_L g965 ( 
.A(n_813),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_910),
.A2(n_710),
.B(n_725),
.Y(n_966)
);

O2A1O1Ixp33_ASAP7_75t_L g967 ( 
.A1(n_768),
.A2(n_654),
.B(n_655),
.C(n_665),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_930),
.B(n_674),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_930),
.B(n_674),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_896),
.B(n_755),
.Y(n_970)
);

A2O1A1Ixp33_ASAP7_75t_L g971 ( 
.A1(n_932),
.A2(n_717),
.B(n_728),
.C(n_733),
.Y(n_971)
);

INVx3_ASAP7_75t_L g972 ( 
.A(n_813),
.Y(n_972)
);

NOR2x1_ASAP7_75t_L g973 ( 
.A(n_801),
.B(n_755),
.Y(n_973)
);

INVx3_ASAP7_75t_L g974 ( 
.A(n_813),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_764),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_L g976 ( 
.A(n_784),
.B(n_751),
.Y(n_976)
);

A2O1A1Ixp33_ASAP7_75t_L g977 ( 
.A1(n_932),
.A2(n_733),
.B(n_750),
.C(n_748),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_L g978 ( 
.A(n_936),
.B(n_751),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_896),
.B(n_928),
.Y(n_979)
);

OAI21xp5_ASAP7_75t_L g980 ( 
.A1(n_904),
.A2(n_750),
.B(n_748),
.Y(n_980)
);

HB1xp67_ASAP7_75t_L g981 ( 
.A(n_776),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_822),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_827),
.B(n_17),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_L g984 ( 
.A(n_928),
.B(n_17),
.Y(n_984)
);

O2A1O1Ixp33_ASAP7_75t_L g985 ( 
.A1(n_895),
.A2(n_724),
.B(n_22),
.C(n_24),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_901),
.B(n_558),
.Y(n_986)
);

AND2x4_ASAP7_75t_L g987 ( 
.A(n_851),
.B(n_480),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_912),
.B(n_558),
.Y(n_988)
);

AND2x6_ASAP7_75t_L g989 ( 
.A(n_766),
.B(n_584),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_922),
.B(n_539),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_818),
.A2(n_539),
.B(n_500),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_761),
.B(n_810),
.Y(n_992)
);

INVx5_ASAP7_75t_L g993 ( 
.A(n_762),
.Y(n_993)
);

OAI22x1_ASAP7_75t_L g994 ( 
.A1(n_929),
.A2(n_20),
.B1(n_22),
.B2(n_24),
.Y(n_994)
);

OR2x2_ASAP7_75t_L g995 ( 
.A(n_786),
.B(n_25),
.Y(n_995)
);

NOR2xp33_ASAP7_75t_L g996 ( 
.A(n_810),
.B(n_805),
.Y(n_996)
);

OAI22xp5_ASAP7_75t_L g997 ( 
.A1(n_889),
.A2(n_500),
.B1(n_480),
.B2(n_584),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_836),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_889),
.B(n_500),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_818),
.A2(n_584),
.B(n_75),
.Y(n_1000)
);

OAI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_904),
.A2(n_584),
.B(n_71),
.Y(n_1001)
);

A2O1A1Ixp33_ASAP7_75t_L g1002 ( 
.A1(n_873),
.A2(n_27),
.B(n_28),
.C(n_34),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_816),
.B(n_80),
.Y(n_1003)
);

BUFx12f_ASAP7_75t_L g1004 ( 
.A(n_907),
.Y(n_1004)
);

OAI22xp5_ASAP7_75t_L g1005 ( 
.A1(n_862),
.A2(n_79),
.B1(n_149),
.B2(n_147),
.Y(n_1005)
);

INVx4_ASAP7_75t_L g1006 ( 
.A(n_821),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_L g1007 ( 
.A(n_805),
.B(n_36),
.Y(n_1007)
);

A2O1A1Ixp33_ASAP7_75t_L g1008 ( 
.A1(n_934),
.A2(n_36),
.B(n_44),
.C(n_45),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_862),
.B(n_44),
.Y(n_1009)
);

A2O1A1Ixp33_ASAP7_75t_L g1010 ( 
.A1(n_855),
.A2(n_834),
.B(n_774),
.C(n_761),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_779),
.A2(n_81),
.B(n_140),
.Y(n_1011)
);

CKINVDCx16_ASAP7_75t_R g1012 ( 
.A(n_909),
.Y(n_1012)
);

INVx2_ASAP7_75t_SL g1013 ( 
.A(n_820),
.Y(n_1013)
);

BUFx2_ASAP7_75t_L g1014 ( 
.A(n_852),
.Y(n_1014)
);

INVx3_ASAP7_75t_L g1015 ( 
.A(n_821),
.Y(n_1015)
);

A2O1A1Ixp33_ASAP7_75t_L g1016 ( 
.A1(n_855),
.A2(n_45),
.B(n_46),
.C(n_49),
.Y(n_1016)
);

INVx3_ASAP7_75t_L g1017 ( 
.A(n_821),
.Y(n_1017)
);

NOR2xp67_ASAP7_75t_L g1018 ( 
.A(n_816),
.B(n_852),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_870),
.B(n_46),
.Y(n_1019)
);

A2O1A1Ixp33_ASAP7_75t_L g1020 ( 
.A1(n_834),
.A2(n_51),
.B(n_54),
.C(n_61),
.Y(n_1020)
);

OAI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_833),
.A2(n_62),
.B1(n_65),
.B2(n_67),
.Y(n_1021)
);

BUFx6f_ASAP7_75t_L g1022 ( 
.A(n_821),
.Y(n_1022)
);

HB1xp67_ASAP7_75t_L g1023 ( 
.A(n_860),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_849),
.B(n_150),
.Y(n_1024)
);

AND2x4_ASAP7_75t_SL g1025 ( 
.A(n_787),
.B(n_98),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_882),
.Y(n_1026)
);

AOI22xp5_ASAP7_75t_L g1027 ( 
.A1(n_771),
.A2(n_100),
.B1(n_104),
.B2(n_108),
.Y(n_1027)
);

BUFx2_ASAP7_75t_L g1028 ( 
.A(n_854),
.Y(n_1028)
);

O2A1O1Ixp33_ASAP7_75t_L g1029 ( 
.A1(n_866),
.A2(n_129),
.B(n_137),
.C(n_868),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_807),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_890),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_858),
.B(n_833),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_891),
.Y(n_1033)
);

NAND2xp33_ASAP7_75t_L g1034 ( 
.A(n_908),
.B(n_762),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_809),
.Y(n_1035)
);

O2A1O1Ixp33_ASAP7_75t_L g1036 ( 
.A1(n_825),
.A2(n_865),
.B(n_795),
.C(n_767),
.Y(n_1036)
);

OAI22x1_ASAP7_75t_L g1037 ( 
.A1(n_854),
.A2(n_778),
.B1(n_920),
.B2(n_771),
.Y(n_1037)
);

A2O1A1Ixp33_ASAP7_75t_L g1038 ( 
.A1(n_769),
.A2(n_783),
.B(n_848),
.C(n_916),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_SL g1039 ( 
.A(n_908),
.B(n_787),
.Y(n_1039)
);

A2O1A1Ixp33_ASAP7_75t_L g1040 ( 
.A1(n_848),
.A2(n_925),
.B(n_913),
.C(n_937),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_847),
.Y(n_1041)
);

BUFx12f_ASAP7_75t_L g1042 ( 
.A(n_806),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_876),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_L g1044 ( 
.A(n_903),
.B(n_914),
.Y(n_1044)
);

OAI22xp5_ASAP7_75t_L g1045 ( 
.A1(n_908),
.A2(n_792),
.B1(n_770),
.B2(n_893),
.Y(n_1045)
);

BUFx3_ASAP7_75t_L g1046 ( 
.A(n_765),
.Y(n_1046)
);

INVx1_ASAP7_75t_SL g1047 ( 
.A(n_871),
.Y(n_1047)
);

A2O1A1Ixp33_ASAP7_75t_L g1048 ( 
.A1(n_925),
.A2(n_913),
.B(n_885),
.C(n_899),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_878),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_918),
.A2(n_931),
.B(n_919),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_823),
.Y(n_1051)
);

OAI22xp5_ASAP7_75t_L g1052 ( 
.A1(n_908),
.A2(n_792),
.B1(n_770),
.B2(n_893),
.Y(n_1052)
);

OAI21x1_ASAP7_75t_L g1053 ( 
.A1(n_923),
.A2(n_874),
.B(n_927),
.Y(n_1053)
);

INVx1_ASAP7_75t_SL g1054 ( 
.A(n_788),
.Y(n_1054)
);

OAI22xp5_ASAP7_75t_L g1055 ( 
.A1(n_905),
.A2(n_924),
.B1(n_840),
.B2(n_880),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_826),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_926),
.A2(n_894),
.B(n_835),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_892),
.A2(n_782),
.B(n_853),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_886),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_840),
.B(n_829),
.Y(n_1060)
);

O2A1O1Ixp5_ASAP7_75t_L g1061 ( 
.A1(n_935),
.A2(n_917),
.B(n_790),
.C(n_831),
.Y(n_1061)
);

AOI21x1_ASAP7_75t_L g1062 ( 
.A1(n_935),
.A2(n_917),
.B(n_831),
.Y(n_1062)
);

AOI22xp5_ASAP7_75t_L g1063 ( 
.A1(n_850),
.A2(n_837),
.B1(n_883),
.B2(n_867),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_838),
.B(n_859),
.Y(n_1064)
);

INVxp67_ASAP7_75t_L g1065 ( 
.A(n_881),
.Y(n_1065)
);

INVx3_ASAP7_75t_SL g1066 ( 
.A(n_802),
.Y(n_1066)
);

OAI22xp5_ASAP7_75t_L g1067 ( 
.A1(n_905),
.A2(n_924),
.B1(n_846),
.B2(n_775),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_L g1068 ( 
.A(n_785),
.B(n_860),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_785),
.B(n_791),
.Y(n_1069)
);

INVx1_ASAP7_75t_SL g1070 ( 
.A(n_897),
.Y(n_1070)
);

AOI221x1_ASAP7_75t_L g1071 ( 
.A1(n_906),
.A2(n_898),
.B1(n_811),
.B2(n_841),
.C(n_863),
.Y(n_1071)
);

INVx1_ASAP7_75t_SL g1072 ( 
.A(n_765),
.Y(n_1072)
);

BUFx6f_ASAP7_75t_L g1073 ( 
.A(n_939),
.Y(n_1073)
);

BUFx3_ASAP7_75t_L g1074 ( 
.A(n_824),
.Y(n_1074)
);

OAI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_812),
.A2(n_857),
.B(n_775),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_SL g1076 ( 
.A(n_802),
.B(n_791),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_869),
.Y(n_1077)
);

NOR2x1_ASAP7_75t_L g1078 ( 
.A(n_824),
.B(n_845),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_L g1079 ( 
.A(n_789),
.B(n_794),
.Y(n_1079)
);

CKINVDCx16_ASAP7_75t_R g1080 ( 
.A(n_884),
.Y(n_1080)
);

OAI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_812),
.A2(n_857),
.B(n_879),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_SL g1082 ( 
.A(n_845),
.B(n_884),
.Y(n_1082)
);

AND2x4_ASAP7_75t_L g1083 ( 
.A(n_802),
.B(n_842),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_887),
.B(n_819),
.Y(n_1084)
);

BUFx6f_ASAP7_75t_L g1085 ( 
.A(n_1066),
.Y(n_1085)
);

AO32x2_ASAP7_75t_L g1086 ( 
.A1(n_1067),
.A2(n_938),
.A3(n_843),
.B1(n_837),
.B2(n_808),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_SL g1087 ( 
.A(n_956),
.B(n_842),
.Y(n_1087)
);

NAND2x1p5_ASAP7_75t_L g1088 ( 
.A(n_993),
.B(n_844),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_1030),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_999),
.A2(n_877),
.B(n_844),
.Y(n_1090)
);

OAI21x1_ASAP7_75t_L g1091 ( 
.A1(n_1053),
.A2(n_798),
.B(n_800),
.Y(n_1091)
);

OAI21x1_ASAP7_75t_L g1092 ( 
.A1(n_963),
.A2(n_815),
.B(n_832),
.Y(n_1092)
);

OAI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_1061),
.A2(n_1010),
.B(n_1048),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_947),
.B(n_837),
.Y(n_1094)
);

OAI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_1061),
.A2(n_843),
.B(n_837),
.Y(n_1095)
);

OAI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_941),
.A2(n_1050),
.B(n_966),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_947),
.B(n_819),
.Y(n_1097)
);

OAI21x1_ASAP7_75t_L g1098 ( 
.A1(n_991),
.A2(n_808),
.B(n_933),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_1050),
.A2(n_803),
.B(n_884),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_951),
.B(n_817),
.Y(n_1100)
);

OAI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_941),
.A2(n_843),
.B(n_804),
.Y(n_1101)
);

OAI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_966),
.A2(n_843),
.B(n_817),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1035),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_L g1104 ( 
.A(n_953),
.B(n_872),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_1034),
.A2(n_803),
.B(n_888),
.Y(n_1105)
);

NOR2x1_ASAP7_75t_L g1106 ( 
.A(n_949),
.B(n_888),
.Y(n_1106)
);

INVx4_ASAP7_75t_L g1107 ( 
.A(n_1066),
.Y(n_1107)
);

OA21x2_ASAP7_75t_L g1108 ( 
.A1(n_1058),
.A2(n_839),
.B(n_864),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_1057),
.A2(n_839),
.B(n_864),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_1051),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_1058),
.A2(n_872),
.B(n_875),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1056),
.Y(n_1112)
);

AND2x4_ASAP7_75t_L g1113 ( 
.A(n_1018),
.B(n_762),
.Y(n_1113)
);

AOI21x1_ASAP7_75t_L g1114 ( 
.A1(n_1062),
.A2(n_875),
.B(n_762),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_L g1115 ( 
.A(n_942),
.B(n_992),
.Y(n_1115)
);

NOR2xp67_ASAP7_75t_R g1116 ( 
.A(n_993),
.B(n_762),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_SL g1117 ( 
.A(n_993),
.B(n_938),
.Y(n_1117)
);

OAI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_977),
.A2(n_952),
.B(n_957),
.Y(n_1118)
);

BUFx3_ASAP7_75t_L g1119 ( 
.A(n_964),
.Y(n_1119)
);

OAI21x1_ASAP7_75t_L g1120 ( 
.A1(n_991),
.A2(n_957),
.B(n_960),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_979),
.B(n_978),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_SL g1122 ( 
.A1(n_1040),
.A2(n_1075),
.B(n_1045),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_1059),
.Y(n_1123)
);

OAI22x1_ASAP7_75t_L g1124 ( 
.A1(n_1069),
.A2(n_1007),
.B1(n_1068),
.B2(n_976),
.Y(n_1124)
);

AO31x2_ASAP7_75t_L g1125 ( 
.A1(n_1038),
.A2(n_1055),
.A3(n_1052),
.B(n_1000),
.Y(n_1125)
);

OAI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_1032),
.A2(n_969),
.B1(n_968),
.B2(n_1009),
.Y(n_1126)
);

AO22x2_ASAP7_75t_L g1127 ( 
.A1(n_1076),
.A2(n_1001),
.B1(n_1047),
.B2(n_995),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_967),
.A2(n_997),
.B(n_958),
.Y(n_1128)
);

AND2x4_ASAP7_75t_L g1129 ( 
.A(n_944),
.B(n_1083),
.Y(n_1129)
);

AO31x2_ASAP7_75t_L g1130 ( 
.A1(n_1000),
.A2(n_976),
.A3(n_1079),
.B(n_971),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_1079),
.B(n_970),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_996),
.B(n_1077),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_996),
.B(n_983),
.Y(n_1133)
);

O2A1O1Ixp33_ASAP7_75t_SL g1134 ( 
.A1(n_1002),
.A2(n_1016),
.B(n_1020),
.C(n_1003),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1064),
.Y(n_1135)
);

OAI21x1_ASAP7_75t_L g1136 ( 
.A1(n_1036),
.A2(n_980),
.B(n_1081),
.Y(n_1136)
);

A2O1A1Ixp33_ASAP7_75t_L g1137 ( 
.A1(n_1063),
.A2(n_1036),
.B(n_967),
.C(n_1029),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_1044),
.B(n_1023),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_1024),
.A2(n_993),
.B(n_986),
.Y(n_1139)
);

AO22x2_ASAP7_75t_L g1140 ( 
.A1(n_1005),
.A2(n_1019),
.B1(n_1054),
.B2(n_1011),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_943),
.Y(n_1141)
);

OAI21x1_ASAP7_75t_L g1142 ( 
.A1(n_1060),
.A2(n_1011),
.B(n_990),
.Y(n_1142)
);

BUFx6f_ASAP7_75t_L g1143 ( 
.A(n_1022),
.Y(n_1143)
);

OAI21x1_ASAP7_75t_L g1144 ( 
.A1(n_988),
.A2(n_1078),
.B(n_1084),
.Y(n_1144)
);

OAI21x1_ASAP7_75t_SL g1145 ( 
.A1(n_985),
.A2(n_1029),
.B(n_1027),
.Y(n_1145)
);

NOR2xp33_ASAP7_75t_L g1146 ( 
.A(n_959),
.B(n_1012),
.Y(n_1146)
);

OR2x2_ASAP7_75t_L g1147 ( 
.A(n_961),
.B(n_981),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_SL g1148 ( 
.A(n_1033),
.B(n_981),
.Y(n_1148)
);

OA21x2_ASAP7_75t_L g1149 ( 
.A1(n_1008),
.A2(n_1041),
.B(n_982),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_984),
.B(n_1044),
.Y(n_1150)
);

NOR3xp33_ASAP7_75t_SL g1151 ( 
.A(n_1080),
.B(n_962),
.C(n_984),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1065),
.B(n_961),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_945),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_948),
.Y(n_1154)
);

OAI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_989),
.A2(n_985),
.B(n_998),
.Y(n_1155)
);

OAI22x1_ASAP7_75t_L g1156 ( 
.A1(n_1014),
.A2(n_1028),
.B1(n_973),
.B2(n_1070),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_1082),
.A2(n_1039),
.B(n_1083),
.Y(n_1157)
);

AO31x2_ASAP7_75t_L g1158 ( 
.A1(n_1037),
.A2(n_1021),
.A3(n_994),
.B(n_1031),
.Y(n_1158)
);

OAI21x1_ASAP7_75t_L g1159 ( 
.A1(n_946),
.A2(n_965),
.B(n_1017),
.Y(n_1159)
);

AND2x2_ASAP7_75t_L g1160 ( 
.A(n_1025),
.B(n_1065),
.Y(n_1160)
);

AND2x2_ASAP7_75t_L g1161 ( 
.A(n_940),
.B(n_1042),
.Y(n_1161)
);

OAI21xp5_ASAP7_75t_SL g1162 ( 
.A1(n_944),
.A2(n_1073),
.B(n_1013),
.Y(n_1162)
);

NOR2x1_ASAP7_75t_SL g1163 ( 
.A(n_940),
.B(n_1022),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_954),
.Y(n_1164)
);

AND2x4_ASAP7_75t_L g1165 ( 
.A(n_1073),
.B(n_987),
.Y(n_1165)
);

AOI221x1_ASAP7_75t_L g1166 ( 
.A1(n_972),
.A2(n_1015),
.B1(n_974),
.B2(n_1049),
.C(n_1043),
.Y(n_1166)
);

OA22x2_ASAP7_75t_L g1167 ( 
.A1(n_940),
.A2(n_1072),
.B1(n_1023),
.B2(n_975),
.Y(n_1167)
);

OA21x2_ASAP7_75t_L g1168 ( 
.A1(n_1026),
.A2(n_989),
.B(n_987),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_1046),
.Y(n_1169)
);

INVx2_ASAP7_75t_L g1170 ( 
.A(n_1074),
.Y(n_1170)
);

BUFx3_ASAP7_75t_L g1171 ( 
.A(n_1004),
.Y(n_1171)
);

OAI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_989),
.A2(n_1006),
.B(n_955),
.Y(n_1172)
);

OAI21xp33_ASAP7_75t_L g1173 ( 
.A1(n_950),
.A2(n_682),
.B(n_523),
.Y(n_1173)
);

A2O1A1Ixp33_ASAP7_75t_L g1174 ( 
.A1(n_976),
.A2(n_772),
.B(n_932),
.C(n_1068),
.Y(n_1174)
);

OAI22xp5_ASAP7_75t_L g1175 ( 
.A1(n_1075),
.A2(n_1067),
.B1(n_915),
.B2(n_771),
.Y(n_1175)
);

NOR2xp33_ASAP7_75t_L g1176 ( 
.A(n_953),
.B(n_312),
.Y(n_1176)
);

OAI21x1_ASAP7_75t_L g1177 ( 
.A1(n_1053),
.A2(n_963),
.B(n_799),
.Y(n_1177)
);

O2A1O1Ixp5_ASAP7_75t_L g1178 ( 
.A1(n_1009),
.A2(n_976),
.B(n_953),
.C(n_1001),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_947),
.B(n_1032),
.Y(n_1179)
);

BUFx2_ASAP7_75t_L g1180 ( 
.A(n_964),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1030),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1030),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_950),
.Y(n_1183)
);

OAI22xp5_ASAP7_75t_L g1184 ( 
.A1(n_1075),
.A2(n_1067),
.B1(n_915),
.B2(n_771),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_999),
.A2(n_1050),
.B(n_921),
.Y(n_1185)
);

AND2x4_ASAP7_75t_L g1186 ( 
.A(n_1018),
.B(n_944),
.Y(n_1186)
);

NOR2xp33_ASAP7_75t_R g1187 ( 
.A(n_1033),
.B(n_501),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_947),
.B(n_1032),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_947),
.B(n_856),
.Y(n_1189)
);

OAI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1061),
.A2(n_1010),
.B(n_1048),
.Y(n_1190)
);

AOI21x1_ASAP7_75t_L g1191 ( 
.A1(n_1057),
.A2(n_894),
.B(n_892),
.Y(n_1191)
);

A2O1A1Ixp33_ASAP7_75t_L g1192 ( 
.A1(n_976),
.A2(n_772),
.B(n_932),
.C(n_1068),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_947),
.B(n_1032),
.Y(n_1193)
);

OA21x2_ASAP7_75t_L g1194 ( 
.A1(n_1071),
.A2(n_1061),
.B(n_1058),
.Y(n_1194)
);

INVx3_ASAP7_75t_L g1195 ( 
.A(n_1083),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_947),
.B(n_856),
.Y(n_1196)
);

AND3x4_ASAP7_75t_L g1197 ( 
.A(n_1018),
.B(n_760),
.C(n_801),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1030),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1030),
.Y(n_1199)
);

INVx3_ASAP7_75t_L g1200 ( 
.A(n_1083),
.Y(n_1200)
);

BUFx12f_ASAP7_75t_L g1201 ( 
.A(n_950),
.Y(n_1201)
);

OAI22xp5_ASAP7_75t_L g1202 ( 
.A1(n_1075),
.A2(n_1067),
.B1(n_915),
.B2(n_771),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_947),
.B(n_856),
.Y(n_1203)
);

NOR2xp67_ASAP7_75t_L g1204 ( 
.A(n_956),
.B(n_467),
.Y(n_1204)
);

OAI22xp5_ASAP7_75t_L g1205 ( 
.A1(n_1075),
.A2(n_1067),
.B1(n_915),
.B2(n_771),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1030),
.Y(n_1206)
);

BUFx3_ASAP7_75t_L g1207 ( 
.A(n_964),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_947),
.B(n_856),
.Y(n_1208)
);

OAI22xp5_ASAP7_75t_L g1209 ( 
.A1(n_1075),
.A2(n_1067),
.B1(n_915),
.B2(n_771),
.Y(n_1209)
);

AO21x2_ASAP7_75t_L g1210 ( 
.A1(n_1058),
.A2(n_1057),
.B(n_1050),
.Y(n_1210)
);

OR2x2_ASAP7_75t_L g1211 ( 
.A(n_956),
.B(n_830),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_SL g1212 ( 
.A1(n_1010),
.A2(n_1040),
.B(n_1075),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_1059),
.Y(n_1213)
);

BUFx3_ASAP7_75t_L g1214 ( 
.A(n_964),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_SL g1215 ( 
.A(n_956),
.B(n_861),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_999),
.A2(n_1050),
.B(n_921),
.Y(n_1216)
);

NOR2xp33_ASAP7_75t_L g1217 ( 
.A(n_953),
.B(n_312),
.Y(n_1217)
);

INVx3_ASAP7_75t_L g1218 ( 
.A(n_1083),
.Y(n_1218)
);

A2O1A1Ixp33_ASAP7_75t_L g1219 ( 
.A1(n_976),
.A2(n_772),
.B(n_932),
.C(n_1068),
.Y(n_1219)
);

AND2x4_ASAP7_75t_L g1220 ( 
.A(n_1018),
.B(n_944),
.Y(n_1220)
);

AOI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_953),
.A2(n_830),
.B1(n_622),
.B2(n_317),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_950),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_947),
.B(n_1032),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1096),
.A2(n_1216),
.B(n_1185),
.Y(n_1224)
);

HB1xp67_ASAP7_75t_L g1225 ( 
.A(n_1147),
.Y(n_1225)
);

OAI22xp33_ASAP7_75t_L g1226 ( 
.A1(n_1175),
.A2(n_1209),
.B1(n_1205),
.B2(n_1202),
.Y(n_1226)
);

OAI21x1_ASAP7_75t_SL g1227 ( 
.A1(n_1163),
.A2(n_1172),
.B(n_1155),
.Y(n_1227)
);

INVx3_ASAP7_75t_L g1228 ( 
.A(n_1129),
.Y(n_1228)
);

BUFx10_ASAP7_75t_L g1229 ( 
.A(n_1146),
.Y(n_1229)
);

OA21x2_ASAP7_75t_L g1230 ( 
.A1(n_1096),
.A2(n_1137),
.B(n_1093),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1212),
.A2(n_1128),
.B(n_1122),
.Y(n_1231)
);

AOI21x1_ASAP7_75t_L g1232 ( 
.A1(n_1191),
.A2(n_1099),
.B(n_1139),
.Y(n_1232)
);

AOI22xp5_ASAP7_75t_L g1233 ( 
.A1(n_1176),
.A2(n_1217),
.B1(n_1205),
.B2(n_1175),
.Y(n_1233)
);

BUFx2_ASAP7_75t_R g1234 ( 
.A(n_1183),
.Y(n_1234)
);

BUFx3_ASAP7_75t_L g1235 ( 
.A(n_1085),
.Y(n_1235)
);

OAI21x1_ASAP7_75t_L g1236 ( 
.A1(n_1120),
.A2(n_1092),
.B(n_1098),
.Y(n_1236)
);

OAI21x1_ASAP7_75t_L g1237 ( 
.A1(n_1102),
.A2(n_1111),
.B(n_1142),
.Y(n_1237)
);

AO31x2_ASAP7_75t_L g1238 ( 
.A1(n_1174),
.A2(n_1192),
.A3(n_1219),
.B(n_1184),
.Y(n_1238)
);

AOI21xp33_ASAP7_75t_SL g1239 ( 
.A1(n_1197),
.A2(n_1173),
.B(n_1215),
.Y(n_1239)
);

OAI21x1_ASAP7_75t_L g1240 ( 
.A1(n_1102),
.A2(n_1109),
.B(n_1095),
.Y(n_1240)
);

OAI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1178),
.A2(n_1202),
.B(n_1184),
.Y(n_1241)
);

OAI21x1_ASAP7_75t_L g1242 ( 
.A1(n_1095),
.A2(n_1101),
.B(n_1118),
.Y(n_1242)
);

OAI21x1_ASAP7_75t_L g1243 ( 
.A1(n_1101),
.A2(n_1118),
.B(n_1114),
.Y(n_1243)
);

BUFx4f_ASAP7_75t_L g1244 ( 
.A(n_1085),
.Y(n_1244)
);

INVx3_ASAP7_75t_L g1245 ( 
.A(n_1129),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1136),
.A2(n_1093),
.B(n_1190),
.Y(n_1246)
);

AO31x2_ASAP7_75t_L g1247 ( 
.A1(n_1209),
.A2(n_1124),
.A3(n_1126),
.B(n_1166),
.Y(n_1247)
);

AOI22xp5_ASAP7_75t_L g1248 ( 
.A1(n_1221),
.A2(n_1204),
.B1(n_1115),
.B2(n_1167),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1089),
.Y(n_1249)
);

AOI22xp33_ASAP7_75t_L g1250 ( 
.A1(n_1127),
.A2(n_1145),
.B1(n_1150),
.B2(n_1190),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_SL g1251 ( 
.A1(n_1172),
.A2(n_1155),
.B(n_1179),
.Y(n_1251)
);

INVx2_ASAP7_75t_SL g1252 ( 
.A(n_1119),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1103),
.Y(n_1253)
);

AND2x4_ASAP7_75t_L g1254 ( 
.A(n_1195),
.B(n_1200),
.Y(n_1254)
);

CKINVDCx16_ASAP7_75t_R g1255 ( 
.A(n_1187),
.Y(n_1255)
);

BUFx2_ASAP7_75t_L g1256 ( 
.A(n_1207),
.Y(n_1256)
);

HB1xp67_ASAP7_75t_L g1257 ( 
.A(n_1180),
.Y(n_1257)
);

A2O1A1Ixp33_ASAP7_75t_L g1258 ( 
.A1(n_1179),
.A2(n_1223),
.B(n_1193),
.C(n_1188),
.Y(n_1258)
);

INVx1_ASAP7_75t_SL g1259 ( 
.A(n_1214),
.Y(n_1259)
);

BUFx4f_ASAP7_75t_L g1260 ( 
.A(n_1085),
.Y(n_1260)
);

NAND3xp33_ASAP7_75t_SL g1261 ( 
.A(n_1121),
.B(n_1189),
.C(n_1203),
.Y(n_1261)
);

INVx2_ASAP7_75t_L g1262 ( 
.A(n_1168),
.Y(n_1262)
);

OAI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1126),
.A2(n_1131),
.B(n_1094),
.Y(n_1263)
);

OAI21x1_ASAP7_75t_SL g1264 ( 
.A1(n_1188),
.A2(n_1223),
.B(n_1193),
.Y(n_1264)
);

OAI21x1_ASAP7_75t_L g1265 ( 
.A1(n_1144),
.A2(n_1090),
.B(n_1105),
.Y(n_1265)
);

AND2x2_ASAP7_75t_L g1266 ( 
.A(n_1133),
.B(n_1211),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1110),
.Y(n_1267)
);

INVx3_ASAP7_75t_L g1268 ( 
.A(n_1195),
.Y(n_1268)
);

AOI22xp33_ASAP7_75t_L g1269 ( 
.A1(n_1127),
.A2(n_1140),
.B1(n_1131),
.B2(n_1208),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_1112),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_1201),
.Y(n_1271)
);

OAI21x1_ASAP7_75t_L g1272 ( 
.A1(n_1194),
.A2(n_1108),
.B(n_1159),
.Y(n_1272)
);

OA21x2_ASAP7_75t_L g1273 ( 
.A1(n_1138),
.A2(n_1104),
.B(n_1097),
.Y(n_1273)
);

AO31x2_ASAP7_75t_L g1274 ( 
.A1(n_1210),
.A2(n_1125),
.A3(n_1156),
.B(n_1138),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_1181),
.Y(n_1275)
);

OAI22xp33_ASAP7_75t_L g1276 ( 
.A1(n_1196),
.A2(n_1117),
.B1(n_1132),
.B2(n_1167),
.Y(n_1276)
);

AOI22xp5_ASAP7_75t_L g1277 ( 
.A1(n_1087),
.A2(n_1151),
.B1(n_1162),
.B2(n_1148),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1182),
.Y(n_1278)
);

BUFx2_ASAP7_75t_L g1279 ( 
.A(n_1160),
.Y(n_1279)
);

OA21x2_ASAP7_75t_L g1280 ( 
.A1(n_1132),
.A2(n_1206),
.B(n_1198),
.Y(n_1280)
);

INVx2_ASAP7_75t_L g1281 ( 
.A(n_1199),
.Y(n_1281)
);

OR2x2_ASAP7_75t_L g1282 ( 
.A(n_1152),
.B(n_1123),
.Y(n_1282)
);

OAI21x1_ASAP7_75t_L g1283 ( 
.A1(n_1149),
.A2(n_1157),
.B(n_1088),
.Y(n_1283)
);

OAI21x1_ASAP7_75t_L g1284 ( 
.A1(n_1088),
.A2(n_1106),
.B(n_1213),
.Y(n_1284)
);

OAI21x1_ASAP7_75t_L g1285 ( 
.A1(n_1164),
.A2(n_1154),
.B(n_1153),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1141),
.Y(n_1286)
);

NOR2xp33_ASAP7_75t_L g1287 ( 
.A(n_1135),
.B(n_1100),
.Y(n_1287)
);

HB1xp67_ASAP7_75t_L g1288 ( 
.A(n_1169),
.Y(n_1288)
);

AOI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1116),
.A2(n_1134),
.B(n_1140),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1130),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_1130),
.Y(n_1291)
);

OAI221xp5_ASAP7_75t_L g1292 ( 
.A1(n_1117),
.A2(n_1162),
.B1(n_1161),
.B2(n_1171),
.C(n_1170),
.Y(n_1292)
);

NAND2x1p5_ASAP7_75t_L g1293 ( 
.A(n_1107),
.B(n_1113),
.Y(n_1293)
);

NAND2x1p5_ASAP7_75t_L g1294 ( 
.A(n_1107),
.B(n_1113),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1143),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_SL g1296 ( 
.A(n_1186),
.B(n_1220),
.Y(n_1296)
);

AOI22xp5_ASAP7_75t_L g1297 ( 
.A1(n_1186),
.A2(n_1220),
.B1(n_1165),
.B2(n_1218),
.Y(n_1297)
);

INVx3_ASAP7_75t_L g1298 ( 
.A(n_1143),
.Y(n_1298)
);

NAND2x1p5_ASAP7_75t_L g1299 ( 
.A(n_1143),
.B(n_1158),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_1086),
.Y(n_1300)
);

OAI21x1_ASAP7_75t_L g1301 ( 
.A1(n_1158),
.A2(n_1177),
.B(n_1053),
.Y(n_1301)
);

OR2x2_ASAP7_75t_L g1302 ( 
.A(n_1158),
.B(n_1222),
.Y(n_1302)
);

O2A1O1Ixp33_ASAP7_75t_SL g1303 ( 
.A1(n_1174),
.A2(n_1002),
.B(n_1219),
.C(n_1192),
.Y(n_1303)
);

BUFx6f_ASAP7_75t_L g1304 ( 
.A(n_1085),
.Y(n_1304)
);

NAND2x1p5_ASAP7_75t_L g1305 ( 
.A(n_1168),
.B(n_993),
.Y(n_1305)
);

AOI221xp5_ASAP7_75t_L g1306 ( 
.A1(n_1175),
.A2(n_1202),
.B1(n_1209),
.B2(n_1205),
.C(n_1184),
.Y(n_1306)
);

OAI22xp5_ASAP7_75t_SL g1307 ( 
.A1(n_1176),
.A2(n_861),
.B1(n_569),
.B2(n_785),
.Y(n_1307)
);

BUFx2_ASAP7_75t_SL g1308 ( 
.A(n_1085),
.Y(n_1308)
);

AOI21xp5_ASAP7_75t_L g1309 ( 
.A1(n_1096),
.A2(n_1216),
.B(n_1185),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1089),
.Y(n_1310)
);

NAND2x1p5_ASAP7_75t_L g1311 ( 
.A(n_1168),
.B(n_993),
.Y(n_1311)
);

CKINVDCx14_ASAP7_75t_R g1312 ( 
.A(n_1187),
.Y(n_1312)
);

BUFx2_ASAP7_75t_SL g1313 ( 
.A(n_1085),
.Y(n_1313)
);

OAI21x1_ASAP7_75t_SL g1314 ( 
.A1(n_1163),
.A2(n_1172),
.B(n_1155),
.Y(n_1314)
);

AND2x4_ASAP7_75t_L g1315 ( 
.A(n_1195),
.B(n_1200),
.Y(n_1315)
);

HB1xp67_ASAP7_75t_L g1316 ( 
.A(n_1147),
.Y(n_1316)
);

OAI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1178),
.A2(n_1192),
.B(n_1174),
.Y(n_1317)
);

AOI22xp33_ASAP7_75t_L g1318 ( 
.A1(n_1175),
.A2(n_1202),
.B1(n_1209),
.B2(n_1184),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1150),
.B(n_1179),
.Y(n_1319)
);

OA21x2_ASAP7_75t_L g1320 ( 
.A1(n_1096),
.A2(n_1137),
.B(n_1093),
.Y(n_1320)
);

OAI22xp5_ASAP7_75t_L g1321 ( 
.A1(n_1221),
.A2(n_861),
.B1(n_915),
.B2(n_771),
.Y(n_1321)
);

OAI21x1_ASAP7_75t_L g1322 ( 
.A1(n_1177),
.A2(n_1053),
.B(n_1091),
.Y(n_1322)
);

BUFx2_ASAP7_75t_L g1323 ( 
.A(n_1119),
.Y(n_1323)
);

OAI22xp5_ASAP7_75t_L g1324 ( 
.A1(n_1221),
.A2(n_861),
.B1(n_915),
.B2(n_771),
.Y(n_1324)
);

OR2x2_ASAP7_75t_L g1325 ( 
.A(n_1211),
.B(n_1133),
.Y(n_1325)
);

AOI22xp33_ASAP7_75t_L g1326 ( 
.A1(n_1175),
.A2(n_1202),
.B1(n_1209),
.B2(n_1184),
.Y(n_1326)
);

OA21x2_ASAP7_75t_L g1327 ( 
.A1(n_1096),
.A2(n_1137),
.B(n_1093),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1150),
.B(n_1179),
.Y(n_1328)
);

A2O1A1Ixp33_ASAP7_75t_L g1329 ( 
.A1(n_1175),
.A2(n_1202),
.B(n_1205),
.C(n_1184),
.Y(n_1329)
);

BUFx2_ASAP7_75t_L g1330 ( 
.A(n_1119),
.Y(n_1330)
);

OAI22xp33_ASAP7_75t_SL g1331 ( 
.A1(n_1175),
.A2(n_1184),
.B1(n_1205),
.B2(n_1202),
.Y(n_1331)
);

AOI22xp33_ASAP7_75t_L g1332 ( 
.A1(n_1175),
.A2(n_1202),
.B1(n_1209),
.B2(n_1184),
.Y(n_1332)
);

NOR2xp33_ASAP7_75t_L g1333 ( 
.A(n_1175),
.B(n_1184),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1089),
.Y(n_1334)
);

AOI22xp5_ASAP7_75t_L g1335 ( 
.A1(n_1176),
.A2(n_312),
.B1(n_322),
.B2(n_317),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1089),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1089),
.Y(n_1337)
);

INVx6_ASAP7_75t_L g1338 ( 
.A(n_1085),
.Y(n_1338)
);

OAI21x1_ASAP7_75t_L g1339 ( 
.A1(n_1177),
.A2(n_1053),
.B(n_1091),
.Y(n_1339)
);

OAI21x1_ASAP7_75t_L g1340 ( 
.A1(n_1177),
.A2(n_1053),
.B(n_1091),
.Y(n_1340)
);

OAI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1178),
.A2(n_1192),
.B(n_1174),
.Y(n_1341)
);

INVx2_ASAP7_75t_SL g1342 ( 
.A(n_1119),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_SL g1343 ( 
.A(n_1174),
.B(n_1192),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1266),
.B(n_1325),
.Y(n_1344)
);

AOI221x1_ASAP7_75t_SL g1345 ( 
.A1(n_1226),
.A2(n_1321),
.B1(n_1324),
.B2(n_1333),
.C(n_1276),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1274),
.B(n_1241),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1274),
.B(n_1318),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1274),
.B(n_1318),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1279),
.B(n_1287),
.Y(n_1349)
);

OAI22xp5_ASAP7_75t_L g1350 ( 
.A1(n_1326),
.A2(n_1332),
.B1(n_1233),
.B2(n_1329),
.Y(n_1350)
);

INVx3_ASAP7_75t_SL g1351 ( 
.A(n_1271),
.Y(n_1351)
);

AOI21xp5_ASAP7_75t_L g1352 ( 
.A1(n_1231),
.A2(n_1309),
.B(n_1224),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1287),
.B(n_1248),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1282),
.B(n_1288),
.Y(n_1354)
);

AOI221xp5_ASAP7_75t_L g1355 ( 
.A1(n_1226),
.A2(n_1331),
.B1(n_1306),
.B2(n_1332),
.C(n_1326),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1225),
.B(n_1316),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1239),
.B(n_1228),
.Y(n_1357)
);

O2A1O1Ixp33_ASAP7_75t_L g1358 ( 
.A1(n_1329),
.A2(n_1333),
.B(n_1303),
.C(n_1343),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1319),
.B(n_1328),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1261),
.B(n_1258),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1228),
.B(n_1245),
.Y(n_1361)
);

OAI22xp5_ASAP7_75t_L g1362 ( 
.A1(n_1307),
.A2(n_1277),
.B1(n_1292),
.B2(n_1250),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1245),
.B(n_1257),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1258),
.B(n_1264),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1286),
.B(n_1250),
.Y(n_1365)
);

OA21x2_ASAP7_75t_L g1366 ( 
.A1(n_1237),
.A2(n_1240),
.B(n_1236),
.Y(n_1366)
);

O2A1O1Ixp33_ASAP7_75t_L g1367 ( 
.A1(n_1303),
.A2(n_1343),
.B(n_1341),
.C(n_1317),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1263),
.B(n_1273),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1274),
.B(n_1273),
.Y(n_1369)
);

INVxp67_ASAP7_75t_L g1370 ( 
.A(n_1256),
.Y(n_1370)
);

HB1xp67_ASAP7_75t_L g1371 ( 
.A(n_1262),
.Y(n_1371)
);

AND2x4_ASAP7_75t_L g1372 ( 
.A(n_1270),
.B(n_1275),
.Y(n_1372)
);

INVx3_ASAP7_75t_L g1373 ( 
.A(n_1305),
.Y(n_1373)
);

OAI22xp5_ASAP7_75t_L g1374 ( 
.A1(n_1269),
.A2(n_1302),
.B1(n_1335),
.B2(n_1297),
.Y(n_1374)
);

OAI22xp5_ASAP7_75t_L g1375 ( 
.A1(n_1276),
.A2(n_1312),
.B1(n_1244),
.B2(n_1260),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1254),
.B(n_1315),
.Y(n_1376)
);

AND2x4_ASAP7_75t_L g1377 ( 
.A(n_1270),
.B(n_1275),
.Y(n_1377)
);

OAI22xp5_ASAP7_75t_L g1378 ( 
.A1(n_1312),
.A2(n_1260),
.B1(n_1244),
.B2(n_1255),
.Y(n_1378)
);

AOI21x1_ASAP7_75t_SL g1379 ( 
.A1(n_1254),
.A2(n_1315),
.B(n_1234),
.Y(n_1379)
);

OAI22xp5_ASAP7_75t_L g1380 ( 
.A1(n_1259),
.A2(n_1296),
.B1(n_1323),
.B2(n_1330),
.Y(n_1380)
);

OR2x2_ASAP7_75t_L g1381 ( 
.A(n_1238),
.B(n_1281),
.Y(n_1381)
);

NAND2x1p5_ASAP7_75t_L g1382 ( 
.A(n_1280),
.B(n_1284),
.Y(n_1382)
);

CKINVDCx5p33_ASAP7_75t_R g1383 ( 
.A(n_1271),
.Y(n_1383)
);

O2A1O1Ixp5_ASAP7_75t_L g1384 ( 
.A1(n_1289),
.A2(n_1290),
.B(n_1291),
.C(n_1232),
.Y(n_1384)
);

CKINVDCx20_ASAP7_75t_R g1385 ( 
.A(n_1235),
.Y(n_1385)
);

NOR2xp67_ASAP7_75t_L g1386 ( 
.A(n_1252),
.B(n_1342),
.Y(n_1386)
);

AOI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1230),
.A2(n_1327),
.B(n_1320),
.Y(n_1387)
);

O2A1O1Ixp33_ASAP7_75t_L g1388 ( 
.A1(n_1251),
.A2(n_1227),
.B(n_1314),
.C(n_1296),
.Y(n_1388)
);

OA21x2_ASAP7_75t_L g1389 ( 
.A1(n_1237),
.A2(n_1240),
.B(n_1236),
.Y(n_1389)
);

O2A1O1Ixp33_ASAP7_75t_L g1390 ( 
.A1(n_1249),
.A2(n_1253),
.B(n_1278),
.C(n_1334),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1238),
.B(n_1327),
.Y(n_1391)
);

AOI21xp5_ASAP7_75t_L g1392 ( 
.A1(n_1230),
.A2(n_1320),
.B(n_1327),
.Y(n_1392)
);

OA21x2_ASAP7_75t_L g1393 ( 
.A1(n_1243),
.A2(n_1301),
.B(n_1272),
.Y(n_1393)
);

INVx3_ASAP7_75t_SL g1394 ( 
.A(n_1338),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1281),
.B(n_1280),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1267),
.Y(n_1396)
);

AOI21xp5_ASAP7_75t_SL g1397 ( 
.A1(n_1230),
.A2(n_1320),
.B(n_1311),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1310),
.Y(n_1398)
);

OR2x2_ASAP7_75t_L g1399 ( 
.A(n_1238),
.B(n_1337),
.Y(n_1399)
);

OAI22xp5_ASAP7_75t_L g1400 ( 
.A1(n_1293),
.A2(n_1294),
.B1(n_1336),
.B2(n_1338),
.Y(n_1400)
);

AOI21xp5_ASAP7_75t_L g1401 ( 
.A1(n_1265),
.A2(n_1311),
.B(n_1305),
.Y(n_1401)
);

OAI22xp5_ASAP7_75t_SL g1402 ( 
.A1(n_1338),
.A2(n_1293),
.B1(n_1294),
.B2(n_1235),
.Y(n_1402)
);

OAI22xp5_ASAP7_75t_L g1403 ( 
.A1(n_1268),
.A2(n_1308),
.B1(n_1313),
.B2(n_1299),
.Y(n_1403)
);

AND2x4_ASAP7_75t_L g1404 ( 
.A(n_1285),
.B(n_1283),
.Y(n_1404)
);

HB1xp67_ASAP7_75t_L g1405 ( 
.A(n_1246),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1229),
.B(n_1285),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1295),
.B(n_1298),
.Y(n_1407)
);

OR2x2_ASAP7_75t_L g1408 ( 
.A(n_1247),
.B(n_1246),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1300),
.B(n_1242),
.Y(n_1409)
);

INVxp67_ASAP7_75t_L g1410 ( 
.A(n_1304),
.Y(n_1410)
);

INVxp33_ASAP7_75t_L g1411 ( 
.A(n_1304),
.Y(n_1411)
);

AND2x4_ASAP7_75t_L g1412 ( 
.A(n_1322),
.B(n_1339),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1340),
.B(n_1266),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1266),
.B(n_1325),
.Y(n_1414)
);

OR2x2_ASAP7_75t_L g1415 ( 
.A(n_1325),
.B(n_1225),
.Y(n_1415)
);

INVx1_ASAP7_75t_SL g1416 ( 
.A(n_1259),
.Y(n_1416)
);

BUFx2_ASAP7_75t_L g1417 ( 
.A(n_1257),
.Y(n_1417)
);

OAI22xp5_ASAP7_75t_L g1418 ( 
.A1(n_1318),
.A2(n_1326),
.B1(n_1332),
.B2(n_1233),
.Y(n_1418)
);

INVx1_ASAP7_75t_SL g1419 ( 
.A(n_1259),
.Y(n_1419)
);

AOI21xp5_ASAP7_75t_L g1420 ( 
.A1(n_1231),
.A2(n_1309),
.B(n_1224),
.Y(n_1420)
);

BUFx3_ASAP7_75t_L g1421 ( 
.A(n_1244),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1266),
.B(n_1325),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1266),
.B(n_1319),
.Y(n_1423)
);

OR2x2_ASAP7_75t_L g1424 ( 
.A(n_1325),
.B(n_1225),
.Y(n_1424)
);

AOI21xp5_ASAP7_75t_L g1425 ( 
.A1(n_1231),
.A2(n_1309),
.B(n_1224),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1266),
.B(n_1319),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1391),
.B(n_1409),
.Y(n_1427)
);

AO21x2_ASAP7_75t_L g1428 ( 
.A1(n_1352),
.A2(n_1425),
.B(n_1420),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_SL g1429 ( 
.A(n_1367),
.B(n_1358),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1391),
.B(n_1409),
.Y(n_1430)
);

INVx3_ASAP7_75t_L g1431 ( 
.A(n_1404),
.Y(n_1431)
);

INVx1_ASAP7_75t_SL g1432 ( 
.A(n_1349),
.Y(n_1432)
);

OA21x2_ASAP7_75t_L g1433 ( 
.A1(n_1387),
.A2(n_1392),
.B(n_1384),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1395),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1413),
.B(n_1368),
.Y(n_1435)
);

AOI22xp33_ASAP7_75t_L g1436 ( 
.A1(n_1350),
.A2(n_1418),
.B1(n_1355),
.B2(n_1362),
.Y(n_1436)
);

OR2x6_ASAP7_75t_L g1437 ( 
.A(n_1397),
.B(n_1401),
.Y(n_1437)
);

OR2x2_ASAP7_75t_L g1438 ( 
.A(n_1408),
.B(n_1369),
.Y(n_1438)
);

OR2x2_ASAP7_75t_L g1439 ( 
.A(n_1369),
.B(n_1346),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1346),
.B(n_1347),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1347),
.B(n_1348),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1371),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1360),
.B(n_1348),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1382),
.Y(n_1444)
);

OAI21xp5_ASAP7_75t_L g1445 ( 
.A1(n_1364),
.A2(n_1374),
.B(n_1353),
.Y(n_1445)
);

BUFx4f_ASAP7_75t_SL g1446 ( 
.A(n_1385),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1405),
.B(n_1381),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1359),
.B(n_1365),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1393),
.Y(n_1449)
);

OR2x2_ASAP7_75t_L g1450 ( 
.A(n_1405),
.B(n_1399),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1393),
.Y(n_1451)
);

INVx3_ASAP7_75t_L g1452 ( 
.A(n_1412),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1396),
.Y(n_1453)
);

OA21x2_ASAP7_75t_L g1454 ( 
.A1(n_1398),
.A2(n_1406),
.B(n_1372),
.Y(n_1454)
);

AO21x2_ASAP7_75t_L g1455 ( 
.A1(n_1388),
.A2(n_1390),
.B(n_1377),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1372),
.Y(n_1456)
);

AOI21x1_ASAP7_75t_L g1457 ( 
.A1(n_1366),
.A2(n_1389),
.B(n_1403),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1377),
.Y(n_1458)
);

INVxp67_ASAP7_75t_R g1459 ( 
.A(n_1402),
.Y(n_1459)
);

INVx1_ASAP7_75t_SL g1460 ( 
.A(n_1415),
.Y(n_1460)
);

INVx4_ASAP7_75t_SL g1461 ( 
.A(n_1394),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1366),
.Y(n_1462)
);

BUFx3_ASAP7_75t_L g1463 ( 
.A(n_1373),
.Y(n_1463)
);

HB1xp67_ASAP7_75t_L g1464 ( 
.A(n_1356),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1354),
.Y(n_1465)
);

AO21x2_ASAP7_75t_L g1466 ( 
.A1(n_1400),
.A2(n_1375),
.B(n_1357),
.Y(n_1466)
);

BUFx3_ASAP7_75t_L g1467 ( 
.A(n_1463),
.Y(n_1467)
);

OR2x2_ASAP7_75t_L g1468 ( 
.A(n_1439),
.B(n_1424),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1427),
.B(n_1344),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1427),
.B(n_1414),
.Y(n_1470)
);

OR2x2_ASAP7_75t_L g1471 ( 
.A(n_1439),
.B(n_1417),
.Y(n_1471)
);

OAI222xp33_ASAP7_75t_L g1472 ( 
.A1(n_1436),
.A2(n_1345),
.B1(n_1426),
.B2(n_1423),
.C1(n_1380),
.C2(n_1422),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1427),
.B(n_1376),
.Y(n_1473)
);

OR2x2_ASAP7_75t_L g1474 ( 
.A(n_1439),
.B(n_1363),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1435),
.B(n_1370),
.Y(n_1475)
);

NOR2xp33_ASAP7_75t_L g1476 ( 
.A(n_1446),
.B(n_1416),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1453),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1453),
.Y(n_1478)
);

NOR2xp33_ASAP7_75t_L g1479 ( 
.A(n_1446),
.B(n_1419),
.Y(n_1479)
);

HB1xp67_ASAP7_75t_L g1480 ( 
.A(n_1454),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1435),
.B(n_1434),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1449),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1434),
.B(n_1407),
.Y(n_1483)
);

AND2x6_ASAP7_75t_L g1484 ( 
.A(n_1456),
.B(n_1361),
.Y(n_1484)
);

AOI22xp33_ASAP7_75t_L g1485 ( 
.A1(n_1436),
.A2(n_1378),
.B1(n_1385),
.B2(n_1421),
.Y(n_1485)
);

INVx2_ASAP7_75t_SL g1486 ( 
.A(n_1452),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_SL g1487 ( 
.A(n_1445),
.B(n_1448),
.Y(n_1487)
);

NAND3xp33_ASAP7_75t_SL g1488 ( 
.A(n_1429),
.B(n_1383),
.C(n_1411),
.Y(n_1488)
);

AO21x1_ASAP7_75t_L g1489 ( 
.A1(n_1429),
.A2(n_1379),
.B(n_1410),
.Y(n_1489)
);

AND2x4_ASAP7_75t_L g1490 ( 
.A(n_1431),
.B(n_1386),
.Y(n_1490)
);

AOI22xp33_ASAP7_75t_L g1491 ( 
.A1(n_1445),
.A2(n_1421),
.B1(n_1351),
.B2(n_1383),
.Y(n_1491)
);

BUFx2_ASAP7_75t_L g1492 ( 
.A(n_1454),
.Y(n_1492)
);

AOI22xp33_ASAP7_75t_L g1493 ( 
.A1(n_1487),
.A2(n_1466),
.B1(n_1443),
.B2(n_1448),
.Y(n_1493)
);

OAI22xp5_ASAP7_75t_L g1494 ( 
.A1(n_1491),
.A2(n_1459),
.B1(n_1443),
.B2(n_1460),
.Y(n_1494)
);

NAND3xp33_ASAP7_75t_L g1495 ( 
.A(n_1491),
.B(n_1485),
.C(n_1475),
.Y(n_1495)
);

AOI31xp33_ASAP7_75t_L g1496 ( 
.A1(n_1489),
.A2(n_1432),
.A3(n_1460),
.B(n_1464),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1475),
.B(n_1464),
.Y(n_1497)
);

OR2x6_ASAP7_75t_L g1498 ( 
.A(n_1489),
.B(n_1437),
.Y(n_1498)
);

HB1xp67_ASAP7_75t_L g1499 ( 
.A(n_1480),
.Y(n_1499)
);

AO21x2_ASAP7_75t_L g1500 ( 
.A1(n_1480),
.A2(n_1462),
.B(n_1457),
.Y(n_1500)
);

AOI221xp5_ASAP7_75t_L g1501 ( 
.A1(n_1472),
.A2(n_1432),
.B1(n_1465),
.B2(n_1434),
.C(n_1466),
.Y(n_1501)
);

AOI222xp33_ASAP7_75t_L g1502 ( 
.A1(n_1472),
.A2(n_1465),
.B1(n_1440),
.B2(n_1441),
.C1(n_1447),
.C2(n_1456),
.Y(n_1502)
);

AND2x6_ASAP7_75t_SL g1503 ( 
.A(n_1476),
.B(n_1351),
.Y(n_1503)
);

AND2x4_ASAP7_75t_L g1504 ( 
.A(n_1490),
.B(n_1467),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1469),
.B(n_1430),
.Y(n_1505)
);

INVxp67_ASAP7_75t_L g1506 ( 
.A(n_1481),
.Y(n_1506)
);

OR2x2_ASAP7_75t_L g1507 ( 
.A(n_1468),
.B(n_1438),
.Y(n_1507)
);

AO21x2_ASAP7_75t_L g1508 ( 
.A1(n_1482),
.A2(n_1462),
.B(n_1457),
.Y(n_1508)
);

INVx5_ASAP7_75t_L g1509 ( 
.A(n_1484),
.Y(n_1509)
);

NAND2xp33_ASAP7_75t_R g1510 ( 
.A(n_1490),
.B(n_1483),
.Y(n_1510)
);

OR2x2_ASAP7_75t_L g1511 ( 
.A(n_1468),
.B(n_1474),
.Y(n_1511)
);

AOI221xp5_ASAP7_75t_L g1512 ( 
.A1(n_1488),
.A2(n_1465),
.B1(n_1466),
.B2(n_1456),
.C(n_1441),
.Y(n_1512)
);

AOI22xp33_ASAP7_75t_SL g1513 ( 
.A1(n_1492),
.A2(n_1455),
.B1(n_1466),
.B2(n_1428),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_1474),
.Y(n_1514)
);

OAI22xp5_ASAP7_75t_L g1515 ( 
.A1(n_1485),
.A2(n_1459),
.B1(n_1394),
.B2(n_1438),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1477),
.Y(n_1516)
);

OR2x2_ASAP7_75t_L g1517 ( 
.A(n_1471),
.B(n_1438),
.Y(n_1517)
);

CKINVDCx5p33_ASAP7_75t_R g1518 ( 
.A(n_1479),
.Y(n_1518)
);

HB1xp67_ASAP7_75t_L g1519 ( 
.A(n_1492),
.Y(n_1519)
);

AOI221xp5_ASAP7_75t_L g1520 ( 
.A1(n_1488),
.A2(n_1466),
.B1(n_1441),
.B2(n_1440),
.C(n_1447),
.Y(n_1520)
);

OR2x2_ASAP7_75t_L g1521 ( 
.A(n_1469),
.B(n_1458),
.Y(n_1521)
);

INVx4_ASAP7_75t_L g1522 ( 
.A(n_1467),
.Y(n_1522)
);

INVx2_ASAP7_75t_SL g1523 ( 
.A(n_1473),
.Y(n_1523)
);

OAI31xp33_ASAP7_75t_L g1524 ( 
.A1(n_1467),
.A2(n_1463),
.A3(n_1444),
.B(n_1450),
.Y(n_1524)
);

AOI221xp5_ASAP7_75t_L g1525 ( 
.A1(n_1483),
.A2(n_1440),
.B1(n_1447),
.B2(n_1455),
.C(n_1442),
.Y(n_1525)
);

NOR2xp33_ASAP7_75t_L g1526 ( 
.A(n_1469),
.B(n_1458),
.Y(n_1526)
);

INVxp67_ASAP7_75t_L g1527 ( 
.A(n_1477),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1478),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1527),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1516),
.Y(n_1530)
);

AOI21xp5_ASAP7_75t_SL g1531 ( 
.A1(n_1496),
.A2(n_1455),
.B(n_1437),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1508),
.Y(n_1532)
);

HB1xp67_ASAP7_75t_L g1533 ( 
.A(n_1527),
.Y(n_1533)
);

OA21x2_ASAP7_75t_L g1534 ( 
.A1(n_1525),
.A2(n_1520),
.B(n_1512),
.Y(n_1534)
);

BUFx6f_ASAP7_75t_L g1535 ( 
.A(n_1509),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1508),
.Y(n_1536)
);

BUFx2_ASAP7_75t_L g1537 ( 
.A(n_1498),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1528),
.Y(n_1538)
);

HB1xp67_ASAP7_75t_L g1539 ( 
.A(n_1499),
.Y(n_1539)
);

AO21x2_ASAP7_75t_L g1540 ( 
.A1(n_1500),
.A2(n_1462),
.B(n_1451),
.Y(n_1540)
);

BUFx2_ASAP7_75t_L g1541 ( 
.A(n_1498),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1500),
.Y(n_1542)
);

AOI21xp5_ASAP7_75t_L g1543 ( 
.A1(n_1498),
.A2(n_1428),
.B(n_1437),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1519),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1506),
.B(n_1470),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1509),
.Y(n_1546)
);

BUFx2_ASAP7_75t_L g1547 ( 
.A(n_1509),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1509),
.Y(n_1548)
);

INVx2_ASAP7_75t_SL g1549 ( 
.A(n_1504),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_SL g1550 ( 
.A(n_1501),
.B(n_1461),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1511),
.Y(n_1551)
);

INVx1_ASAP7_75t_SL g1552 ( 
.A(n_1503),
.Y(n_1552)
);

NAND3xp33_ASAP7_75t_L g1553 ( 
.A(n_1501),
.B(n_1433),
.C(n_1437),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1507),
.Y(n_1554)
);

NOR2xp33_ASAP7_75t_L g1555 ( 
.A(n_1495),
.B(n_1470),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1514),
.Y(n_1556)
);

INVx3_ASAP7_75t_L g1557 ( 
.A(n_1504),
.Y(n_1557)
);

INVx4_ASAP7_75t_SL g1558 ( 
.A(n_1523),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1533),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1555),
.B(n_1493),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1537),
.B(n_1505),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1537),
.B(n_1522),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1537),
.B(n_1526),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1540),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1540),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1541),
.B(n_1513),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1533),
.Y(n_1567)
);

NOR2xp33_ASAP7_75t_L g1568 ( 
.A(n_1552),
.B(n_1518),
.Y(n_1568)
);

OR2x2_ASAP7_75t_L g1569 ( 
.A(n_1554),
.B(n_1517),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1538),
.Y(n_1570)
);

AND2x2_ASAP7_75t_SL g1571 ( 
.A(n_1534),
.B(n_1520),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1555),
.B(n_1497),
.Y(n_1572)
);

INVx1_ASAP7_75t_SL g1573 ( 
.A(n_1552),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1541),
.B(n_1513),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1541),
.B(n_1470),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1529),
.B(n_1525),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1538),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1557),
.B(n_1512),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_SL g1579 ( 
.A(n_1535),
.B(n_1502),
.Y(n_1579)
);

AND2x4_ASAP7_75t_L g1580 ( 
.A(n_1558),
.B(n_1486),
.Y(n_1580)
);

OR2x2_ASAP7_75t_L g1581 ( 
.A(n_1554),
.B(n_1521),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1538),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1530),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1558),
.B(n_1524),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1530),
.Y(n_1585)
);

NOR2x1_ASAP7_75t_L g1586 ( 
.A(n_1531),
.B(n_1494),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1529),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1539),
.Y(n_1588)
);

HB1xp67_ASAP7_75t_L g1589 ( 
.A(n_1539),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1540),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1551),
.B(n_1473),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1540),
.Y(n_1592)
);

HB1xp67_ASAP7_75t_L g1593 ( 
.A(n_1544),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1551),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1544),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1557),
.B(n_1473),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1573),
.B(n_1545),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1573),
.B(n_1550),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1571),
.B(n_1550),
.Y(n_1599)
);

OAI22xp5_ASAP7_75t_L g1600 ( 
.A1(n_1586),
.A2(n_1553),
.B1(n_1534),
.B2(n_1459),
.Y(n_1600)
);

INVxp67_ASAP7_75t_L g1601 ( 
.A(n_1568),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1589),
.Y(n_1602)
);

INVx3_ASAP7_75t_L g1603 ( 
.A(n_1580),
.Y(n_1603)
);

OAI22xp33_ASAP7_75t_SL g1604 ( 
.A1(n_1586),
.A2(n_1547),
.B1(n_1549),
.B2(n_1557),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1562),
.B(n_1557),
.Y(n_1605)
);

AND2x4_ASAP7_75t_L g1606 ( 
.A(n_1562),
.B(n_1558),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1589),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1587),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1596),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1571),
.B(n_1556),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1587),
.Y(n_1611)
);

HB1xp67_ASAP7_75t_L g1612 ( 
.A(n_1588),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1583),
.Y(n_1613)
);

OR2x2_ASAP7_75t_L g1614 ( 
.A(n_1588),
.B(n_1534),
.Y(n_1614)
);

AND2x4_ASAP7_75t_L g1615 ( 
.A(n_1575),
.B(n_1558),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_SL g1616 ( 
.A(n_1571),
.B(n_1535),
.Y(n_1616)
);

NOR2xp33_ASAP7_75t_L g1617 ( 
.A(n_1560),
.B(n_1549),
.Y(n_1617)
);

INVx2_ASAP7_75t_SL g1618 ( 
.A(n_1593),
.Y(n_1618)
);

BUFx2_ASAP7_75t_L g1619 ( 
.A(n_1559),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1560),
.B(n_1556),
.Y(n_1620)
);

HB1xp67_ASAP7_75t_L g1621 ( 
.A(n_1559),
.Y(n_1621)
);

OAI21xp5_ASAP7_75t_SL g1622 ( 
.A1(n_1579),
.A2(n_1553),
.B(n_1515),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1583),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1572),
.B(n_1549),
.Y(n_1624)
);

AOI21xp5_ASAP7_75t_L g1625 ( 
.A1(n_1576),
.A2(n_1534),
.B(n_1543),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1572),
.B(n_1534),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1585),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1575),
.B(n_1534),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1585),
.Y(n_1629)
);

HB1xp67_ASAP7_75t_L g1630 ( 
.A(n_1567),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1570),
.Y(n_1631)
);

INVxp67_ASAP7_75t_L g1632 ( 
.A(n_1616),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1619),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1605),
.B(n_1561),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1605),
.B(n_1561),
.Y(n_1635)
);

AOI22xp33_ASAP7_75t_L g1636 ( 
.A1(n_1600),
.A2(n_1566),
.B1(n_1574),
.B2(n_1576),
.Y(n_1636)
);

OR2x2_ASAP7_75t_L g1637 ( 
.A(n_1597),
.B(n_1567),
.Y(n_1637)
);

INVx1_ASAP7_75t_SL g1638 ( 
.A(n_1616),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1601),
.B(n_1563),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_1618),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1618),
.Y(n_1641)
);

INVx1_ASAP7_75t_SL g1642 ( 
.A(n_1598),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1617),
.B(n_1563),
.Y(n_1643)
);

INVx1_ASAP7_75t_SL g1644 ( 
.A(n_1619),
.Y(n_1644)
);

AND2x4_ASAP7_75t_L g1645 ( 
.A(n_1607),
.B(n_1558),
.Y(n_1645)
);

AOI222xp33_ASAP7_75t_L g1646 ( 
.A1(n_1622),
.A2(n_1566),
.B1(n_1574),
.B2(n_1578),
.C1(n_1584),
.C2(n_1594),
.Y(n_1646)
);

OR2x2_ASAP7_75t_L g1647 ( 
.A(n_1614),
.B(n_1594),
.Y(n_1647)
);

NOR2xp33_ASAP7_75t_L g1648 ( 
.A(n_1599),
.B(n_1591),
.Y(n_1648)
);

OR2x2_ASAP7_75t_L g1649 ( 
.A(n_1614),
.B(n_1602),
.Y(n_1649)
);

NOR2xp33_ASAP7_75t_L g1650 ( 
.A(n_1617),
.B(n_1591),
.Y(n_1650)
);

INVxp67_ASAP7_75t_L g1651 ( 
.A(n_1621),
.Y(n_1651)
);

INVx1_ASAP7_75t_SL g1652 ( 
.A(n_1610),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1630),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1625),
.B(n_1566),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1603),
.Y(n_1655)
);

NOR2xp33_ASAP7_75t_L g1656 ( 
.A(n_1620),
.B(n_1569),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1633),
.Y(n_1657)
);

INVx2_ASAP7_75t_SL g1658 ( 
.A(n_1634),
.Y(n_1658)
);

AO22x1_ASAP7_75t_L g1659 ( 
.A1(n_1654),
.A2(n_1607),
.B1(n_1574),
.B2(n_1626),
.Y(n_1659)
);

NAND3xp33_ASAP7_75t_SL g1660 ( 
.A(n_1646),
.B(n_1628),
.C(n_1624),
.Y(n_1660)
);

OAI322xp33_ASAP7_75t_L g1661 ( 
.A1(n_1651),
.A2(n_1612),
.A3(n_1608),
.B1(n_1611),
.B2(n_1623),
.C1(n_1613),
.C2(n_1627),
.Y(n_1661)
);

OR2x2_ASAP7_75t_L g1662 ( 
.A(n_1639),
.B(n_1643),
.Y(n_1662)
);

NAND2x1p5_ASAP7_75t_L g1663 ( 
.A(n_1638),
.B(n_1535),
.Y(n_1663)
);

HB1xp67_ASAP7_75t_L g1664 ( 
.A(n_1644),
.Y(n_1664)
);

OAI22xp33_ASAP7_75t_L g1665 ( 
.A1(n_1632),
.A2(n_1535),
.B1(n_1557),
.B2(n_1510),
.Y(n_1665)
);

OR2x2_ASAP7_75t_L g1666 ( 
.A(n_1652),
.B(n_1609),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1633),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1644),
.Y(n_1668)
);

OR2x2_ASAP7_75t_L g1669 ( 
.A(n_1642),
.B(n_1609),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1634),
.B(n_1596),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1649),
.Y(n_1671)
);

AOI221xp5_ASAP7_75t_L g1672 ( 
.A1(n_1636),
.A2(n_1604),
.B1(n_1650),
.B2(n_1656),
.C(n_1648),
.Y(n_1672)
);

AOI22xp5_ASAP7_75t_L g1673 ( 
.A1(n_1653),
.A2(n_1640),
.B1(n_1641),
.B2(n_1578),
.Y(n_1673)
);

OAI211xp5_ASAP7_75t_L g1674 ( 
.A1(n_1653),
.A2(n_1543),
.B(n_1629),
.C(n_1631),
.Y(n_1674)
);

O2A1O1Ixp5_ASAP7_75t_L g1675 ( 
.A1(n_1640),
.A2(n_1603),
.B(n_1606),
.C(n_1584),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1664),
.B(n_1641),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1658),
.B(n_1635),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1671),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1670),
.B(n_1635),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1668),
.B(n_1637),
.Y(n_1680)
);

OAI221xp5_ASAP7_75t_L g1681 ( 
.A1(n_1672),
.A2(n_1637),
.B1(n_1649),
.B2(n_1655),
.C(n_1647),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1673),
.B(n_1655),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1673),
.B(n_1659),
.Y(n_1683)
);

NOR2xp33_ASAP7_75t_L g1684 ( 
.A(n_1662),
.B(n_1660),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1669),
.B(n_1666),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1657),
.B(n_1647),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1667),
.Y(n_1687)
);

OAI22xp5_ASAP7_75t_L g1688 ( 
.A1(n_1684),
.A2(n_1663),
.B1(n_1665),
.B2(n_1606),
.Y(n_1688)
);

AOI222xp33_ASAP7_75t_L g1689 ( 
.A1(n_1683),
.A2(n_1674),
.B1(n_1661),
.B2(n_1542),
.C1(n_1584),
.C2(n_1593),
.Y(n_1689)
);

OAI221xp5_ASAP7_75t_L g1690 ( 
.A1(n_1681),
.A2(n_1675),
.B1(n_1603),
.B2(n_1547),
.C(n_1546),
.Y(n_1690)
);

NOR3xp33_ASAP7_75t_L g1691 ( 
.A(n_1676),
.B(n_1661),
.C(n_1645),
.Y(n_1691)
);

NOR3xp33_ASAP7_75t_L g1692 ( 
.A(n_1676),
.B(n_1645),
.C(n_1595),
.Y(n_1692)
);

AOI21xp5_ASAP7_75t_L g1693 ( 
.A1(n_1680),
.A2(n_1685),
.B(n_1686),
.Y(n_1693)
);

AOI221x1_ASAP7_75t_L g1694 ( 
.A1(n_1687),
.A2(n_1678),
.B1(n_1682),
.B2(n_1686),
.C(n_1677),
.Y(n_1694)
);

NAND4xp75_ASAP7_75t_L g1695 ( 
.A(n_1679),
.B(n_1595),
.C(n_1546),
.D(n_1548),
.Y(n_1695)
);

OAI21xp33_ASAP7_75t_L g1696 ( 
.A1(n_1684),
.A2(n_1645),
.B(n_1606),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1694),
.Y(n_1697)
);

OAI21xp33_ASAP7_75t_SL g1698 ( 
.A1(n_1689),
.A2(n_1582),
.B(n_1577),
.Y(n_1698)
);

CKINVDCx5p33_ASAP7_75t_R g1699 ( 
.A(n_1693),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1691),
.B(n_1615),
.Y(n_1700)
);

OAI22xp33_ASAP7_75t_SL g1701 ( 
.A1(n_1690),
.A2(n_1547),
.B1(n_1615),
.B2(n_1548),
.Y(n_1701)
);

OR2x2_ASAP7_75t_L g1702 ( 
.A(n_1697),
.B(n_1699),
.Y(n_1702)
);

AOI21xp33_ASAP7_75t_SL g1703 ( 
.A1(n_1699),
.A2(n_1688),
.B(n_1696),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1700),
.B(n_1692),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1701),
.Y(n_1705)
);

NOR2x1_ASAP7_75t_L g1706 ( 
.A(n_1698),
.B(n_1695),
.Y(n_1706)
);

OR2x2_ASAP7_75t_L g1707 ( 
.A(n_1697),
.B(n_1569),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1707),
.Y(n_1708)
);

AOI22xp33_ASAP7_75t_L g1709 ( 
.A1(n_1705),
.A2(n_1535),
.B1(n_1615),
.B2(n_1542),
.Y(n_1709)
);

O2A1O1Ixp33_ASAP7_75t_L g1710 ( 
.A1(n_1703),
.A2(n_1542),
.B(n_1592),
.C(n_1564),
.Y(n_1710)
);

OAI21xp5_ASAP7_75t_L g1711 ( 
.A1(n_1706),
.A2(n_1546),
.B(n_1548),
.Y(n_1711)
);

OR2x2_ASAP7_75t_L g1712 ( 
.A(n_1702),
.B(n_1581),
.Y(n_1712)
);

NAND3xp33_ASAP7_75t_SL g1713 ( 
.A(n_1708),
.B(n_1704),
.C(n_1548),
.Y(n_1713)
);

NAND4xp25_ASAP7_75t_L g1714 ( 
.A(n_1709),
.B(n_1546),
.C(n_1592),
.D(n_1565),
.Y(n_1714)
);

NAND4xp25_ASAP7_75t_L g1715 ( 
.A(n_1712),
.B(n_1565),
.C(n_1592),
.D(n_1590),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1713),
.Y(n_1716)
);

A2O1A1Ixp33_ASAP7_75t_L g1717 ( 
.A1(n_1716),
.A2(n_1711),
.B(n_1710),
.C(n_1714),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1717),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1718),
.Y(n_1719)
);

O2A1O1Ixp33_ASAP7_75t_L g1720 ( 
.A1(n_1719),
.A2(n_1715),
.B(n_1564),
.C(n_1565),
.Y(n_1720)
);

AOI21xp33_ASAP7_75t_SL g1721 ( 
.A1(n_1720),
.A2(n_1564),
.B(n_1590),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1720),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1722),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1721),
.Y(n_1724)
);

AOI21xp5_ASAP7_75t_L g1725 ( 
.A1(n_1723),
.A2(n_1590),
.B(n_1577),
.Y(n_1725)
);

AND2x4_ASAP7_75t_L g1726 ( 
.A(n_1724),
.B(n_1570),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1726),
.Y(n_1727)
);

AOI22xp33_ASAP7_75t_SL g1728 ( 
.A1(n_1725),
.A2(n_1542),
.B1(n_1582),
.B2(n_1535),
.Y(n_1728)
);

AOI22xp33_ASAP7_75t_SL g1729 ( 
.A1(n_1727),
.A2(n_1535),
.B1(n_1532),
.B2(n_1536),
.Y(n_1729)
);

AOI211xp5_ASAP7_75t_L g1730 ( 
.A1(n_1729),
.A2(n_1728),
.B(n_1535),
.C(n_1532),
.Y(n_1730)
);


endmodule