module fake_jpeg_26531_n_299 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_299);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_299;

wire n_159;
wire n_117;
wire n_286;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_270;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_282;
wire n_258;
wire n_96;

BUFx3_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx6f_ASAP7_75t_SL g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_28),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_37),
.Y(n_46)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

CKINVDCx5p33_ASAP7_75t_R g37 ( 
.A(n_27),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_38),
.B(n_24),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_20),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_41),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx3_ASAP7_75t_SL g65 ( 
.A(n_40),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_20),
.B(n_0),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_53),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_35),
.A2(n_19),
.B1(n_26),
.B2(n_22),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_45),
.B(n_60),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_41),
.Y(n_48)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_48),
.B(n_50),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_28),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_38),
.A2(n_22),
.B1(n_26),
.B2(n_21),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_51),
.A2(n_52),
.B1(n_62),
.B2(n_43),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_43),
.A2(n_18),
.B1(n_24),
.B2(n_23),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_36),
.A2(n_43),
.B1(n_33),
.B2(n_29),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_56),
.A2(n_64),
.B1(n_36),
.B2(n_38),
.Y(n_95)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_58),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_25),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_47),
.Y(n_69)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_43),
.A2(n_29),
.B1(n_33),
.B2(n_34),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_36),
.A2(n_34),
.B1(n_31),
.B2(n_21),
.Y(n_64)
);

A2O1A1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_48),
.A2(n_35),
.B(n_31),
.C(n_38),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_68),
.A2(n_9),
.B(n_16),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_69),
.B(n_17),
.Y(n_125)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_70),
.B(n_76),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_25),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_71),
.B(n_79),
.Y(n_98)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_73),
.Y(n_104)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g115 ( 
.A(n_77),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_57),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_78),
.Y(n_100)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_80),
.B(n_83),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_82),
.B(n_24),
.Y(n_113)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_46),
.B(n_25),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_84),
.B(n_89),
.Y(n_123)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_85),
.B(n_87),
.Y(n_103)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_86),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_50),
.B(n_25),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_49),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_90),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_47),
.B(n_30),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_30),
.Y(n_108)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_93),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_45),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_94),
.Y(n_102)
);

O2A1O1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_95),
.A2(n_65),
.B(n_75),
.C(n_93),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_44),
.B(n_23),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_96),
.B(n_97),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_53),
.B(n_23),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_85),
.A2(n_59),
.B1(n_54),
.B2(n_52),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_101),
.A2(n_70),
.B1(n_75),
.B2(n_88),
.Y(n_128)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_72),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_105),
.B(n_107),
.Y(n_126)
);

BUFx5_ASAP7_75t_L g107 ( 
.A(n_73),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_108),
.B(n_125),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_69),
.B(n_42),
.C(n_30),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_110),
.B(n_121),
.C(n_42),
.Y(n_138)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_72),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_111),
.B(n_78),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_76),
.A2(n_54),
.B1(n_55),
.B2(n_65),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_112),
.A2(n_92),
.B1(n_67),
.B2(n_83),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_113),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_91),
.B(n_30),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_114),
.B(n_120),
.Y(n_148)
);

OAI22x1_ASAP7_75t_L g151 ( 
.A1(n_116),
.A2(n_37),
.B1(n_42),
.B2(n_80),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_74),
.B(n_66),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_66),
.B(n_42),
.C(n_32),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_124),
.A2(n_88),
.B(n_102),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_127),
.A2(n_125),
.B(n_121),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_128),
.A2(n_134),
.B1(n_135),
.B2(n_147),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_100),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_130),
.Y(n_167)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_115),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_131),
.B(n_136),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_106),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_132),
.B(n_133),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_120),
.B(n_74),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_99),
.A2(n_88),
.B1(n_79),
.B2(n_67),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_100),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_112),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_137),
.B(n_142),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_138),
.B(n_149),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_119),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_139),
.B(n_141),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_103),
.B(n_68),
.Y(n_140)
);

BUFx24_ASAP7_75t_SL g168 ( 
.A(n_140),
.Y(n_168)
);

BUFx5_ASAP7_75t_L g141 ( 
.A(n_115),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_99),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_98),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_143),
.B(n_144),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_123),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_145),
.B(n_153),
.Y(n_173)
);

AO21x1_ASAP7_75t_L g146 ( 
.A1(n_124),
.A2(n_37),
.B(n_42),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_146),
.A2(n_151),
.B(n_154),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_113),
.A2(n_90),
.B1(n_81),
.B2(n_77),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_110),
.B(n_114),
.Y(n_149)
);

OA22x2_ASAP7_75t_L g150 ( 
.A1(n_116),
.A2(n_37),
.B1(n_86),
.B2(n_81),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_150),
.B(n_115),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_113),
.A2(n_42),
.B1(n_17),
.B2(n_32),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_152),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_179)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_119),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_102),
.A2(n_32),
.B(n_17),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_125),
.B(n_7),
.C(n_15),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_155),
.B(n_12),
.C(n_15),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_156),
.A2(n_109),
.B1(n_117),
.B2(n_122),
.Y(n_165)
);

AND2x4_ASAP7_75t_L g157 ( 
.A(n_151),
.B(n_103),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_157),
.A2(n_162),
.B(n_176),
.Y(n_189)
);

NAND3xp33_ASAP7_75t_L g159 ( 
.A(n_148),
.B(n_108),
.C(n_118),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_159),
.B(n_165),
.Y(n_191)
);

AO21x1_ASAP7_75t_L g211 ( 
.A1(n_160),
.A2(n_131),
.B(n_141),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_127),
.A2(n_118),
.B(n_101),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_137),
.A2(n_105),
.B1(n_111),
.B2(n_117),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_163),
.A2(n_175),
.B1(n_182),
.B2(n_185),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_166),
.B(n_155),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_148),
.A2(n_122),
.B1(n_104),
.B2(n_109),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_149),
.B(n_104),
.C(n_115),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_177),
.B(n_184),
.C(n_152),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_130),
.B(n_107),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_178),
.B(n_183),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_179),
.A2(n_181),
.B(n_154),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_138),
.B(n_7),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_180),
.B(n_186),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_129),
.A2(n_1),
.B(n_3),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_147),
.A2(n_8),
.B1(n_4),
.B2(n_5),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_136),
.B(n_143),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_142),
.B(n_8),
.C(n_4),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_150),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_134),
.B(n_5),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_150),
.A2(n_6),
.B1(n_11),
.B2(n_13),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_187),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_157),
.B(n_150),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_188),
.A2(n_199),
.B(n_212),
.Y(n_215)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_170),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_190),
.B(n_207),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_169),
.B(n_160),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_194),
.B(n_169),
.C(n_162),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_158),
.B(n_139),
.Y(n_195)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_195),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_SL g232 ( 
.A(n_196),
.B(n_198),
.C(n_211),
.Y(n_232)
);

BUFx2_ASAP7_75t_L g197 ( 
.A(n_171),
.Y(n_197)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_197),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_176),
.A2(n_146),
.B(n_144),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_167),
.B(n_126),
.Y(n_201)
);

CKINVDCx14_ASAP7_75t_R g229 ( 
.A(n_201),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_167),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_202),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_203),
.B(n_177),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_158),
.B(n_153),
.Y(n_204)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_204),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_173),
.B(n_135),
.Y(n_206)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_206),
.Y(n_227)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_163),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_172),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_208),
.B(n_210),
.Y(n_218)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_175),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_209),
.B(n_164),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_161),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_176),
.A2(n_6),
.B(n_11),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_157),
.Y(n_213)
);

CKINVDCx14_ASAP7_75t_R g230 ( 
.A(n_213),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_192),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_216),
.B(n_235),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_207),
.A2(n_164),
.B1(n_157),
.B2(n_187),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_219),
.A2(n_200),
.B1(n_191),
.B2(n_182),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_220),
.B(n_193),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_209),
.A2(n_205),
.B1(n_200),
.B2(n_188),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_221),
.A2(n_213),
.B1(n_211),
.B2(n_189),
.Y(n_243)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_223),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_224),
.B(n_233),
.C(n_234),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_195),
.B(n_186),
.Y(n_225)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_225),
.Y(n_241)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_204),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_228),
.B(n_188),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_194),
.B(n_180),
.C(n_174),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_193),
.B(n_174),
.C(n_184),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_206),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_231),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_237),
.B(n_247),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_238),
.A2(n_243),
.B1(n_219),
.B2(n_185),
.Y(n_262)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_242),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_214),
.A2(n_230),
.B(n_221),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_244),
.A2(n_248),
.B(n_215),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_231),
.B(n_190),
.Y(n_245)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_245),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_218),
.B(n_205),
.Y(n_246)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_246),
.Y(n_260)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_214),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_215),
.A2(n_189),
.B(n_199),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_249),
.B(n_239),
.Y(n_261)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_223),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_250),
.B(n_251),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_217),
.B(n_181),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_224),
.B(n_203),
.C(n_198),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_252),
.B(n_220),
.C(n_233),
.Y(n_259)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_242),
.Y(n_254)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_254),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_256),
.B(n_261),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_259),
.B(n_239),
.C(n_252),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_263),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_243),
.A2(n_232),
.B1(n_227),
.B2(n_229),
.Y(n_263)
);

NAND4xp25_ASAP7_75t_L g264 ( 
.A(n_237),
.B(n_232),
.C(n_225),
.D(n_197),
.Y(n_264)
);

NOR2xp67_ASAP7_75t_SL g276 ( 
.A(n_264),
.B(n_248),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_251),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_265),
.B(n_227),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_266),
.B(n_267),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_261),
.B(n_249),
.C(n_234),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_257),
.B(n_222),
.C(n_240),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_268),
.B(n_270),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_259),
.B(n_222),
.C(n_244),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_260),
.B(n_241),
.C(n_247),
.Y(n_271)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_271),
.Y(n_280)
);

NAND2xp33_ASAP7_75t_SL g284 ( 
.A(n_272),
.B(n_228),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_263),
.B(n_241),
.C(n_250),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_274),
.B(n_273),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_276),
.A2(n_256),
.B(n_265),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_277),
.A2(n_284),
.B(n_226),
.Y(n_286)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_278),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_275),
.B(n_255),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_282),
.B(n_269),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_272),
.A2(n_262),
.B1(n_258),
.B2(n_217),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_283),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_286),
.B(n_290),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_287),
.B(n_288),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_282),
.B(n_253),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_279),
.B(n_168),
.Y(n_290)
);

AOI322xp5_ASAP7_75t_L g291 ( 
.A1(n_285),
.A2(n_281),
.A3(n_280),
.B1(n_278),
.B2(n_284),
.C1(n_236),
.C2(n_196),
.Y(n_291)
);

NOR4xp25_ASAP7_75t_L g295 ( 
.A(n_291),
.B(n_293),
.C(n_11),
.D(n_15),
.Y(n_295)
);

AOI322xp5_ASAP7_75t_L g293 ( 
.A1(n_285),
.A2(n_236),
.A3(n_226),
.B1(n_212),
.B2(n_179),
.C1(n_166),
.C2(n_16),
.Y(n_293)
);

OR2x2_ASAP7_75t_L g297 ( 
.A(n_295),
.B(n_296),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_294),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_297),
.A2(n_292),
.B(n_289),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_298),
.B(n_16),
.Y(n_299)
);


endmodule