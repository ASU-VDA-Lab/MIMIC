module fake_jpeg_30256_n_100 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_100);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_100;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

INVx3_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_9),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx14_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g18 ( 
.A(n_3),
.B(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_23),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_18),
.B(n_0),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_26),
.B(n_32),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

CKINVDCx6p67_ASAP7_75t_R g45 ( 
.A(n_30),
.Y(n_45)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

INVx4_ASAP7_75t_SL g44 ( 
.A(n_31),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_0),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_34),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g34 ( 
.A(n_11),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_16),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_24),
.A2(n_29),
.B1(n_30),
.B2(n_33),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_40),
.A2(n_30),
.B1(n_31),
.B2(n_13),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_34),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_42),
.B(n_46),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_28),
.B(n_17),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_48),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_17),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_49),
.B(n_55),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_47),
.A2(n_27),
.B1(n_25),
.B2(n_35),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_50),
.A2(n_53),
.B1(n_57),
.B2(n_44),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_13),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_56),
.Y(n_69)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_14),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_14),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_38),
.A2(n_15),
.B1(n_19),
.B2(n_20),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_45),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_60),
.B(n_45),
.Y(n_63)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_15),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_62),
.B(n_20),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_67),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_66),
.A2(n_53),
.B1(n_52),
.B2(n_54),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_19),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_68),
.A2(n_40),
.B(n_61),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_1),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_2),
.Y(n_79)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_72),
.Y(n_73)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_73),
.Y(n_80)
);

HAxp5_ASAP7_75t_SL g74 ( 
.A(n_69),
.B(n_51),
.CON(n_74),
.SN(n_74)
);

NOR3xp33_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_68),
.C(n_66),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_65),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_75),
.B(n_76),
.Y(n_83)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_78),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_79),
.A2(n_64),
.B(n_65),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_84),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_82),
.B(n_77),
.C(n_74),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_88),
.C(n_71),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_83),
.A2(n_76),
.B1(n_57),
.B2(n_73),
.Y(n_86)
);

AOI322xp5_ASAP7_75t_L g91 ( 
.A1(n_86),
.A2(n_59),
.A3(n_71),
.B1(n_37),
.B2(n_39),
.C1(n_38),
.C2(n_5),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_80),
.B(n_78),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_87),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_84),
.B(n_50),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_91),
.B(n_89),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_92),
.A2(n_87),
.B(n_39),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_93),
.B(n_90),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_94),
.B(n_5),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_95),
.B(n_96),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_97),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_6),
.C(n_95),
.Y(n_99)
);

BUFx24_ASAP7_75t_SL g100 ( 
.A(n_99),
.Y(n_100)
);


endmodule