module fake_jpeg_2282_n_710 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_710);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_710;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_696;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_686;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_699;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_701;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_688;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_689;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_704;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_698;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_694;
wire n_692;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_697;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_691;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_709;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_708;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_690;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_693;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_703;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_695;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_702;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_687;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_707;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_705;
wire n_665;
wire n_706;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_700;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx24_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_18),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_12),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_14),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx4f_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_19),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

BUFx10_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

INVx11_ASAP7_75t_SL g53 ( 
.A(n_4),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_14),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_4),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_16),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_0),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_9),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_62),
.B(n_63),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_10),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_10),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_64),
.B(n_70),
.Y(n_166)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g146 ( 
.A(n_65),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_41),
.A2(n_8),
.B(n_17),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g175 ( 
.A(n_66),
.B(n_81),
.Y(n_175)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_67),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g149 ( 
.A(n_68),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_69),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_43),
.B(n_46),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g168 ( 
.A(n_71),
.Y(n_168)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_72),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_46),
.B(n_8),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_73),
.B(n_77),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_74),
.Y(n_155)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g207 ( 
.A(n_75),
.Y(n_207)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_76),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_57),
.B(n_18),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_26),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_78),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_34),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_79),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_34),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_80),
.Y(n_196)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_57),
.B(n_18),
.Y(n_81)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_23),
.Y(n_82)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_82),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_34),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_83),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_22),
.B(n_16),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g184 ( 
.A(n_84),
.B(n_97),
.Y(n_184)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_85),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_86),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_23),
.Y(n_87)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_87),
.Y(n_177)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

INVx2_ASAP7_75t_SL g205 ( 
.A(n_88),
.Y(n_205)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_89),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

INVx6_ASAP7_75t_L g190 ( 
.A(n_90),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

INVx8_ASAP7_75t_L g161 ( 
.A(n_91),
.Y(n_161)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

INVxp67_ASAP7_75t_SL g218 ( 
.A(n_92),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

INVx8_ASAP7_75t_L g208 ( 
.A(n_93),
.Y(n_208)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_94),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_95),
.Y(n_197)
);

BUFx4f_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_96),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_22),
.B(n_15),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_98),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_37),
.Y(n_99)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_99),
.Y(n_140)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_100),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_48),
.Y(n_101)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_101),
.Y(n_152)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_102),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_103),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_56),
.B(n_15),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_104),
.B(n_120),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_50),
.Y(n_105)
);

INVx5_ASAP7_75t_L g212 ( 
.A(n_105),
.Y(n_212)
);

INVx13_ASAP7_75t_L g106 ( 
.A(n_23),
.Y(n_106)
);

INVx6_ASAP7_75t_SL g156 ( 
.A(n_106),
.Y(n_156)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_55),
.Y(n_107)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_107),
.Y(n_214)
);

BUFx5_ASAP7_75t_L g108 ( 
.A(n_23),
.Y(n_108)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_108),
.Y(n_206)
);

BUFx12_ASAP7_75t_L g109 ( 
.A(n_21),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g198 ( 
.A(n_109),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_31),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_110),
.Y(n_158)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_31),
.Y(n_111)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_111),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_55),
.Y(n_112)
);

INVx5_ASAP7_75t_L g220 ( 
.A(n_112),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_30),
.B(n_15),
.Y(n_113)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_113),
.Y(n_147)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_33),
.Y(n_114)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_114),
.Y(n_173)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_33),
.Y(n_115)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_115),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_55),
.Y(n_116)
);

INVx5_ASAP7_75t_L g221 ( 
.A(n_116),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_58),
.Y(n_117)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_117),
.Y(n_170)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_25),
.Y(n_118)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_118),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_58),
.Y(n_119)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_119),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_30),
.B(n_39),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_58),
.Y(n_121)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_121),
.Y(n_174)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_47),
.Y(n_122)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_122),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_27),
.Y(n_123)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_123),
.Y(n_178)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_25),
.Y(n_124)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_124),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_27),
.Y(n_125)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_125),
.Y(n_187)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_25),
.Y(n_126)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_126),
.Y(n_211)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_27),
.Y(n_127)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_127),
.Y(n_193)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_33),
.Y(n_128)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_128),
.Y(n_160)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_41),
.Y(n_129)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_129),
.Y(n_200)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_20),
.Y(n_130)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_130),
.Y(n_163)
);

BUFx4f_ASAP7_75t_L g131 ( 
.A(n_49),
.Y(n_131)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_131),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_28),
.Y(n_132)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_132),
.Y(n_204)
);

BUFx12f_ASAP7_75t_SL g133 ( 
.A(n_21),
.Y(n_133)
);

HAxp5_ASAP7_75t_SL g209 ( 
.A(n_133),
.B(n_52),
.CON(n_209),
.SN(n_209)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_88),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_136),
.B(n_141),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_123),
.A2(n_49),
.B1(n_41),
.B2(n_28),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_139),
.A2(n_154),
.B1(n_199),
.B2(n_202),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_92),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_96),
.A2(n_49),
.B1(n_61),
.B2(n_54),
.Y(n_151)
);

OA22x2_ASAP7_75t_L g284 ( 
.A1(n_151),
.A2(n_157),
.B1(n_189),
.B2(n_191),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_125),
.A2(n_132),
.B1(n_86),
.B2(n_105),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_96),
.A2(n_61),
.B1(n_41),
.B2(n_38),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_69),
.A2(n_95),
.B1(n_74),
.B2(n_79),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_159),
.A2(n_180),
.B1(n_181),
.B2(n_183),
.Y(n_238)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_131),
.Y(n_164)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_164),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_78),
.A2(n_45),
.B1(n_28),
.B2(n_38),
.Y(n_180)
);

OAI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_80),
.A2(n_38),
.B1(n_40),
.B2(n_39),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_131),
.Y(n_182)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_182),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_81),
.A2(n_45),
.B1(n_36),
.B2(n_40),
.Y(n_183)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_118),
.Y(n_188)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_188),
.Y(n_265)
);

OA22x2_ASAP7_75t_L g189 ( 
.A1(n_133),
.A2(n_45),
.B1(n_59),
.B2(n_20),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_124),
.A2(n_59),
.B1(n_29),
.B2(n_32),
.Y(n_191)
);

INVx6_ASAP7_75t_SL g195 ( 
.A(n_106),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_195),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_83),
.A2(n_29),
.B1(n_32),
.B2(n_36),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_90),
.A2(n_52),
.B1(n_21),
.B2(n_35),
.Y(n_202)
);

OR2x2_ASAP7_75t_L g283 ( 
.A(n_209),
.B(n_210),
.Y(n_283)
);

HAxp5_ASAP7_75t_SL g210 ( 
.A(n_109),
.B(n_52),
.CON(n_210),
.SN(n_210)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_126),
.Y(n_213)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_213),
.Y(n_266)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_72),
.Y(n_216)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_216),
.Y(n_242)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_114),
.Y(n_217)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_217),
.Y(n_273)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_75),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_219),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_127),
.A2(n_52),
.B1(n_21),
.B2(n_60),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_222),
.A2(n_121),
.B1(n_119),
.B2(n_117),
.Y(n_251)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_91),
.Y(n_224)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_224),
.Y(n_268)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_67),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_225),
.Y(n_281)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_65),
.Y(n_226)
);

BUFx2_ASAP7_75t_L g277 ( 
.A(n_226),
.Y(n_277)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_82),
.Y(n_227)
);

INVx4_ASAP7_75t_L g290 ( 
.A(n_227),
.Y(n_290)
);

INVx8_ASAP7_75t_L g228 ( 
.A(n_156),
.Y(n_228)
);

BUFx2_ASAP7_75t_L g363 ( 
.A(n_228),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_138),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_229),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_137),
.B(n_203),
.Y(n_230)
);

CKINVDCx14_ASAP7_75t_R g337 ( 
.A(n_230),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_147),
.B(n_153),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_232),
.B(n_233),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_166),
.B(n_68),
.Y(n_233)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_135),
.Y(n_235)
);

INVx4_ASAP7_75t_L g317 ( 
.A(n_235),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_158),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_236),
.B(n_241),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_138),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_237),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_223),
.B(n_13),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_239),
.B(n_276),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_209),
.A2(n_89),
.B1(n_76),
.B2(n_99),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_240),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_184),
.B(n_215),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_158),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_245),
.B(n_246),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_184),
.B(n_71),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_140),
.Y(n_247)
);

INVx5_ASAP7_75t_L g318 ( 
.A(n_247),
.Y(n_318)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_193),
.Y(n_248)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_248),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_142),
.B(n_122),
.Y(n_249)
);

AND2x2_ASAP7_75t_SL g324 ( 
.A(n_249),
.B(n_252),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_223),
.B(n_103),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_250),
.B(n_309),
.C(n_201),
.Y(n_354)
);

OA22x2_ASAP7_75t_L g336 ( 
.A1(n_251),
.A2(n_307),
.B1(n_285),
.B2(n_256),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_145),
.B(n_85),
.Y(n_252)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_165),
.Y(n_253)
);

INVx4_ASAP7_75t_L g345 ( 
.A(n_253),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_155),
.Y(n_254)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_254),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_181),
.A2(n_116),
.B1(n_112),
.B2(n_101),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_256),
.B(n_282),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_146),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_257),
.B(n_267),
.Y(n_349)
);

INVx5_ASAP7_75t_L g258 ( 
.A(n_161),
.Y(n_258)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_258),
.Y(n_358)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_205),
.A2(n_107),
.B1(n_102),
.B2(n_93),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g316 ( 
.A1(n_259),
.A2(n_280),
.B1(n_294),
.B2(n_177),
.Y(n_316)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_214),
.Y(n_260)
);

INVx2_ASAP7_75t_SL g315 ( 
.A(n_260),
.Y(n_315)
);

BUFx12_ASAP7_75t_L g261 ( 
.A(n_198),
.Y(n_261)
);

INVx13_ASAP7_75t_L g326 ( 
.A(n_261),
.Y(n_326)
);

BUFx3_ASAP7_75t_L g262 ( 
.A(n_149),
.Y(n_262)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_262),
.Y(n_347)
);

INVx5_ASAP7_75t_L g263 ( 
.A(n_161),
.Y(n_263)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_263),
.Y(n_310)
);

INVx5_ASAP7_75t_L g264 ( 
.A(n_208),
.Y(n_264)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_264),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_163),
.B(n_107),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_146),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_269),
.B(n_296),
.Y(n_355)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_186),
.Y(n_271)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_271),
.Y(n_321)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_200),
.Y(n_272)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_272),
.Y(n_330)
);

INVx5_ASAP7_75t_L g274 ( 
.A(n_208),
.Y(n_274)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_274),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_175),
.A2(n_102),
.B1(n_109),
.B2(n_52),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_275),
.A2(n_210),
.B1(n_189),
.B2(n_206),
.Y(n_323)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_144),
.Y(n_276)
);

BUFx2_ASAP7_75t_L g278 ( 
.A(n_205),
.Y(n_278)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_278),
.Y(n_333)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_143),
.Y(n_279)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_279),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_218),
.A2(n_60),
.B1(n_35),
.B2(n_24),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_175),
.A2(n_21),
.B1(n_24),
.B2(n_35),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_149),
.A2(n_24),
.B1(n_14),
.B2(n_13),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_285),
.B(n_306),
.Y(n_351)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_178),
.Y(n_286)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_286),
.Y(n_339)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_207),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_287),
.B(n_298),
.Y(n_334)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_170),
.Y(n_288)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_288),
.Y(n_350)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_162),
.Y(n_289)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_289),
.Y(n_364)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_187),
.Y(n_291)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_291),
.Y(n_369)
);

AOI22xp33_ASAP7_75t_L g292 ( 
.A1(n_199),
.A2(n_13),
.B1(n_12),
.B2(n_11),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_292),
.A2(n_303),
.B1(n_139),
.B2(n_191),
.Y(n_312)
);

INVx4_ASAP7_75t_L g293 ( 
.A(n_179),
.Y(n_293)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_293),
.Y(n_372)
);

AOI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_218),
.A2(n_168),
.B1(n_207),
.B2(n_169),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_155),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_295),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_167),
.A2(n_12),
.B(n_11),
.Y(n_296)
);

INVx8_ASAP7_75t_L g297 ( 
.A(n_198),
.Y(n_297)
);

INVx13_ASAP7_75t_L g341 ( 
.A(n_297),
.Y(n_341)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_176),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_168),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_299),
.B(n_300),
.Y(n_343)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_194),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_150),
.B(n_0),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_301),
.B(n_305),
.Y(n_371)
);

INVx6_ASAP7_75t_L g302 ( 
.A(n_185),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_302),
.Y(n_365)
);

AOI22xp33_ASAP7_75t_L g303 ( 
.A1(n_154),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_303)
);

BUFx2_ASAP7_75t_L g304 ( 
.A(n_151),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_304),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_160),
.B(n_1),
.Y(n_305)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_211),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_189),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_148),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_308),
.B(n_3),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_173),
.B(n_1),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_L g402 ( 
.A1(n_312),
.A2(n_274),
.B1(n_264),
.B2(n_258),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_238),
.A2(n_157),
.B1(n_190),
.B2(n_134),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_314),
.A2(n_361),
.B1(n_368),
.B2(n_263),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g386 ( 
.A(n_316),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_238),
.A2(n_204),
.B1(n_174),
.B2(n_171),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_322),
.A2(n_323),
.B1(n_342),
.B2(n_249),
.Y(n_373)
);

INVx6_ASAP7_75t_SL g332 ( 
.A(n_270),
.Y(n_332)
);

BUFx2_ASAP7_75t_SL g394 ( 
.A(n_332),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_336),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_251),
.A2(n_134),
.B1(n_201),
.B2(n_196),
.Y(n_342)
);

AOI22xp33_ASAP7_75t_SL g344 ( 
.A1(n_304),
.A2(n_221),
.B1(n_220),
.B2(n_212),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_344),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_250),
.B(n_172),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_348),
.B(n_356),
.Y(n_384)
);

AND2x6_ASAP7_75t_L g352 ( 
.A(n_283),
.B(n_197),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_352),
.B(n_297),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_354),
.B(n_357),
.Y(n_375)
);

A2O1A1Ixp33_ASAP7_75t_L g356 ( 
.A1(n_283),
.A2(n_152),
.B(n_192),
.C(n_185),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_309),
.B(n_192),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_231),
.B(n_196),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_359),
.B(n_278),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_360),
.Y(n_421)
);

AOI22xp33_ASAP7_75t_L g361 ( 
.A1(n_243),
.A2(n_284),
.B1(n_307),
.B2(n_255),
.Y(n_361)
);

INVx13_ASAP7_75t_L g362 ( 
.A(n_228),
.Y(n_362)
);

INVx5_ASAP7_75t_L g406 ( 
.A(n_362),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_309),
.B(n_3),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_366),
.B(n_357),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_243),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_368)
);

AOI22xp33_ASAP7_75t_SL g370 ( 
.A1(n_275),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_370),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_373),
.B(n_407),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_314),
.A2(n_284),
.B1(n_282),
.B2(n_252),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_374),
.A2(n_387),
.B1(n_402),
.B2(n_403),
.Y(n_427)
);

OR2x2_ASAP7_75t_L g376 ( 
.A(n_323),
.B(n_284),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_L g423 ( 
.A1(n_376),
.A2(n_410),
.B(n_353),
.Y(n_423)
);

INVx3_ASAP7_75t_L g377 ( 
.A(n_317),
.Y(n_377)
);

INVx2_ASAP7_75t_SL g440 ( 
.A(n_377),
.Y(n_440)
);

OAI21xp5_ASAP7_75t_L g378 ( 
.A1(n_355),
.A2(n_284),
.B(n_244),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_SL g438 ( 
.A1(n_378),
.A2(n_379),
.B(n_343),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_L g379 ( 
.A1(n_353),
.A2(n_273),
.B(n_266),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_327),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g451 ( 
.A(n_380),
.Y(n_451)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_339),
.Y(n_381)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_381),
.Y(n_429)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_339),
.Y(n_382)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_382),
.Y(n_434)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_315),
.Y(n_383)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_383),
.Y(n_437)
);

OAI22xp33_ASAP7_75t_SL g385 ( 
.A1(n_368),
.A2(n_271),
.B1(n_235),
.B2(n_277),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_385),
.A2(n_392),
.B1(n_396),
.B2(n_337),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_322),
.A2(n_249),
.B1(n_252),
.B2(n_291),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_332),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_388),
.B(n_390),
.Y(n_428)
);

OAI32xp33_ASAP7_75t_L g389 ( 
.A1(n_313),
.A2(n_265),
.A3(n_272),
.B1(n_248),
.B2(n_230),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_389),
.B(n_391),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_393),
.B(n_397),
.Y(n_439)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_369),
.Y(n_395)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_395),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_346),
.A2(n_302),
.B1(n_286),
.B2(n_268),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_319),
.B(n_306),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_319),
.B(n_300),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_398),
.B(n_415),
.Y(n_446)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_369),
.Y(n_399)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_399),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_354),
.B(n_230),
.C(n_242),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_400),
.B(n_414),
.C(n_321),
.Y(n_452)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_330),
.Y(n_401)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_401),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_346),
.A2(n_298),
.B1(n_277),
.B2(n_237),
.Y(n_403)
);

FAx1_ASAP7_75t_SL g405 ( 
.A(n_348),
.B(n_281),
.CI(n_234),
.CON(n_405),
.SN(n_405)
);

OAI32xp33_ASAP7_75t_L g426 ( 
.A1(n_405),
.A2(n_351),
.A3(n_328),
.B1(n_352),
.B2(n_324),
.Y(n_426)
);

AO22x2_ASAP7_75t_L g407 ( 
.A1(n_312),
.A2(n_289),
.B1(n_234),
.B2(n_279),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_371),
.B(n_290),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_409),
.B(n_412),
.Y(n_433)
);

OR2x2_ASAP7_75t_L g410 ( 
.A(n_329),
.B(n_290),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_346),
.A2(n_295),
.B1(n_254),
.B2(n_229),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_411),
.A2(n_416),
.B1(n_419),
.B2(n_363),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_371),
.B(n_366),
.Y(n_412)
);

INVx3_ASAP7_75t_L g413 ( 
.A(n_317),
.Y(n_413)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_413),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_324),
.B(n_247),
.C(n_260),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_363),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_356),
.A2(n_293),
.B1(n_262),
.B2(n_253),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_359),
.B(n_4),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_417),
.B(n_418),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_349),
.B(n_5),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_342),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_330),
.Y(n_420)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_420),
.Y(n_462)
);

OAI21xp5_ASAP7_75t_SL g492 ( 
.A1(n_423),
.A2(n_438),
.B(n_445),
.Y(n_492)
);

INVx1_ASAP7_75t_SL g477 ( 
.A(n_424),
.Y(n_477)
);

INVxp67_ASAP7_75t_L g466 ( 
.A(n_426),
.Y(n_466)
);

NOR2x1_ASAP7_75t_L g430 ( 
.A(n_378),
.B(n_351),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_SL g475 ( 
.A1(n_430),
.A2(n_405),
.B(n_389),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_404),
.A2(n_351),
.B1(n_367),
.B2(n_336),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_431),
.A2(n_449),
.B1(n_407),
.B2(n_408),
.Y(n_480)
);

AOI21xp5_ASAP7_75t_SL g432 ( 
.A1(n_404),
.A2(n_367),
.B(n_343),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_L g486 ( 
.A1(n_432),
.A2(n_383),
.B(n_333),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_406),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_435),
.B(n_388),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_436),
.A2(n_464),
.B1(n_396),
.B2(n_415),
.Y(n_465)
);

NAND2x1_ASAP7_75t_L g441 ( 
.A(n_376),
.B(n_324),
.Y(n_441)
);

XNOR2x1_ASAP7_75t_L g481 ( 
.A(n_441),
.B(n_452),
.Y(n_481)
);

NOR2x1_ASAP7_75t_R g443 ( 
.A(n_405),
.B(n_324),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g499 ( 
.A(n_443),
.Y(n_499)
);

OAI21xp5_ASAP7_75t_L g445 ( 
.A1(n_384),
.A2(n_334),
.B(n_363),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_374),
.A2(n_336),
.B1(n_365),
.B2(n_325),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_391),
.B(n_365),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_454),
.B(n_460),
.Y(n_487)
);

AOI22xp33_ASAP7_75t_SL g455 ( 
.A1(n_386),
.A2(n_358),
.B1(n_325),
.B2(n_315),
.Y(n_455)
);

OAI21xp33_ASAP7_75t_SL g490 ( 
.A1(n_455),
.A2(n_358),
.B(n_347),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_375),
.B(n_400),
.C(n_414),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_456),
.B(n_457),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_375),
.B(n_334),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_L g458 ( 
.A1(n_379),
.A2(n_321),
.B(n_315),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_L g483 ( 
.A1(n_458),
.A2(n_382),
.B(n_395),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_412),
.B(n_336),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_459),
.B(n_456),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_417),
.B(n_331),
.Y(n_460)
);

AOI21xp5_ASAP7_75t_L g461 ( 
.A1(n_408),
.A2(n_345),
.B(n_372),
.Y(n_461)
);

AOI21xp5_ASAP7_75t_L g497 ( 
.A1(n_461),
.A2(n_345),
.B(n_326),
.Y(n_497)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_381),
.Y(n_463)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_463),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_373),
.A2(n_320),
.B1(n_331),
.B2(n_310),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_465),
.B(n_480),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_L g467 ( 
.A1(n_453),
.A2(n_416),
.B1(n_411),
.B2(n_419),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_467),
.A2(n_468),
.B1(n_490),
.B2(n_495),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_453),
.A2(n_386),
.B1(n_407),
.B2(n_403),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_469),
.B(n_472),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_SL g471 ( 
.A(n_433),
.B(n_409),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_471),
.B(n_482),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_460),
.B(n_421),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_429),
.Y(n_473)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_473),
.Y(n_524)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_429),
.Y(n_474)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_474),
.Y(n_506)
);

OAI21xp5_ASAP7_75t_SL g518 ( 
.A1(n_475),
.A2(n_486),
.B(n_497),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_453),
.A2(n_422),
.B1(n_410),
.B2(n_407),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_SL g519 ( 
.A1(n_476),
.A2(n_485),
.B1(n_496),
.B2(n_501),
.Y(n_519)
);

OAI32xp33_ASAP7_75t_L g478 ( 
.A1(n_425),
.A2(n_387),
.A3(n_421),
.B1(n_422),
.B2(n_401),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_478),
.B(n_479),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_433),
.B(n_418),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_SL g482 ( 
.A(n_447),
.B(n_420),
.Y(n_482)
);

INVx1_ASAP7_75t_SL g525 ( 
.A(n_483),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_453),
.A2(n_407),
.B1(n_394),
.B2(n_399),
.Y(n_485)
);

CKINVDCx16_ASAP7_75t_R g488 ( 
.A(n_446),
.Y(n_488)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_488),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_454),
.B(n_413),
.Y(n_489)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_489),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_428),
.B(n_446),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_SL g504 ( 
.A(n_491),
.B(n_500),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_SL g517 ( 
.A(n_493),
.B(n_441),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_447),
.B(n_377),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_494),
.B(n_498),
.Y(n_536)
);

OAI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_425),
.A2(n_340),
.B1(n_380),
.B2(n_310),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_449),
.A2(n_427),
.B1(n_436),
.B2(n_459),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_428),
.B(n_320),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_SL g500 ( 
.A(n_439),
.B(n_406),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_427),
.A2(n_340),
.B1(n_380),
.B2(n_338),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_439),
.B(n_438),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_502),
.B(n_503),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_458),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_SL g508 ( 
.A(n_502),
.B(n_457),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_508),
.B(n_526),
.Y(n_562)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_489),
.Y(n_511)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_511),
.Y(n_545)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_473),
.Y(n_513)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_513),
.Y(n_546)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_477),
.A2(n_464),
.B1(n_423),
.B2(n_445),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_SL g555 ( 
.A1(n_514),
.A2(n_516),
.B1(n_522),
.B2(n_534),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_484),
.B(n_452),
.C(n_441),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_515),
.B(n_520),
.C(n_538),
.Y(n_543)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_477),
.A2(n_424),
.B1(n_431),
.B2(n_461),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g551 ( 
.A(n_517),
.B(n_529),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_484),
.B(n_443),
.C(n_430),
.Y(n_520)
);

OAI22xp5_ASAP7_75t_SL g521 ( 
.A1(n_496),
.A2(n_443),
.B1(n_455),
.B2(n_426),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g561 ( 
.A1(n_521),
.A2(n_542),
.B1(n_476),
.B2(n_467),
.Y(n_561)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_477),
.A2(n_430),
.B1(n_432),
.B2(n_444),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_470),
.Y(n_523)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_523),
.Y(n_554)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_498),
.Y(n_526)
);

XOR2xp5_ASAP7_75t_L g529 ( 
.A(n_484),
.B(n_432),
.Y(n_529)
);

XOR2x2_ASAP7_75t_SL g530 ( 
.A(n_481),
.B(n_463),
.Y(n_530)
);

A2O1A1O1Ixp25_ASAP7_75t_L g552 ( 
.A1(n_530),
.A2(n_491),
.B(n_486),
.C(n_483),
.D(n_475),
.Y(n_552)
);

AOI21xp5_ASAP7_75t_L g531 ( 
.A1(n_492),
.A2(n_435),
.B(n_450),
.Y(n_531)
);

OAI21xp5_ASAP7_75t_SL g566 ( 
.A1(n_531),
.A2(n_541),
.B(n_437),
.Y(n_566)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_470),
.Y(n_532)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_532),
.Y(n_556)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_474),
.Y(n_533)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_533),
.Y(n_558)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_480),
.A2(n_462),
.B1(n_442),
.B2(n_434),
.Y(n_534)
);

XOR2xp5_ASAP7_75t_L g535 ( 
.A(n_493),
.B(n_462),
.Y(n_535)
);

XOR2xp5_ASAP7_75t_L g569 ( 
.A(n_535),
.B(n_478),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_SL g537 ( 
.A(n_472),
.B(n_444),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_537),
.B(n_539),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_493),
.B(n_448),
.C(n_434),
.Y(n_538)
);

CKINVDCx16_ASAP7_75t_R g539 ( 
.A(n_469),
.Y(n_539)
);

AOI21xp5_ASAP7_75t_L g541 ( 
.A1(n_492),
.A2(n_450),
.B(n_448),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_SL g542 ( 
.A1(n_466),
.A2(n_442),
.B1(n_437),
.B2(n_440),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_512),
.B(n_487),
.Y(n_544)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_544),
.Y(n_586)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_535),
.B(n_481),
.C(n_503),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g585 ( 
.A(n_547),
.B(n_577),
.C(n_529),
.Y(n_585)
);

NOR4xp25_ASAP7_75t_L g548 ( 
.A(n_512),
.B(n_499),
.C(n_487),
.D(n_481),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_L g605 ( 
.A1(n_548),
.A2(n_564),
.B1(n_318),
.B2(n_364),
.Y(n_605)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_536),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_549),
.B(n_550),
.Y(n_595)
);

CKINVDCx20_ASAP7_75t_R g550 ( 
.A(n_536),
.Y(n_550)
);

XNOR2xp5_ASAP7_75t_SL g599 ( 
.A(n_552),
.B(n_572),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_510),
.B(n_494),
.Y(n_553)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_553),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_510),
.B(n_488),
.Y(n_557)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_557),
.Y(n_589)
);

INVxp67_ASAP7_75t_L g559 ( 
.A(n_531),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_559),
.B(n_563),
.Y(n_604)
);

O2A1O1Ixp33_ASAP7_75t_L g560 ( 
.A1(n_540),
.A2(n_486),
.B(n_468),
.C(n_475),
.Y(n_560)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_560),
.Y(n_596)
);

OAI22xp5_ASAP7_75t_SL g592 ( 
.A1(n_561),
.A2(n_509),
.B1(n_514),
.B2(n_516),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_504),
.B(n_482),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_L g564 ( 
.A1(n_505),
.A2(n_485),
.B1(n_465),
.B2(n_471),
.Y(n_564)
);

AOI21xp5_ASAP7_75t_L g565 ( 
.A1(n_518),
.A2(n_497),
.B(n_495),
.Y(n_565)
);

CKINVDCx20_ASAP7_75t_R g581 ( 
.A(n_565),
.Y(n_581)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_566),
.Y(n_602)
);

OR2x2_ASAP7_75t_L g568 ( 
.A(n_525),
.B(n_500),
.Y(n_568)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_568),
.Y(n_606)
);

XOR2xp5_ASAP7_75t_L g584 ( 
.A(n_569),
.B(n_551),
.Y(n_584)
);

OAI22xp5_ASAP7_75t_SL g570 ( 
.A1(n_505),
.A2(n_501),
.B1(n_479),
.B2(n_490),
.Y(n_570)
);

AOI22xp5_ASAP7_75t_L g583 ( 
.A1(n_570),
.A2(n_519),
.B1(n_509),
.B2(n_542),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_507),
.B(n_440),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_571),
.B(n_573),
.Y(n_582)
);

XNOR2xp5_ASAP7_75t_SL g572 ( 
.A(n_517),
.B(n_335),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_507),
.B(n_440),
.Y(n_573)
);

INVx1_ASAP7_75t_SL g574 ( 
.A(n_524),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_574),
.B(n_575),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_511),
.B(n_451),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_538),
.B(n_335),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_SL g578 ( 
.A(n_576),
.B(n_525),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g577 ( 
.A(n_515),
.B(n_364),
.C(n_372),
.Y(n_577)
);

INVxp67_ASAP7_75t_L g608 ( 
.A(n_578),
.Y(n_608)
);

BUFx24_ASAP7_75t_SL g580 ( 
.A(n_562),
.Y(n_580)
);

BUFx24_ASAP7_75t_SL g607 ( 
.A(n_580),
.Y(n_607)
);

OAI22xp5_ASAP7_75t_SL g609 ( 
.A1(n_583),
.A2(n_565),
.B1(n_568),
.B2(n_545),
.Y(n_609)
);

XOR2xp5_ASAP7_75t_L g612 ( 
.A(n_584),
.B(n_603),
.Y(n_612)
);

XNOR2xp5_ASAP7_75t_L g625 ( 
.A(n_585),
.B(n_572),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_567),
.B(n_527),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_SL g610 ( 
.A(n_587),
.B(n_594),
.Y(n_610)
);

MAJIxp5_ASAP7_75t_L g590 ( 
.A(n_577),
.B(n_530),
.C(n_541),
.Y(n_590)
);

MAJIxp5_ASAP7_75t_L g611 ( 
.A(n_590),
.B(n_585),
.C(n_543),
.Y(n_611)
);

AOI22xp5_ASAP7_75t_L g591 ( 
.A1(n_555),
.A2(n_519),
.B1(n_509),
.B2(n_521),
.Y(n_591)
);

OAI22xp5_ASAP7_75t_L g614 ( 
.A1(n_591),
.A2(n_598),
.B1(n_600),
.B2(n_601),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_592),
.Y(n_615)
);

OAI22xp5_ASAP7_75t_SL g593 ( 
.A1(n_561),
.A2(n_527),
.B1(n_540),
.B2(n_522),
.Y(n_593)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_593),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_SL g594 ( 
.A(n_563),
.B(n_528),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_569),
.B(n_533),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_SL g631 ( 
.A(n_597),
.B(n_558),
.Y(n_631)
);

OAI22xp5_ASAP7_75t_SL g598 ( 
.A1(n_568),
.A2(n_534),
.B1(n_518),
.B2(n_506),
.Y(n_598)
);

AOI22xp5_ASAP7_75t_L g600 ( 
.A1(n_555),
.A2(n_520),
.B1(n_513),
.B2(n_532),
.Y(n_600)
);

AOI22xp5_ASAP7_75t_L g601 ( 
.A1(n_564),
.A2(n_506),
.B1(n_523),
.B2(n_524),
.Y(n_601)
);

XNOR2xp5_ASAP7_75t_SL g603 ( 
.A(n_551),
.B(n_326),
.Y(n_603)
);

OAI22xp5_ASAP7_75t_L g617 ( 
.A1(n_605),
.A2(n_549),
.B1(n_550),
.B2(n_557),
.Y(n_617)
);

AOI22xp5_ASAP7_75t_L g646 ( 
.A1(n_609),
.A2(n_617),
.B1(n_618),
.B2(n_621),
.Y(n_646)
);

AOI21xp33_ASAP7_75t_SL g638 ( 
.A1(n_611),
.A2(n_599),
.B(n_603),
.Y(n_638)
);

BUFx24_ASAP7_75t_SL g613 ( 
.A(n_604),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_613),
.B(n_616),
.Y(n_643)
);

CKINVDCx20_ASAP7_75t_R g616 ( 
.A(n_595),
.Y(n_616)
);

OAI22xp5_ASAP7_75t_SL g618 ( 
.A1(n_583),
.A2(n_591),
.B1(n_606),
.B2(n_604),
.Y(n_618)
);

MAJIxp5_ASAP7_75t_L g619 ( 
.A(n_600),
.B(n_543),
.C(n_590),
.Y(n_619)
);

MAJIxp5_ASAP7_75t_L g634 ( 
.A(n_619),
.B(n_620),
.C(n_626),
.Y(n_634)
);

MAJIxp5_ASAP7_75t_L g620 ( 
.A(n_584),
.B(n_547),
.C(n_559),
.Y(n_620)
);

OAI22xp5_ASAP7_75t_SL g621 ( 
.A1(n_606),
.A2(n_545),
.B1(n_544),
.B2(n_553),
.Y(n_621)
);

OAI22xp5_ASAP7_75t_L g623 ( 
.A1(n_601),
.A2(n_546),
.B1(n_554),
.B2(n_556),
.Y(n_623)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_623),
.Y(n_636)
);

OAI21xp5_ASAP7_75t_SL g624 ( 
.A1(n_581),
.A2(n_566),
.B(n_552),
.Y(n_624)
);

CKINVDCx14_ASAP7_75t_R g650 ( 
.A(n_624),
.Y(n_650)
);

XNOR2xp5_ASAP7_75t_L g640 ( 
.A(n_625),
.B(n_630),
.Y(n_640)
);

MAJIxp5_ASAP7_75t_L g626 ( 
.A(n_602),
.B(n_575),
.C(n_570),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_582),
.Y(n_627)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_627),
.Y(n_642)
);

MAJIxp5_ASAP7_75t_L g628 ( 
.A(n_602),
.B(n_546),
.C(n_573),
.Y(n_628)
);

MAJIxp5_ASAP7_75t_L g635 ( 
.A(n_628),
.B(n_629),
.C(n_588),
.Y(n_635)
);

MAJIxp5_ASAP7_75t_L g629 ( 
.A(n_581),
.B(n_571),
.C(n_574),
.Y(n_629)
);

XNOR2xp5_ASAP7_75t_L g630 ( 
.A(n_593),
.B(n_560),
.Y(n_630)
);

XNOR2xp5_ASAP7_75t_L g641 ( 
.A(n_631),
.B(n_588),
.Y(n_641)
);

OAI22xp5_ASAP7_75t_SL g632 ( 
.A1(n_615),
.A2(n_596),
.B1(n_595),
.B2(n_589),
.Y(n_632)
);

AOI22xp5_ASAP7_75t_L g668 ( 
.A1(n_632),
.A2(n_651),
.B1(n_636),
.B2(n_639),
.Y(n_668)
);

OAI21xp5_ASAP7_75t_SL g633 ( 
.A1(n_624),
.A2(n_596),
.B(n_548),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_633),
.B(n_649),
.Y(n_659)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_635),
.Y(n_663)
);

MAJIxp5_ASAP7_75t_L g637 ( 
.A(n_619),
.B(n_592),
.C(n_598),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_637),
.B(n_644),
.Y(n_656)
);

XNOR2xp5_ASAP7_75t_L g653 ( 
.A(n_638),
.B(n_625),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_629),
.B(n_589),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_639),
.B(n_648),
.Y(n_662)
);

OR2x2_ASAP7_75t_L g661 ( 
.A(n_641),
.B(n_652),
.Y(n_661)
);

XNOR2xp5_ASAP7_75t_L g644 ( 
.A(n_611),
.B(n_599),
.Y(n_644)
);

AOI21xp5_ASAP7_75t_L g645 ( 
.A1(n_608),
.A2(n_579),
.B(n_586),
.Y(n_645)
);

OAI21x1_ASAP7_75t_SL g655 ( 
.A1(n_645),
.A2(n_647),
.B(n_622),
.Y(n_655)
);

AOI21xp5_ASAP7_75t_L g647 ( 
.A1(n_608),
.A2(n_586),
.B(n_558),
.Y(n_647)
);

XNOR2xp5_ASAP7_75t_L g648 ( 
.A(n_626),
.B(n_556),
.Y(n_648)
);

MAJIxp5_ASAP7_75t_L g649 ( 
.A(n_620),
.B(n_554),
.C(n_347),
.Y(n_649)
);

OAI22xp5_ASAP7_75t_SL g651 ( 
.A1(n_615),
.A2(n_327),
.B1(n_338),
.B2(n_318),
.Y(n_651)
);

FAx1_ASAP7_75t_SL g652 ( 
.A(n_621),
.B(n_362),
.CI(n_341),
.CON(n_652),
.SN(n_652)
);

MAJx2_ASAP7_75t_L g677 ( 
.A(n_653),
.B(n_665),
.C(n_640),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_SL g654 ( 
.A(n_643),
.B(n_607),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_654),
.B(n_658),
.Y(n_680)
);

AOI21x1_ASAP7_75t_L g684 ( 
.A1(n_655),
.A2(n_326),
.B(n_362),
.Y(n_684)
);

MAJIxp5_ASAP7_75t_L g657 ( 
.A(n_634),
.B(n_614),
.C(n_618),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_657),
.B(n_660),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_SL g658 ( 
.A(n_642),
.B(n_610),
.Y(n_658)
);

MAJIxp5_ASAP7_75t_L g660 ( 
.A(n_634),
.B(n_622),
.C(n_628),
.Y(n_660)
);

XNOR2xp5_ASAP7_75t_L g664 ( 
.A(n_649),
.B(n_630),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_664),
.B(n_666),
.Y(n_679)
);

OAI21xp5_ASAP7_75t_SL g665 ( 
.A1(n_646),
.A2(n_609),
.B(n_612),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_635),
.B(n_338),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_641),
.Y(n_667)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_667),
.Y(n_675)
);

INVxp67_ASAP7_75t_L g676 ( 
.A(n_668),
.Y(n_676)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_639),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_669),
.B(n_350),
.Y(n_683)
);

MAJIxp5_ASAP7_75t_L g670 ( 
.A(n_637),
.B(n_612),
.C(n_327),
.Y(n_670)
);

AOI21xp5_ASAP7_75t_L g682 ( 
.A1(n_670),
.A2(n_652),
.B(n_350),
.Y(n_682)
);

OAI21xp5_ASAP7_75t_SL g671 ( 
.A1(n_656),
.A2(n_650),
.B(n_646),
.Y(n_671)
);

AOI21xp5_ASAP7_75t_SL g687 ( 
.A1(n_671),
.A2(n_683),
.B(n_661),
.Y(n_687)
);

AOI22xp5_ASAP7_75t_SL g673 ( 
.A1(n_663),
.A2(n_632),
.B1(n_651),
.B2(n_644),
.Y(n_673)
);

OAI21xp5_ASAP7_75t_L g692 ( 
.A1(n_673),
.A2(n_674),
.B(n_681),
.Y(n_692)
);

AOI21xp5_ASAP7_75t_SL g674 ( 
.A1(n_665),
.A2(n_648),
.B(n_640),
.Y(n_674)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_677),
.Y(n_689)
);

XOR2xp5_ASAP7_75t_L g678 ( 
.A(n_664),
.B(n_652),
.Y(n_678)
);

MAJIxp5_ASAP7_75t_L g685 ( 
.A(n_678),
.B(n_670),
.C(n_662),
.Y(n_685)
);

AOI22xp5_ASAP7_75t_SL g681 ( 
.A1(n_659),
.A2(n_662),
.B1(n_657),
.B2(n_660),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_682),
.B(n_653),
.Y(n_688)
);

OAI21xp5_ASAP7_75t_SL g686 ( 
.A1(n_684),
.A2(n_661),
.B(n_341),
.Y(n_686)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_685),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_686),
.B(n_687),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_688),
.B(n_691),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_672),
.B(n_676),
.Y(n_690)
);

AOI21xp5_ASAP7_75t_SL g696 ( 
.A1(n_690),
.A2(n_694),
.B(n_680),
.Y(n_696)
);

MAJIxp5_ASAP7_75t_L g691 ( 
.A(n_674),
.B(n_677),
.C(n_679),
.Y(n_691)
);

MAJIxp5_ASAP7_75t_L g693 ( 
.A(n_676),
.B(n_668),
.C(n_311),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_SL g698 ( 
.A(n_693),
.B(n_690),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_675),
.B(n_678),
.Y(n_694)
);

XOR2xp5_ASAP7_75t_L g702 ( 
.A(n_696),
.B(n_700),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_698),
.B(n_694),
.Y(n_701)
);

OAI21xp5_ASAP7_75t_SL g699 ( 
.A1(n_692),
.A2(n_341),
.B(n_333),
.Y(n_699)
);

AOI21xp5_ASAP7_75t_L g703 ( 
.A1(n_699),
.A2(n_689),
.B(n_311),
.Y(n_703)
);

MAJIxp5_ASAP7_75t_L g704 ( 
.A(n_701),
.B(n_702),
.C(n_703),
.Y(n_704)
);

MAJIxp5_ASAP7_75t_L g705 ( 
.A(n_702),
.B(n_697),
.C(n_695),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_705),
.Y(n_706)
);

OAI21xp5_ASAP7_75t_SL g707 ( 
.A1(n_706),
.A2(n_704),
.B(n_261),
.Y(n_707)
);

AO21x1_ASAP7_75t_L g708 ( 
.A1(n_707),
.A2(n_261),
.B(n_7),
.Y(n_708)
);

MAJIxp5_ASAP7_75t_L g709 ( 
.A(n_708),
.B(n_7),
.C(n_270),
.Y(n_709)
);

BUFx24_ASAP7_75t_SL g710 ( 
.A(n_709),
.Y(n_710)
);


endmodule