module fake_aes_2315_n_597 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_597);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_597;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_593;
wire n_554;
wire n_447;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_415;
wire n_482;
wire n_394;
wire n_243;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_446;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_285;
wire n_370;
wire n_589;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_395;
wire n_132;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
BUFx2_ASAP7_75t_SL g78 ( .A(n_34), .Y(n_78) );
NOR2xp67_ASAP7_75t_L g79 ( .A(n_63), .B(n_39), .Y(n_79) );
INVxp67_ASAP7_75t_SL g80 ( .A(n_1), .Y(n_80) );
INVxp67_ASAP7_75t_L g81 ( .A(n_53), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_4), .Y(n_82) );
CKINVDCx16_ASAP7_75t_R g83 ( .A(n_69), .Y(n_83) );
INVxp67_ASAP7_75t_L g84 ( .A(n_58), .Y(n_84) );
CKINVDCx5p33_ASAP7_75t_R g85 ( .A(n_67), .Y(n_85) );
CKINVDCx20_ASAP7_75t_R g86 ( .A(n_13), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_12), .Y(n_87) );
INVxp67_ASAP7_75t_SL g88 ( .A(n_28), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_38), .Y(n_89) );
INVx2_ASAP7_75t_L g90 ( .A(n_55), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_61), .Y(n_91) );
INVx3_ASAP7_75t_L g92 ( .A(n_20), .Y(n_92) );
INVxp67_ASAP7_75t_SL g93 ( .A(n_8), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_18), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_49), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_13), .Y(n_96) );
INVx2_ASAP7_75t_L g97 ( .A(n_56), .Y(n_97) );
CKINVDCx14_ASAP7_75t_R g98 ( .A(n_29), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_52), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_15), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_33), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_23), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_41), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_51), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_6), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_2), .Y(n_106) );
CKINVDCx14_ASAP7_75t_R g107 ( .A(n_8), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_36), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_27), .Y(n_109) );
CKINVDCx16_ASAP7_75t_R g110 ( .A(n_77), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_21), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_26), .Y(n_112) );
INVxp67_ASAP7_75t_SL g113 ( .A(n_7), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_68), .Y(n_114) );
OR2x2_ASAP7_75t_L g115 ( .A(n_10), .B(n_35), .Y(n_115) );
INVx2_ASAP7_75t_SL g116 ( .A(n_12), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_22), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_20), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_73), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_70), .Y(n_120) );
INVxp67_ASAP7_75t_L g121 ( .A(n_64), .Y(n_121) );
INVxp33_ASAP7_75t_SL g122 ( .A(n_50), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_40), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_62), .Y(n_124) );
INVx1_ASAP7_75t_SL g125 ( .A(n_26), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_32), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_90), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_116), .B(n_0), .Y(n_128) );
AND2x6_ASAP7_75t_L g129 ( .A(n_89), .B(n_31), .Y(n_129) );
HB1xp67_ASAP7_75t_L g130 ( .A(n_107), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_108), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_92), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_92), .Y(n_133) );
CKINVDCx20_ASAP7_75t_R g134 ( .A(n_86), .Y(n_134) );
CKINVDCx20_ASAP7_75t_R g135 ( .A(n_112), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_92), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_89), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_91), .Y(n_138) );
INVx5_ASAP7_75t_L g139 ( .A(n_90), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g140 ( .A(n_83), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_97), .Y(n_141) );
AND2x4_ASAP7_75t_L g142 ( .A(n_116), .B(n_0), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_110), .Y(n_143) );
INVx3_ASAP7_75t_L g144 ( .A(n_82), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_97), .Y(n_145) );
AND2x2_ASAP7_75t_L g146 ( .A(n_98), .B(n_1), .Y(n_146) );
CKINVDCx5p33_ASAP7_75t_R g147 ( .A(n_122), .Y(n_147) );
INVx2_ASAP7_75t_SL g148 ( .A(n_114), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_91), .Y(n_149) );
INVx3_ASAP7_75t_L g150 ( .A(n_95), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g151 ( .A(n_85), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_95), .Y(n_152) );
NOR2xp33_ASAP7_75t_L g153 ( .A(n_99), .B(n_2), .Y(n_153) );
AND2x6_ASAP7_75t_L g154 ( .A(n_99), .B(n_42), .Y(n_154) );
CKINVDCx20_ASAP7_75t_R g155 ( .A(n_125), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_114), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_101), .Y(n_157) );
CKINVDCx5p33_ASAP7_75t_R g158 ( .A(n_126), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_101), .Y(n_159) );
CKINVDCx20_ASAP7_75t_R g160 ( .A(n_115), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_103), .Y(n_161) );
NOR2xp33_ASAP7_75t_L g162 ( .A(n_103), .B(n_3), .Y(n_162) );
CKINVDCx20_ASAP7_75t_R g163 ( .A(n_115), .Y(n_163) );
CKINVDCx5p33_ASAP7_75t_R g164 ( .A(n_78), .Y(n_164) );
INVx3_ASAP7_75t_L g165 ( .A(n_104), .Y(n_165) );
NAND2xp5_ASAP7_75t_SL g166 ( .A(n_104), .B(n_3), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g167 ( .A(n_124), .B(n_4), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_109), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_109), .Y(n_169) );
OAI22xp5_ASAP7_75t_L g170 ( .A1(n_82), .A2(n_5), .B1(n_6), .B2(n_7), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_119), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_119), .B(n_5), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_142), .Y(n_173) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_150), .B(n_124), .Y(n_174) );
CKINVDCx20_ASAP7_75t_R g175 ( .A(n_134), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_142), .Y(n_176) );
CKINVDCx5p33_ASAP7_75t_R g177 ( .A(n_140), .Y(n_177) );
AO22x2_ASAP7_75t_L g178 ( .A1(n_142), .A2(n_100), .B1(n_94), .B2(n_87), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_142), .Y(n_179) );
AND2x4_ASAP7_75t_L g180 ( .A(n_132), .B(n_100), .Y(n_180) );
AND2x6_ASAP7_75t_L g181 ( .A(n_146), .B(n_123), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_164), .B(n_121), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_150), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_150), .Y(n_184) );
AND2x2_ASAP7_75t_SL g185 ( .A(n_146), .B(n_123), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_150), .B(n_120), .Y(n_186) );
BUFx3_ASAP7_75t_L g187 ( .A(n_129), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_130), .B(n_81), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_165), .Y(n_189) );
AND2x4_ASAP7_75t_L g190 ( .A(n_132), .B(n_96), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_144), .Y(n_191) );
AND2x4_ASAP7_75t_L g192 ( .A(n_133), .B(n_96), .Y(n_192) );
OAI221xp5_ASAP7_75t_L g193 ( .A1(n_137), .A2(n_94), .B1(n_118), .B2(n_117), .C(n_87), .Y(n_193) );
BUFx2_ASAP7_75t_L g194 ( .A(n_155), .Y(n_194) );
OAI22xp5_ASAP7_75t_L g195 ( .A1(n_160), .A2(n_102), .B1(n_118), .B2(n_117), .Y(n_195) );
BUFx6f_ASAP7_75t_L g196 ( .A(n_129), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_137), .B(n_84), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_144), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_144), .Y(n_199) );
AND2x4_ASAP7_75t_L g200 ( .A(n_133), .B(n_102), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_136), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_136), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_128), .Y(n_203) );
BUFx3_ASAP7_75t_L g204 ( .A(n_129), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_165), .B(n_120), .Y(n_205) );
BUFx4f_ASAP7_75t_L g206 ( .A(n_129), .Y(n_206) );
AND2x6_ASAP7_75t_L g207 ( .A(n_165), .B(n_111), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_165), .B(n_79), .Y(n_208) );
INVx2_ASAP7_75t_SL g209 ( .A(n_139), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_138), .B(n_88), .Y(n_210) );
BUFx6f_ASAP7_75t_L g211 ( .A(n_129), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_138), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_149), .B(n_78), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_149), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_152), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_152), .Y(n_216) );
NAND2x1p5_ASAP7_75t_L g217 ( .A(n_166), .B(n_111), .Y(n_217) );
NOR2x1p5_ASAP7_75t_L g218 ( .A(n_131), .B(n_113), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_157), .B(n_159), .Y(n_219) );
AND2x2_ASAP7_75t_L g220 ( .A(n_143), .B(n_105), .Y(n_220) );
AND2x4_ASAP7_75t_L g221 ( .A(n_148), .B(n_106), .Y(n_221) );
AND2x4_ASAP7_75t_L g222 ( .A(n_148), .B(n_106), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_157), .B(n_105), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_159), .Y(n_224) );
INVx2_ASAP7_75t_SL g225 ( .A(n_139), .Y(n_225) );
AOI22xp33_ASAP7_75t_L g226 ( .A1(n_129), .A2(n_93), .B1(n_80), .B2(n_11), .Y(n_226) );
INVx4_ASAP7_75t_L g227 ( .A(n_129), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_161), .Y(n_228) );
BUFx2_ASAP7_75t_L g229 ( .A(n_151), .Y(n_229) );
OAI21xp33_ASAP7_75t_SL g230 ( .A1(n_161), .A2(n_9), .B(n_10), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_168), .B(n_9), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_168), .B(n_11), .Y(n_232) );
NOR3xp33_ASAP7_75t_SL g233 ( .A(n_177), .B(n_147), .C(n_170), .Y(n_233) );
AOI22xp33_ASAP7_75t_L g234 ( .A1(n_178), .A2(n_154), .B1(n_171), .B2(n_169), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_183), .Y(n_235) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_227), .B(n_158), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_203), .B(n_171), .Y(n_237) );
BUFx6f_ASAP7_75t_L g238 ( .A(n_196), .Y(n_238) );
OR2x2_ASAP7_75t_SL g239 ( .A(n_188), .B(n_135), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_183), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_184), .Y(n_241) );
BUFx2_ASAP7_75t_L g242 ( .A(n_178), .Y(n_242) );
BUFx6f_ASAP7_75t_L g243 ( .A(n_196), .Y(n_243) );
CKINVDCx5p33_ASAP7_75t_R g244 ( .A(n_175), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_184), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_197), .B(n_169), .Y(n_246) );
INVx5_ASAP7_75t_L g247 ( .A(n_207), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_189), .Y(n_248) );
INVx2_ASAP7_75t_L g249 ( .A(n_189), .Y(n_249) );
BUFx6f_ASAP7_75t_L g250 ( .A(n_196), .Y(n_250) );
OR2x6_ASAP7_75t_L g251 ( .A(n_178), .B(n_172), .Y(n_251) );
BUFx2_ASAP7_75t_L g252 ( .A(n_181), .Y(n_252) );
NAND2xp5_ASAP7_75t_SL g253 ( .A(n_227), .B(n_167), .Y(n_253) );
BUFx3_ASAP7_75t_L g254 ( .A(n_187), .Y(n_254) );
INVx1_ASAP7_75t_SL g255 ( .A(n_194), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_191), .Y(n_256) );
HB1xp67_ASAP7_75t_L g257 ( .A(n_229), .Y(n_257) );
INVx3_ASAP7_75t_L g258 ( .A(n_207), .Y(n_258) );
AOI22xp5_ASAP7_75t_L g259 ( .A1(n_185), .A2(n_153), .B1(n_162), .B2(n_163), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_198), .Y(n_260) );
NOR2xp33_ASAP7_75t_L g261 ( .A(n_182), .B(n_156), .Y(n_261) );
NOR2xp33_ASAP7_75t_R g262 ( .A(n_177), .B(n_154), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_199), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_212), .B(n_154), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_173), .Y(n_265) );
BUFx3_ASAP7_75t_L g266 ( .A(n_187), .Y(n_266) );
INVx2_ASAP7_75t_L g267 ( .A(n_196), .Y(n_267) );
BUFx2_ASAP7_75t_L g268 ( .A(n_181), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_176), .Y(n_269) );
BUFx6f_ASAP7_75t_L g270 ( .A(n_211), .Y(n_270) );
INVx2_ASAP7_75t_SL g271 ( .A(n_207), .Y(n_271) );
BUFx3_ASAP7_75t_L g272 ( .A(n_204), .Y(n_272) );
AND2x4_ASAP7_75t_L g273 ( .A(n_180), .B(n_154), .Y(n_273) );
HB1xp67_ASAP7_75t_L g274 ( .A(n_181), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_211), .Y(n_275) );
OAI22xp5_ASAP7_75t_L g276 ( .A1(n_185), .A2(n_226), .B1(n_193), .B2(n_179), .Y(n_276) );
INVx2_ASAP7_75t_SL g277 ( .A(n_207), .Y(n_277) );
HB1xp67_ASAP7_75t_L g278 ( .A(n_181), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_201), .Y(n_279) );
INVx4_ASAP7_75t_L g280 ( .A(n_207), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_211), .Y(n_281) );
CKINVDCx5p33_ASAP7_75t_R g282 ( .A(n_175), .Y(n_282) );
OR2x2_ASAP7_75t_SL g283 ( .A(n_218), .B(n_156), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_202), .Y(n_284) );
INVxp67_ASAP7_75t_SL g285 ( .A(n_211), .Y(n_285) );
BUFx3_ASAP7_75t_L g286 ( .A(n_204), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_214), .Y(n_287) );
INVxp67_ASAP7_75t_L g288 ( .A(n_195), .Y(n_288) );
INVx3_ASAP7_75t_L g289 ( .A(n_180), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_215), .B(n_154), .Y(n_290) );
BUFx6f_ASAP7_75t_L g291 ( .A(n_227), .Y(n_291) );
CKINVDCx5p33_ASAP7_75t_R g292 ( .A(n_220), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_216), .Y(n_293) );
INVx3_ASAP7_75t_L g294 ( .A(n_180), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_224), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_228), .Y(n_296) );
NAND2xp5_ASAP7_75t_SL g297 ( .A(n_206), .B(n_139), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_209), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_190), .B(n_145), .Y(n_299) );
AOI22xp33_ASAP7_75t_L g300 ( .A1(n_181), .A2(n_154), .B1(n_145), .B2(n_141), .Y(n_300) );
BUFx3_ASAP7_75t_L g301 ( .A(n_291), .Y(n_301) );
INVx1_ASAP7_75t_SL g302 ( .A(n_255), .Y(n_302) );
A2O1A1Ixp33_ASAP7_75t_L g303 ( .A1(n_287), .A2(n_219), .B(n_213), .C(n_210), .Y(n_303) );
AOI22xp33_ASAP7_75t_SL g304 ( .A1(n_242), .A2(n_230), .B1(n_222), .B2(n_221), .Y(n_304) );
INVxp67_ASAP7_75t_SL g305 ( .A(n_242), .Y(n_305) );
HB1xp67_ASAP7_75t_L g306 ( .A(n_255), .Y(n_306) );
INVx1_ASAP7_75t_SL g307 ( .A(n_257), .Y(n_307) );
AND2x4_ASAP7_75t_L g308 ( .A(n_280), .B(n_200), .Y(n_308) );
AND2x4_ASAP7_75t_L g309 ( .A(n_280), .B(n_200), .Y(n_309) );
BUFx3_ASAP7_75t_L g310 ( .A(n_291), .Y(n_310) );
AOI21xp5_ASAP7_75t_L g311 ( .A1(n_264), .A2(n_206), .B(n_174), .Y(n_311) );
AOI21xp5_ASAP7_75t_L g312 ( .A1(n_264), .A2(n_206), .B(n_174), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_287), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_237), .B(n_219), .Y(n_314) );
NOR2xp33_ASAP7_75t_L g315 ( .A(n_288), .B(n_182), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_249), .Y(n_316) );
BUFx12f_ASAP7_75t_L g317 ( .A(n_251), .Y(n_317) );
OAI21xp33_ASAP7_75t_L g318 ( .A1(n_237), .A2(n_210), .B(n_213), .Y(n_318) );
AO22x1_ASAP7_75t_L g319 ( .A1(n_252), .A2(n_154), .B1(n_222), .B2(n_221), .Y(n_319) );
NOR3xp33_ASAP7_75t_L g320 ( .A(n_276), .B(n_232), .C(n_231), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_296), .Y(n_321) );
AND2x4_ASAP7_75t_L g322 ( .A(n_280), .B(n_200), .Y(n_322) );
BUFx3_ASAP7_75t_L g323 ( .A(n_291), .Y(n_323) );
CKINVDCx5p33_ASAP7_75t_R g324 ( .A(n_244), .Y(n_324) );
INVxp67_ASAP7_75t_SL g325 ( .A(n_280), .Y(n_325) );
BUFx2_ASAP7_75t_SL g326 ( .A(n_247), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_296), .B(n_222), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_279), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_251), .B(n_190), .Y(n_329) );
BUFx2_ASAP7_75t_L g330 ( .A(n_251), .Y(n_330) );
BUFx6f_ASAP7_75t_L g331 ( .A(n_291), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_249), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_251), .B(n_190), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_279), .B(n_221), .Y(n_334) );
BUFx6f_ASAP7_75t_L g335 ( .A(n_291), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_249), .Y(n_336) );
AOI22xp33_ASAP7_75t_L g337 ( .A1(n_251), .A2(n_192), .B1(n_186), .B2(n_205), .Y(n_337) );
INVx3_ASAP7_75t_L g338 ( .A(n_258), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_293), .Y(n_339) );
NAND2xp33_ASAP7_75t_L g340 ( .A(n_247), .B(n_225), .Y(n_340) );
BUFx3_ASAP7_75t_L g341 ( .A(n_291), .Y(n_341) );
NOR2x1_ASAP7_75t_L g342 ( .A(n_289), .B(n_205), .Y(n_342) );
AOI22xp33_ASAP7_75t_L g343 ( .A1(n_276), .A2(n_192), .B1(n_186), .B2(n_208), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_284), .Y(n_344) );
BUFx12f_ASAP7_75t_L g345 ( .A(n_292), .Y(n_345) );
INVx4_ASAP7_75t_L g346 ( .A(n_247), .Y(n_346) );
NOR2x1_ASAP7_75t_L g347 ( .A(n_289), .B(n_294), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_284), .Y(n_348) );
INVx2_ASAP7_75t_SL g349 ( .A(n_289), .Y(n_349) );
AOI21xp5_ASAP7_75t_L g350 ( .A1(n_290), .A2(n_225), .B(n_209), .Y(n_350) );
INVxp67_ASAP7_75t_SL g351 ( .A(n_254), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_256), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_293), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_293), .Y(n_354) );
NOR2xp33_ASAP7_75t_L g355 ( .A(n_259), .B(n_217), .Y(n_355) );
AOI221xp5_ASAP7_75t_L g356 ( .A1(n_246), .A2(n_223), .B1(n_192), .B2(n_208), .C(n_141), .Y(n_356) );
HB1xp67_ASAP7_75t_L g357 ( .A(n_282), .Y(n_357) );
AOI21xp5_ASAP7_75t_L g358 ( .A1(n_290), .A2(n_217), .B(n_127), .Y(n_358) );
A2O1A1Ixp33_ASAP7_75t_L g359 ( .A1(n_320), .A2(n_261), .B(n_269), .C(n_265), .Y(n_359) );
INVx3_ASAP7_75t_L g360 ( .A(n_346), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_314), .B(n_265), .Y(n_361) );
OAI21x1_ASAP7_75t_L g362 ( .A1(n_350), .A2(n_234), .B(n_300), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_339), .Y(n_363) );
OAI22xp33_ASAP7_75t_L g364 ( .A1(n_302), .A2(n_259), .B1(n_252), .B2(n_268), .Y(n_364) );
OAI21x1_ASAP7_75t_L g365 ( .A1(n_358), .A2(n_295), .B(n_236), .Y(n_365) );
AOI21xp5_ASAP7_75t_L g366 ( .A1(n_303), .A2(n_253), .B(n_273), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_314), .B(n_269), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_313), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_313), .B(n_289), .Y(n_369) );
AO21x2_ASAP7_75t_L g370 ( .A1(n_321), .A2(n_344), .B(n_328), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_339), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_339), .Y(n_372) );
AOI22xp33_ASAP7_75t_SL g373 ( .A1(n_317), .A2(n_268), .B1(n_262), .B2(n_278), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_353), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_321), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_328), .B(n_294), .Y(n_376) );
AOI22xp33_ASAP7_75t_L g377 ( .A1(n_355), .A2(n_294), .B1(n_274), .B2(n_273), .Y(n_377) );
AO31x2_ASAP7_75t_L g378 ( .A1(n_330), .A2(n_295), .A3(n_127), .B(n_256), .Y(n_378) );
AOI22xp33_ASAP7_75t_L g379 ( .A1(n_315), .A2(n_294), .B1(n_273), .B2(n_299), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_344), .Y(n_380) );
AOI22xp33_ASAP7_75t_L g381 ( .A1(n_329), .A2(n_273), .B1(n_299), .B2(n_260), .Y(n_381) );
OR2x6_ASAP7_75t_L g382 ( .A(n_317), .B(n_271), .Y(n_382) );
OAI22xp5_ASAP7_75t_L g383 ( .A1(n_304), .A2(n_295), .B1(n_260), .B2(n_235), .Y(n_383) );
OAI221xp5_ASAP7_75t_L g384 ( .A1(n_318), .A2(n_233), .B1(n_263), .B2(n_235), .C(n_240), .Y(n_384) );
AOI332xp33_ASAP7_75t_L g385 ( .A1(n_343), .A2(n_239), .A3(n_283), .B1(n_240), .B2(n_241), .B3(n_245), .C1(n_248), .C2(n_21), .Y(n_385) );
OAI21x1_ASAP7_75t_L g386 ( .A1(n_311), .A2(n_281), .B(n_275), .Y(n_386) );
AND2x4_ASAP7_75t_L g387 ( .A(n_308), .B(n_247), .Y(n_387) );
OAI22xp5_ASAP7_75t_L g388 ( .A1(n_348), .A2(n_248), .B1(n_245), .B2(n_241), .Y(n_388) );
OAI221xp5_ASAP7_75t_L g389 ( .A1(n_318), .A2(n_263), .B1(n_139), .B2(n_271), .C(n_277), .Y(n_389) );
OAI22xp33_ASAP7_75t_L g390 ( .A1(n_302), .A2(n_247), .B1(n_239), .B2(n_258), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_348), .Y(n_391) );
CKINVDCx5p33_ASAP7_75t_R g392 ( .A(n_324), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_353), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g394 ( .A1(n_329), .A2(n_263), .B1(n_258), .B2(n_277), .Y(n_394) );
CKINVDCx20_ASAP7_75t_R g395 ( .A(n_306), .Y(n_395) );
INVx3_ASAP7_75t_L g396 ( .A(n_387), .Y(n_396) );
AOI22xp33_ASAP7_75t_SL g397 ( .A1(n_395), .A2(n_317), .B1(n_307), .B2(n_345), .Y(n_397) );
OAI22xp33_ASAP7_75t_L g398 ( .A1(n_361), .A2(n_307), .B1(n_345), .B2(n_330), .Y(n_398) );
OAI22xp33_ASAP7_75t_L g399 ( .A1(n_361), .A2(n_345), .B1(n_305), .B2(n_334), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_368), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_368), .Y(n_401) );
BUFx6f_ASAP7_75t_L g402 ( .A(n_363), .Y(n_402) );
AOI22xp33_ASAP7_75t_L g403 ( .A1(n_384), .A2(n_333), .B1(n_357), .B2(n_356), .Y(n_403) );
INVx4_ASAP7_75t_SL g404 ( .A(n_378), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_367), .B(n_353), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_363), .Y(n_406) );
OAI222xp33_ASAP7_75t_L g407 ( .A1(n_383), .A2(n_333), .B1(n_352), .B2(n_354), .C1(n_334), .C2(n_327), .Y(n_407) );
AOI22xp33_ASAP7_75t_L g408 ( .A1(n_384), .A2(n_356), .B1(n_352), .B2(n_327), .Y(n_408) );
AND2x4_ASAP7_75t_L g409 ( .A(n_367), .B(n_308), .Y(n_409) );
AOI221xp5_ASAP7_75t_L g410 ( .A1(n_383), .A2(n_337), .B1(n_354), .B2(n_319), .C(n_349), .Y(n_410) );
AOI221xp5_ASAP7_75t_L g411 ( .A1(n_364), .A2(n_354), .B1(n_319), .B2(n_349), .C(n_308), .Y(n_411) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_390), .A2(n_322), .B1(n_309), .B2(n_308), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_379), .A2(n_322), .B1(n_309), .B2(n_347), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_375), .Y(n_414) );
AO31x2_ASAP7_75t_L g415 ( .A1(n_359), .A2(n_316), .A3(n_336), .B(n_332), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_381), .A2(n_322), .B1(n_309), .B2(n_347), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_375), .Y(n_417) );
OR2x2_ASAP7_75t_L g418 ( .A(n_363), .B(n_316), .Y(n_418) );
OAI22xp5_ASAP7_75t_L g419 ( .A1(n_388), .A2(n_316), .B1(n_332), .B2(n_336), .Y(n_419) );
AOI22xp5_ASAP7_75t_L g420 ( .A1(n_377), .A2(n_322), .B1(n_309), .B2(n_342), .Y(n_420) );
AOI22xp33_ASAP7_75t_L g421 ( .A1(n_380), .A2(n_342), .B1(n_338), .B2(n_332), .Y(n_421) );
OAI321xp33_ASAP7_75t_L g422 ( .A1(n_388), .A2(n_336), .A3(n_297), .B1(n_312), .B2(n_298), .C(n_351), .Y(n_422) );
OAI221xp5_ASAP7_75t_L g423 ( .A1(n_366), .A2(n_283), .B1(n_325), .B2(n_338), .C(n_258), .Y(n_423) );
OAI221xp5_ASAP7_75t_SL g424 ( .A1(n_385), .A2(n_338), .B1(n_301), .B2(n_310), .C(n_323), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_380), .Y(n_425) );
OAI332xp33_ASAP7_75t_L g426 ( .A1(n_398), .A2(n_385), .A3(n_391), .B1(n_369), .B2(n_374), .B3(n_372), .C1(n_371), .C2(n_393), .Y(n_426) );
NAND3xp33_ASAP7_75t_L g427 ( .A(n_424), .B(n_366), .C(n_393), .Y(n_427) );
OAI33xp33_ASAP7_75t_L g428 ( .A1(n_399), .A2(n_391), .A3(n_369), .B1(n_392), .B2(n_393), .B3(n_374), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_406), .Y(n_429) );
OAI33xp33_ASAP7_75t_L g430 ( .A1(n_400), .A2(n_374), .A3(n_372), .B1(n_371), .B2(n_17), .B3(n_18), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_405), .B(n_376), .Y(n_431) );
AOI221xp5_ASAP7_75t_L g432 ( .A1(n_403), .A2(n_376), .B1(n_370), .B2(n_371), .C(n_372), .Y(n_432) );
BUFx2_ASAP7_75t_L g433 ( .A(n_404), .Y(n_433) );
INVxp67_ASAP7_75t_L g434 ( .A(n_405), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_406), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_402), .Y(n_436) );
AOI21xp5_ASAP7_75t_SL g437 ( .A1(n_419), .A2(n_410), .B(n_411), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_400), .Y(n_438) );
OR2x2_ASAP7_75t_L g439 ( .A(n_418), .B(n_378), .Y(n_439) );
BUFx2_ASAP7_75t_L g440 ( .A(n_404), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_401), .B(n_370), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_402), .Y(n_442) );
INVxp67_ASAP7_75t_L g443 ( .A(n_418), .Y(n_443) );
INVx1_ASAP7_75t_SL g444 ( .A(n_402), .Y(n_444) );
OAI33xp33_ASAP7_75t_L g445 ( .A1(n_414), .A2(n_14), .A3(n_15), .B1(n_16), .B2(n_17), .B3(n_19), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_414), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_409), .B(n_370), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g448 ( .A1(n_409), .A2(n_370), .B1(n_382), .B2(n_373), .Y(n_448) );
AOI221xp5_ASAP7_75t_L g449 ( .A1(n_407), .A2(n_394), .B1(n_389), .B2(n_139), .C(n_360), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_417), .B(n_378), .Y(n_450) );
AOI21xp5_ASAP7_75t_SL g451 ( .A1(n_402), .A2(n_389), .B(n_382), .Y(n_451) );
AOI221xp5_ASAP7_75t_L g452 ( .A1(n_425), .A2(n_139), .B1(n_360), .B2(n_387), .C(n_373), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_415), .Y(n_453) );
AOI322xp5_ASAP7_75t_L g454 ( .A1(n_397), .A2(n_416), .A3(n_413), .B1(n_408), .B2(n_412), .C1(n_420), .C2(n_396), .Y(n_454) );
AOI22xp5_ASAP7_75t_L g455 ( .A1(n_423), .A2(n_382), .B1(n_387), .B2(n_360), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_396), .B(n_378), .Y(n_456) );
AO21x2_ASAP7_75t_L g457 ( .A1(n_422), .A2(n_386), .B(n_365), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_447), .B(n_404), .Y(n_458) );
AOI221xp5_ASAP7_75t_L g459 ( .A1(n_426), .A2(n_421), .B1(n_396), .B2(n_360), .C(n_387), .Y(n_459) );
INVxp67_ASAP7_75t_L g460 ( .A(n_439), .Y(n_460) );
INVx2_ASAP7_75t_SL g461 ( .A(n_433), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_447), .B(n_404), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_441), .B(n_378), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_441), .B(n_378), .Y(n_464) );
NAND3xp33_ASAP7_75t_L g465 ( .A(n_454), .B(n_382), .C(n_331), .Y(n_465) );
INVx2_ASAP7_75t_SL g466 ( .A(n_440), .Y(n_466) );
OR2x2_ASAP7_75t_L g467 ( .A(n_450), .B(n_415), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_434), .B(n_415), .Y(n_468) );
INVx6_ASAP7_75t_L g469 ( .A(n_456), .Y(n_469) );
NAND2xp33_ASAP7_75t_SL g470 ( .A(n_440), .B(n_346), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_438), .Y(n_471) );
INVxp67_ASAP7_75t_SL g472 ( .A(n_443), .Y(n_472) );
HB1xp67_ASAP7_75t_L g473 ( .A(n_429), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_456), .B(n_415), .Y(n_474) );
OAI21xp5_ASAP7_75t_L g475 ( .A1(n_454), .A2(n_362), .B(n_365), .Y(n_475) );
OR2x2_ASAP7_75t_L g476 ( .A(n_450), .B(n_415), .Y(n_476) );
AND2x4_ASAP7_75t_L g477 ( .A(n_436), .B(n_386), .Y(n_477) );
OR2x2_ASAP7_75t_L g478 ( .A(n_446), .B(n_14), .Y(n_478) );
OAI33xp33_ASAP7_75t_L g479 ( .A1(n_446), .A2(n_16), .A3(n_19), .B1(n_22), .B2(n_23), .B3(n_24), .Y(n_479) );
OR2x2_ASAP7_75t_L g480 ( .A(n_429), .B(n_24), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_435), .Y(n_481) );
AO211x2_ASAP7_75t_L g482 ( .A1(n_426), .A2(n_25), .B(n_382), .C(n_37), .Y(n_482) );
OR2x2_ASAP7_75t_L g483 ( .A(n_435), .B(n_25), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_453), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_436), .Y(n_485) );
NAND2x1p5_ASAP7_75t_L g486 ( .A(n_444), .B(n_335), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_442), .Y(n_487) );
OR2x2_ASAP7_75t_L g488 ( .A(n_431), .B(n_382), .Y(n_488) );
AOI211xp5_ASAP7_75t_L g489 ( .A1(n_428), .A2(n_340), .B(n_331), .C(n_335), .Y(n_489) );
NOR2xp33_ASAP7_75t_L g490 ( .A(n_472), .B(n_445), .Y(n_490) );
NAND5xp2_ASAP7_75t_SL g491 ( .A(n_459), .B(n_448), .C(n_455), .D(n_452), .E(n_449), .Y(n_491) );
AND2x4_ASAP7_75t_L g492 ( .A(n_458), .B(n_457), .Y(n_492) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_479), .B(n_430), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_460), .B(n_432), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_474), .B(n_457), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_474), .B(n_457), .Y(n_496) );
OR2x2_ASAP7_75t_L g497 ( .A(n_463), .B(n_427), .Y(n_497) );
AOI221xp5_ASAP7_75t_L g498 ( .A1(n_465), .A2(n_437), .B1(n_427), .B2(n_451), .C(n_455), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_463), .B(n_451), .Y(n_499) );
INVx2_ASAP7_75t_SL g500 ( .A(n_461), .Y(n_500) );
OAI22xp5_ASAP7_75t_L g501 ( .A1(n_465), .A2(n_437), .B1(n_301), .B2(n_341), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_471), .Y(n_502) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_478), .B(n_30), .Y(n_503) );
BUFx2_ASAP7_75t_L g504 ( .A(n_461), .Y(n_504) );
NOR3xp33_ASAP7_75t_SL g505 ( .A(n_470), .B(n_43), .C(n_44), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_464), .B(n_331), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_464), .B(n_45), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_469), .B(n_46), .Y(n_508) );
INVx2_ASAP7_75t_SL g509 ( .A(n_466), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_469), .B(n_47), .Y(n_510) );
AND2x4_ASAP7_75t_L g511 ( .A(n_458), .B(n_48), .Y(n_511) );
INVx2_ASAP7_75t_SL g512 ( .A(n_466), .Y(n_512) );
HB1xp67_ASAP7_75t_L g513 ( .A(n_473), .Y(n_513) );
AND2x4_ASAP7_75t_L g514 ( .A(n_462), .B(n_54), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_469), .B(n_57), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_484), .Y(n_516) );
AND2x4_ASAP7_75t_L g517 ( .A(n_484), .B(n_59), .Y(n_517) );
INVx4_ASAP7_75t_L g518 ( .A(n_480), .Y(n_518) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_488), .B(n_60), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_488), .B(n_335), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_483), .Y(n_521) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_489), .B(n_247), .Y(n_522) );
INVx2_ASAP7_75t_SL g523 ( .A(n_481), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_485), .Y(n_524) );
AOI22xp5_ASAP7_75t_L g525 ( .A1(n_490), .A2(n_482), .B1(n_468), .B2(n_489), .Y(n_525) );
OAI211xp5_ASAP7_75t_L g526 ( .A1(n_498), .A2(n_475), .B(n_467), .C(n_476), .Y(n_526) );
OAI22xp5_ASAP7_75t_L g527 ( .A1(n_518), .A2(n_476), .B1(n_482), .B2(n_487), .Y(n_527) );
INVxp67_ASAP7_75t_L g528 ( .A(n_504), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_502), .Y(n_529) );
INVx2_ASAP7_75t_L g530 ( .A(n_513), .Y(n_530) );
INVx2_ASAP7_75t_L g531 ( .A(n_523), .Y(n_531) );
INVxp33_ASAP7_75t_SL g532 ( .A(n_507), .Y(n_532) );
AOI322xp5_ASAP7_75t_L g533 ( .A1(n_493), .A2(n_477), .A3(n_341), .B1(n_323), .B2(n_310), .C1(n_301), .C2(n_486), .Y(n_533) );
NOR3xp33_ASAP7_75t_L g534 ( .A(n_503), .B(n_338), .C(n_323), .Y(n_534) );
OAI22xp5_ASAP7_75t_L g535 ( .A1(n_518), .A2(n_341), .B1(n_310), .B2(n_326), .Y(n_535) );
OAI21xp33_ASAP7_75t_L g536 ( .A1(n_499), .A2(n_298), .B(n_66), .Y(n_536) );
AOI33xp33_ASAP7_75t_L g537 ( .A1(n_495), .A2(n_298), .A3(n_71), .B1(n_72), .B2(n_74), .B3(n_75), .Y(n_537) );
OAI22xp33_ASAP7_75t_SL g538 ( .A1(n_500), .A2(n_65), .B1(n_76), .B2(n_286), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_523), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_516), .Y(n_540) );
INVx1_ASAP7_75t_SL g541 ( .A(n_509), .Y(n_541) );
OAI32xp33_ASAP7_75t_L g542 ( .A1(n_518), .A2(n_286), .A3(n_254), .B1(n_266), .B2(n_272), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_524), .Y(n_543) );
INVx1_ASAP7_75t_SL g544 ( .A(n_512), .Y(n_544) );
OAI22xp33_ASAP7_75t_SL g545 ( .A1(n_512), .A2(n_266), .B1(n_272), .B2(n_285), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_521), .Y(n_546) );
AOI22xp5_ASAP7_75t_L g547 ( .A1(n_519), .A2(n_267), .B1(n_275), .B2(n_281), .Y(n_547) );
O2A1O1Ixp33_ASAP7_75t_L g548 ( .A1(n_491), .A2(n_267), .B(n_243), .C(n_250), .Y(n_548) );
OAI32xp33_ASAP7_75t_L g549 ( .A1(n_497), .A2(n_238), .A3(n_243), .B1(n_250), .B2(n_270), .Y(n_549) );
AOI22xp5_ASAP7_75t_L g550 ( .A1(n_494), .A2(n_238), .B1(n_243), .B2(n_250), .Y(n_550) );
OR2x2_ASAP7_75t_L g551 ( .A(n_506), .B(n_238), .Y(n_551) );
AOI22xp33_ASAP7_75t_SL g552 ( .A1(n_511), .A2(n_238), .B1(n_243), .B2(n_250), .Y(n_552) );
AOI21xp33_ASAP7_75t_SL g553 ( .A1(n_511), .A2(n_238), .B(n_243), .Y(n_553) );
AOI221xp5_ASAP7_75t_L g554 ( .A1(n_527), .A2(n_495), .B1(n_496), .B2(n_501), .C(n_507), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_530), .Y(n_555) );
AOI22xp5_ASAP7_75t_L g556 ( .A1(n_527), .A2(n_496), .B1(n_514), .B2(n_492), .Y(n_556) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_532), .A2(n_514), .B1(n_492), .B2(n_520), .Y(n_557) );
INVx3_ASAP7_75t_SL g558 ( .A(n_541), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_546), .B(n_525), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g560 ( .A(n_528), .B(n_522), .Y(n_560) );
A2O1A1Ixp33_ASAP7_75t_L g561 ( .A1(n_534), .A2(n_514), .B(n_505), .C(n_510), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_529), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_540), .Y(n_563) );
AOI22xp5_ASAP7_75t_L g564 ( .A1(n_526), .A2(n_515), .B1(n_508), .B2(n_517), .Y(n_564) );
INVx3_ASAP7_75t_SL g565 ( .A(n_541), .Y(n_565) );
INVx1_ASAP7_75t_SL g566 ( .A(n_544), .Y(n_566) );
HB1xp67_ASAP7_75t_L g567 ( .A(n_544), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_543), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_531), .B(n_270), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_539), .B(n_270), .Y(n_570) );
NAND3xp33_ASAP7_75t_L g571 ( .A(n_533), .B(n_250), .C(n_270), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_559), .B(n_551), .Y(n_572) );
INVxp67_ASAP7_75t_L g573 ( .A(n_567), .Y(n_573) );
OAI22xp5_ASAP7_75t_L g574 ( .A1(n_557), .A2(n_535), .B1(n_553), .B2(n_536), .Y(n_574) );
NOR3xp33_ASAP7_75t_L g575 ( .A(n_554), .B(n_538), .C(n_537), .Y(n_575) );
AOI22xp5_ASAP7_75t_L g576 ( .A1(n_556), .A2(n_560), .B1(n_564), .B2(n_557), .Y(n_576) );
BUFx3_ASAP7_75t_L g577 ( .A(n_558), .Y(n_577) );
OAI22xp33_ASAP7_75t_L g578 ( .A1(n_565), .A2(n_547), .B1(n_550), .B2(n_552), .Y(n_578) );
AOI21xp5_ASAP7_75t_L g579 ( .A1(n_561), .A2(n_545), .B(n_542), .Y(n_579) );
NAND3xp33_ASAP7_75t_L g580 ( .A(n_560), .B(n_548), .C(n_549), .Y(n_580) );
BUFx3_ASAP7_75t_L g581 ( .A(n_566), .Y(n_581) );
NOR3xp33_ASAP7_75t_L g582 ( .A(n_571), .B(n_561), .C(n_555), .Y(n_582) );
INVx2_ASAP7_75t_SL g583 ( .A(n_577), .Y(n_583) );
NAND3xp33_ASAP7_75t_L g584 ( .A(n_582), .B(n_562), .C(n_563), .Y(n_584) );
NOR2x1_ASAP7_75t_L g585 ( .A(n_578), .B(n_568), .Y(n_585) );
AOI211xp5_ASAP7_75t_SL g586 ( .A1(n_579), .A2(n_569), .B(n_570), .C(n_575), .Y(n_586) );
CKINVDCx20_ASAP7_75t_R g587 ( .A(n_581), .Y(n_587) );
OAI22xp5_ASAP7_75t_L g588 ( .A1(n_573), .A2(n_574), .B1(n_572), .B2(n_580), .Y(n_588) );
OAI221xp5_ASAP7_75t_R g589 ( .A1(n_576), .A2(n_556), .B1(n_582), .B2(n_575), .C(n_557), .Y(n_589) );
CKINVDCx5p33_ASAP7_75t_R g590 ( .A(n_587), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_585), .B(n_586), .Y(n_591) );
BUFx2_ASAP7_75t_L g592 ( .A(n_583), .Y(n_592) );
AOI22xp33_ASAP7_75t_SL g593 ( .A1(n_591), .A2(n_588), .B1(n_589), .B2(n_584), .Y(n_593) );
XNOR2xp5_ASAP7_75t_L g594 ( .A(n_593), .B(n_590), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_594), .Y(n_595) );
AOI22xp5_ASAP7_75t_SL g596 ( .A1(n_595), .A2(n_591), .B1(n_592), .B2(n_593), .Y(n_596) );
UNKNOWN g597 ( );
endmodule