module real_jpeg_14335_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx10_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx4f_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_2),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_3),
.A2(n_28),
.B1(n_29),
.B2(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_3),
.A2(n_34),
.B1(n_47),
.B2(n_48),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_3),
.A2(n_34),
.B1(n_66),
.B2(n_67),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_3),
.A2(n_34),
.B1(n_61),
.B2(n_63),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_4),
.A2(n_61),
.B1(n_63),
.B2(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_4),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_4),
.A2(n_66),
.B1(n_67),
.B2(n_71),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_4),
.A2(n_47),
.B1(n_48),
.B2(n_71),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_4),
.A2(n_28),
.B1(n_29),
.B2(n_71),
.Y(n_215)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_6),
.A2(n_28),
.B1(n_29),
.B2(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

OAI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_6),
.A2(n_39),
.B1(n_47),
.B2(n_48),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_6),
.A2(n_39),
.B1(n_66),
.B2(n_67),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g269 ( 
.A1(n_6),
.A2(n_39),
.B1(n_61),
.B2(n_63),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_7),
.A2(n_61),
.B1(n_63),
.B2(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_7),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_7),
.A2(n_66),
.B1(n_67),
.B2(n_112),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_7),
.A2(n_47),
.B1(n_48),
.B2(n_112),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_7),
.A2(n_28),
.B1(n_29),
.B2(n_112),
.Y(n_221)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_8),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_9),
.A2(n_61),
.B1(n_63),
.B2(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_9),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_9),
.A2(n_66),
.B1(n_67),
.B2(n_69),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_9),
.A2(n_47),
.B1(n_48),
.B2(n_69),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_9),
.A2(n_28),
.B1(n_29),
.B2(n_69),
.Y(n_213)
);

BUFx12_ASAP7_75t_L g76 ( 
.A(n_10),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_11),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_11),
.B(n_127),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_11),
.B(n_29),
.C(n_45),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_11),
.A2(n_47),
.B1(n_48),
.B2(n_102),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_11),
.A2(n_26),
.B1(n_37),
.B2(n_221),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_11),
.B(n_108),
.Y(n_232)
);

BUFx8_ASAP7_75t_L g60 ( 
.A(n_12),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_13),
.A2(n_66),
.B1(n_67),
.B2(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_13),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_13),
.A2(n_28),
.B1(n_29),
.B2(n_80),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_13),
.A2(n_61),
.B1(n_63),
.B2(n_80),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_13),
.A2(n_47),
.B1(n_48),
.B2(n_80),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_14),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_46)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_14),
.A2(n_28),
.B1(n_29),
.B2(n_49),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_14),
.A2(n_49),
.B1(n_66),
.B2(n_67),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_14),
.A2(n_49),
.B1(n_61),
.B2(n_63),
.Y(n_285)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_329),
.Y(n_16)
);

AOI21xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_317),
.B(n_328),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_279),
.B(n_314),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_256),
.B(n_278),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_138),
.B(n_255),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_113),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_22),
.B(n_113),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_83),
.C(n_93),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_23),
.B(n_83),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_55),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_24),
.B(n_56),
.C(n_73),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_40),
.Y(n_24)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_25),
.B(n_40),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_32),
.B(n_35),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_26),
.A2(n_37),
.B(n_133),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_26),
.A2(n_37),
.B1(n_213),
.B2(n_221),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_26),
.A2(n_88),
.B(n_215),
.Y(n_235)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_27),
.B(n_87),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_27),
.A2(n_31),
.B1(n_33),
.B2(n_98),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_27),
.A2(n_36),
.B(n_89),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_27),
.A2(n_31),
.B1(n_212),
.B2(n_214),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_31),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_28),
.A2(n_29),
.B1(n_43),
.B2(n_45),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_28),
.B(n_219),
.Y(n_218)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_29),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_31),
.B(n_89),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_33),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_38),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_37),
.A2(n_86),
.B(n_99),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_37),
.B(n_102),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_38),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_46),
.B(n_50),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_41),
.A2(n_46),
.B1(n_53),
.B2(n_92),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_41),
.A2(n_53),
.B1(n_209),
.B2(n_210),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_41),
.B(n_102),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_41),
.A2(n_53),
.B1(n_185),
.B2(n_210),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_41),
.A2(n_53),
.B(n_149),
.Y(n_292)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_42),
.B(n_51),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_42),
.A2(n_52),
.B1(n_184),
.B2(n_186),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_42),
.B(n_196),
.Y(n_195)
);

CKINVDCx14_ASAP7_75t_SL g45 ( 
.A(n_43),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_43),
.A2(n_45),
.B1(n_47),
.B2(n_48),
.Y(n_54)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OA22x2_ASAP7_75t_SL g78 ( 
.A1(n_47),
.A2(n_48),
.B1(n_76),
.B2(n_77),
.Y(n_78)
);

NAND3xp33_ASAP7_75t_L g181 ( 
.A(n_47),
.B(n_67),
.C(n_77),
.Y(n_181)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

A2O1A1Ixp33_ASAP7_75t_L g179 ( 
.A1(n_48),
.A2(n_76),
.B(n_180),
.C(n_181),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_48),
.B(n_206),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_50),
.B(n_195),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_52),
.Y(n_50)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_53),
.A2(n_92),
.B(n_135),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_53),
.A2(n_135),
.B(n_149),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_53),
.A2(n_194),
.B(n_195),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_56),
.A2(n_57),
.B1(n_72),
.B2(n_73),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_65),
.B1(n_68),
.B2(n_70),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_58),
.A2(n_65),
.B1(n_68),
.B2(n_110),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_58),
.A2(n_70),
.B(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_58),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_58),
.B(n_269),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_65),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_61),
.B1(n_63),
.B2(n_64),
.Y(n_59)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_60),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_60),
.A2(n_64),
.B1(n_66),
.B2(n_67),
.Y(n_65)
);

A2O1A1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_60),
.A2(n_67),
.B(n_101),
.C(n_103),
.Y(n_100)
);

INVx3_ASAP7_75t_SL g63 ( 
.A(n_61),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

HAxp5_ASAP7_75t_SL g101 ( 
.A(n_63),
.B(n_102),
.CON(n_101),
.SN(n_101)
);

NAND3xp33_ASAP7_75t_L g103 ( 
.A(n_63),
.B(n_64),
.C(n_66),
.Y(n_103)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_65),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_65),
.B(n_269),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_66),
.A2(n_67),
.B1(n_76),
.B2(n_77),
.Y(n_75)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

HAxp5_ASAP7_75t_SL g180 ( 
.A(n_67),
.B(n_102),
.CON(n_180),
.SN(n_180)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_79),
.B(n_81),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_74),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_74),
.B(n_124),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_74),
.A2(n_108),
.B1(n_157),
.B2(n_180),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_74),
.A2(n_108),
.B1(n_274),
.B2(n_275),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_74),
.A2(n_79),
.B(n_108),
.Y(n_324)
);

AND2x2_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_78),
.Y(n_74)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_76),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_78),
.B(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_78),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_78),
.A2(n_122),
.B(n_123),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_78),
.A2(n_105),
.B1(n_106),
.B2(n_147),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_78),
.A2(n_106),
.B1(n_147),
.B2(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_79),
.B(n_108),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_81),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_82),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_85),
.B1(n_90),
.B2(n_91),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_84),
.B(n_91),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_88),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_89),
.Y(n_133)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_93),
.B(n_253),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_104),
.C(n_109),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_94),
.A2(n_95),
.B1(n_163),
.B2(n_164),
.Y(n_162)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_100),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_96),
.A2(n_97),
.B1(n_100),
.B2(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_100),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_101),
.A2(n_111),
.B1(n_127),
.B2(n_143),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_104),
.B(n_109),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_106),
.B(n_107),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_106),
.A2(n_290),
.B(n_291),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_107),
.B(n_123),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_137),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_115),
.A2(n_116),
.B1(n_129),
.B2(n_130),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_115),
.B(n_130),
.C(n_137),
.Y(n_277)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_118),
.B1(n_119),
.B2(n_120),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_117),
.B(n_121),
.C(n_125),
.Y(n_259)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_125),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_122),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_126),
.B(n_332),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_128),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_127),
.A2(n_285),
.B(n_286),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_127),
.A2(n_143),
.B1(n_285),
.B2(n_303),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_128),
.A2(n_143),
.B(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_132),
.B1(n_134),
.B2(n_136),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_131),
.A2(n_132),
.B1(n_266),
.B2(n_267),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_132),
.B(n_134),
.Y(n_264)
);

AOI21xp33_ASAP7_75t_L g296 ( 
.A1(n_132),
.A2(n_264),
.B(n_267),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_134),
.Y(n_136)
);

O2A1O1Ixp33_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_168),
.B(n_250),
.C(n_254),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_161),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_140),
.B(n_161),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_151),
.C(n_154),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_141),
.B(n_246),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_144),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_142),
.B(n_145),
.C(n_150),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_143),
.A2(n_268),
.B(n_303),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_146),
.B1(n_148),
.B2(n_150),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_148),
.Y(n_150)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_149),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_151),
.A2(n_152),
.B1(n_154),
.B2(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_154),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_158),
.C(n_160),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g188 ( 
.A(n_155),
.B(n_189),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_158),
.A2(n_159),
.B1(n_160),
.B2(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_160),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_165),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_162),
.B(n_166),
.C(n_167),
.Y(n_251)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_163),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_171),
.A2(n_244),
.B(n_249),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_199),
.B(n_243),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_187),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_173),
.B(n_187),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_182),
.C(n_183),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_174),
.A2(n_175),
.B1(n_239),
.B2(n_240),
.Y(n_238)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_177),
.B1(n_178),
.B2(n_179),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_176),
.B(n_179),
.Y(n_192)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_182),
.B(n_183),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

CKINVDCx14_ASAP7_75t_R g194 ( 
.A(n_186),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_191),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_188),
.B(n_193),
.C(n_197),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_192),
.A2(n_193),
.B1(n_197),
.B2(n_198),
.Y(n_191)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_192),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_193),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_237),
.B(n_242),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_227),
.B(n_236),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_216),
.B(n_226),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_211),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_203),
.B(n_211),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_207),
.B2(n_208),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_205),
.B(n_207),
.Y(n_228)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

CKINVDCx14_ASAP7_75t_R g214 ( 
.A(n_215),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_222),
.B(n_225),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_220),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_223),
.B(n_224),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_228),
.B(n_229),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_235),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_232),
.B1(n_233),
.B2(n_234),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_231),
.B(n_234),
.C(n_235),
.Y(n_241)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_238),
.B(n_241),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_238),
.B(n_241),
.Y(n_242)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_245),
.B(n_248),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_245),
.B(n_248),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_251),
.B(n_252),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_257),
.B(n_277),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_257),
.B(n_277),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_259),
.B1(n_260),
.B2(n_261),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_258),
.B(n_262),
.C(n_271),
.Y(n_310)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_262),
.A2(n_263),
.B1(n_270),
.B2(n_271),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

CKINVDCx14_ASAP7_75t_R g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_272),
.A2(n_273),
.B(n_276),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_272),
.B(n_273),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_275),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_276),
.B(n_282),
.C(n_296),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_276),
.A2(n_282),
.B1(n_283),
.B2(n_313),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_276),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_280),
.B(n_309),
.Y(n_279)
);

AOI21xp33_ASAP7_75t_L g314 ( 
.A1(n_280),
.A2(n_315),
.B(n_316),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_297),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_281),
.B(n_297),
.Y(n_316)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_287),
.B1(n_294),
.B2(n_295),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_284),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_284),
.B(n_289),
.C(n_292),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_284),
.A2(n_294),
.B1(n_301),
.B2(n_307),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_286),
.Y(n_332)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_287),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_289),
.B1(n_292),
.B2(n_293),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_289),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_292),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_292),
.A2(n_293),
.B1(n_305),
.B2(n_306),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_292),
.B(n_302),
.C(n_306),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_294),
.B(n_298),
.C(n_307),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_296),
.B(n_312),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_298),
.A2(n_299),
.B1(n_300),
.B2(n_308),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_300),
.Y(n_308)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_301),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_304),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_306),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_310),
.B(n_311),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_318),
.B(n_319),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_318),
.B(n_319),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_320),
.A2(n_325),
.B1(n_326),
.B2(n_327),
.Y(n_319)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_320),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_321),
.A2(n_322),
.B1(n_323),
.B2(n_324),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_322),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_322),
.B(n_323),
.C(n_325),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_324),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_326),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_335),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_333),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_331),
.Y(n_336)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_336),
.Y(n_335)
);


endmodule