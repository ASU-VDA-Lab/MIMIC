module fake_jpeg_2778_n_308 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_308);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_308;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx8_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx24_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

INVx11_ASAP7_75t_SL g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_1),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_13),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_10),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_0),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_15),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_10),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_5),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_2),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_52),
.Y(n_131)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_53),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_54),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

INVx4_ASAP7_75t_SL g121 ( 
.A(n_55),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_56),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_1),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_57),
.B(n_58),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_28),
.B(n_47),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_59),
.Y(n_150)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_60),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_41),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_61),
.B(n_64),
.Y(n_109)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_62),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_63),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_41),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_65),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_66),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_1),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_67),
.B(n_68),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_18),
.B(n_33),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_18),
.B(n_3),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_69),
.B(n_71),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_17),
.Y(n_70)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_70),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_19),
.B(n_4),
.Y(n_71)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_26),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g151 ( 
.A(n_72),
.Y(n_151)
);

OR2x2_ASAP7_75t_SL g73 ( 
.A(n_50),
.B(n_51),
.Y(n_73)
);

NAND2xp33_ASAP7_75t_SL g132 ( 
.A(n_73),
.B(n_97),
.Y(n_132)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_74),
.Y(n_140)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_30),
.Y(n_75)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_75),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_26),
.Y(n_76)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_76),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_19),
.B(n_4),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_77),
.B(n_78),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_21),
.B(n_4),
.Y(n_78)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_26),
.Y(n_79)
);

INVx8_ASAP7_75t_L g139 ( 
.A(n_79),
.Y(n_139)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_26),
.Y(n_80)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_80),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_50),
.A2(n_7),
.B1(n_10),
.B2(n_12),
.Y(n_81)
);

OA22x2_ASAP7_75t_L g118 ( 
.A1(n_81),
.A2(n_12),
.B1(n_14),
.B2(n_36),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_21),
.B(n_7),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_82),
.B(n_87),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_31),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g130 ( 
.A(n_83),
.Y(n_130)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_32),
.Y(n_85)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_85),
.Y(n_155)
);

BUFx4f_ASAP7_75t_SL g86 ( 
.A(n_32),
.Y(n_86)
);

INVx5_ASAP7_75t_SL g144 ( 
.A(n_86),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_24),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_40),
.Y(n_88)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_88),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_40),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_89),
.B(n_90),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_24),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_25),
.Y(n_91)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_91),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_27),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_92),
.B(n_101),
.Y(n_122)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_25),
.Y(n_93)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_48),
.Y(n_94)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_94),
.Y(n_115)
);

BUFx12_ASAP7_75t_L g95 ( 
.A(n_25),
.Y(n_95)
);

CKINVDCx12_ASAP7_75t_R g126 ( 
.A(n_95),
.Y(n_126)
);

BUFx4f_ASAP7_75t_L g96 ( 
.A(n_48),
.Y(n_96)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_96),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

INVx2_ASAP7_75t_SL g98 ( 
.A(n_49),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_98),
.B(n_100),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_51),
.Y(n_99)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_99),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_27),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_33),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_34),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_102),
.B(n_104),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_34),
.B(n_7),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_58),
.Y(n_124)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_35),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_91),
.A2(n_39),
.B1(n_45),
.B2(n_35),
.Y(n_105)
);

OA22x2_ASAP7_75t_L g166 ( 
.A1(n_105),
.A2(n_80),
.B1(n_79),
.B2(n_63),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_39),
.C(n_45),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_111),
.B(n_138),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_83),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_112),
.B(n_124),
.Y(n_172)
);

AOI21xp33_ASAP7_75t_L g188 ( 
.A1(n_118),
.A2(n_126),
.B(n_144),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_82),
.A2(n_38),
.B1(n_44),
.B2(n_36),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_127),
.A2(n_128),
.B1(n_129),
.B2(n_105),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_54),
.A2(n_42),
.B1(n_44),
.B2(n_37),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_103),
.B(n_37),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_137),
.B(n_147),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_100),
.B(n_38),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_100),
.B(n_42),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_152),
.B(n_86),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_94),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_154),
.B(n_72),
.Y(n_171)
);

OR2x4_ASAP7_75t_L g156 ( 
.A(n_132),
.B(n_81),
.Y(n_156)
);

OA21x2_ASAP7_75t_L g196 ( 
.A1(n_156),
.A2(n_178),
.B(n_195),
.Y(n_196)
);

A2O1A1Ixp33_ASAP7_75t_L g157 ( 
.A1(n_116),
.A2(n_43),
.B(n_47),
.C(n_98),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_157),
.B(n_158),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_134),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_128),
.A2(n_96),
.B1(n_56),
.B2(n_99),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_159),
.A2(n_188),
.B1(n_192),
.B2(n_194),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_148),
.A2(n_43),
.B1(n_76),
.B2(n_66),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_160),
.B(n_161),
.Y(n_208)
);

OAI21xp33_ASAP7_75t_L g161 ( 
.A1(n_134),
.A2(n_95),
.B(n_14),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_141),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_162),
.Y(n_221)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_107),
.Y(n_163)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_163),
.Y(n_203)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_115),
.Y(n_164)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_164),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_120),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_165),
.B(n_181),
.Y(n_201)
);

OAI21xp33_ASAP7_75t_SL g212 ( 
.A1(n_166),
.A2(n_174),
.B(n_179),
.Y(n_212)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_135),
.Y(n_168)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_168),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_169),
.B(n_170),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_108),
.B(n_12),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_171),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_113),
.A2(n_70),
.B(n_55),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_173),
.B(n_176),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_148),
.A2(n_125),
.B1(n_110),
.B2(n_123),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_141),
.Y(n_175)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_175),
.Y(n_216)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_106),
.Y(n_177)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_177),
.Y(n_218)
);

OR2x4_ASAP7_75t_L g178 ( 
.A(n_108),
.B(n_129),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_119),
.B(n_155),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_180),
.B(n_182),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_122),
.B(n_153),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_121),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_109),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_183),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_150),
.B(n_114),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_184),
.B(n_185),
.Y(n_207)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_151),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_151),
.Y(n_186)
);

INVxp33_ASAP7_75t_L g202 ( 
.A(n_186),
.Y(n_202)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_145),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_187),
.B(n_189),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_121),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_145),
.B(n_130),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_190),
.B(n_182),
.Y(n_220)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_139),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_191),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_118),
.A2(n_143),
.B1(n_123),
.B2(n_139),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_144),
.B(n_117),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_193),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_140),
.A2(n_130),
.B1(n_146),
.B2(n_133),
.Y(n_194)
);

BUFx12f_ASAP7_75t_SL g195 ( 
.A(n_130),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_176),
.B(n_136),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_197),
.B(n_219),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_156),
.A2(n_118),
.B1(n_136),
.B2(n_142),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_204),
.A2(n_210),
.B1(n_217),
.B2(n_198),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_192),
.A2(n_142),
.B1(n_149),
.B2(n_133),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_178),
.B(n_149),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_211),
.B(n_166),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_160),
.A2(n_131),
.B1(n_140),
.B2(n_166),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_157),
.B(n_131),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_220),
.B(n_161),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_207),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_225),
.B(n_226),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_214),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_227),
.B(n_231),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_201),
.B(n_167),
.Y(n_228)
);

NAND3xp33_ASAP7_75t_L g249 ( 
.A(n_228),
.B(n_232),
.C(n_233),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_197),
.A2(n_166),
.B1(n_180),
.B2(n_187),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_229),
.A2(n_227),
.B1(n_240),
.B2(n_238),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_221),
.Y(n_230)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_230),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_211),
.B(n_172),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_214),
.B(n_180),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_209),
.B(n_189),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_216),
.Y(n_234)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_234),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_235),
.B(n_196),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_223),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_236),
.Y(n_251)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_216),
.Y(n_237)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_237),
.Y(n_261)
);

OR2x4_ASAP7_75t_L g239 ( 
.A(n_196),
.B(n_195),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_239),
.A2(n_240),
.B(n_246),
.Y(n_254)
);

AND2x4_ASAP7_75t_L g240 ( 
.A(n_222),
.B(n_191),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_241),
.A2(n_243),
.B1(n_244),
.B2(n_245),
.Y(n_260)
);

INVx13_ASAP7_75t_L g242 ( 
.A(n_202),
.Y(n_242)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_242),
.Y(n_252)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_205),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_205),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_206),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_219),
.A2(n_186),
.B(n_163),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_239),
.A2(n_217),
.B(n_224),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_247),
.A2(n_256),
.B(n_208),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g269 ( 
.A(n_255),
.B(n_240),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_238),
.A2(n_196),
.B(n_246),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_241),
.A2(n_212),
.B1(n_208),
.B2(n_220),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_257),
.B(n_240),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_259),
.A2(n_262),
.B1(n_236),
.B2(n_209),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_229),
.A2(n_199),
.B1(n_208),
.B2(n_215),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_251),
.B(n_225),
.Y(n_263)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_263),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_248),
.B(n_231),
.C(n_199),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_264),
.B(n_273),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_265),
.A2(n_268),
.B(n_272),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_250),
.Y(n_266)
);

OAI322xp33_ASAP7_75t_L g283 ( 
.A1(n_266),
.A2(n_271),
.A3(n_274),
.B1(n_213),
.B2(n_252),
.C1(n_265),
.C2(n_261),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_254),
.Y(n_267)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_267),
.Y(n_276)
);

XNOR2x1_ASAP7_75t_L g275 ( 
.A(n_269),
.B(n_270),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_249),
.B(n_226),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_254),
.A2(n_200),
.B(n_222),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_248),
.B(n_222),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_258),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_268),
.A2(n_259),
.B1(n_247),
.B2(n_262),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_279),
.A2(n_281),
.B1(n_264),
.B2(n_269),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_267),
.A2(n_257),
.B1(n_260),
.B2(n_255),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_273),
.B(n_256),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_282),
.B(n_277),
.C(n_275),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_283),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_278),
.B(n_252),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_284),
.B(n_286),
.Y(n_292)
);

OA21x2_ASAP7_75t_L g294 ( 
.A1(n_285),
.A2(n_288),
.B(n_289),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_279),
.B(n_200),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_282),
.A2(n_272),
.B(n_243),
.Y(n_289)
);

BUFx24_ASAP7_75t_SL g290 ( 
.A(n_277),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_290),
.B(n_275),
.C(n_276),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_291),
.B(n_293),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_287),
.B(n_276),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_286),
.B(n_280),
.C(n_281),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_295),
.B(n_280),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_292),
.B(n_253),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_296),
.B(n_298),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_294),
.A2(n_245),
.B(n_244),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_299),
.B(n_237),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_297),
.B(n_293),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_300),
.B(n_302),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_301),
.A2(n_253),
.B(n_234),
.Y(n_303)
);

AOI322xp5_ASAP7_75t_L g306 ( 
.A1(n_303),
.A2(n_230),
.A3(n_221),
.B1(n_203),
.B2(n_162),
.C1(n_218),
.C2(n_168),
.Y(n_306)
);

A2O1A1O1Ixp25_ASAP7_75t_L g305 ( 
.A1(n_304),
.A2(n_203),
.B(n_242),
.C(n_206),
.D(n_202),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_305),
.A2(n_306),
.B1(n_175),
.B2(n_218),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_307),
.B(n_164),
.Y(n_308)
);


endmodule