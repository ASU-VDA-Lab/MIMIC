module fake_ariane_1580_n_430 (n_8, n_7, n_1, n_6, n_13, n_20, n_17, n_4, n_2, n_18, n_9, n_11, n_3, n_14, n_0, n_19, n_16, n_5, n_12, n_15, n_10, n_430);

input n_8;
input n_7;
input n_1;
input n_6;
input n_13;
input n_20;
input n_17;
input n_4;
input n_2;
input n_18;
input n_9;
input n_11;
input n_3;
input n_14;
input n_0;
input n_19;
input n_16;
input n_5;
input n_12;
input n_15;
input n_10;

output n_430;

wire n_295;
wire n_356;
wire n_170;
wire n_190;
wire n_160;
wire n_64;
wire n_180;
wire n_119;
wire n_124;
wire n_386;
wire n_307;
wire n_332;
wire n_294;
wire n_197;
wire n_176;
wire n_34;
wire n_404;
wire n_172;
wire n_347;
wire n_423;
wire n_183;
wire n_373;
wire n_299;
wire n_133;
wire n_66;
wire n_205;
wire n_341;
wire n_71;
wire n_109;
wire n_245;
wire n_421;
wire n_96;
wire n_319;
wire n_49;
wire n_416;
wire n_283;
wire n_50;
wire n_187;
wire n_367;
wire n_345;
wire n_374;
wire n_318;
wire n_103;
wire n_244;
wire n_226;
wire n_220;
wire n_261;
wire n_36;
wire n_370;
wire n_189;
wire n_286;
wire n_72;
wire n_57;
wire n_424;
wire n_387;
wire n_406;
wire n_117;
wire n_139;
wire n_85;
wire n_130;
wire n_349;
wire n_391;
wire n_346;
wire n_214;
wire n_348;
wire n_32;
wire n_410;
wire n_379;
wire n_138;
wire n_162;
wire n_264;
wire n_137;
wire n_122;
wire n_198;
wire n_232;
wire n_52;
wire n_385;
wire n_73;
wire n_327;
wire n_77;
wire n_372;
wire n_377;
wire n_396;
wire n_23;
wire n_399;
wire n_87;
wire n_279;
wire n_207;
wire n_363;
wire n_354;
wire n_41;
wire n_140;
wire n_419;
wire n_151;
wire n_28;
wire n_146;
wire n_230;
wire n_270;
wire n_194;
wire n_154;
wire n_338;
wire n_142;
wire n_285;
wire n_186;
wire n_202;
wire n_145;
wire n_193;
wire n_59;
wire n_336;
wire n_315;
wire n_311;
wire n_239;
wire n_402;
wire n_35;
wire n_272;
wire n_54;
wire n_339;
wire n_167;
wire n_90;
wire n_38;
wire n_422;
wire n_47;
wire n_153;
wire n_269;
wire n_75;
wire n_158;
wire n_69;
wire n_259;
wire n_95;
wire n_143;
wire n_152;
wire n_405;
wire n_120;
wire n_169;
wire n_106;
wire n_173;
wire n_242;
wire n_331;
wire n_320;
wire n_115;
wire n_309;
wire n_401;
wire n_267;
wire n_335;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_398;
wire n_62;
wire n_210;
wire n_200;
wire n_166;
wire n_253;
wire n_218;
wire n_79;
wire n_271;
wire n_247;
wire n_91;
wire n_240;
wire n_369;
wire n_128;
wire n_224;
wire n_44;
wire n_82;
wire n_31;
wire n_420;
wire n_222;
wire n_256;
wire n_326;
wire n_227;
wire n_48;
wire n_188;
wire n_323;
wire n_330;
wire n_400;
wire n_129;
wire n_126;
wire n_282;
wire n_328;
wire n_368;
wire n_277;
wire n_301;
wire n_248;
wire n_293;
wire n_228;
wire n_325;
wire n_276;
wire n_93;
wire n_427;
wire n_108;
wire n_303;
wire n_168;
wire n_81;
wire n_206;
wire n_352;
wire n_238;
wire n_365;
wire n_429;
wire n_136;
wire n_334;
wire n_192;
wire n_300;
wire n_163;
wire n_88;
wire n_141;
wire n_390;
wire n_104;
wire n_314;
wire n_273;
wire n_305;
wire n_312;
wire n_233;
wire n_56;
wire n_60;
wire n_388;
wire n_333;
wire n_413;
wire n_392;
wire n_376;
wire n_221;
wire n_321;
wire n_86;
wire n_361;
wire n_89;
wire n_149;
wire n_383;
wire n_237;
wire n_175;
wire n_74;
wire n_40;
wire n_181;
wire n_53;
wire n_362;
wire n_260;
wire n_310;
wire n_236;
wire n_281;
wire n_24;
wire n_209;
wire n_262;
wire n_225;
wire n_235;
wire n_297;
wire n_290;
wire n_46;
wire n_84;
wire n_371;
wire n_199;
wire n_107;
wire n_217;
wire n_178;
wire n_42;
wire n_308;
wire n_417;
wire n_201;
wire n_70;
wire n_343;
wire n_414;
wire n_287;
wire n_302;
wire n_380;
wire n_94;
wire n_284;
wire n_249;
wire n_58;
wire n_37;
wire n_65;
wire n_123;
wire n_212;
wire n_355;
wire n_278;
wire n_255;
wire n_257;
wire n_148;
wire n_135;
wire n_409;
wire n_171;
wire n_384;
wire n_61;
wire n_102;
wire n_182;
wire n_316;
wire n_196;
wire n_125;
wire n_43;
wire n_407;
wire n_27;
wire n_254;
wire n_219;
wire n_55;
wire n_231;
wire n_366;
wire n_234;
wire n_280;
wire n_215;
wire n_252;
wire n_161;
wire n_298;
wire n_68;
wire n_415;
wire n_78;
wire n_63;
wire n_99;
wire n_216;
wire n_418;
wire n_223;
wire n_403;
wire n_25;
wire n_83;
wire n_389;
wire n_288;
wire n_179;
wire n_395;
wire n_195;
wire n_213;
wire n_110;
wire n_304;
wire n_67;
wire n_306;
wire n_313;
wire n_92;
wire n_203;
wire n_378;
wire n_150;
wire n_98;
wire n_375;
wire n_113;
wire n_114;
wire n_33;
wire n_324;
wire n_337;
wire n_111;
wire n_21;
wire n_274;
wire n_296;
wire n_265;
wire n_208;
wire n_156;
wire n_292;
wire n_174;
wire n_275;
wire n_100;
wire n_132;
wire n_147;
wire n_204;
wire n_51;
wire n_76;
wire n_342;
wire n_26;
wire n_246;
wire n_428;
wire n_159;
wire n_358;
wire n_105;
wire n_30;
wire n_131;
wire n_263;
wire n_360;
wire n_229;
wire n_394;
wire n_250;
wire n_165;
wire n_144;
wire n_317;
wire n_101;
wire n_243;
wire n_134;
wire n_329;
wire n_185;
wire n_340;
wire n_289;
wire n_112;
wire n_45;
wire n_268;
wire n_266;
wire n_164;
wire n_157;
wire n_184;
wire n_177;
wire n_364;
wire n_258;
wire n_425;
wire n_118;
wire n_121;
wire n_411;
wire n_353;
wire n_22;
wire n_241;
wire n_29;
wire n_357;
wire n_412;
wire n_191;
wire n_382;
wire n_80;
wire n_211;
wire n_97;
wire n_408;
wire n_322;
wire n_251;
wire n_116;
wire n_397;
wire n_351;
wire n_39;
wire n_393;
wire n_359;
wire n_155;
wire n_127;

CKINVDCx5p33_ASAP7_75t_R g21 ( 
.A(n_18),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

CKINVDCx5p33_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx8_ASAP7_75t_SL g26 ( 
.A(n_16),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVxp67_ASAP7_75t_SL g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVxp67_ASAP7_75t_SL g35 ( 
.A(n_16),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_11),
.B(n_1),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVxp33_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_1),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_39),
.B(n_0),
.Y(n_42)
);

CKINVDCx5p33_ASAP7_75t_R g43 ( 
.A(n_26),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_2),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_3),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_3),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_5),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_39),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_43),
.Y(n_56)
);

BUFx10_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_48),
.B(n_23),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_49),
.B(n_23),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_51),
.B(n_28),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_51),
.B(n_28),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_L g68 ( 
.A1(n_51),
.A2(n_41),
.B1(n_22),
.B2(n_30),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_51),
.A2(n_28),
.B1(n_34),
.B2(n_40),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_68),
.A2(n_34),
.B1(n_50),
.B2(n_46),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_68),
.A2(n_30),
.B1(n_35),
.B2(n_32),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_70),
.A2(n_34),
.B1(n_44),
.B2(n_35),
.Y(n_75)
);

BUFx6f_ASAP7_75t_SL g76 ( 
.A(n_57),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_54),
.B(n_52),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_54),
.B(n_39),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_53),
.Y(n_80)
);

NOR2x1_ASAP7_75t_L g81 ( 
.A(n_58),
.B(n_52),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_53),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_55),
.B(n_39),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_53),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_47),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_70),
.B(n_52),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_63),
.B(n_52),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_63),
.B(n_52),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_63),
.B(n_47),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_60),
.Y(n_93)
);

AND2x4_ASAP7_75t_L g94 ( 
.A(n_61),
.B(n_32),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_64),
.A2(n_21),
.B1(n_25),
.B2(n_36),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

NAND3xp33_ASAP7_75t_SL g97 ( 
.A(n_56),
.B(n_36),
.C(n_37),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_69),
.A2(n_40),
.B1(n_37),
.B2(n_33),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_63),
.B(n_47),
.Y(n_99)
);

INVx2_ASAP7_75t_SL g100 ( 
.A(n_65),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_60),
.B(n_33),
.Y(n_101)
);

AND3x1_ASAP7_75t_L g102 ( 
.A(n_62),
.B(n_31),
.C(n_29),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_78),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_78),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g105 ( 
.A(n_74),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_78),
.B(n_69),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_72),
.B(n_79),
.Y(n_107)
);

AND3x1_ASAP7_75t_SL g108 ( 
.A(n_97),
.B(n_31),
.C(n_29),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_79),
.A2(n_62),
.B(n_67),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_74),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_72),
.B(n_67),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_96),
.B(n_57),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_82),
.Y(n_113)
);

O2A1O1Ixp33_ASAP7_75t_L g114 ( 
.A1(n_97),
.A2(n_27),
.B(n_7),
.C(n_11),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_67),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_84),
.A2(n_67),
.B(n_27),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_100),
.B(n_57),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_87),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_94),
.B(n_57),
.Y(n_119)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_76),
.Y(n_120)
);

OAI21x1_ASAP7_75t_L g121 ( 
.A1(n_80),
.A2(n_67),
.B(n_7),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_96),
.B(n_67),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_84),
.A2(n_77),
.B(n_82),
.Y(n_123)
);

AND2x6_ASAP7_75t_L g124 ( 
.A(n_88),
.B(n_96),
.Y(n_124)
);

OA22x2_ASAP7_75t_L g125 ( 
.A1(n_95),
.A2(n_73),
.B1(n_94),
.B2(n_88),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_92),
.A2(n_6),
.B(n_12),
.Y(n_126)
);

A2O1A1Ixp33_ASAP7_75t_L g127 ( 
.A1(n_73),
.A2(n_6),
.B(n_13),
.C(n_14),
.Y(n_127)
);

AND2x6_ASAP7_75t_L g128 ( 
.A(n_88),
.B(n_13),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_82),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_94),
.B(n_15),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_77),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_87),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_89),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_75),
.A2(n_15),
.B1(n_18),
.B2(n_19),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_75),
.A2(n_19),
.B1(n_102),
.B2(n_76),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_101),
.Y(n_136)
);

NOR2xp67_ASAP7_75t_L g137 ( 
.A(n_100),
.B(n_95),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_94),
.B(n_81),
.Y(n_138)
);

INVx1_ASAP7_75t_SL g139 ( 
.A(n_101),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_96),
.B(n_102),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_92),
.A2(n_99),
.B(n_80),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_99),
.B(n_89),
.Y(n_142)
);

AO32x1_ASAP7_75t_L g143 ( 
.A1(n_89),
.A2(n_93),
.A3(n_100),
.B1(n_90),
.B2(n_91),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_81),
.B(n_93),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_141),
.A2(n_83),
.B(n_85),
.Y(n_145)
);

OAI22x1_ASAP7_75t_L g146 ( 
.A1(n_105),
.A2(n_98),
.B1(n_90),
.B2(n_91),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_118),
.A2(n_132),
.B1(n_104),
.B2(n_103),
.Y(n_147)
);

O2A1O1Ixp33_ASAP7_75t_L g148 ( 
.A1(n_134),
.A2(n_93),
.B(n_98),
.C(n_85),
.Y(n_148)
);

HB1xp67_ASAP7_75t_L g149 ( 
.A(n_110),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_142),
.A2(n_86),
.B(n_83),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_139),
.B(n_119),
.Y(n_151)
);

A2O1A1Ixp33_ASAP7_75t_L g152 ( 
.A1(n_117),
.A2(n_76),
.B(n_86),
.C(n_137),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_142),
.A2(n_106),
.B(n_136),
.Y(n_153)
);

NOR2x1_ASAP7_75t_R g154 ( 
.A(n_130),
.B(n_76),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_124),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_122),
.A2(n_76),
.B(n_131),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_135),
.A2(n_125),
.B1(n_117),
.B2(n_128),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_124),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_113),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_125),
.A2(n_128),
.B1(n_107),
.B2(n_124),
.Y(n_160)
);

O2A1O1Ixp33_ASAP7_75t_SL g161 ( 
.A1(n_112),
.A2(n_140),
.B(n_122),
.C(n_127),
.Y(n_161)
);

INVx3_ASAP7_75t_SL g162 ( 
.A(n_128),
.Y(n_162)
);

A2O1A1Ixp33_ASAP7_75t_L g163 ( 
.A1(n_114),
.A2(n_127),
.B(n_140),
.C(n_131),
.Y(n_163)
);

A2O1A1Ixp33_ASAP7_75t_L g164 ( 
.A1(n_123),
.A2(n_133),
.B(n_116),
.C(n_111),
.Y(n_164)
);

O2A1O1Ixp33_ASAP7_75t_SL g165 ( 
.A1(n_126),
.A2(n_112),
.B(n_133),
.C(n_144),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_128),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_113),
.A2(n_109),
.B(n_129),
.Y(n_167)
);

A2O1A1Ixp33_ASAP7_75t_L g168 ( 
.A1(n_138),
.A2(n_115),
.B(n_129),
.C(n_121),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_128),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_124),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_129),
.A2(n_143),
.B(n_121),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_124),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_129),
.B(n_120),
.Y(n_173)
);

OA21x2_ASAP7_75t_L g174 ( 
.A1(n_143),
.A2(n_108),
.B(n_120),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_120),
.B(n_143),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_143),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_118),
.Y(n_177)
);

O2A1O1Ixp33_ASAP7_75t_SL g178 ( 
.A1(n_127),
.A2(n_114),
.B(n_126),
.C(n_112),
.Y(n_178)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_124),
.Y(n_179)
);

OAI22x1_ASAP7_75t_L g180 ( 
.A1(n_105),
.A2(n_74),
.B1(n_110),
.B2(n_73),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_145),
.A2(n_165),
.B(n_153),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_151),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_149),
.Y(n_183)
);

OA21x2_ASAP7_75t_L g184 ( 
.A1(n_171),
.A2(n_175),
.B(n_176),
.Y(n_184)
);

AO22x2_ASAP7_75t_L g185 ( 
.A1(n_160),
.A2(n_157),
.B1(n_166),
.B2(n_147),
.Y(n_185)
);

OR2x2_ASAP7_75t_L g186 ( 
.A(n_149),
.B(n_177),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_180),
.B(n_163),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_162),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_165),
.A2(n_150),
.B(n_167),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_158),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_164),
.A2(n_168),
.B(n_152),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_160),
.B(n_155),
.Y(n_192)
);

NOR2x1_ASAP7_75t_SL g193 ( 
.A(n_179),
.B(n_158),
.Y(n_193)
);

AO21x2_ASAP7_75t_L g194 ( 
.A1(n_156),
.A2(n_161),
.B(n_178),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_159),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_179),
.A2(n_162),
.B1(n_155),
.B2(n_158),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_179),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_158),
.B(n_179),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_170),
.Y(n_199)
);

OR2x2_ASAP7_75t_L g200 ( 
.A(n_172),
.B(n_146),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_169),
.A2(n_173),
.B1(n_148),
.B2(n_174),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_174),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_174),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_173),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_178),
.A2(n_73),
.B1(n_22),
.B2(n_41),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_154),
.A2(n_145),
.B(n_165),
.Y(n_206)
);

NAND2x1p5_ASAP7_75t_L g207 ( 
.A(n_179),
.B(n_158),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_151),
.B(n_139),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_151),
.B(n_74),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_159),
.Y(n_210)
);

AOI222xp33_ASAP7_75t_L g211 ( 
.A1(n_180),
.A2(n_68),
.B1(n_97),
.B2(n_127),
.C1(n_22),
.C2(n_41),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_149),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_159),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_159),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_151),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_145),
.A2(n_165),
.B(n_153),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_211),
.A2(n_205),
.B1(n_187),
.B2(n_185),
.Y(n_217)
);

OA21x2_ASAP7_75t_L g218 ( 
.A1(n_181),
.A2(n_216),
.B(n_191),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_204),
.B(n_192),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_192),
.B(n_185),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_199),
.Y(n_221)
);

BUFx8_ASAP7_75t_SL g222 ( 
.A(n_208),
.Y(n_222)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_207),
.Y(n_223)
);

AOI21x1_ASAP7_75t_L g224 ( 
.A1(n_189),
.A2(n_206),
.B(n_201),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_183),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_202),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_199),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_200),
.A2(n_202),
.B(n_203),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_205),
.A2(n_186),
.B1(n_185),
.B2(n_212),
.Y(n_229)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_207),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_202),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_195),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_195),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_210),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_209),
.B(n_182),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_200),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_210),
.Y(n_237)
);

OR2x6_ASAP7_75t_L g238 ( 
.A(n_185),
.B(n_207),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_213),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_203),
.A2(n_184),
.B(n_204),
.Y(n_240)
);

NAND4xp25_ASAP7_75t_L g241 ( 
.A(n_211),
.B(n_186),
.C(n_215),
.D(n_182),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_213),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_215),
.B(n_188),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_214),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_220),
.B(n_226),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_220),
.B(n_203),
.Y(n_246)
);

OAI211xp5_ASAP7_75t_L g247 ( 
.A1(n_217),
.A2(n_188),
.B(n_184),
.C(n_190),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_238),
.Y(n_248)
);

AND2x4_ASAP7_75t_L g249 ( 
.A(n_238),
.B(n_194),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_240),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_231),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_231),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g253 ( 
.A(n_238),
.Y(n_253)
);

AND2x4_ASAP7_75t_L g254 ( 
.A(n_238),
.B(n_194),
.Y(n_254)
);

OR2x2_ASAP7_75t_L g255 ( 
.A(n_240),
.B(n_184),
.Y(n_255)
);

AND2x4_ASAP7_75t_SL g256 ( 
.A(n_238),
.B(n_197),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_231),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_220),
.B(n_184),
.Y(n_258)
);

AOI221xp5_ASAP7_75t_L g259 ( 
.A1(n_241),
.A2(n_194),
.B1(n_196),
.B2(n_214),
.C(n_198),
.Y(n_259)
);

AND2x4_ASAP7_75t_L g260 ( 
.A(n_238),
.B(n_197),
.Y(n_260)
);

INVxp67_ASAP7_75t_SL g261 ( 
.A(n_218),
.Y(n_261)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_224),
.Y(n_262)
);

OR2x2_ASAP7_75t_L g263 ( 
.A(n_226),
.B(n_197),
.Y(n_263)
);

AO21x2_ASAP7_75t_L g264 ( 
.A1(n_224),
.A2(n_193),
.B(n_198),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_226),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_226),
.B(n_193),
.Y(n_266)
);

OAI31xp33_ASAP7_75t_L g267 ( 
.A1(n_229),
.A2(n_241),
.A3(n_217),
.B(n_235),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_224),
.A2(n_218),
.B(n_227),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_258),
.B(n_236),
.Y(n_269)
);

OR2x2_ASAP7_75t_L g270 ( 
.A(n_258),
.B(n_236),
.Y(n_270)
);

OR2x2_ASAP7_75t_L g271 ( 
.A(n_258),
.B(n_228),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_265),
.Y(n_272)
);

OR2x2_ASAP7_75t_L g273 ( 
.A(n_258),
.B(n_228),
.Y(n_273)
);

OR2x2_ASAP7_75t_L g274 ( 
.A(n_246),
.B(n_219),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_246),
.B(n_219),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_266),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_251),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g278 ( 
.A(n_266),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_246),
.B(n_238),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_246),
.B(n_227),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_265),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_266),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_250),
.B(n_221),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_251),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_245),
.B(n_221),
.Y(n_285)
);

OR2x2_ASAP7_75t_L g286 ( 
.A(n_245),
.B(n_225),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_251),
.Y(n_287)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_255),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_245),
.B(n_225),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_252),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_245),
.B(n_249),
.Y(n_291)
);

BUFx2_ASAP7_75t_L g292 ( 
.A(n_255),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_252),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_283),
.B(n_250),
.Y(n_294)
);

OR2x2_ASAP7_75t_L g295 ( 
.A(n_292),
.B(n_255),
.Y(n_295)
);

AND2x2_ASAP7_75t_SL g296 ( 
.A(n_279),
.B(n_249),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_293),
.Y(n_297)
);

AND2x4_ASAP7_75t_L g298 ( 
.A(n_291),
.B(n_249),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_291),
.B(n_254),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_272),
.Y(n_300)
);

OR2x2_ASAP7_75t_L g301 ( 
.A(n_292),
.B(n_270),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_272),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_285),
.B(n_288),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_293),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_285),
.B(n_254),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_286),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_288),
.B(n_254),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_283),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_288),
.B(n_254),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_277),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_286),
.B(n_222),
.Y(n_311)
);

INVxp67_ASAP7_75t_SL g312 ( 
.A(n_288),
.Y(n_312)
);

OR2x2_ASAP7_75t_L g313 ( 
.A(n_270),
.B(n_255),
.Y(n_313)
);

OR2x2_ASAP7_75t_L g314 ( 
.A(n_269),
.B(n_250),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_289),
.B(n_222),
.Y(n_315)
);

OR2x2_ASAP7_75t_L g316 ( 
.A(n_269),
.B(n_254),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_289),
.B(n_261),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_290),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_280),
.B(n_261),
.Y(n_319)
);

OR2x2_ASAP7_75t_L g320 ( 
.A(n_301),
.B(n_271),
.Y(n_320)
);

NAND2xp67_ASAP7_75t_L g321 ( 
.A(n_294),
.B(n_272),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_308),
.B(n_280),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_311),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_297),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_297),
.Y(n_325)
);

OR2x2_ASAP7_75t_L g326 ( 
.A(n_301),
.B(n_271),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_304),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_299),
.B(n_278),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_304),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_310),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_300),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_315),
.A2(n_259),
.B1(n_229),
.B2(n_247),
.Y(n_332)
);

OR2x2_ASAP7_75t_L g333 ( 
.A(n_306),
.B(n_273),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_299),
.B(n_278),
.Y(n_334)
);

INVx1_ASAP7_75t_SL g335 ( 
.A(n_306),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_310),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_318),
.Y(n_337)
);

OAI22xp33_ASAP7_75t_L g338 ( 
.A1(n_316),
.A2(n_259),
.B1(n_253),
.B2(n_248),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_314),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g340 ( 
.A(n_303),
.B(n_276),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_308),
.B(n_273),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_318),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_325),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_323),
.B(n_314),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_332),
.A2(n_294),
.B(n_247),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_325),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_335),
.B(n_319),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_327),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_327),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_339),
.B(n_319),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_328),
.B(n_303),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_322),
.B(n_317),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_328),
.B(n_298),
.Y(n_353)
);

OAI22xp33_ASAP7_75t_L g354 ( 
.A1(n_338),
.A2(n_316),
.B1(n_295),
.B2(n_313),
.Y(n_354)
);

INVx1_ASAP7_75t_SL g355 ( 
.A(n_333),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_331),
.Y(n_356)
);

AOI211xp5_ASAP7_75t_SL g357 ( 
.A1(n_341),
.A2(n_312),
.B(n_247),
.C(n_295),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_334),
.B(n_298),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_324),
.Y(n_359)
);

OR2x2_ASAP7_75t_L g360 ( 
.A(n_333),
.B(n_313),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_320),
.B(n_317),
.Y(n_361)
);

AOI31xp33_ASAP7_75t_L g362 ( 
.A1(n_320),
.A2(n_259),
.A3(n_309),
.B(n_307),
.Y(n_362)
);

HB1xp67_ASAP7_75t_L g363 ( 
.A(n_321),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_345),
.B(n_321),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_354),
.A2(n_296),
.B1(n_235),
.B2(n_298),
.Y(n_365)
);

AOI21xp33_ASAP7_75t_L g366 ( 
.A1(n_362),
.A2(n_342),
.B(n_330),
.Y(n_366)
);

OAI221xp5_ASAP7_75t_L g367 ( 
.A1(n_357),
.A2(n_267),
.B1(n_326),
.B2(n_331),
.C(n_337),
.Y(n_367)
);

OAI221xp5_ASAP7_75t_SL g368 ( 
.A1(n_355),
.A2(n_267),
.B1(n_326),
.B2(n_305),
.C(n_334),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_344),
.B(n_336),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_SL g370 ( 
.A1(n_362),
.A2(n_267),
.B(n_340),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_359),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_360),
.A2(n_298),
.B1(n_296),
.B2(n_340),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_363),
.A2(n_296),
.B1(n_275),
.B2(n_243),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_352),
.B(n_329),
.Y(n_374)
);

OAI221xp5_ASAP7_75t_L g375 ( 
.A1(n_355),
.A2(n_275),
.B1(n_274),
.B2(n_243),
.C(n_282),
.Y(n_375)
);

AOI222xp33_ASAP7_75t_L g376 ( 
.A1(n_347),
.A2(n_249),
.B1(n_254),
.B2(n_279),
.C1(n_248),
.C2(n_253),
.Y(n_376)
);

AOI221xp5_ASAP7_75t_L g377 ( 
.A1(n_350),
.A2(n_305),
.B1(n_261),
.B2(n_300),
.C(n_302),
.Y(n_377)
);

OAI211xp5_ASAP7_75t_L g378 ( 
.A1(n_361),
.A2(n_268),
.B(n_262),
.C(n_309),
.Y(n_378)
);

NAND4xp25_ASAP7_75t_L g379 ( 
.A(n_359),
.B(n_268),
.C(n_262),
.D(n_307),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_360),
.A2(n_254),
.B1(n_249),
.B2(n_274),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_SL g381 ( 
.A(n_353),
.B(n_249),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_L g382 ( 
.A1(n_343),
.A2(n_302),
.B(n_300),
.Y(n_382)
);

AOI211xp5_ASAP7_75t_L g383 ( 
.A1(n_366),
.A2(n_343),
.B(n_346),
.C(n_348),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_370),
.A2(n_356),
.B1(n_348),
.B2(n_346),
.Y(n_384)
);

AOI221xp5_ASAP7_75t_L g385 ( 
.A1(n_368),
.A2(n_349),
.B1(n_356),
.B2(n_351),
.C(n_249),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_374),
.B(n_349),
.Y(n_386)
);

AOI221xp5_ASAP7_75t_L g387 ( 
.A1(n_364),
.A2(n_351),
.B1(n_358),
.B2(n_353),
.C(n_268),
.Y(n_387)
);

AOI211xp5_ASAP7_75t_SL g388 ( 
.A1(n_378),
.A2(n_358),
.B(n_262),
.C(n_290),
.Y(n_388)
);

AOI211x1_ASAP7_75t_SL g389 ( 
.A1(n_379),
.A2(n_302),
.B(n_281),
.C(n_262),
.Y(n_389)
);

AOI221xp5_ASAP7_75t_L g390 ( 
.A1(n_367),
.A2(n_287),
.B1(n_284),
.B2(n_277),
.C(n_253),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_L g391 ( 
.A1(n_365),
.A2(n_287),
.B(n_284),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_377),
.A2(n_374),
.B(n_369),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_371),
.B(n_262),
.Y(n_393)
);

AOI211xp5_ASAP7_75t_L g394 ( 
.A1(n_372),
.A2(n_262),
.B(n_253),
.C(n_248),
.Y(n_394)
);

O2A1O1Ixp33_ASAP7_75t_L g395 ( 
.A1(n_375),
.A2(n_262),
.B(n_218),
.C(n_264),
.Y(n_395)
);

INVx1_ASAP7_75t_SL g396 ( 
.A(n_373),
.Y(n_396)
);

NOR2xp67_ASAP7_75t_L g397 ( 
.A(n_384),
.B(n_382),
.Y(n_397)
);

AOI221xp5_ASAP7_75t_SL g398 ( 
.A1(n_392),
.A2(n_381),
.B1(n_376),
.B2(n_380),
.C(n_281),
.Y(n_398)
);

NAND5xp2_ASAP7_75t_L g399 ( 
.A(n_388),
.B(n_266),
.C(n_244),
.D(n_232),
.E(n_234),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_386),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_396),
.B(n_281),
.Y(n_401)
);

NAND3xp33_ASAP7_75t_L g402 ( 
.A(n_383),
.B(n_218),
.C(n_242),
.Y(n_402)
);

OAI211xp5_ASAP7_75t_SL g403 ( 
.A1(n_389),
.A2(n_242),
.B(n_244),
.C(n_239),
.Y(n_403)
);

NAND3xp33_ASAP7_75t_SL g404 ( 
.A(n_385),
.B(n_263),
.C(n_239),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_401),
.Y(n_405)
);

XOR2x2_ASAP7_75t_L g406 ( 
.A(n_398),
.B(n_390),
.Y(n_406)
);

NOR3xp33_ASAP7_75t_L g407 ( 
.A(n_402),
.B(n_395),
.C(n_387),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_397),
.A2(n_391),
.B1(n_394),
.B2(n_393),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_400),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_403),
.Y(n_410)
);

OAI211xp5_ASAP7_75t_SL g411 ( 
.A1(n_399),
.A2(n_237),
.B(n_234),
.C(n_233),
.Y(n_411)
);

NOR3xp33_ASAP7_75t_L g412 ( 
.A(n_404),
.B(n_237),
.C(n_233),
.Y(n_412)
);

INVx3_ASAP7_75t_L g413 ( 
.A(n_409),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_406),
.A2(n_253),
.B1(n_248),
.B2(n_260),
.Y(n_414)
);

AND3x4_ASAP7_75t_L g415 ( 
.A(n_407),
.B(n_248),
.C(n_260),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_410),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_412),
.Y(n_417)
);

OR3x1_ASAP7_75t_L g418 ( 
.A(n_411),
.B(n_232),
.C(n_257),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_413),
.B(n_408),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_416),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_416),
.Y(n_421)
);

INVx4_ASAP7_75t_L g422 ( 
.A(n_417),
.Y(n_422)
);

OR2x2_ASAP7_75t_L g423 ( 
.A(n_422),
.B(n_419),
.Y(n_423)
);

OAI22x1_ASAP7_75t_L g424 ( 
.A1(n_422),
.A2(n_414),
.B1(n_415),
.B2(n_405),
.Y(n_424)
);

OAI22x1_ASAP7_75t_L g425 ( 
.A1(n_420),
.A2(n_418),
.B1(n_218),
.B2(n_260),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_423),
.B(n_421),
.Y(n_426)
);

OAI21x1_ASAP7_75t_L g427 ( 
.A1(n_424),
.A2(n_230),
.B(n_223),
.Y(n_427)
);

OAI21xp33_ASAP7_75t_L g428 ( 
.A1(n_426),
.A2(n_425),
.B(n_256),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_428),
.Y(n_429)
);

AOI22xp33_ASAP7_75t_SL g430 ( 
.A1(n_429),
.A2(n_427),
.B1(n_264),
.B2(n_256),
.Y(n_430)
);


endmodule