module fake_jpeg_14935_n_355 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_355);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_355;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_20),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_5),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_9),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_11),
.Y(n_45)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx6_ASAP7_75t_SL g48 ( 
.A(n_22),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_48),
.B(n_26),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_11),
.Y(n_49)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_0),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_50),
.B(n_40),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_57),
.A2(n_37),
.B1(n_32),
.B2(n_28),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_62),
.A2(n_85),
.B1(n_59),
.B2(n_37),
.Y(n_92)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_66),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_57),
.A2(n_44),
.B1(n_43),
.B2(n_25),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_69),
.A2(n_33),
.B1(n_39),
.B2(n_23),
.Y(n_101)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_45),
.B(n_29),
.C(n_42),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_73),
.B(n_88),
.Y(n_107)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_55),
.Y(n_94)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_84),
.B(n_50),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_59),
.A2(n_37),
.B1(n_33),
.B2(n_39),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_86),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_49),
.B(n_61),
.C(n_60),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_89),
.B(n_109),
.Y(n_127)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_91),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_92),
.A2(n_93),
.B1(n_105),
.B2(n_116),
.Y(n_152)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_94),
.Y(n_134)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_96),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_63),
.A2(n_56),
.B1(n_54),
.B2(n_46),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_97),
.A2(n_112),
.B1(n_120),
.B2(n_34),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_65),
.B(n_40),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_99),
.B(n_106),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_33),
.Y(n_100)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_100),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_104),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_102),
.B(n_110),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_68),
.A2(n_36),
.B1(n_23),
.B2(n_41),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_68),
.A2(n_39),
.B1(n_54),
.B2(n_46),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_79),
.B(n_51),
.Y(n_106)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_70),
.Y(n_108)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_108),
.Y(n_149)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_83),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_77),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_73),
.B(n_51),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_111),
.B(n_31),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_64),
.A2(n_48),
.B1(n_47),
.B2(n_36),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_74),
.Y(n_113)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_113),
.Y(n_125)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_74),
.Y(n_114)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_114),
.Y(n_144)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_87),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_115),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_81),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_64),
.B(n_41),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_117),
.B(n_121),
.Y(n_140)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_70),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_118),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_72),
.A2(n_47),
.B1(n_31),
.B2(n_43),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_71),
.B(n_35),
.Y(n_121)
);

INVx2_ASAP7_75t_SL g122 ( 
.A(n_96),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_122),
.Y(n_172)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_119),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_123),
.Y(n_171)
);

OAI22xp33_ASAP7_75t_L g124 ( 
.A1(n_111),
.A2(n_71),
.B1(n_82),
.B2(n_76),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_124),
.A2(n_112),
.B1(n_90),
.B2(n_120),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_130),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_100),
.A2(n_21),
.B(n_44),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_131),
.A2(n_133),
.B(n_137),
.Y(n_173)
);

BUFx24_ASAP7_75t_SL g132 ( 
.A(n_89),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_132),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_104),
.Y(n_133)
);

MAJx2_ASAP7_75t_L g135 ( 
.A(n_107),
.B(n_42),
.C(n_81),
.Y(n_135)
);

MAJx2_ASAP7_75t_L g170 ( 
.A(n_135),
.B(n_29),
.C(n_42),
.Y(n_170)
);

OAI21xp33_ASAP7_75t_L g137 ( 
.A1(n_99),
.A2(n_31),
.B(n_35),
.Y(n_137)
);

INVx3_ASAP7_75t_SL g138 ( 
.A(n_93),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_138),
.A2(n_139),
.B1(n_146),
.B2(n_147),
.Y(n_174)
);

INVx4_ASAP7_75t_SL g139 ( 
.A(n_108),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_95),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_141),
.B(n_121),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_107),
.B(n_30),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_142),
.B(n_153),
.C(n_94),
.Y(n_157)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_119),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_118),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_150),
.B(n_101),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_107),
.B(n_75),
.C(n_67),
.Y(n_153)
);

XOR2x2_ASAP7_75t_L g154 ( 
.A(n_135),
.B(n_107),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_154),
.A2(n_170),
.B(n_134),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_151),
.A2(n_97),
.B1(n_106),
.B2(n_108),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_155),
.A2(n_159),
.B1(n_160),
.B2(n_163),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_157),
.B(n_162),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_158),
.B(n_166),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_150),
.A2(n_109),
.B1(n_103),
.B2(n_95),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_153),
.A2(n_103),
.B1(n_114),
.B2(n_113),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_136),
.A2(n_90),
.B1(n_96),
.B2(n_98),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_136),
.A2(n_91),
.B1(n_119),
.B2(n_117),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_164),
.A2(n_165),
.B1(n_168),
.B2(n_149),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_152),
.A2(n_91),
.B1(n_93),
.B2(n_76),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_142),
.B(n_115),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_167),
.B(n_169),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_124),
.A2(n_116),
.B1(n_75),
.B2(n_25),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_127),
.B(n_31),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_154),
.A2(n_129),
.B(n_131),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_175),
.A2(n_187),
.B(n_192),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_166),
.B(n_140),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_176),
.B(n_193),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_178),
.A2(n_179),
.B(n_183),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_154),
.A2(n_149),
.B(n_147),
.Y(n_179)
);

AO22x1_ASAP7_75t_L g180 ( 
.A1(n_161),
.A2(n_130),
.B1(n_122),
.B2(n_123),
.Y(n_180)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_180),
.Y(n_212)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_172),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_181),
.B(n_185),
.Y(n_204)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_172),
.Y(n_184)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_184),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_169),
.Y(n_185)
);

A2O1A1Ixp33_ASAP7_75t_SL g186 ( 
.A1(n_155),
.A2(n_145),
.B(n_129),
.C(n_139),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_186),
.A2(n_171),
.B(n_172),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_161),
.A2(n_146),
.B1(n_143),
.B2(n_148),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_174),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_190),
.B(n_168),
.Y(n_215)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_159),
.Y(n_191)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_191),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_173),
.A2(n_143),
.B(n_148),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_162),
.B(n_167),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_162),
.B(n_128),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_194),
.B(n_164),
.Y(n_209)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_174),
.Y(n_195)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_195),
.Y(n_219)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_174),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_196),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_182),
.B(n_157),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_198),
.B(n_203),
.C(n_211),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_195),
.A2(n_196),
.B1(n_191),
.B2(n_177),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_200),
.A2(n_201),
.B1(n_206),
.B2(n_220),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_177),
.A2(n_157),
.B1(n_160),
.B2(n_170),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_182),
.B(n_170),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_186),
.A2(n_158),
.B1(n_165),
.B2(n_173),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_184),
.Y(n_207)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_207),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_209),
.B(n_220),
.Y(n_242)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_187),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_210),
.B(n_214),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_183),
.B(n_163),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_176),
.B(n_156),
.Y(n_214)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_215),
.Y(n_228)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_216),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_187),
.Y(n_217)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_217),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_193),
.B(n_122),
.C(n_126),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_218),
.B(n_223),
.C(n_192),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_186),
.A2(n_125),
.B1(n_144),
.B2(n_128),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_188),
.B(n_144),
.Y(n_221)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_221),
.Y(n_234)
);

OA21x2_ASAP7_75t_L g222 ( 
.A1(n_186),
.A2(n_125),
.B(n_138),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_222),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_179),
.B(n_30),
.Y(n_223)
);

NAND3xp33_ASAP7_75t_L g226 ( 
.A(n_205),
.B(n_185),
.C(n_175),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_226),
.B(n_213),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_221),
.B(n_188),
.Y(n_229)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_229),
.Y(n_250)
);

INVx2_ASAP7_75t_SL g231 ( 
.A(n_207),
.Y(n_231)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_231),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_222),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_233),
.B(n_227),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_203),
.B(n_194),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_237),
.B(n_240),
.C(n_241),
.Y(n_255)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_204),
.Y(n_238)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_238),
.Y(n_265)
);

BUFx2_ASAP7_75t_L g239 ( 
.A(n_197),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_239),
.B(n_181),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_198),
.B(n_175),
.C(n_189),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_242),
.B(n_180),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_218),
.B(n_189),
.C(n_178),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_243),
.B(n_245),
.C(n_247),
.Y(n_267)
);

INVx2_ASAP7_75t_SL g244 ( 
.A(n_222),
.Y(n_244)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_244),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_201),
.B(n_178),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_202),
.Y(n_246)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_246),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_211),
.B(n_186),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_223),
.B(n_186),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_248),
.B(n_180),
.C(n_181),
.Y(n_271)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_202),
.Y(n_249)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_249),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_251),
.A2(n_254),
.B1(n_261),
.B2(n_247),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_225),
.B(n_205),
.Y(n_252)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_252),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_213),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_253),
.B(n_257),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_244),
.A2(n_212),
.B1(n_210),
.B2(n_209),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_235),
.B(n_216),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_230),
.A2(n_212),
.B1(n_199),
.B2(n_219),
.Y(n_258)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_258),
.Y(n_278)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_259),
.Y(n_282)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_260),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_233),
.A2(n_208),
.B1(n_206),
.B2(n_200),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_229),
.B(n_180),
.Y(n_262)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_262),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_234),
.B(n_228),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_263),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_264),
.B(n_271),
.Y(n_291)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_231),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_270),
.B(n_239),
.Y(n_280)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_224),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_272),
.B(n_248),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_266),
.A2(n_232),
.B(n_236),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_274),
.A2(n_283),
.B(n_254),
.Y(n_293)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_275),
.Y(n_301)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_279),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_280),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_255),
.B(n_237),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_281),
.B(n_288),
.C(n_290),
.Y(n_296)
);

XOR2x2_ASAP7_75t_L g283 ( 
.A(n_264),
.B(n_242),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_265),
.B(n_243),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_285),
.B(n_257),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_269),
.A2(n_241),
.B1(n_245),
.B2(n_236),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_286),
.A2(n_271),
.B1(n_262),
.B2(n_260),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_250),
.B(n_240),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_287),
.B(n_263),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_255),
.B(n_30),
.C(n_26),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_267),
.B(n_26),
.Y(n_290)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_292),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_293),
.A2(n_294),
.B1(n_297),
.B2(n_34),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_284),
.A2(n_269),
.B1(n_268),
.B2(n_256),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_281),
.B(n_267),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_295),
.B(n_253),
.C(n_258),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_282),
.B(n_277),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_299),
.B(n_302),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_278),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_300),
.B(n_250),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_276),
.B(n_272),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_304),
.B(n_307),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_287),
.B(n_273),
.C(n_291),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_305),
.B(n_306),
.C(n_296),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_273),
.B(n_291),
.C(n_290),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_286),
.B(n_261),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_308),
.B(n_312),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_301),
.A2(n_283),
.B1(n_278),
.B2(n_289),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_309),
.B(n_314),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_297),
.A2(n_294),
.B(n_274),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_310),
.A2(n_306),
.B1(n_298),
.B2(n_27),
.Y(n_322)
);

OR2x2_ASAP7_75t_L g312 ( 
.A(n_303),
.B(n_279),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_295),
.B(n_288),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_313),
.B(n_317),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_305),
.A2(n_256),
.B(n_21),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_318),
.A2(n_319),
.B1(n_316),
.B2(n_314),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_296),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_320),
.B(n_0),
.Y(n_330)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_322),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_315),
.B(n_156),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_323),
.B(n_325),
.Y(n_334)
);

OR2x2_ASAP7_75t_L g339 ( 
.A(n_324),
.B(n_328),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_311),
.A2(n_27),
.B1(n_11),
.B2(n_12),
.Y(n_325)
);

AOI21x1_ASAP7_75t_L g328 ( 
.A1(n_312),
.A2(n_10),
.B(n_19),
.Y(n_328)
);

OAI21x1_ASAP7_75t_SL g329 ( 
.A1(n_309),
.A2(n_10),
.B(n_19),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_329),
.A2(n_330),
.B(n_12),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_319),
.B(n_320),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_331),
.B(n_13),
.Y(n_335)
);

OAI321xp33_ASAP7_75t_L g341 ( 
.A1(n_332),
.A2(n_340),
.A3(n_8),
.B1(n_20),
.B2(n_17),
.C(n_4),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_321),
.B(n_9),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_333),
.B(n_338),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_335),
.B(n_336),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_324),
.B(n_13),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_327),
.B(n_328),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_326),
.A2(n_13),
.B(n_18),
.Y(n_340)
);

OAI321xp33_ASAP7_75t_L g348 ( 
.A1(n_341),
.A2(n_345),
.A3(n_4),
.B1(n_5),
.B2(n_15),
.C(n_20),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_333),
.B(n_326),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_342),
.A2(n_344),
.B1(n_343),
.B2(n_5),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_337),
.A2(n_8),
.B(n_17),
.Y(n_345)
);

AOI31xp33_ASAP7_75t_L g346 ( 
.A1(n_339),
.A2(n_6),
.A3(n_17),
.B(n_16),
.Y(n_346)
);

AOI31xp33_ASAP7_75t_L g347 ( 
.A1(n_346),
.A2(n_334),
.A3(n_6),
.B(n_14),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_347),
.B(n_348),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_349),
.B(n_4),
.Y(n_350)
);

OAI321xp33_ASAP7_75t_L g352 ( 
.A1(n_350),
.A2(n_1),
.A3(n_2),
.B1(n_3),
.B2(n_15),
.C(n_351),
.Y(n_352)
);

OAI221xp5_ASAP7_75t_L g353 ( 
.A1(n_352),
.A2(n_1),
.B1(n_3),
.B2(n_351),
.C(n_328),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_353),
.B(n_1),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_354),
.B(n_1),
.Y(n_355)
);


endmodule