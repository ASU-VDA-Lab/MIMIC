module fake_ibex_674_n_944 (n_151, n_147, n_85, n_167, n_128, n_84, n_64, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_177, n_148, n_2, n_76, n_8, n_118, n_67, n_9, n_164, n_38, n_124, n_37, n_110, n_47, n_169, n_108, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_172, n_49, n_40, n_66, n_17, n_74, n_90, n_176, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_166, n_163, n_26, n_114, n_34, n_97, n_102, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_156, n_126, n_1, n_154, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_50, n_11, n_92, n_144, n_170, n_101, n_113, n_138, n_96, n_68, n_117, n_79, n_81, n_35, n_159, n_158, n_132, n_174, n_157, n_160, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_944);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_177;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_67;
input n_9;
input n_164;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_169;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_172;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_176;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_166;
input n_163;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_1;
input n_154;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_50;
input n_11;
input n_92;
input n_144;
input n_170;
input n_101;
input n_113;
input n_138;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_159;
input n_158;
input n_132;
input n_174;
input n_157;
input n_160;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_944;

wire n_599;
wire n_822;
wire n_778;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_707;
wire n_273;
wire n_309;
wire n_330;
wire n_926;
wire n_328;
wire n_372;
wire n_293;
wire n_341;
wire n_256;
wire n_418;
wire n_193;
wire n_510;
wire n_845;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_790;
wire n_920;
wire n_452;
wire n_664;
wire n_255;
wire n_586;
wire n_773;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_191;
wire n_873;
wire n_593;
wire n_862;
wire n_545;
wire n_909;
wire n_583;
wire n_887;
wire n_678;
wire n_663;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_357;
wire n_457;
wire n_412;
wire n_494;
wire n_226;
wire n_930;
wire n_336;
wire n_258;
wire n_861;
wire n_449;
wire n_547;
wire n_727;
wire n_216;
wire n_915;
wire n_911;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_698;
wire n_280;
wire n_317;
wire n_340;
wire n_375;
wire n_708;
wire n_901;
wire n_187;
wire n_667;
wire n_884;
wire n_682;
wire n_850;
wire n_182;
wire n_196;
wire n_326;
wire n_327;
wire n_879;
wire n_723;
wire n_270;
wire n_383;
wire n_346;
wire n_886;
wire n_840;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_859;
wire n_259;
wire n_339;
wire n_276;
wire n_470;
wire n_770;
wire n_210;
wire n_348;
wire n_220;
wire n_875;
wire n_941;
wire n_674;
wire n_481;
wire n_243;
wire n_497;
wire n_287;
wire n_671;
wire n_228;
wire n_711;
wire n_876;
wire n_552;
wire n_384;
wire n_251;
wire n_632;
wire n_373;
wire n_854;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_936;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_939;
wire n_453;
wire n_591;
wire n_898;
wire n_655;
wire n_333;
wire n_928;
wire n_400;
wire n_306;
wire n_550;
wire n_736;
wire n_673;
wire n_732;
wire n_798;
wire n_832;
wire n_278;
wire n_242;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_914;
wire n_835;
wire n_526;
wire n_785;
wire n_824;
wire n_929;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_923;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_933;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_938;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_281;
wire n_758;
wire n_594;
wire n_636;
wire n_720;
wire n_710;
wire n_490;
wire n_407;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_543;
wire n_420;
wire n_483;
wire n_580;
wire n_769;
wire n_487;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_765;
wire n_849;
wire n_857;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_917;
wire n_185;
wire n_388;
wire n_625;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_931;
wire n_666;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_207;
wire n_922;
wire n_438;
wire n_851;
wire n_689;
wire n_793;
wire n_676;
wire n_937;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_488;
wire n_514;
wire n_705;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_635;
wire n_844;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_847;
wire n_830;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_826;
wire n_299;
wire n_433;
wire n_439;
wire n_262;
wire n_704;
wire n_924;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_696;
wire n_837;
wire n_796;
wire n_797;
wire n_477;
wire n_640;
wire n_363;
wire n_402;
wire n_725;
wire n_180;
wire n_369;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_935;
wire n_869;
wire n_925;
wire n_718;
wire n_801;
wire n_918;
wire n_672;
wire n_722;
wire n_401;
wire n_554;
wire n_553;
wire n_735;
wire n_305;
wire n_882;
wire n_942;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_605;
wire n_539;
wire n_354;
wire n_206;
wire n_392;
wire n_630;
wire n_516;
wire n_548;
wire n_567;
wire n_943;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_940;
wire n_188;
wire n_200;
wire n_444;
wire n_506;
wire n_562;
wire n_564;
wire n_868;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_927;
wire n_934;
wire n_658;
wire n_512;
wire n_615;
wire n_685;
wire n_283;
wire n_366;
wire n_397;
wire n_894;
wire n_803;
wire n_692;
wire n_627;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_757;
wire n_248;
wire n_702;
wire n_451;
wire n_712;
wire n_190;
wire n_906;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_818;
wire n_653;
wire n_214;
wire n_238;
wire n_579;
wire n_899;
wire n_843;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_919;
wire n_780;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_288;
wire n_285;
wire n_247;
wire n_320;
wire n_379;
wire n_551;
wire n_612;
wire n_318;
wire n_291;
wire n_819;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_858;
wire n_342;
wire n_233;
wire n_414;
wire n_385;
wire n_430;
wire n_741;
wire n_729;
wire n_603;
wire n_378;
wire n_486;
wire n_422;
wire n_264;
wire n_198;
wire n_616;
wire n_782;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_820;
wire n_670;
wire n_805;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_808;
wire n_250;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_903;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_885;
wire n_513;
wire n_212;
wire n_588;
wire n_877;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_896;
wire n_197;
wire n_528;
wire n_181;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_794;
wire n_836;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_572;
wire n_867;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_897;
wire n_889;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_697;
wire n_874;
wire n_816;
wire n_890;
wire n_912;
wire n_921;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_213;
wire n_424;
wire n_565;
wire n_916;
wire n_823;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_394;
wire n_364;
wire n_687;
wire n_895;
wire n_298;
wire n_202;
wire n_231;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_932;
wire n_657;
wire n_764;
wire n_184;
wire n_492;
wire n_649;
wire n_855;
wire n_812;
wire n_232;
wire n_380;
wire n_749;
wire n_866;
wire n_559;
wire n_425;

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_178),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_168),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_61),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_169),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_114),
.Y(n_184)
);

BUFx2_ASAP7_75t_L g185 ( 
.A(n_72),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_131),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_76),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_167),
.Y(n_188)
);

NOR2xp67_ASAP7_75t_L g189 ( 
.A(n_89),
.B(n_173),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_16),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_137),
.Y(n_191)
);

INVx2_ASAP7_75t_SL g192 ( 
.A(n_117),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_95),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_60),
.Y(n_194)
);

INVxp33_ASAP7_75t_L g195 ( 
.A(n_106),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_133),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_26),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_62),
.B(n_148),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_47),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_123),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_113),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_165),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_115),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_3),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_30),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_138),
.Y(n_206)
);

INVxp67_ASAP7_75t_SL g207 ( 
.A(n_150),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_166),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_139),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_25),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_26),
.Y(n_211)
);

INVxp33_ASAP7_75t_SL g212 ( 
.A(n_34),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_81),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_145),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_109),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_177),
.Y(n_216)
);

INVxp67_ASAP7_75t_SL g217 ( 
.A(n_55),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_155),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_110),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_102),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_172),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_90),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_40),
.Y(n_223)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_136),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_158),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_68),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_157),
.Y(n_227)
);

NOR2xp67_ASAP7_75t_L g228 ( 
.A(n_39),
.B(n_111),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_126),
.Y(n_229)
);

OR2x2_ASAP7_75t_L g230 ( 
.A(n_156),
.B(n_49),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_96),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_163),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_57),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_7),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_121),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_105),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_130),
.Y(n_237)
);

NOR2xp67_ASAP7_75t_L g238 ( 
.A(n_143),
.B(n_84),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_77),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_103),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_107),
.Y(n_241)
);

NOR2xp67_ASAP7_75t_L g242 ( 
.A(n_170),
.B(n_104),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g243 ( 
.A(n_63),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_128),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_48),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_52),
.Y(n_246)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_45),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_19),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_8),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_152),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_119),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_116),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_41),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_162),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_3),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_65),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_18),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_127),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_12),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_174),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_175),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_100),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_36),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_80),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_171),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_88),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_93),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_9),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_8),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_161),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_159),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_118),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_59),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_179),
.Y(n_274)
);

INVxp67_ASAP7_75t_SL g275 ( 
.A(n_9),
.Y(n_275)
);

INVxp67_ASAP7_75t_SL g276 ( 
.A(n_98),
.Y(n_276)
);

AND2x4_ASAP7_75t_L g277 ( 
.A(n_67),
.B(n_134),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_124),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_132),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_10),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_160),
.Y(n_281)
);

INVxp67_ASAP7_75t_SL g282 ( 
.A(n_82),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_53),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_5),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_140),
.Y(n_285)
);

BUFx3_ASAP7_75t_L g286 ( 
.A(n_176),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_149),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_13),
.Y(n_288)
);

BUFx3_ASAP7_75t_L g289 ( 
.A(n_122),
.Y(n_289)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_31),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_74),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_87),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_125),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_92),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_135),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_112),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_54),
.Y(n_297)
);

INVx2_ASAP7_75t_SL g298 ( 
.A(n_17),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_142),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_1),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_22),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_25),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_2),
.Y(n_303)
);

BUFx2_ASAP7_75t_SL g304 ( 
.A(n_99),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_31),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_79),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_56),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_85),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_27),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_94),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_108),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_129),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_91),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_153),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_272),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_224),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_204),
.B(n_0),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_224),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_224),
.Y(n_319)
);

AND2x4_ASAP7_75t_L g320 ( 
.A(n_290),
.B(n_247),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_195),
.B(n_0),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_288),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_322)
);

BUFx8_ASAP7_75t_L g323 ( 
.A(n_185),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_195),
.B(n_4),
.Y(n_324)
);

BUFx2_ASAP7_75t_L g325 ( 
.A(n_290),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_290),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_247),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_247),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_209),
.B(n_6),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_184),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_184),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_244),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_272),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_222),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_267),
.Y(n_335)
);

CKINVDCx6p67_ASAP7_75t_R g336 ( 
.A(n_261),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_272),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_244),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_298),
.B(n_11),
.Y(n_339)
);

AND2x4_ASAP7_75t_L g340 ( 
.A(n_257),
.B(n_11),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_272),
.Y(n_341)
);

INVx3_ASAP7_75t_L g342 ( 
.A(n_257),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_268),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_268),
.Y(n_344)
);

AND2x6_ASAP7_75t_L g345 ( 
.A(n_277),
.B(n_69),
.Y(n_345)
);

AND2x4_ASAP7_75t_L g346 ( 
.A(n_192),
.B(n_13),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_183),
.Y(n_347)
);

CKINVDCx11_ASAP7_75t_R g348 ( 
.A(n_248),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_190),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_197),
.Y(n_350)
);

INVx6_ASAP7_75t_L g351 ( 
.A(n_277),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_205),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_210),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_186),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_243),
.Y(n_355)
);

BUFx3_ASAP7_75t_L g356 ( 
.A(n_243),
.Y(n_356)
);

HB1xp67_ASAP7_75t_L g357 ( 
.A(n_288),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_212),
.B(n_14),
.Y(n_358)
);

AND2x4_ASAP7_75t_L g359 ( 
.A(n_277),
.B(n_15),
.Y(n_359)
);

HB1xp67_ASAP7_75t_L g360 ( 
.A(n_300),
.Y(n_360)
);

INVx3_ASAP7_75t_L g361 ( 
.A(n_211),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_212),
.B(n_252),
.Y(n_362)
);

HB1xp67_ASAP7_75t_L g363 ( 
.A(n_302),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_270),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_302),
.B(n_15),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_186),
.A2(n_16),
.B1(n_17),
.B2(n_19),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_215),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_270),
.B(n_20),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_234),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_249),
.B(n_255),
.Y(n_370)
);

INVx3_ASAP7_75t_L g371 ( 
.A(n_259),
.Y(n_371)
);

AND2x4_ASAP7_75t_L g372 ( 
.A(n_246),
.B(n_286),
.Y(n_372)
);

AND2x2_ASAP7_75t_SL g373 ( 
.A(n_230),
.B(n_75),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_263),
.Y(n_374)
);

INVx3_ASAP7_75t_L g375 ( 
.A(n_280),
.Y(n_375)
);

BUFx12f_ASAP7_75t_L g376 ( 
.A(n_180),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_284),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_246),
.B(n_21),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_289),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_248),
.Y(n_380)
);

AOI22xp33_ASAP7_75t_SL g381 ( 
.A1(n_269),
.A2(n_23),
.B1(n_24),
.B2(n_27),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_289),
.B(n_23),
.Y(n_382)
);

AND2x4_ASAP7_75t_L g383 ( 
.A(n_285),
.B(n_24),
.Y(n_383)
);

AND2x4_ASAP7_75t_L g384 ( 
.A(n_297),
.B(n_28),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_297),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_301),
.B(n_29),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_181),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_182),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_303),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_305),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.Y(n_390)
);

AND2x4_ASAP7_75t_L g391 ( 
.A(n_309),
.B(n_32),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_187),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_215),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_180),
.B(n_33),
.Y(n_394)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_202),
.B(n_34),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_188),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_191),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_193),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_194),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_196),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_199),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_200),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_201),
.B(n_35),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_203),
.Y(n_404)
);

AND2x4_ASAP7_75t_L g405 ( 
.A(n_206),
.B(n_35),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_213),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_214),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_216),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_366),
.A2(n_269),
.B1(n_314),
.B2(n_236),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_340),
.Y(n_410)
);

BUFx4f_ASAP7_75t_L g411 ( 
.A(n_359),
.Y(n_411)
);

INVxp67_ASAP7_75t_SL g412 ( 
.A(n_321),
.Y(n_412)
);

OR2x6_ASAP7_75t_L g413 ( 
.A(n_376),
.B(n_304),
.Y(n_413)
);

INVxp67_ASAP7_75t_SL g414 ( 
.A(n_321),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_325),
.B(n_202),
.Y(n_415)
);

INVxp33_ASAP7_75t_L g416 ( 
.A(n_357),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_383),
.Y(n_417)
);

AND2x6_ASAP7_75t_L g418 ( 
.A(n_359),
.B(n_198),
.Y(n_418)
);

INVx4_ASAP7_75t_L g419 ( 
.A(n_345),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_334),
.B(n_335),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_347),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_383),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_336),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_320),
.B(n_218),
.Y(n_424)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_320),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_383),
.Y(n_426)
);

OR2x6_ASAP7_75t_L g427 ( 
.A(n_376),
.B(n_189),
.Y(n_427)
);

INVx4_ASAP7_75t_L g428 ( 
.A(n_345),
.Y(n_428)
);

NOR2x1p5_ASAP7_75t_L g429 ( 
.A(n_336),
.B(n_275),
.Y(n_429)
);

BUFx2_ASAP7_75t_L g430 ( 
.A(n_360),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_326),
.B(n_219),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_398),
.B(n_399),
.Y(n_432)
);

INVx3_ASAP7_75t_L g433 ( 
.A(n_384),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_384),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_372),
.B(n_208),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_346),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_347),
.Y(n_437)
);

NAND2xp33_ASAP7_75t_L g438 ( 
.A(n_345),
.B(n_237),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_346),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_346),
.Y(n_440)
);

NAND2xp33_ASAP7_75t_SL g441 ( 
.A(n_324),
.B(n_232),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_315),
.Y(n_442)
);

INVx5_ASAP7_75t_L g443 ( 
.A(n_359),
.Y(n_443)
);

NAND3xp33_ASAP7_75t_L g444 ( 
.A(n_362),
.B(n_391),
.C(n_386),
.Y(n_444)
);

INVx6_ASAP7_75t_L g445 ( 
.A(n_391),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_351),
.B(n_221),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_347),
.Y(n_447)
);

BUFx10_ASAP7_75t_L g448 ( 
.A(n_362),
.Y(n_448)
);

INVx2_ASAP7_75t_SL g449 ( 
.A(n_363),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_316),
.B(n_225),
.Y(n_450)
);

INVx4_ASAP7_75t_L g451 ( 
.A(n_345),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_316),
.B(n_226),
.Y(n_452)
);

AOI22xp33_ASAP7_75t_L g453 ( 
.A1(n_391),
.A2(n_271),
.B1(n_313),
.B2(n_312),
.Y(n_453)
);

AND2x4_ASAP7_75t_L g454 ( 
.A(n_372),
.B(n_227),
.Y(n_454)
);

HB1xp67_ASAP7_75t_L g455 ( 
.A(n_365),
.Y(n_455)
);

BUFx6f_ASAP7_75t_SL g456 ( 
.A(n_373),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_339),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_354),
.Y(n_458)
);

AOI22xp33_ASAP7_75t_L g459 ( 
.A1(n_324),
.A2(n_231),
.B1(n_311),
.B2(n_310),
.Y(n_459)
);

BUFx3_ASAP7_75t_L g460 ( 
.A(n_356),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_318),
.B(n_229),
.Y(n_461)
);

INVx4_ASAP7_75t_SL g462 ( 
.A(n_345),
.Y(n_462)
);

INVx2_ASAP7_75t_SL g463 ( 
.A(n_323),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_405),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_380),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_380),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_SL g467 ( 
.A(n_373),
.B(n_232),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_318),
.B(n_233),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_361),
.B(n_239),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_361),
.B(n_240),
.Y(n_470)
);

OR2x2_ASAP7_75t_L g471 ( 
.A(n_370),
.B(n_220),
.Y(n_471)
);

OR2x2_ASAP7_75t_L g472 ( 
.A(n_349),
.B(n_223),
.Y(n_472)
);

INVx3_ASAP7_75t_L g473 ( 
.A(n_405),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_361),
.B(n_245),
.Y(n_474)
);

BUFx6f_ASAP7_75t_L g475 ( 
.A(n_333),
.Y(n_475)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_387),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_354),
.Y(n_477)
);

INVx3_ASAP7_75t_L g478 ( 
.A(n_387),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_319),
.B(n_327),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_319),
.B(n_250),
.Y(n_480)
);

INVx1_ASAP7_75t_SL g481 ( 
.A(n_329),
.Y(n_481)
);

INVx1_ASAP7_75t_SL g482 ( 
.A(n_394),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_L g483 ( 
.A1(n_367),
.A2(n_314),
.B1(n_236),
.B2(n_296),
.Y(n_483)
);

OR2x2_ASAP7_75t_L g484 ( 
.A(n_350),
.B(n_235),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_327),
.B(n_251),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_371),
.B(n_253),
.Y(n_486)
);

AND2x2_ASAP7_75t_SL g487 ( 
.A(n_394),
.B(n_254),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_358),
.A2(n_296),
.B1(n_241),
.B2(n_274),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_333),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_328),
.Y(n_490)
);

INVx4_ASAP7_75t_L g491 ( 
.A(n_345),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_355),
.Y(n_492)
);

INVx5_ASAP7_75t_L g493 ( 
.A(n_355),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_358),
.A2(n_241),
.B1(n_274),
.B2(n_281),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_393),
.Y(n_495)
);

INVx6_ASAP7_75t_L g496 ( 
.A(n_387),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_378),
.Y(n_497)
);

BUFx8_ASAP7_75t_SL g498 ( 
.A(n_348),
.Y(n_498)
);

OAI22xp33_ASAP7_75t_L g499 ( 
.A1(n_317),
.A2(n_278),
.B1(n_265),
.B2(n_266),
.Y(n_499)
);

BUFx6f_ASAP7_75t_L g500 ( 
.A(n_333),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_337),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_337),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_378),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_402),
.Y(n_504)
);

AND2x4_ASAP7_75t_L g505 ( 
.A(n_371),
.B(n_256),
.Y(n_505)
);

NAND2xp33_ASAP7_75t_SL g506 ( 
.A(n_395),
.B(n_266),
.Y(n_506)
);

BUFx2_ASAP7_75t_L g507 ( 
.A(n_323),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_355),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_382),
.Y(n_509)
);

BUFx4f_ASAP7_75t_L g510 ( 
.A(n_402),
.Y(n_510)
);

INVx2_ASAP7_75t_SL g511 ( 
.A(n_395),
.Y(n_511)
);

BUFx3_ASAP7_75t_L g512 ( 
.A(n_355),
.Y(n_512)
);

INVx1_ASAP7_75t_SL g513 ( 
.A(n_348),
.Y(n_513)
);

CKINVDCx16_ASAP7_75t_R g514 ( 
.A(n_322),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_352),
.B(n_353),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_375),
.Y(n_516)
);

AND2x4_ASAP7_75t_L g517 ( 
.A(n_375),
.B(n_258),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_419),
.B(n_279),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_L g519 ( 
.A1(n_482),
.A2(n_381),
.B1(n_389),
.B2(n_369),
.Y(n_519)
);

AOI22xp33_ASAP7_75t_L g520 ( 
.A1(n_436),
.A2(n_408),
.B1(n_392),
.B2(n_406),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_457),
.B(n_375),
.Y(n_521)
);

OR2x6_ASAP7_75t_L g522 ( 
.A(n_413),
.B(n_390),
.Y(n_522)
);

INVx1_ASAP7_75t_SL g523 ( 
.A(n_430),
.Y(n_523)
);

INVx2_ASAP7_75t_SL g524 ( 
.A(n_471),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_498),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_412),
.B(n_374),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_414),
.B(n_377),
.Y(n_527)
);

NAND2x1p5_ASAP7_75t_L g528 ( 
.A(n_482),
.B(n_403),
.Y(n_528)
);

INVx3_ASAP7_75t_L g529 ( 
.A(n_425),
.Y(n_529)
);

INVx2_ASAP7_75t_SL g530 ( 
.A(n_472),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_505),
.B(n_388),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_517),
.B(n_388),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_496),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_496),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_512),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_445),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_516),
.Y(n_537)
);

NOR2xp67_ASAP7_75t_L g538 ( 
.A(n_463),
.B(n_392),
.Y(n_538)
);

INVx3_ASAP7_75t_L g539 ( 
.A(n_445),
.Y(n_539)
);

OR2x2_ASAP7_75t_L g540 ( 
.A(n_416),
.B(n_343),
.Y(n_540)
);

AO22x1_ASAP7_75t_L g541 ( 
.A1(n_507),
.A2(n_291),
.B1(n_299),
.B2(n_283),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_479),
.Y(n_542)
);

OR2x6_ASAP7_75t_L g543 ( 
.A(n_413),
.B(n_368),
.Y(n_543)
);

AOI22xp33_ASAP7_75t_L g544 ( 
.A1(n_439),
.A2(n_396),
.B1(n_404),
.B2(n_397),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_484),
.B(n_397),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_435),
.B(n_415),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_432),
.B(n_400),
.Y(n_547)
);

AOI22xp33_ASAP7_75t_L g548 ( 
.A1(n_440),
.A2(n_433),
.B1(n_422),
.B2(n_426),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_454),
.B(n_401),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_479),
.Y(n_550)
);

AOI22xp5_ASAP7_75t_L g551 ( 
.A1(n_487),
.A2(n_283),
.B1(n_291),
.B2(n_293),
.Y(n_551)
);

AOI21xp5_ASAP7_75t_L g552 ( 
.A1(n_438),
.A2(n_364),
.B(n_332),
.Y(n_552)
);

NOR2x1p5_ASAP7_75t_L g553 ( 
.A(n_423),
.B(n_342),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_455),
.B(n_344),
.Y(n_554)
);

NAND2x1p5_ASAP7_75t_L g555 ( 
.A(n_411),
.B(n_330),
.Y(n_555)
);

OR2x6_ASAP7_75t_L g556 ( 
.A(n_413),
.B(n_331),
.Y(n_556)
);

AND2x6_ASAP7_75t_SL g557 ( 
.A(n_427),
.B(n_260),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_497),
.B(n_307),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_503),
.B(n_308),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_509),
.B(n_332),
.Y(n_560)
);

NAND2x1_ASAP7_75t_L g561 ( 
.A(n_418),
.B(n_338),
.Y(n_561)
);

OAI21xp5_ASAP7_75t_L g562 ( 
.A1(n_444),
.A2(n_292),
.B(n_287),
.Y(n_562)
);

A2O1A1Ixp33_ASAP7_75t_L g563 ( 
.A1(n_464),
.A2(n_294),
.B(n_273),
.C(n_295),
.Y(n_563)
);

BUFx8_ASAP7_75t_SL g564 ( 
.A(n_465),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_490),
.Y(n_565)
);

INVx2_ASAP7_75t_SL g566 ( 
.A(n_448),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_424),
.B(n_407),
.Y(n_567)
);

AO22x1_ASAP7_75t_L g568 ( 
.A1(n_458),
.A2(n_207),
.B1(n_217),
.B2(n_276),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_460),
.Y(n_569)
);

HB1xp67_ASAP7_75t_L g570 ( 
.A(n_481),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_420),
.B(n_282),
.Y(n_571)
);

OR2x2_ASAP7_75t_L g572 ( 
.A(n_481),
.B(n_407),
.Y(n_572)
);

AOI22xp33_ASAP7_75t_L g573 ( 
.A1(n_417),
.A2(n_407),
.B1(n_402),
.B2(n_385),
.Y(n_573)
);

AND2x6_ASAP7_75t_SL g574 ( 
.A(n_427),
.B(n_264),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_453),
.B(n_306),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_511),
.B(n_262),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_476),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_428),
.B(n_379),
.Y(n_578)
);

AOI22xp33_ASAP7_75t_SL g579 ( 
.A1(n_456),
.A2(n_385),
.B1(n_341),
.B2(n_337),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_449),
.B(n_36),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_473),
.Y(n_581)
);

A2O1A1Ixp33_ASAP7_75t_L g582 ( 
.A1(n_434),
.A2(n_242),
.B(n_238),
.C(n_228),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_446),
.B(n_341),
.Y(n_583)
);

INVx4_ASAP7_75t_L g584 ( 
.A(n_443),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_476),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_410),
.Y(n_586)
);

INVx4_ASAP7_75t_L g587 ( 
.A(n_443),
.Y(n_587)
);

AOI22xp5_ASAP7_75t_L g588 ( 
.A1(n_506),
.A2(n_341),
.B1(n_337),
.B2(n_37),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_478),
.Y(n_589)
);

AOI22xp33_ASAP7_75t_L g590 ( 
.A1(n_418),
.A2(n_37),
.B1(n_38),
.B2(n_42),
.Y(n_590)
);

AOI21xp5_ASAP7_75t_L g591 ( 
.A1(n_428),
.A2(n_101),
.B(n_43),
.Y(n_591)
);

AOI22xp33_ASAP7_75t_SL g592 ( 
.A1(n_409),
.A2(n_38),
.B1(n_44),
.B2(n_46),
.Y(n_592)
);

AOI21xp5_ASAP7_75t_L g593 ( 
.A1(n_451),
.A2(n_50),
.B(n_51),
.Y(n_593)
);

NAND2x1p5_ASAP7_75t_L g594 ( 
.A(n_429),
.B(n_58),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_478),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_515),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_504),
.Y(n_597)
);

HB1xp67_ASAP7_75t_L g598 ( 
.A(n_462),
.Y(n_598)
);

AOI22xp33_ASAP7_75t_L g599 ( 
.A1(n_418),
.A2(n_491),
.B1(n_451),
.B2(n_470),
.Y(n_599)
);

AOI22xp33_ASAP7_75t_L g600 ( 
.A1(n_491),
.A2(n_64),
.B1(n_66),
.B2(n_70),
.Y(n_600)
);

NOR2x1p5_ASAP7_75t_L g601 ( 
.A(n_477),
.B(n_71),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_542),
.B(n_459),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_550),
.Y(n_603)
);

OAI22xp5_ASAP7_75t_L g604 ( 
.A1(n_548),
.A2(n_494),
.B1(n_488),
.B2(n_514),
.Y(n_604)
);

A2O1A1Ixp33_ASAP7_75t_L g605 ( 
.A1(n_562),
.A2(n_469),
.B(n_474),
.C(n_486),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_524),
.B(n_499),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_561),
.Y(n_607)
);

AND2x4_ASAP7_75t_L g608 ( 
.A(n_556),
.B(n_462),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_581),
.Y(n_609)
);

INVx8_ASAP7_75t_L g610 ( 
.A(n_556),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_566),
.B(n_523),
.Y(n_611)
);

AND2x4_ASAP7_75t_L g612 ( 
.A(n_556),
.B(n_538),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_530),
.B(n_441),
.Y(n_613)
);

AOI21xp5_ASAP7_75t_L g614 ( 
.A1(n_552),
.A2(n_521),
.B(n_546),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_529),
.Y(n_615)
);

HB1xp67_ASAP7_75t_L g616 ( 
.A(n_570),
.Y(n_616)
);

NOR3xp33_ASAP7_75t_SL g617 ( 
.A(n_525),
.B(n_483),
.C(n_409),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_526),
.B(n_494),
.Y(n_618)
);

O2A1O1Ixp33_ASAP7_75t_L g619 ( 
.A1(n_519),
.A2(n_483),
.B(n_431),
.C(n_452),
.Y(n_619)
);

AOI21xp5_ASAP7_75t_L g620 ( 
.A1(n_578),
.A2(n_485),
.B(n_480),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_527),
.B(n_431),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_551),
.B(n_495),
.Y(n_622)
);

HB1xp67_ASAP7_75t_L g623 ( 
.A(n_540),
.Y(n_623)
);

OAI21xp33_ASAP7_75t_L g624 ( 
.A1(n_571),
.A2(n_488),
.B(n_450),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_529),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_547),
.B(n_468),
.Y(n_626)
);

OAI21xp5_ASAP7_75t_L g627 ( 
.A1(n_591),
.A2(n_468),
.B(n_461),
.Y(n_627)
);

AOI21xp5_ASAP7_75t_L g628 ( 
.A1(n_518),
.A2(n_461),
.B(n_510),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_572),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_545),
.B(n_427),
.Y(n_630)
);

BUFx2_ASAP7_75t_L g631 ( 
.A(n_564),
.Y(n_631)
);

OAI22xp5_ASAP7_75t_L g632 ( 
.A1(n_548),
.A2(n_513),
.B1(n_466),
.B2(n_504),
.Y(n_632)
);

OR2x2_ASAP7_75t_L g633 ( 
.A(n_554),
.B(n_508),
.Y(n_633)
);

AOI22xp5_ASAP7_75t_L g634 ( 
.A1(n_522),
.A2(n_421),
.B1(n_437),
.B2(n_447),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_560),
.Y(n_635)
);

INVx1_ASAP7_75t_SL g636 ( 
.A(n_580),
.Y(n_636)
);

AOI21xp5_ASAP7_75t_L g637 ( 
.A1(n_586),
.A2(n_492),
.B(n_493),
.Y(n_637)
);

AND2x4_ASAP7_75t_L g638 ( 
.A(n_553),
.B(n_73),
.Y(n_638)
);

AND2x4_ASAP7_75t_L g639 ( 
.A(n_543),
.B(n_78),
.Y(n_639)
);

NAND2xp33_ASAP7_75t_SL g640 ( 
.A(n_601),
.B(n_502),
.Y(n_640)
);

OAI21xp5_ASAP7_75t_L g641 ( 
.A1(n_591),
.A2(n_502),
.B(n_501),
.Y(n_641)
);

OAI22xp5_ASAP7_75t_L g642 ( 
.A1(n_599),
.A2(n_501),
.B1(n_500),
.B2(n_489),
.Y(n_642)
);

OAI22xp5_ASAP7_75t_L g643 ( 
.A1(n_599),
.A2(n_549),
.B1(n_544),
.B2(n_520),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_537),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_565),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_SL g646 ( 
.A(n_598),
.B(n_475),
.Y(n_646)
);

O2A1O1Ixp33_ASAP7_75t_L g647 ( 
.A1(n_563),
.A2(n_83),
.B(n_86),
.C(n_97),
.Y(n_647)
);

BUFx6f_ASAP7_75t_SL g648 ( 
.A(n_522),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_SL g649 ( 
.A(n_594),
.B(n_593),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_543),
.B(n_120),
.Y(n_650)
);

NOR3xp33_ASAP7_75t_SL g651 ( 
.A(n_575),
.B(n_582),
.C(n_576),
.Y(n_651)
);

INVxp67_ASAP7_75t_L g652 ( 
.A(n_541),
.Y(n_652)
);

INVx3_ASAP7_75t_L g653 ( 
.A(n_584),
.Y(n_653)
);

BUFx12f_ASAP7_75t_L g654 ( 
.A(n_557),
.Y(n_654)
);

INVx2_ASAP7_75t_SL g655 ( 
.A(n_543),
.Y(n_655)
);

O2A1O1Ixp33_ASAP7_75t_L g656 ( 
.A1(n_531),
.A2(n_141),
.B(n_144),
.C(n_146),
.Y(n_656)
);

BUFx2_ASAP7_75t_L g657 ( 
.A(n_555),
.Y(n_657)
);

OAI22xp5_ASAP7_75t_L g658 ( 
.A1(n_520),
.A2(n_442),
.B1(n_151),
.B2(n_154),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_532),
.B(n_147),
.Y(n_659)
);

HB1xp67_ASAP7_75t_L g660 ( 
.A(n_555),
.Y(n_660)
);

AOI21xp5_ASAP7_75t_L g661 ( 
.A1(n_558),
.A2(n_559),
.B(n_567),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_583),
.Y(n_662)
);

INVxp67_ASAP7_75t_L g663 ( 
.A(n_528),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_544),
.B(n_164),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_536),
.B(n_539),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_596),
.B(n_568),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_SL g667 ( 
.A(n_584),
.B(n_587),
.Y(n_667)
);

AOI21xp5_ASAP7_75t_L g668 ( 
.A1(n_577),
.A2(n_589),
.B(n_585),
.Y(n_668)
);

AOI21xp5_ASAP7_75t_L g669 ( 
.A1(n_595),
.A2(n_597),
.B(n_535),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_587),
.Y(n_670)
);

NAND2x1p5_ASAP7_75t_L g671 ( 
.A(n_569),
.B(n_588),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_579),
.B(n_592),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_579),
.B(n_590),
.Y(n_673)
);

INVxp67_ASAP7_75t_L g674 ( 
.A(n_592),
.Y(n_674)
);

BUFx2_ASAP7_75t_L g675 ( 
.A(n_574),
.Y(n_675)
);

OR2x6_ASAP7_75t_SL g676 ( 
.A(n_590),
.B(n_533),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_534),
.Y(n_677)
);

AOI22xp33_ASAP7_75t_L g678 ( 
.A1(n_604),
.A2(n_573),
.B1(n_600),
.B2(n_674),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_618),
.B(n_600),
.Y(n_679)
);

OAI22xp5_ASAP7_75t_L g680 ( 
.A1(n_635),
.A2(n_573),
.B1(n_603),
.B2(n_626),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_623),
.B(n_616),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_611),
.B(n_652),
.Y(n_682)
);

O2A1O1Ixp33_ASAP7_75t_L g683 ( 
.A1(n_619),
.A2(n_606),
.B(n_624),
.C(n_672),
.Y(n_683)
);

INVx1_ASAP7_75t_SL g684 ( 
.A(n_610),
.Y(n_684)
);

OAI21xp5_ASAP7_75t_L g685 ( 
.A1(n_614),
.A2(n_661),
.B(n_627),
.Y(n_685)
);

AO32x2_ASAP7_75t_L g686 ( 
.A1(n_643),
.A2(n_642),
.A3(n_655),
.B1(n_676),
.B2(n_658),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_617),
.B(n_613),
.Y(n_687)
);

OAI22xp5_ASAP7_75t_L g688 ( 
.A1(n_602),
.A2(n_636),
.B1(n_629),
.B2(n_645),
.Y(n_688)
);

O2A1O1Ixp33_ASAP7_75t_L g689 ( 
.A1(n_630),
.A2(n_632),
.B(n_673),
.C(n_651),
.Y(n_689)
);

NAND3xp33_ASAP7_75t_L g690 ( 
.A(n_649),
.B(n_641),
.C(n_647),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_644),
.Y(n_691)
);

AOI22xp5_ASAP7_75t_L g692 ( 
.A1(n_648),
.A2(n_639),
.B1(n_622),
.B2(n_636),
.Y(n_692)
);

CKINVDCx12_ASAP7_75t_R g693 ( 
.A(n_631),
.Y(n_693)
);

OR2x2_ASAP7_75t_L g694 ( 
.A(n_610),
.B(n_666),
.Y(n_694)
);

OAI22xp5_ASAP7_75t_L g695 ( 
.A1(n_639),
.A2(n_633),
.B1(n_663),
.B2(n_608),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_648),
.B(n_612),
.Y(n_696)
);

NOR2xp67_ASAP7_75t_L g697 ( 
.A(n_608),
.B(n_650),
.Y(n_697)
);

OAI21xp5_ASAP7_75t_L g698 ( 
.A1(n_620),
.A2(n_662),
.B(n_664),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_609),
.Y(n_699)
);

AOI21xp5_ASAP7_75t_L g700 ( 
.A1(n_668),
.A2(n_669),
.B(n_659),
.Y(n_700)
);

BUFx8_ASAP7_75t_L g701 ( 
.A(n_654),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_660),
.B(n_657),
.Y(n_702)
);

A2O1A1Ixp33_ASAP7_75t_L g703 ( 
.A1(n_640),
.A2(n_628),
.B(n_634),
.C(n_656),
.Y(n_703)
);

INVx1_ASAP7_75t_SL g704 ( 
.A(n_638),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_670),
.Y(n_705)
);

INVx1_ASAP7_75t_SL g706 ( 
.A(n_638),
.Y(n_706)
);

BUFx8_ASAP7_75t_L g707 ( 
.A(n_675),
.Y(n_707)
);

BUFx6f_ASAP7_75t_L g708 ( 
.A(n_607),
.Y(n_708)
);

A2O1A1Ixp33_ASAP7_75t_L g709 ( 
.A1(n_637),
.A2(n_615),
.B(n_625),
.C(n_677),
.Y(n_709)
);

BUFx10_ASAP7_75t_L g710 ( 
.A(n_665),
.Y(n_710)
);

AOI21xp5_ASAP7_75t_L g711 ( 
.A1(n_646),
.A2(n_667),
.B(n_671),
.Y(n_711)
);

BUFx2_ASAP7_75t_L g712 ( 
.A(n_653),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_604),
.B(n_523),
.Y(n_713)
);

A2O1A1Ixp33_ASAP7_75t_L g714 ( 
.A1(n_661),
.A2(n_614),
.B(n_674),
.C(n_605),
.Y(n_714)
);

OAI21xp5_ASAP7_75t_L g715 ( 
.A1(n_614),
.A2(n_661),
.B(n_627),
.Y(n_715)
);

BUFx3_ASAP7_75t_L g716 ( 
.A(n_631),
.Y(n_716)
);

HB1xp67_ASAP7_75t_L g717 ( 
.A(n_616),
.Y(n_717)
);

NOR2xp67_ASAP7_75t_SL g718 ( 
.A(n_623),
.B(n_566),
.Y(n_718)
);

INVx2_ASAP7_75t_SL g719 ( 
.A(n_610),
.Y(n_719)
);

BUFx12f_ASAP7_75t_L g720 ( 
.A(n_631),
.Y(n_720)
);

NOR2x1_ASAP7_75t_R g721 ( 
.A(n_631),
.B(n_348),
.Y(n_721)
);

NAND3xp33_ASAP7_75t_L g722 ( 
.A(n_651),
.B(n_674),
.C(n_582),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_616),
.Y(n_723)
);

CKINVDCx6p67_ASAP7_75t_R g724 ( 
.A(n_631),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_603),
.Y(n_725)
);

NAND4xp25_ASAP7_75t_L g726 ( 
.A(n_604),
.B(n_618),
.C(n_619),
.D(n_467),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_603),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_604),
.B(n_523),
.Y(n_728)
);

INVx3_ASAP7_75t_L g729 ( 
.A(n_608),
.Y(n_729)
);

OAI21xp5_ASAP7_75t_L g730 ( 
.A1(n_614),
.A2(n_661),
.B(n_627),
.Y(n_730)
);

NAND2x1p5_ASAP7_75t_L g731 ( 
.A(n_608),
.B(n_523),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_616),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_616),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_604),
.B(n_523),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_616),
.Y(n_735)
);

BUFx6f_ASAP7_75t_L g736 ( 
.A(n_608),
.Y(n_736)
);

A2O1A1Ixp33_ASAP7_75t_L g737 ( 
.A1(n_661),
.A2(n_614),
.B(n_674),
.C(n_605),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_621),
.B(n_603),
.Y(n_738)
);

AOI22xp33_ASAP7_75t_L g739 ( 
.A1(n_604),
.A2(n_456),
.B1(n_467),
.B2(n_674),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_616),
.Y(n_740)
);

O2A1O1Ixp33_ASAP7_75t_L g741 ( 
.A1(n_674),
.A2(n_519),
.B(n_619),
.C(n_604),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_604),
.B(n_523),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_621),
.B(n_603),
.Y(n_743)
);

BUFx12f_ASAP7_75t_L g744 ( 
.A(n_631),
.Y(n_744)
);

BUFx6f_ASAP7_75t_L g745 ( 
.A(n_608),
.Y(n_745)
);

HB1xp67_ASAP7_75t_L g746 ( 
.A(n_616),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_603),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_621),
.B(n_603),
.Y(n_748)
);

BUFx6f_ASAP7_75t_L g749 ( 
.A(n_608),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_621),
.B(n_603),
.Y(n_750)
);

AOI22xp33_ASAP7_75t_L g751 ( 
.A1(n_604),
.A2(n_456),
.B1(n_467),
.B2(n_674),
.Y(n_751)
);

BUFx3_ASAP7_75t_L g752 ( 
.A(n_631),
.Y(n_752)
);

A2O1A1Ixp33_ASAP7_75t_L g753 ( 
.A1(n_661),
.A2(n_614),
.B(n_674),
.C(n_605),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_611),
.B(n_566),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_603),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_623),
.B(n_570),
.Y(n_756)
);

BUFx2_ASAP7_75t_SL g757 ( 
.A(n_631),
.Y(n_757)
);

AOI22xp33_ASAP7_75t_L g758 ( 
.A1(n_604),
.A2(n_456),
.B1(n_467),
.B2(n_674),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_604),
.B(n_523),
.Y(n_759)
);

NOR2xp67_ASAP7_75t_SL g760 ( 
.A(n_623),
.B(n_566),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_621),
.B(n_603),
.Y(n_761)
);

OAI21xp5_ASAP7_75t_L g762 ( 
.A1(n_614),
.A2(n_661),
.B(n_627),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_604),
.B(n_523),
.Y(n_763)
);

BUFx2_ASAP7_75t_L g764 ( 
.A(n_616),
.Y(n_764)
);

NOR2xp67_ASAP7_75t_L g765 ( 
.A(n_603),
.B(n_635),
.Y(n_765)
);

CKINVDCx20_ASAP7_75t_R g766 ( 
.A(n_631),
.Y(n_766)
);

AOI221xp5_ASAP7_75t_SL g767 ( 
.A1(n_674),
.A2(n_619),
.B1(n_614),
.B2(n_624),
.C(n_605),
.Y(n_767)
);

OAI21xp5_ASAP7_75t_L g768 ( 
.A1(n_614),
.A2(n_661),
.B(n_627),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_725),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_738),
.B(n_743),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_727),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_691),
.Y(n_772)
);

BUFx4f_ASAP7_75t_SL g773 ( 
.A(n_701),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_747),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_755),
.Y(n_775)
);

AO21x2_ASAP7_75t_L g776 ( 
.A1(n_685),
.A2(n_768),
.B(n_715),
.Y(n_776)
);

OAI21x1_ASAP7_75t_SL g777 ( 
.A1(n_711),
.A2(n_695),
.B(n_692),
.Y(n_777)
);

AOI21xp5_ASAP7_75t_L g778 ( 
.A1(n_714),
.A2(n_737),
.B(n_753),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_748),
.B(n_750),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_723),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_732),
.Y(n_781)
);

AOI21xp5_ASAP7_75t_L g782 ( 
.A1(n_730),
.A2(n_762),
.B(n_690),
.Y(n_782)
);

OAI21xp5_ASAP7_75t_L g783 ( 
.A1(n_679),
.A2(n_683),
.B(n_767),
.Y(n_783)
);

AOI22xp5_ASAP7_75t_L g784 ( 
.A1(n_713),
.A2(n_759),
.B1(n_734),
.B2(n_742),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_699),
.Y(n_785)
);

AOI21xp5_ASAP7_75t_L g786 ( 
.A1(n_700),
.A2(n_698),
.B(n_703),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_701),
.Y(n_787)
);

A2O1A1Ixp33_ASAP7_75t_L g788 ( 
.A1(n_741),
.A2(n_689),
.B(n_765),
.C(n_726),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_720),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_SL g790 ( 
.A(n_704),
.B(n_706),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_733),
.Y(n_791)
);

AO31x2_ASAP7_75t_L g792 ( 
.A1(n_688),
.A2(n_709),
.A3(n_680),
.B(n_728),
.Y(n_792)
);

INVx3_ASAP7_75t_L g793 ( 
.A(n_736),
.Y(n_793)
);

AOI22xp5_ASAP7_75t_L g794 ( 
.A1(n_763),
.A2(n_739),
.B1(n_751),
.B2(n_758),
.Y(n_794)
);

A2O1A1Ixp33_ASAP7_75t_L g795 ( 
.A1(n_722),
.A2(n_761),
.B(n_687),
.C(n_678),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_735),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_740),
.Y(n_797)
);

AOI22xp33_ASAP7_75t_L g798 ( 
.A1(n_722),
.A2(n_692),
.B1(n_764),
.B2(n_756),
.Y(n_798)
);

AND3x2_ASAP7_75t_L g799 ( 
.A(n_721),
.B(n_696),
.C(n_746),
.Y(n_799)
);

AO21x1_ASAP7_75t_L g800 ( 
.A1(n_682),
.A2(n_694),
.B(n_686),
.Y(n_800)
);

AOI21xp5_ASAP7_75t_L g801 ( 
.A1(n_705),
.A2(n_697),
.B(n_681),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_717),
.B(n_702),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_731),
.B(n_684),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_708),
.Y(n_804)
);

AOI21xp5_ASAP7_75t_L g805 ( 
.A1(n_697),
.A2(n_754),
.B(n_708),
.Y(n_805)
);

AOI22xp5_ASAP7_75t_L g806 ( 
.A1(n_718),
.A2(n_760),
.B1(n_766),
.B2(n_757),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_710),
.B(n_708),
.Y(n_807)
);

CKINVDCx6p67_ASAP7_75t_R g808 ( 
.A(n_693),
.Y(n_808)
);

OAI22xp33_ASAP7_75t_L g809 ( 
.A1(n_724),
.A2(n_752),
.B1(n_716),
.B2(n_719),
.Y(n_809)
);

AOI22xp33_ASAP7_75t_L g810 ( 
.A1(n_710),
.A2(n_712),
.B1(n_729),
.B2(n_745),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_744),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_749),
.B(n_721),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_707),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_707),
.Y(n_814)
);

AOI21xp33_ASAP7_75t_L g815 ( 
.A1(n_683),
.A2(n_741),
.B(n_689),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_701),
.Y(n_816)
);

AOI221xp5_ASAP7_75t_L g817 ( 
.A1(n_741),
.A2(n_604),
.B1(n_713),
.B2(n_734),
.C(n_728),
.Y(n_817)
);

AOI21xp5_ASAP7_75t_SL g818 ( 
.A1(n_695),
.A2(n_639),
.B(n_711),
.Y(n_818)
);

OAI21xp5_ASAP7_75t_L g819 ( 
.A1(n_679),
.A2(n_737),
.B(n_714),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_692),
.B(n_695),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_738),
.B(n_743),
.Y(n_821)
);

OA21x2_ASAP7_75t_L g822 ( 
.A1(n_685),
.A2(n_730),
.B(n_715),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_691),
.Y(n_823)
);

OR2x2_ASAP7_75t_L g824 ( 
.A(n_681),
.B(n_523),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_738),
.B(n_743),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_692),
.B(n_695),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_738),
.B(n_743),
.Y(n_827)
);

HB1xp67_ASAP7_75t_L g828 ( 
.A(n_764),
.Y(n_828)
);

AOI22xp5_ASAP7_75t_L g829 ( 
.A1(n_713),
.A2(n_467),
.B1(n_380),
.B2(n_393),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_738),
.B(n_743),
.Y(n_830)
);

AOI22xp33_ASAP7_75t_L g831 ( 
.A1(n_713),
.A2(n_728),
.B1(n_742),
.B2(n_734),
.Y(n_831)
);

HB1xp67_ASAP7_75t_L g832 ( 
.A(n_776),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_822),
.Y(n_833)
);

OA21x2_ASAP7_75t_L g834 ( 
.A1(n_786),
.A2(n_778),
.B(n_782),
.Y(n_834)
);

HB1xp67_ASAP7_75t_L g835 ( 
.A(n_776),
.Y(n_835)
);

INVxp67_ASAP7_75t_L g836 ( 
.A(n_770),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_819),
.B(n_783),
.Y(n_837)
);

OAI31xp33_ASAP7_75t_SL g838 ( 
.A1(n_820),
.A2(n_826),
.A3(n_817),
.B(n_809),
.Y(n_838)
);

OAI22xp33_ASAP7_75t_L g839 ( 
.A1(n_794),
.A2(n_784),
.B1(n_770),
.B2(n_830),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_819),
.B(n_783),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_779),
.B(n_821),
.Y(n_841)
);

INVxp67_ASAP7_75t_SL g842 ( 
.A(n_779),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_772),
.Y(n_843)
);

AND2x6_ASAP7_75t_L g844 ( 
.A(n_818),
.B(n_804),
.Y(n_844)
);

OR2x6_ASAP7_75t_L g845 ( 
.A(n_777),
.B(n_801),
.Y(n_845)
);

OAI21xp5_ASAP7_75t_L g846 ( 
.A1(n_795),
.A2(n_788),
.B(n_815),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_823),
.Y(n_847)
);

INVxp67_ASAP7_75t_L g848 ( 
.A(n_821),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_SL g849 ( 
.A1(n_825),
.A2(n_830),
.B(n_827),
.Y(n_849)
);

BUFx2_ASAP7_75t_L g850 ( 
.A(n_792),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_817),
.B(n_831),
.Y(n_851)
);

OAI21xp5_ASAP7_75t_L g852 ( 
.A1(n_825),
.A2(n_827),
.B(n_805),
.Y(n_852)
);

AND2x4_ASAP7_75t_SL g853 ( 
.A(n_769),
.B(n_771),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_833),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_837),
.B(n_792),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_837),
.B(n_800),
.Y(n_856)
);

INVxp67_ASAP7_75t_SL g857 ( 
.A(n_842),
.Y(n_857)
);

AND2x2_ASAP7_75t_L g858 ( 
.A(n_837),
.B(n_798),
.Y(n_858)
);

INVx4_ASAP7_75t_L g859 ( 
.A(n_853),
.Y(n_859)
);

NOR2x1_ASAP7_75t_L g860 ( 
.A(n_849),
.B(n_807),
.Y(n_860)
);

AND2x4_ASAP7_75t_L g861 ( 
.A(n_840),
.B(n_805),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_840),
.B(n_850),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_834),
.B(n_785),
.Y(n_863)
);

INVx5_ASAP7_75t_L g864 ( 
.A(n_844),
.Y(n_864)
);

INVxp67_ASAP7_75t_L g865 ( 
.A(n_841),
.Y(n_865)
);

OR2x2_ASAP7_75t_L g866 ( 
.A(n_836),
.B(n_824),
.Y(n_866)
);

OR2x2_ASAP7_75t_L g867 ( 
.A(n_836),
.B(n_828),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_851),
.B(n_774),
.Y(n_868)
);

AND2x4_ASAP7_75t_L g869 ( 
.A(n_845),
.B(n_793),
.Y(n_869)
);

OR2x2_ASAP7_75t_L g870 ( 
.A(n_848),
.B(n_775),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_858),
.B(n_851),
.Y(n_871)
);

AND2x2_ASAP7_75t_L g872 ( 
.A(n_862),
.B(n_832),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_858),
.B(n_839),
.Y(n_873)
);

AND2x4_ASAP7_75t_L g874 ( 
.A(n_864),
.B(n_861),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_858),
.B(n_839),
.Y(n_875)
);

OR2x2_ASAP7_75t_L g876 ( 
.A(n_862),
.B(n_857),
.Y(n_876)
);

INVxp67_ASAP7_75t_SL g877 ( 
.A(n_857),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_854),
.Y(n_878)
);

AND2x4_ASAP7_75t_L g879 ( 
.A(n_864),
.B(n_845),
.Y(n_879)
);

INVx1_ASAP7_75t_SL g880 ( 
.A(n_870),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_862),
.B(n_832),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_855),
.B(n_835),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_882),
.B(n_863),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_878),
.Y(n_884)
);

AND2x4_ASAP7_75t_L g885 ( 
.A(n_874),
.B(n_864),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_878),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_882),
.B(n_863),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_880),
.B(n_865),
.Y(n_888)
);

AND2x4_ASAP7_75t_L g889 ( 
.A(n_879),
.B(n_864),
.Y(n_889)
);

AND2x4_ASAP7_75t_L g890 ( 
.A(n_879),
.B(n_864),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_872),
.B(n_863),
.Y(n_891)
);

NOR2xp33_ASAP7_75t_SL g892 ( 
.A(n_885),
.B(n_773),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_884),
.Y(n_893)
);

AOI22xp5_ASAP7_75t_L g894 ( 
.A1(n_888),
.A2(n_875),
.B1(n_873),
.B2(n_871),
.Y(n_894)
);

INVx1_ASAP7_75t_SL g895 ( 
.A(n_891),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_L g896 ( 
.A(n_891),
.B(n_873),
.Y(n_896)
);

OR2x2_ASAP7_75t_L g897 ( 
.A(n_883),
.B(n_876),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_883),
.B(n_880),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_884),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_886),
.Y(n_900)
);

INVx1_ASAP7_75t_SL g901 ( 
.A(n_887),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_887),
.B(n_875),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_885),
.B(n_872),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_886),
.B(n_871),
.Y(n_904)
);

NOR2xp33_ASAP7_75t_L g905 ( 
.A(n_896),
.B(n_813),
.Y(n_905)
);

AND2x2_ASAP7_75t_L g906 ( 
.A(n_903),
.B(n_874),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_893),
.Y(n_907)
);

NOR3xp33_ASAP7_75t_L g908 ( 
.A(n_904),
.B(n_860),
.C(n_814),
.Y(n_908)
);

AOI22xp5_ASAP7_75t_L g909 ( 
.A1(n_892),
.A2(n_860),
.B1(n_881),
.B2(n_856),
.Y(n_909)
);

AOI21xp33_ASAP7_75t_L g910 ( 
.A1(n_894),
.A2(n_838),
.B(n_867),
.Y(n_910)
);

OAI22xp33_ASAP7_75t_SL g911 ( 
.A1(n_897),
.A2(n_876),
.B1(n_877),
.B2(n_885),
.Y(n_911)
);

NAND3xp33_ASAP7_75t_SL g912 ( 
.A(n_895),
.B(n_816),
.C(n_787),
.Y(n_912)
);

OAI22xp5_ASAP7_75t_L g913 ( 
.A1(n_901),
.A2(n_890),
.B1(n_889),
.B2(n_885),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_899),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_896),
.B(n_902),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_907),
.Y(n_916)
);

OAI22xp33_ASAP7_75t_L g917 ( 
.A1(n_909),
.A2(n_897),
.B1(n_859),
.B2(n_864),
.Y(n_917)
);

AOI21xp33_ASAP7_75t_L g918 ( 
.A1(n_905),
.A2(n_838),
.B(n_867),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_914),
.Y(n_919)
);

AOI222xp33_ASAP7_75t_L g920 ( 
.A1(n_912),
.A2(n_848),
.B1(n_865),
.B2(n_898),
.C1(n_856),
.C2(n_900),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_911),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_915),
.B(n_908),
.Y(n_922)
);

OAI22xp5_ASAP7_75t_SL g923 ( 
.A1(n_921),
.A2(n_912),
.B1(n_811),
.B2(n_789),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_916),
.Y(n_924)
);

OAI31xp33_ASAP7_75t_L g925 ( 
.A1(n_917),
.A2(n_913),
.A3(n_910),
.B(n_906),
.Y(n_925)
);

AOI22xp5_ASAP7_75t_L g926 ( 
.A1(n_920),
.A2(n_903),
.B1(n_856),
.B2(n_889),
.Y(n_926)
);

OAI22xp5_ASAP7_75t_L g927 ( 
.A1(n_922),
.A2(n_890),
.B1(n_889),
.B2(n_859),
.Y(n_927)
);

AOI31xp33_ASAP7_75t_L g928 ( 
.A1(n_918),
.A2(n_806),
.A3(n_808),
.B(n_812),
.Y(n_928)
);

NOR3xp33_ASAP7_75t_SL g929 ( 
.A(n_923),
.B(n_925),
.C(n_927),
.Y(n_929)
);

NAND3xp33_ASAP7_75t_SL g930 ( 
.A(n_926),
.B(n_829),
.C(n_846),
.Y(n_930)
);

OAI311xp33_ASAP7_75t_L g931 ( 
.A1(n_928),
.A2(n_919),
.A3(n_866),
.B1(n_852),
.C1(n_868),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_924),
.B(n_890),
.Y(n_932)
);

OR5x1_ASAP7_75t_L g933 ( 
.A(n_929),
.B(n_799),
.C(n_917),
.D(n_866),
.E(n_864),
.Y(n_933)
);

HB1xp67_ASAP7_75t_L g934 ( 
.A(n_932),
.Y(n_934)
);

AOI211xp5_ASAP7_75t_L g935 ( 
.A1(n_931),
.A2(n_852),
.B(n_868),
.C(n_802),
.Y(n_935)
);

XNOR2x1_ASAP7_75t_L g936 ( 
.A(n_933),
.B(n_930),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_934),
.Y(n_937)
);

XOR2xp5_ASAP7_75t_L g938 ( 
.A(n_935),
.B(n_870),
.Y(n_938)
);

AOI22xp33_ASAP7_75t_L g939 ( 
.A1(n_937),
.A2(n_861),
.B1(n_874),
.B2(n_869),
.Y(n_939)
);

BUFx2_ASAP7_75t_L g940 ( 
.A(n_939),
.Y(n_940)
);

AOI221xp5_ASAP7_75t_L g941 ( 
.A1(n_940),
.A2(n_938),
.B1(n_936),
.B2(n_781),
.C(n_780),
.Y(n_941)
);

AOI21xp33_ASAP7_75t_L g942 ( 
.A1(n_941),
.A2(n_791),
.B(n_796),
.Y(n_942)
);

OAI22xp5_ASAP7_75t_L g943 ( 
.A1(n_942),
.A2(n_810),
.B1(n_847),
.B2(n_843),
.Y(n_943)
);

AOI22xp5_ASAP7_75t_L g944 ( 
.A1(n_943),
.A2(n_790),
.B1(n_803),
.B2(n_797),
.Y(n_944)
);


endmodule