module fake_ariane_2173_n_2222 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_213, n_47, n_110, n_153, n_18, n_197, n_221, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_208, n_96, n_156, n_209, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_200, n_51, n_166, n_76, n_218, n_103, n_79, n_26, n_3, n_46, n_220, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_217, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_222, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_214, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_29, n_41, n_219, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_211, n_194, n_97, n_154, n_215, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_216, n_16, n_5, n_155, n_127, n_223, n_35, n_54, n_25, n_2222);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_221;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_96;
input n_156;
input n_209;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_200;
input n_51;
input n_166;
input n_76;
input n_218;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_220;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_217;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_222;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_214;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_29;
input n_41;
input n_219;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_211;
input n_194;
input n_97;
input n_154;
input n_215;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_216;
input n_16;
input n_5;
input n_155;
input n_127;
input n_223;
input n_35;
input n_54;
input n_25;

output n_2222;

wire n_913;
wire n_1681;
wire n_2163;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_2131;
wire n_423;
wire n_1383;
wire n_2182;
wire n_603;
wire n_373;
wire n_2135;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_2207;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_2084;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_945;
wire n_279;
wire n_958;
wire n_813;
wire n_419;
wire n_1985;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_2221;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_2200;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_238;
wire n_365;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_2098;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1654;
wire n_1560;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_2043;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_2116;
wire n_2145;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_2166;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_2185;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_306;
wire n_436;
wire n_324;
wire n_2087;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_967;
wire n_274;
wire n_337;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_2155;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_2172;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_2167;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_976;
wire n_712;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_964;
wire n_1627;
wire n_2220;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_2213;
wire n_1447;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2142;
wire n_1633;
wire n_404;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_2144;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_2120;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_2168;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_2099;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2129;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_2059;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_2122;
wire n_320;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_2195;
wire n_502;
wire n_2194;
wire n_1467;
wire n_247;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_677;
wire n_604;
wire n_439;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_2075;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_2118;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_2125;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_2184;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_2217;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_2211;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_1400;
wire n_342;
wire n_2035;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_2137;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_2032;
wire n_2090;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_2022;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2143;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_2203;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_2158;
wire n_1288;
wire n_1201;
wire n_858;
wire n_1185;
wire n_2173;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_2070;
wire n_2136;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_689;
wire n_400;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_2177;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_2196;
wire n_1038;
wire n_1978;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_2154;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_540;
wire n_692;
wire n_2054;
wire n_1857;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_2189;
wire n_395;
wire n_621;
wire n_1587;
wire n_2093;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_2204;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_2199;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_2180;
wire n_580;
wire n_1579;
wire n_494;
wire n_2181;
wire n_434;
wire n_2014;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_2197;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_2165;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_2169;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_663;
wire n_1720;
wire n_443;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_2096;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_2212;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_2111;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_784;
wire n_648;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_2103;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_2062;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_2153;
wire n_1510;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_2206;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_2101;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_2088;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2108;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2191;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_2085;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_1768;
wire n_2193;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_252;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_415;
wire n_1967;
wire n_2179;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_537;
wire n_1063;
wire n_991;
wire n_2183;
wire n_2205;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_2209;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_2081;
wire n_265;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2152;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_484;
wire n_411;
wire n_849;
wire n_2095;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_2208;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

BUFx8_ASAP7_75t_SL g224 ( 
.A(n_187),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_93),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_101),
.Y(n_226)
);

BUFx5_ASAP7_75t_L g227 ( 
.A(n_151),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_2),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_156),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_222),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_103),
.Y(n_231)
);

BUFx2_ASAP7_75t_L g232 ( 
.A(n_118),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_180),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_97),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_4),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_25),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_203),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_16),
.Y(n_238)
);

BUFx2_ASAP7_75t_L g239 ( 
.A(n_57),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_42),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_141),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_60),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_136),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_53),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_125),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_37),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_186),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_24),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_185),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_105),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_109),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_113),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_10),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_130),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_40),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_207),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_190),
.Y(n_257)
);

BUFx2_ASAP7_75t_SL g258 ( 
.A(n_2),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_91),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_71),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_179),
.Y(n_261)
);

BUFx2_ASAP7_75t_SL g262 ( 
.A(n_39),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_143),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_178),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_223),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_65),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_123),
.Y(n_267)
);

BUFx5_ASAP7_75t_L g268 ( 
.A(n_149),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_64),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_37),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_98),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_211),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_74),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_171),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_83),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_35),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_59),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_131),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_104),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_5),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_20),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_183),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_73),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_81),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_107),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_119),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_63),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_191),
.Y(n_288)
);

INVx2_ASAP7_75t_SL g289 ( 
.A(n_11),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_154),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_100),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_64),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_117),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_92),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_175),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_50),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_58),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_128),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_69),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_39),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_60),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_24),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_159),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_124),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_87),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_169),
.Y(n_306)
);

BUFx3_ASAP7_75t_L g307 ( 
.A(n_36),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_62),
.Y(n_308)
);

BUFx5_ASAP7_75t_L g309 ( 
.A(n_146),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_114),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_121),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_38),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_61),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_26),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_85),
.Y(n_315)
);

BUFx8_ASAP7_75t_SL g316 ( 
.A(n_198),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_194),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_38),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_193),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_116),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_43),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_215),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_102),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_19),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_150),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_192),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_218),
.Y(n_327)
);

BUFx10_ASAP7_75t_L g328 ( 
.A(n_140),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_217),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_86),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_195),
.Y(n_331)
);

INVx1_ASAP7_75t_SL g332 ( 
.A(n_188),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_51),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_202),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_19),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_61),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_152),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_20),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_68),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_54),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_7),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_164),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_112),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_29),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_162),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_68),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_205),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_158),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_88),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_3),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_165),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_86),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_209),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_96),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_78),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_4),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_29),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_44),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_67),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_219),
.Y(n_360)
);

BUFx3_ASAP7_75t_L g361 ( 
.A(n_163),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_51),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_78),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_167),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_213),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_9),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_65),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_170),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_122),
.Y(n_369)
);

BUFx8_ASAP7_75t_SL g370 ( 
.A(n_6),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_85),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_36),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_22),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_14),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_83),
.Y(n_375)
);

BUFx3_ASAP7_75t_L g376 ( 
.A(n_18),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_76),
.Y(n_377)
);

INVx1_ASAP7_75t_SL g378 ( 
.A(n_210),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_221),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_120),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_127),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_95),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_17),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_142),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_52),
.Y(n_385)
);

BUFx10_ASAP7_75t_L g386 ( 
.A(n_47),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_174),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_73),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_212),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_138),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_14),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_200),
.Y(n_392)
);

BUFx10_ASAP7_75t_L g393 ( 
.A(n_99),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_9),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_8),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_173),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_23),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_184),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_139),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_56),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_25),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_94),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_135),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_42),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_137),
.Y(n_405)
);

INVx1_ASAP7_75t_SL g406 ( 
.A(n_160),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_16),
.Y(n_407)
);

INVx2_ASAP7_75t_SL g408 ( 
.A(n_89),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_47),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_49),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_28),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_58),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_176),
.Y(n_413)
);

INVx2_ASAP7_75t_SL g414 ( 
.A(n_189),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_126),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_144),
.Y(n_416)
);

BUFx3_ASAP7_75t_L g417 ( 
.A(n_62),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_110),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_66),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_82),
.Y(n_420)
);

INVx1_ASAP7_75t_SL g421 ( 
.A(n_27),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_26),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_177),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_10),
.Y(n_424)
);

BUFx3_ASAP7_75t_L g425 ( 
.A(n_134),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_35),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_115),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_1),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_74),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_197),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_157),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_22),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_72),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_40),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_53),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_7),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_18),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_111),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_34),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_17),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_370),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_248),
.Y(n_442)
);

INVxp33_ASAP7_75t_SL g443 ( 
.A(n_239),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_257),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_224),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_225),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_316),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_225),
.Y(n_448)
);

INVxp67_ASAP7_75t_SL g449 ( 
.A(n_248),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_264),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_334),
.Y(n_451)
);

INVxp67_ASAP7_75t_SL g452 ( 
.A(n_307),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_226),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_384),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_242),
.Y(n_455)
);

INVxp67_ASAP7_75t_L g456 ( 
.A(n_239),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_226),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_398),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_402),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_228),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_276),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_232),
.B(n_0),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_240),
.Y(n_463)
);

INVxp67_ASAP7_75t_L g464 ( 
.A(n_258),
.Y(n_464)
);

INVxp67_ASAP7_75t_SL g465 ( 
.A(n_307),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_234),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_234),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_232),
.B(n_0),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_246),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_243),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_312),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_243),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_249),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_249),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_314),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_260),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_269),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_250),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_273),
.Y(n_479)
);

CKINVDCx16_ASAP7_75t_R g480 ( 
.A(n_386),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_275),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_250),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_251),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_277),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_376),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_376),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_417),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_417),
.Y(n_488)
);

INVxp67_ASAP7_75t_L g489 ( 
.A(n_258),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_372),
.B(n_1),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_251),
.Y(n_491)
);

NOR2xp67_ASAP7_75t_L g492 ( 
.A(n_289),
.B(n_3),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g493 ( 
.A(n_280),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_259),
.B(n_5),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_259),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_394),
.Y(n_496)
);

CKINVDCx16_ASAP7_75t_R g497 ( 
.A(n_386),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_261),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_404),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_261),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_274),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_274),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_282),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_281),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_282),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_410),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_328),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_288),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_288),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_291),
.Y(n_510)
);

INVxp67_ASAP7_75t_SL g511 ( 
.A(n_235),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_291),
.Y(n_512)
);

INVxp67_ASAP7_75t_SL g513 ( 
.A(n_235),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_294),
.Y(n_514)
);

HB1xp67_ASAP7_75t_L g515 ( 
.A(n_283),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_294),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_298),
.B(n_6),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_298),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_311),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_284),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_311),
.Y(n_521)
);

HB1xp67_ASAP7_75t_L g522 ( 
.A(n_287),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_292),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_326),
.Y(n_524)
);

INVxp33_ASAP7_75t_SL g525 ( 
.A(n_262),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_326),
.Y(n_526)
);

HB1xp67_ASAP7_75t_L g527 ( 
.A(n_296),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_297),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_329),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_300),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_329),
.B(n_8),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_353),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_353),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_354),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_354),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_328),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_301),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_302),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_328),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_308),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_328),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_368),
.Y(n_542)
);

INVxp67_ASAP7_75t_L g543 ( 
.A(n_262),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_361),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_324),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_368),
.Y(n_546)
);

INVxp67_ASAP7_75t_SL g547 ( 
.A(n_236),
.Y(n_547)
);

CKINVDCx20_ASAP7_75t_R g548 ( 
.A(n_393),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_393),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_390),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_338),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_341),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_390),
.Y(n_553)
);

INVxp67_ASAP7_75t_L g554 ( 
.A(n_236),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_346),
.Y(n_555)
);

BUFx2_ASAP7_75t_L g556 ( 
.A(n_289),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_403),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_403),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_446),
.B(n_405),
.Y(n_559)
);

HB1xp67_ASAP7_75t_L g560 ( 
.A(n_456),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_483),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_483),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_446),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_448),
.Y(n_564)
);

NAND2xp33_ASAP7_75t_SL g565 ( 
.A(n_507),
.B(n_356),
.Y(n_565)
);

BUFx2_ASAP7_75t_L g566 ( 
.A(n_455),
.Y(n_566)
);

INVx5_ASAP7_75t_L g567 ( 
.A(n_544),
.Y(n_567)
);

BUFx2_ASAP7_75t_L g568 ( 
.A(n_460),
.Y(n_568)
);

OA21x2_ASAP7_75t_L g569 ( 
.A1(n_448),
.A2(n_431),
.B(n_405),
.Y(n_569)
);

AOI22xp5_ASAP7_75t_L g570 ( 
.A1(n_443),
.A2(n_421),
.B1(n_238),
.B2(n_359),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_453),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_453),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_457),
.B(n_431),
.Y(n_573)
);

AND2x4_ASAP7_75t_L g574 ( 
.A(n_457),
.B(n_466),
.Y(n_574)
);

HB1xp67_ASAP7_75t_L g575 ( 
.A(n_463),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_466),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_467),
.Y(n_577)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_467),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_470),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_470),
.Y(n_580)
);

HB1xp67_ASAP7_75t_L g581 ( 
.A(n_469),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_472),
.Y(n_582)
);

AND2x4_ASAP7_75t_L g583 ( 
.A(n_472),
.B(n_330),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_473),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_473),
.Y(n_585)
);

CKINVDCx8_ASAP7_75t_R g586 ( 
.A(n_445),
.Y(n_586)
);

AND2x4_ASAP7_75t_L g587 ( 
.A(n_474),
.B(n_478),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_474),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_478),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_482),
.B(n_290),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_482),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_458),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_491),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_491),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_480),
.B(n_393),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_495),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_495),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_498),
.B(n_408),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_498),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_500),
.Y(n_600)
);

BUFx8_ASAP7_75t_L g601 ( 
.A(n_556),
.Y(n_601)
);

OR2x2_ASAP7_75t_SL g602 ( 
.A(n_497),
.B(n_330),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_500),
.Y(n_603)
);

AND2x4_ASAP7_75t_L g604 ( 
.A(n_501),
.B(n_366),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_501),
.B(n_408),
.Y(n_605)
);

OAI21x1_ASAP7_75t_L g606 ( 
.A1(n_517),
.A2(n_304),
.B(n_265),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_502),
.Y(n_607)
);

BUFx3_ASAP7_75t_L g608 ( 
.A(n_544),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_502),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_503),
.B(n_366),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_503),
.Y(n_611)
);

BUFx2_ASAP7_75t_L g612 ( 
.A(n_476),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_505),
.Y(n_613)
);

CKINVDCx16_ASAP7_75t_R g614 ( 
.A(n_536),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_505),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_508),
.Y(n_616)
);

AND2x4_ASAP7_75t_L g617 ( 
.A(n_508),
.B(n_373),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_509),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_477),
.B(n_393),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_509),
.Y(n_620)
);

INVx3_ASAP7_75t_L g621 ( 
.A(n_510),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_510),
.Y(n_622)
);

OA21x2_ASAP7_75t_L g623 ( 
.A1(n_512),
.A2(n_304),
.B(n_265),
.Y(n_623)
);

BUFx6f_ASAP7_75t_L g624 ( 
.A(n_512),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_514),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_514),
.Y(n_626)
);

BUFx2_ASAP7_75t_L g627 ( 
.A(n_479),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_525),
.B(n_414),
.Y(n_628)
);

BUFx2_ASAP7_75t_L g629 ( 
.A(n_481),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_516),
.Y(n_630)
);

NAND2xp33_ASAP7_75t_SL g631 ( 
.A(n_539),
.B(n_541),
.Y(n_631)
);

INVx3_ASAP7_75t_L g632 ( 
.A(n_516),
.Y(n_632)
);

AND2x4_ASAP7_75t_L g633 ( 
.A(n_518),
.B(n_373),
.Y(n_633)
);

OA21x2_ASAP7_75t_L g634 ( 
.A1(n_518),
.A2(n_345),
.B(n_319),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_519),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_519),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_521),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_521),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_524),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_464),
.B(n_414),
.Y(n_640)
);

BUFx2_ASAP7_75t_L g641 ( 
.A(n_484),
.Y(n_641)
);

HB1xp67_ASAP7_75t_L g642 ( 
.A(n_504),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_524),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_526),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_526),
.B(n_377),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_529),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_529),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_532),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_532),
.B(n_332),
.Y(n_649)
);

AND2x4_ASAP7_75t_L g650 ( 
.A(n_533),
.B(n_377),
.Y(n_650)
);

AND2x4_ASAP7_75t_L g651 ( 
.A(n_608),
.B(n_511),
.Y(n_651)
);

OR2x2_ASAP7_75t_L g652 ( 
.A(n_560),
.B(n_493),
.Y(n_652)
);

BUFx2_ASAP7_75t_L g653 ( 
.A(n_566),
.Y(n_653)
);

BUFx2_ASAP7_75t_L g654 ( 
.A(n_566),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_572),
.Y(n_655)
);

BUFx10_ASAP7_75t_L g656 ( 
.A(n_628),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_568),
.B(n_520),
.Y(n_657)
);

BUFx6f_ASAP7_75t_L g658 ( 
.A(n_572),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_568),
.B(n_523),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_572),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_572),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_612),
.B(n_528),
.Y(n_662)
);

AOI22xp5_ASAP7_75t_L g663 ( 
.A1(n_640),
.A2(n_468),
.B1(n_462),
.B2(n_619),
.Y(n_663)
);

BUFx3_ASAP7_75t_L g664 ( 
.A(n_608),
.Y(n_664)
);

AND2x4_ASAP7_75t_L g665 ( 
.A(n_608),
.B(n_513),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_572),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_572),
.Y(n_667)
);

AND2x6_ASAP7_75t_L g668 ( 
.A(n_574),
.B(n_319),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_572),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_578),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_612),
.B(n_530),
.Y(n_671)
);

INVx2_ASAP7_75t_SL g672 ( 
.A(n_574),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_578),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_592),
.Y(n_674)
);

AND2x2_ASAP7_75t_SL g675 ( 
.A(n_627),
.B(n_494),
.Y(n_675)
);

OAI22xp5_ASAP7_75t_L g676 ( 
.A1(n_570),
.A2(n_489),
.B1(n_543),
.B2(n_560),
.Y(n_676)
);

AND2x6_ASAP7_75t_L g677 ( 
.A(n_574),
.B(n_345),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_578),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_595),
.B(n_537),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_578),
.Y(n_680)
);

NOR3xp33_ASAP7_75t_L g681 ( 
.A(n_627),
.B(n_531),
.C(n_395),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_578),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_578),
.Y(n_683)
);

INVx3_ASAP7_75t_L g684 ( 
.A(n_578),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_649),
.B(n_538),
.Y(n_685)
);

AOI22xp5_ASAP7_75t_L g686 ( 
.A1(n_570),
.A2(n_540),
.B1(n_551),
.B2(n_545),
.Y(n_686)
);

INVx3_ASAP7_75t_L g687 ( 
.A(n_584),
.Y(n_687)
);

BUFx2_ASAP7_75t_L g688 ( 
.A(n_629),
.Y(n_688)
);

INVx2_ASAP7_75t_SL g689 ( 
.A(n_574),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_584),
.Y(n_690)
);

NAND3xp33_ASAP7_75t_L g691 ( 
.A(n_649),
.B(n_555),
.C(n_552),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_571),
.B(n_515),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_584),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_574),
.B(n_533),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_629),
.B(n_447),
.Y(n_695)
);

BUFx2_ASAP7_75t_L g696 ( 
.A(n_641),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_587),
.B(n_449),
.Y(n_697)
);

INVx3_ASAP7_75t_L g698 ( 
.A(n_584),
.Y(n_698)
);

INVx4_ASAP7_75t_L g699 ( 
.A(n_567),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_584),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_571),
.B(n_522),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_584),
.Y(n_702)
);

AOI22xp5_ASAP7_75t_L g703 ( 
.A1(n_641),
.A2(n_492),
.B1(n_549),
.B2(n_548),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_584),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_577),
.Y(n_705)
);

XOR2xp5_ASAP7_75t_R g706 ( 
.A(n_601),
.B(n_490),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_577),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_600),
.Y(n_708)
);

AOI22xp33_ASAP7_75t_L g709 ( 
.A1(n_623),
.A2(n_556),
.B1(n_535),
.B2(n_542),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_587),
.B(n_527),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_600),
.Y(n_711)
);

INVx3_ASAP7_75t_L g712 ( 
.A(n_600),
.Y(n_712)
);

INVx1_ASAP7_75t_SL g713 ( 
.A(n_575),
.Y(n_713)
);

AOI22xp5_ASAP7_75t_L g714 ( 
.A1(n_575),
.A2(n_547),
.B1(n_465),
.B2(n_452),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_580),
.B(n_534),
.Y(n_715)
);

AND2x2_ASAP7_75t_L g716 ( 
.A(n_587),
.B(n_534),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_587),
.B(n_535),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_587),
.B(n_542),
.Y(n_718)
);

AOI22xp5_ASAP7_75t_L g719 ( 
.A1(n_581),
.A2(n_554),
.B1(n_362),
.B2(n_363),
.Y(n_719)
);

AND2x6_ASAP7_75t_L g720 ( 
.A(n_580),
.B(n_387),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_581),
.B(n_546),
.Y(n_721)
);

INVx4_ASAP7_75t_L g722 ( 
.A(n_567),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_576),
.B(n_546),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_582),
.B(n_550),
.Y(n_724)
);

NAND3xp33_ASAP7_75t_L g725 ( 
.A(n_642),
.B(n_558),
.C(n_553),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_600),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_610),
.B(n_550),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_600),
.Y(n_728)
);

BUFx6f_ASAP7_75t_L g729 ( 
.A(n_600),
.Y(n_729)
);

NAND2xp33_ASAP7_75t_L g730 ( 
.A(n_600),
.B(n_227),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_582),
.Y(n_731)
);

BUFx8_ASAP7_75t_SL g732 ( 
.A(n_586),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_611),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_611),
.Y(n_734)
);

BUFx2_ASAP7_75t_L g735 ( 
.A(n_601),
.Y(n_735)
);

INVx4_ASAP7_75t_L g736 ( 
.A(n_567),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_611),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_611),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_611),
.Y(n_739)
);

AO22x2_ASAP7_75t_L g740 ( 
.A1(n_601),
.A2(n_553),
.B1(n_558),
.B2(n_557),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_642),
.B(n_557),
.Y(n_741)
);

BUFx3_ASAP7_75t_L g742 ( 
.A(n_567),
.Y(n_742)
);

INVx3_ASAP7_75t_L g743 ( 
.A(n_611),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_611),
.Y(n_744)
);

AOI22xp33_ASAP7_75t_L g745 ( 
.A1(n_623),
.A2(n_424),
.B1(n_428),
.B2(n_391),
.Y(n_745)
);

INVx4_ASAP7_75t_L g746 ( 
.A(n_567),
.Y(n_746)
);

NAND3xp33_ASAP7_75t_L g747 ( 
.A(n_585),
.B(n_367),
.C(n_358),
.Y(n_747)
);

AO21x2_ASAP7_75t_L g748 ( 
.A1(n_606),
.A2(n_427),
.B(n_387),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_585),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_624),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_624),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_576),
.B(n_621),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_601),
.B(n_386),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_624),
.Y(n_754)
);

OR2x6_ASAP7_75t_L g755 ( 
.A(n_610),
.B(n_442),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_624),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_624),
.Y(n_757)
);

INVx4_ASAP7_75t_L g758 ( 
.A(n_567),
.Y(n_758)
);

OR2x2_ASAP7_75t_L g759 ( 
.A(n_602),
.B(n_485),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_624),
.Y(n_760)
);

NAND2xp33_ASAP7_75t_L g761 ( 
.A(n_624),
.B(n_227),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_643),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_643),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_643),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_L g765 ( 
.A(n_588),
.B(n_486),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_588),
.B(n_487),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_576),
.B(n_488),
.Y(n_767)
);

BUFx2_ASAP7_75t_L g768 ( 
.A(n_601),
.Y(n_768)
);

BUFx6f_ASAP7_75t_L g769 ( 
.A(n_643),
.Y(n_769)
);

AOI22xp5_ASAP7_75t_L g770 ( 
.A1(n_565),
.A2(n_374),
.B1(n_375),
.B2(n_371),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_643),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_643),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_610),
.B(n_386),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_643),
.Y(n_774)
);

INVx3_ASAP7_75t_L g775 ( 
.A(n_576),
.Y(n_775)
);

INVx3_ASAP7_75t_L g776 ( 
.A(n_621),
.Y(n_776)
);

AND2x6_ASAP7_75t_L g777 ( 
.A(n_591),
.B(n_427),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_621),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_621),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_632),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_632),
.B(n_378),
.Y(n_781)
);

INVx1_ASAP7_75t_SL g782 ( 
.A(n_631),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_632),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_563),
.Y(n_784)
);

AO21x2_ASAP7_75t_L g785 ( 
.A1(n_606),
.A2(n_253),
.B(n_244),
.Y(n_785)
);

AND2x2_ASAP7_75t_L g786 ( 
.A(n_645),
.B(n_244),
.Y(n_786)
);

NOR3xp33_ASAP7_75t_L g787 ( 
.A(n_614),
.B(n_255),
.C(n_253),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_563),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_632),
.B(n_591),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_593),
.B(n_406),
.Y(n_790)
);

AOI21x1_ASAP7_75t_L g791 ( 
.A1(n_606),
.A2(n_266),
.B(n_255),
.Y(n_791)
);

OR2x6_ASAP7_75t_L g792 ( 
.A(n_645),
.B(n_391),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_563),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_593),
.B(n_229),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_594),
.Y(n_795)
);

INVx3_ASAP7_75t_L g796 ( 
.A(n_564),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_594),
.B(n_230),
.Y(n_797)
);

AND2x2_ASAP7_75t_SL g798 ( 
.A(n_569),
.B(n_424),
.Y(n_798)
);

OAI22xp33_ASAP7_75t_L g799 ( 
.A1(n_598),
.A2(n_383),
.B1(n_385),
.B2(n_397),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_564),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_596),
.Y(n_801)
);

AOI22xp33_ASAP7_75t_L g802 ( 
.A1(n_623),
.A2(n_428),
.B1(n_357),
.B2(n_318),
.Y(n_802)
);

OAI22xp33_ASAP7_75t_L g803 ( 
.A1(n_598),
.A2(n_605),
.B1(n_590),
.B2(n_573),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_564),
.Y(n_804)
);

INVx5_ASAP7_75t_L g805 ( 
.A(n_567),
.Y(n_805)
);

INVx1_ASAP7_75t_SL g806 ( 
.A(n_614),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_596),
.B(n_231),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_645),
.B(n_266),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_685),
.B(n_599),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_784),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_803),
.B(n_599),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_716),
.B(n_603),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_716),
.B(n_603),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_672),
.B(n_607),
.Y(n_814)
);

OR2x2_ASAP7_75t_L g815 ( 
.A(n_713),
.B(n_602),
.Y(n_815)
);

A2O1A1Ixp33_ASAP7_75t_L g816 ( 
.A1(n_672),
.A2(n_573),
.B(n_559),
.C(n_579),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_689),
.B(n_607),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_689),
.B(n_613),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_784),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_697),
.B(n_613),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_697),
.B(n_618),
.Y(n_821)
);

BUFx3_ASAP7_75t_L g822 ( 
.A(n_664),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_778),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_675),
.B(n_618),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_788),
.Y(n_825)
);

INVx8_ASAP7_75t_L g826 ( 
.A(n_732),
.Y(n_826)
);

INVx2_ASAP7_75t_SL g827 ( 
.A(n_653),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_778),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_788),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_727),
.B(n_620),
.Y(n_830)
);

INVxp67_ASAP7_75t_L g831 ( 
.A(n_653),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_727),
.B(n_620),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_651),
.B(n_626),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_651),
.B(n_626),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_688),
.B(n_696),
.Y(n_835)
);

AOI21xp5_ASAP7_75t_L g836 ( 
.A1(n_752),
.A2(n_605),
.B(n_559),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_651),
.B(n_630),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_793),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_793),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_779),
.Y(n_840)
);

NAND2xp33_ASAP7_75t_SL g841 ( 
.A(n_674),
.B(n_630),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_800),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_665),
.B(n_635),
.Y(n_843)
);

NAND2xp33_ASAP7_75t_L g844 ( 
.A(n_668),
.B(n_635),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_800),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_675),
.B(n_636),
.Y(n_846)
);

OAI22xp5_ASAP7_75t_L g847 ( 
.A1(n_663),
.A2(n_636),
.B1(n_639),
.B2(n_638),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_688),
.B(n_586),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_798),
.B(n_638),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_665),
.B(n_639),
.Y(n_850)
);

NOR3xp33_ASAP7_75t_L g851 ( 
.A(n_696),
.B(n_299),
.C(n_270),
.Y(n_851)
);

INVx5_ASAP7_75t_L g852 ( 
.A(n_668),
.Y(n_852)
);

NAND2x1p5_ASAP7_75t_L g853 ( 
.A(n_735),
.B(n_579),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_798),
.B(n_646),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_796),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_665),
.B(n_646),
.Y(n_856)
);

O2A1O1Ixp33_ASAP7_75t_L g857 ( 
.A1(n_694),
.A2(n_647),
.B(n_589),
.C(n_597),
.Y(n_857)
);

BUFx2_ASAP7_75t_L g858 ( 
.A(n_654),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_775),
.B(n_776),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_656),
.B(n_679),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_796),
.Y(n_861)
);

INVxp67_ASAP7_75t_L g862 ( 
.A(n_654),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_796),
.Y(n_863)
);

AOI22xp33_ASAP7_75t_L g864 ( 
.A1(n_740),
.A2(n_623),
.B1(n_634),
.B2(n_569),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_775),
.B(n_647),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_779),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_775),
.B(n_579),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_780),
.Y(n_868)
);

AOI22xp5_ASAP7_75t_L g869 ( 
.A1(n_668),
.A2(n_590),
.B1(n_597),
.B2(n_589),
.Y(n_869)
);

INVx2_ASAP7_75t_SL g870 ( 
.A(n_773),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_780),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_773),
.B(n_589),
.Y(n_872)
);

AND2x2_ASAP7_75t_L g873 ( 
.A(n_652),
.B(n_586),
.Y(n_873)
);

NAND2xp33_ASAP7_75t_L g874 ( 
.A(n_668),
.B(n_597),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_776),
.B(n_609),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_804),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_776),
.B(n_609),
.Y(n_877)
);

OAI22xp5_ASAP7_75t_L g878 ( 
.A1(n_705),
.A2(n_615),
.B1(n_616),
.B2(n_609),
.Y(n_878)
);

HB1xp67_ASAP7_75t_L g879 ( 
.A(n_652),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_658),
.B(n_615),
.Y(n_880)
);

NAND2xp33_ASAP7_75t_L g881 ( 
.A(n_668),
.B(n_615),
.Y(n_881)
);

NOR2x1p5_ASAP7_75t_L g882 ( 
.A(n_674),
.B(n_441),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_L g883 ( 
.A(n_656),
.B(n_444),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_692),
.B(n_616),
.Y(n_884)
);

BUFx5_ASAP7_75t_L g885 ( 
.A(n_668),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_783),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_658),
.B(n_729),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_701),
.B(n_616),
.Y(n_888)
);

INVx2_ASAP7_75t_SL g889 ( 
.A(n_759),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_804),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_715),
.B(n_622),
.Y(n_891)
);

BUFx6f_ASAP7_75t_SL g892 ( 
.A(n_732),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_SL g893 ( 
.A(n_658),
.B(n_622),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_724),
.B(n_709),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_783),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_707),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_658),
.B(n_622),
.Y(n_897)
);

INVxp33_ASAP7_75t_L g898 ( 
.A(n_686),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_731),
.Y(n_899)
);

INVxp33_ASAP7_75t_L g900 ( 
.A(n_676),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_661),
.Y(n_901)
);

NAND3xp33_ASAP7_75t_L g902 ( 
.A(n_725),
.B(n_490),
.C(n_625),
.Y(n_902)
);

NOR2xp67_ASAP7_75t_L g903 ( 
.A(n_691),
.B(n_625),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_661),
.Y(n_904)
);

OAI22xp33_ASAP7_75t_L g905 ( 
.A1(n_755),
.A2(n_625),
.B1(n_648),
.B2(n_644),
.Y(n_905)
);

AO22x2_ASAP7_75t_L g906 ( 
.A1(n_753),
.A2(n_435),
.B1(n_299),
.B2(n_313),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_790),
.B(n_637),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_656),
.B(n_450),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_666),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_781),
.B(n_637),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_749),
.Y(n_911)
);

NAND2xp33_ASAP7_75t_SL g912 ( 
.A(n_735),
.B(n_637),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_795),
.B(n_801),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_789),
.Y(n_914)
);

AOI22xp5_ASAP7_75t_L g915 ( 
.A1(n_677),
.A2(n_644),
.B1(n_648),
.B2(n_650),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_666),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_SL g917 ( 
.A(n_658),
.B(n_644),
.Y(n_917)
);

BUFx5_ASAP7_75t_L g918 ( 
.A(n_677),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_755),
.B(n_451),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_690),
.Y(n_920)
);

INVx2_ASAP7_75t_SL g921 ( 
.A(n_759),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_755),
.B(n_454),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_717),
.B(n_648),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_SL g924 ( 
.A(n_729),
.B(n_583),
.Y(n_924)
);

BUFx6f_ASAP7_75t_L g925 ( 
.A(n_729),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_767),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_723),
.Y(n_927)
);

INVx2_ASAP7_75t_SL g928 ( 
.A(n_786),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_718),
.Y(n_929)
);

INVxp67_ASAP7_75t_SL g930 ( 
.A(n_664),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_690),
.Y(n_931)
);

INVx2_ASAP7_75t_SL g932 ( 
.A(n_786),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_721),
.B(n_741),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_SL g934 ( 
.A(n_729),
.B(n_583),
.Y(n_934)
);

BUFx3_ASAP7_75t_L g935 ( 
.A(n_768),
.Y(n_935)
);

AOI22xp33_ASAP7_75t_L g936 ( 
.A1(n_740),
.A2(n_634),
.B1(n_623),
.B2(n_569),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_700),
.Y(n_937)
);

INVxp67_ASAP7_75t_L g938 ( 
.A(n_806),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_765),
.B(n_583),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_766),
.B(n_583),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_729),
.B(n_583),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_808),
.B(n_604),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_808),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_657),
.B(n_459),
.Y(n_944)
);

AND2x4_ASAP7_75t_L g945 ( 
.A(n_792),
.B(n_604),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_794),
.B(n_604),
.Y(n_946)
);

AND2x6_ASAP7_75t_SL g947 ( 
.A(n_755),
.B(n_270),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_655),
.Y(n_948)
);

NAND2xp33_ASAP7_75t_SL g949 ( 
.A(n_768),
.B(n_313),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_655),
.A2(n_569),
.B(n_634),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_L g951 ( 
.A(n_659),
.B(n_662),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_797),
.B(n_604),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_807),
.B(n_792),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_700),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_660),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_769),
.B(n_604),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_792),
.B(n_617),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_SL g958 ( 
.A(n_769),
.B(n_617),
.Y(n_958)
);

AOI22xp5_ASAP7_75t_L g959 ( 
.A1(n_677),
.A2(n_650),
.B1(n_633),
.B2(n_617),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_769),
.B(n_617),
.Y(n_960)
);

NAND2xp33_ASAP7_75t_L g961 ( 
.A(n_677),
.B(n_401),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_660),
.A2(n_569),
.B(n_634),
.Y(n_962)
);

BUFx4_ASAP7_75t_L g963 ( 
.A(n_706),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_792),
.B(n_617),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_671),
.B(n_461),
.Y(n_965)
);

NOR2x1p5_ASAP7_75t_L g966 ( 
.A(n_706),
.B(n_411),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_L g967 ( 
.A(n_714),
.B(n_471),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_677),
.B(n_633),
.Y(n_968)
);

AOI22xp33_ASAP7_75t_L g969 ( 
.A1(n_740),
.A2(n_634),
.B1(n_650),
.B2(n_633),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_SL g970 ( 
.A(n_769),
.B(n_633),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_702),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_677),
.B(n_633),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_667),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_L g974 ( 
.A(n_710),
.B(n_475),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_802),
.B(n_650),
.Y(n_975)
);

BUFx6f_ASAP7_75t_L g976 ( 
.A(n_769),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_799),
.B(n_650),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_745),
.B(n_561),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_681),
.B(n_561),
.Y(n_979)
);

BUFx8_ASAP7_75t_L g980 ( 
.A(n_720),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_SL g981 ( 
.A(n_684),
.B(n_562),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_667),
.Y(n_982)
);

NOR2xp33_ASAP7_75t_L g983 ( 
.A(n_860),
.B(n_496),
.Y(n_983)
);

OAI21xp5_ASAP7_75t_L g984 ( 
.A1(n_950),
.A2(n_670),
.B(n_669),
.Y(n_984)
);

AOI22xp5_ASAP7_75t_L g985 ( 
.A1(n_900),
.A2(n_740),
.B1(n_719),
.B2(n_782),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_914),
.B(n_684),
.Y(n_986)
);

OR2x2_ASAP7_75t_L g987 ( 
.A(n_879),
.B(n_703),
.Y(n_987)
);

NOR2x1_ASAP7_75t_L g988 ( 
.A(n_848),
.B(n_935),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_887),
.A2(n_670),
.B(n_669),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_SL g990 ( 
.A(n_873),
.B(n_841),
.Y(n_990)
);

BUFx6f_ASAP7_75t_L g991 ( 
.A(n_925),
.Y(n_991)
);

BUFx4f_ASAP7_75t_L g992 ( 
.A(n_826),
.Y(n_992)
);

NOR3xp33_ASAP7_75t_L g993 ( 
.A(n_841),
.B(n_695),
.C(n_747),
.Y(n_993)
);

OAI21xp33_ASAP7_75t_L g994 ( 
.A1(n_809),
.A2(n_770),
.B(n_419),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_895),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_927),
.B(n_684),
.Y(n_996)
);

AOI22xp5_ASAP7_75t_L g997 ( 
.A1(n_900),
.A2(n_777),
.B1(n_720),
.B2(n_787),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_887),
.A2(n_836),
.B(n_859),
.Y(n_998)
);

NOR2x1_ASAP7_75t_R g999 ( 
.A(n_858),
.B(n_412),
.Y(n_999)
);

NOR2xp33_ASAP7_75t_L g1000 ( 
.A(n_898),
.B(n_499),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_859),
.A2(n_678),
.B(n_673),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_926),
.B(n_687),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_849),
.A2(n_678),
.B(n_673),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_895),
.Y(n_1004)
);

OAI221xp5_ASAP7_75t_L g1005 ( 
.A1(n_870),
.A2(n_420),
.B1(n_422),
.B2(n_429),
.C(n_433),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_823),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_828),
.Y(n_1007)
);

BUFx6f_ASAP7_75t_L g1008 ( 
.A(n_925),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_840),
.Y(n_1009)
);

BUFx6f_ASAP7_75t_L g1010 ( 
.A(n_925),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_849),
.A2(n_682),
.B(n_680),
.Y(n_1011)
);

NOR2x1_ASAP7_75t_R g1012 ( 
.A(n_827),
.B(n_434),
.Y(n_1012)
);

AND2x2_ASAP7_75t_L g1013 ( 
.A(n_835),
.B(n_506),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_884),
.B(n_720),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_888),
.B(n_720),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_928),
.B(n_932),
.Y(n_1016)
);

O2A1O1Ixp33_ASAP7_75t_L g1017 ( 
.A1(n_824),
.A2(n_318),
.B(n_321),
.C(n_315),
.Y(n_1017)
);

BUFx6f_ASAP7_75t_L g1018 ( 
.A(n_925),
.Y(n_1018)
);

AND2x4_ASAP7_75t_L g1019 ( 
.A(n_945),
.B(n_935),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_854),
.A2(n_682),
.B(n_680),
.Y(n_1020)
);

AOI21x1_ASAP7_75t_L g1021 ( 
.A1(n_854),
.A2(n_791),
.B(n_693),
.Y(n_1021)
);

NOR2x1p5_ASAP7_75t_SL g1022 ( 
.A(n_885),
.B(n_791),
.Y(n_1022)
);

INVx3_ASAP7_75t_L g1023 ( 
.A(n_822),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_810),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_872),
.B(n_720),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_810),
.Y(n_1026)
);

BUFx6f_ASAP7_75t_L g1027 ( 
.A(n_976),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_811),
.A2(n_693),
.B(n_683),
.Y(n_1028)
);

NOR2x1_ASAP7_75t_L g1029 ( 
.A(n_822),
.B(n_562),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_812),
.B(n_687),
.Y(n_1030)
);

NAND2x1p5_ASAP7_75t_L g1031 ( 
.A(n_852),
.B(n_687),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_813),
.B(n_698),
.Y(n_1032)
);

AO21x1_ASAP7_75t_L g1033 ( 
.A1(n_824),
.A2(n_711),
.B(n_683),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_817),
.A2(n_726),
.B(n_711),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_SL g1035 ( 
.A(n_852),
.B(n_698),
.Y(n_1035)
);

A2O1A1Ixp33_ASAP7_75t_L g1036 ( 
.A1(n_933),
.A2(n_712),
.B(n_698),
.C(n_743),
.Y(n_1036)
);

AOI22xp33_ASAP7_75t_L g1037 ( 
.A1(n_898),
.A2(n_720),
.B1(n_777),
.B2(n_733),
.Y(n_1037)
);

INVx3_ASAP7_75t_L g1038 ( 
.A(n_976),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_L g1039 ( 
.A(n_831),
.B(n_712),
.Y(n_1039)
);

OAI22xp5_ASAP7_75t_L g1040 ( 
.A1(n_814),
.A2(n_712),
.B1(n_743),
.B2(n_726),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_817),
.A2(n_737),
.B(n_728),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_819),
.Y(n_1042)
);

AND2x4_ASAP7_75t_L g1043 ( 
.A(n_945),
.B(n_777),
.Y(n_1043)
);

OAI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_962),
.A2(n_737),
.B(n_728),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_SL g1045 ( 
.A(n_852),
.B(n_743),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_820),
.B(n_738),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_821),
.B(n_738),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_907),
.B(n_754),
.Y(n_1048)
);

AOI22xp5_ASAP7_75t_L g1049 ( 
.A1(n_846),
.A2(n_777),
.B1(n_754),
.B2(n_760),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_876),
.B(n_760),
.Y(n_1050)
);

O2A1O1Ixp33_ASAP7_75t_L g1051 ( 
.A1(n_846),
.A2(n_315),
.B(n_321),
.C(n_333),
.Y(n_1051)
);

BUFx2_ASAP7_75t_L g1052 ( 
.A(n_862),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_866),
.Y(n_1053)
);

BUFx4f_ASAP7_75t_L g1054 ( 
.A(n_826),
.Y(n_1054)
);

OAI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_816),
.A2(n_764),
.B(n_763),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_891),
.A2(n_764),
.B(n_763),
.Y(n_1056)
);

AND2x2_ASAP7_75t_L g1057 ( 
.A(n_974),
.B(n_333),
.Y(n_1057)
);

BUFx3_ASAP7_75t_L g1058 ( 
.A(n_826),
.Y(n_1058)
);

OAI22xp5_ASAP7_75t_L g1059 ( 
.A1(n_818),
.A2(n_756),
.B1(n_733),
.B2(n_774),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_867),
.A2(n_704),
.B(n_702),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_867),
.A2(n_708),
.B(n_704),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_852),
.B(n_885),
.Y(n_1062)
);

AOI21x1_ASAP7_75t_L g1063 ( 
.A1(n_880),
.A2(n_734),
.B(n_708),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_875),
.A2(n_739),
.B(n_734),
.Y(n_1064)
);

AOI21x1_ASAP7_75t_L g1065 ( 
.A1(n_880),
.A2(n_744),
.B(n_739),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_875),
.A2(n_750),
.B(n_744),
.Y(n_1066)
);

AOI22xp5_ASAP7_75t_L g1067 ( 
.A1(n_951),
.A2(n_777),
.B1(n_751),
.B2(n_750),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_876),
.B(n_751),
.Y(n_1068)
);

OAI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_816),
.A2(n_757),
.B(n_756),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_943),
.B(n_777),
.Y(n_1070)
);

AOI22xp5_ASAP7_75t_L g1071 ( 
.A1(n_949),
.A2(n_762),
.B1(n_757),
.B2(n_774),
.Y(n_1071)
);

NOR2x1_ASAP7_75t_L g1072 ( 
.A(n_882),
.B(n_762),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_819),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_877),
.A2(n_772),
.B(n_771),
.Y(n_1074)
);

AO21x1_ASAP7_75t_L g1075 ( 
.A1(n_905),
.A2(n_761),
.B(n_730),
.Y(n_1075)
);

A2O1A1Ixp33_ASAP7_75t_L g1076 ( 
.A1(n_953),
.A2(n_772),
.B(n_771),
.C(n_730),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_877),
.A2(n_761),
.B(n_785),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_910),
.A2(n_785),
.B(n_748),
.Y(n_1078)
);

BUFx3_ASAP7_75t_L g1079 ( 
.A(n_919),
.Y(n_1079)
);

AOI21xp33_ASAP7_75t_L g1080 ( 
.A1(n_967),
.A2(n_748),
.B(n_439),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_893),
.A2(n_785),
.B(n_748),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_890),
.B(n_699),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_890),
.B(n_699),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_868),
.Y(n_1084)
);

NOR2xp33_ASAP7_75t_SL g1085 ( 
.A(n_892),
.B(n_436),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_894),
.B(n_699),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_893),
.A2(n_736),
.B(n_722),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_833),
.B(n_722),
.Y(n_1088)
);

NOR2xp33_ASAP7_75t_L g1089 ( 
.A(n_883),
.B(n_335),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_871),
.Y(n_1090)
);

OAI21xp33_ASAP7_75t_L g1091 ( 
.A1(n_830),
.A2(n_336),
.B(n_335),
.Y(n_1091)
);

OAI22xp5_ASAP7_75t_L g1092 ( 
.A1(n_832),
.A2(n_336),
.B1(n_339),
.B2(n_340),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_897),
.A2(n_736),
.B(n_722),
.Y(n_1093)
);

OAI22xp5_ASAP7_75t_L g1094 ( 
.A1(n_913),
.A2(n_339),
.B1(n_340),
.B2(n_344),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_834),
.B(n_736),
.Y(n_1095)
);

O2A1O1Ixp33_ASAP7_75t_L g1096 ( 
.A1(n_942),
.A2(n_344),
.B(n_350),
.C(n_352),
.Y(n_1096)
);

INVx3_ASAP7_75t_L g1097 ( 
.A(n_976),
.Y(n_1097)
);

NOR2x1_ASAP7_75t_L g1098 ( 
.A(n_908),
.B(n_361),
.Y(n_1098)
);

INVx4_ASAP7_75t_L g1099 ( 
.A(n_892),
.Y(n_1099)
);

AND2x2_ASAP7_75t_L g1100 ( 
.A(n_889),
.B(n_350),
.Y(n_1100)
);

AO21x1_ASAP7_75t_L g1101 ( 
.A1(n_847),
.A2(n_355),
.B(n_352),
.Y(n_1101)
);

OAI22xp5_ASAP7_75t_L g1102 ( 
.A1(n_837),
.A2(n_355),
.B1(n_357),
.B2(n_388),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_825),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_843),
.B(n_850),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_897),
.A2(n_758),
.B(n_746),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_856),
.B(n_746),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_896),
.B(n_746),
.Y(n_1107)
);

CKINVDCx20_ASAP7_75t_R g1108 ( 
.A(n_938),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_899),
.B(n_758),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_825),
.Y(n_1110)
);

AND2x4_ASAP7_75t_L g1111 ( 
.A(n_945),
.B(n_742),
.Y(n_1111)
);

INVx3_ASAP7_75t_L g1112 ( 
.A(n_976),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_911),
.B(n_758),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_917),
.A2(n_742),
.B(n_805),
.Y(n_1114)
);

OAI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_865),
.A2(n_805),
.B(n_400),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_917),
.A2(n_805),
.B(n_237),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_865),
.A2(n_805),
.B(n_241),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_946),
.A2(n_805),
.B(n_245),
.Y(n_1118)
);

A2O1A1Ixp33_ASAP7_75t_L g1119 ( 
.A1(n_886),
.A2(n_440),
.B(n_388),
.C(n_437),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_923),
.Y(n_1120)
);

NOR2xp33_ASAP7_75t_L g1121 ( 
.A(n_815),
.B(n_400),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_SL g1122 ( 
.A(n_885),
.B(n_233),
.Y(n_1122)
);

OAI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_952),
.A2(n_409),
.B(n_407),
.Y(n_1123)
);

AND2x2_ASAP7_75t_L g1124 ( 
.A(n_921),
.B(n_407),
.Y(n_1124)
);

INVxp67_ASAP7_75t_L g1125 ( 
.A(n_922),
.Y(n_1125)
);

OAI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_857),
.A2(n_426),
.B(n_409),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_939),
.B(n_426),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_981),
.A2(n_861),
.B(n_855),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_940),
.B(n_432),
.Y(n_1129)
);

OAI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_948),
.A2(n_440),
.B(n_432),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_979),
.B(n_435),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_929),
.B(n_957),
.Y(n_1132)
);

AND2x2_ASAP7_75t_L g1133 ( 
.A(n_965),
.B(n_944),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_964),
.B(n_437),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_930),
.B(n_247),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_981),
.A2(n_438),
.B(n_430),
.Y(n_1136)
);

AND2x2_ASAP7_75t_L g1137 ( 
.A(n_851),
.B(n_425),
.Y(n_1137)
);

NOR2xp33_ASAP7_75t_SL g1138 ( 
.A(n_980),
.B(n_252),
.Y(n_1138)
);

AOI22xp5_ASAP7_75t_L g1139 ( 
.A1(n_949),
.A2(n_331),
.B1(n_254),
.B2(n_418),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_855),
.A2(n_327),
.B(n_267),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_861),
.A2(n_337),
.B(n_271),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_863),
.A2(n_342),
.B(n_272),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_863),
.A2(n_343),
.B(n_278),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_SL g1144 ( 
.A(n_885),
.B(n_256),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_R g1145 ( 
.A(n_912),
.B(n_263),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_959),
.B(n_279),
.Y(n_1146)
);

AOI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_906),
.A2(n_874),
.B1(n_881),
.B2(n_844),
.Y(n_1147)
);

NOR2xp33_ASAP7_75t_L g1148 ( 
.A(n_902),
.B(n_285),
.Y(n_1148)
);

NAND2x1p5_ASAP7_75t_L g1149 ( 
.A(n_924),
.B(n_425),
.Y(n_1149)
);

AOI22xp5_ASAP7_75t_L g1150 ( 
.A1(n_906),
.A2(n_349),
.B1(n_416),
.B2(n_415),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_955),
.A2(n_347),
.B(n_413),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_906),
.B(n_286),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_973),
.A2(n_348),
.B(n_399),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_982),
.A2(n_325),
.B(n_396),
.Y(n_1154)
);

AOI22xp5_ASAP7_75t_L g1155 ( 
.A1(n_968),
.A2(n_323),
.B1(n_392),
.B2(n_389),
.Y(n_1155)
);

INVx1_ASAP7_75t_SL g1156 ( 
.A(n_963),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_901),
.A2(n_320),
.B(n_382),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_901),
.A2(n_317),
.B(n_381),
.Y(n_1158)
);

O2A1O1Ixp33_ASAP7_75t_L g1159 ( 
.A1(n_924),
.A2(n_11),
.B(n_12),
.C(n_13),
.Y(n_1159)
);

AND2x4_ASAP7_75t_L g1160 ( 
.A(n_972),
.B(n_12),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_904),
.A2(n_310),
.B(n_380),
.Y(n_1161)
);

INVx1_ASAP7_75t_SL g1162 ( 
.A(n_947),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_904),
.A2(n_909),
.B(n_916),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_829),
.B(n_227),
.Y(n_1164)
);

NOR2xp33_ASAP7_75t_L g1165 ( 
.A(n_853),
.B(n_293),
.Y(n_1165)
);

INVxp67_ASAP7_75t_L g1166 ( 
.A(n_903),
.Y(n_1166)
);

A2O1A1Ixp33_ASAP7_75t_L g1167 ( 
.A1(n_869),
.A2(n_351),
.B(n_379),
.C(n_369),
.Y(n_1167)
);

INVx2_ASAP7_75t_SL g1168 ( 
.A(n_966),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_909),
.A2(n_306),
.B(n_365),
.Y(n_1169)
);

INVxp67_ASAP7_75t_SL g1170 ( 
.A(n_980),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_916),
.A2(n_305),
.B(n_364),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_829),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_920),
.A2(n_303),
.B(n_360),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_838),
.B(n_839),
.Y(n_1174)
);

NAND3xp33_ASAP7_75t_L g1175 ( 
.A(n_934),
.B(n_322),
.C(n_295),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_920),
.A2(n_423),
.B(n_309),
.Y(n_1176)
);

INVx6_ASAP7_75t_L g1177 ( 
.A(n_1019),
.Y(n_1177)
);

O2A1O1Ixp33_ASAP7_75t_L g1178 ( 
.A1(n_1089),
.A2(n_878),
.B(n_977),
.C(n_956),
.Y(n_1178)
);

NOR2xp33_ASAP7_75t_SL g1179 ( 
.A(n_1108),
.B(n_980),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_SL g1180 ( 
.A(n_1133),
.B(n_885),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_998),
.A2(n_961),
.B(n_941),
.Y(n_1181)
);

AOI22xp5_ASAP7_75t_L g1182 ( 
.A1(n_983),
.A2(n_885),
.B1(n_918),
.B2(n_915),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_SL g1183 ( 
.A(n_1019),
.B(n_885),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_1004),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1104),
.B(n_853),
.Y(n_1185)
);

NAND2xp33_ASAP7_75t_L g1186 ( 
.A(n_991),
.B(n_918),
.Y(n_1186)
);

BUFx6f_ASAP7_75t_L g1187 ( 
.A(n_991),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1104),
.B(n_918),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_1046),
.A2(n_956),
.B(n_934),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_995),
.Y(n_1190)
);

A2O1A1Ixp33_ASAP7_75t_SL g1191 ( 
.A1(n_1039),
.A2(n_937),
.B(n_931),
.C(n_971),
.Y(n_1191)
);

OAI21x1_ASAP7_75t_L g1192 ( 
.A1(n_984),
.A2(n_842),
.B(n_838),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1120),
.B(n_918),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1024),
.Y(n_1194)
);

NOR2xp33_ASAP7_75t_SL g1195 ( 
.A(n_1156),
.B(n_1099),
.Y(n_1195)
);

OR2x6_ASAP7_75t_L g1196 ( 
.A(n_1043),
.B(n_975),
.Y(n_1196)
);

OAI22xp5_ASAP7_75t_L g1197 ( 
.A1(n_1147),
.A2(n_969),
.B1(n_941),
.B2(n_970),
.Y(n_1197)
);

OAI21xp33_ASAP7_75t_L g1198 ( 
.A1(n_994),
.A2(n_970),
.B(n_960),
.Y(n_1198)
);

INVx5_ASAP7_75t_L g1199 ( 
.A(n_991),
.Y(n_1199)
);

NOR2xp33_ASAP7_75t_L g1200 ( 
.A(n_990),
.B(n_958),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1006),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1046),
.A2(n_958),
.B(n_960),
.Y(n_1202)
);

NOR2xp33_ASAP7_75t_L g1203 ( 
.A(n_1052),
.B(n_931),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1047),
.A2(n_971),
.B(n_954),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1047),
.A2(n_954),
.B(n_937),
.Y(n_1205)
);

INVx4_ASAP7_75t_L g1206 ( 
.A(n_992),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1057),
.B(n_839),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1007),
.Y(n_1208)
);

NOR2xp33_ASAP7_75t_L g1209 ( 
.A(n_1000),
.B(n_842),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_SL g1210 ( 
.A(n_997),
.B(n_987),
.Y(n_1210)
);

NOR2xp33_ASAP7_75t_L g1211 ( 
.A(n_1013),
.B(n_845),
.Y(n_1211)
);

OAI22xp5_ASAP7_75t_L g1212 ( 
.A1(n_1123),
.A2(n_936),
.B1(n_864),
.B2(n_978),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1009),
.Y(n_1213)
);

A2O1A1Ixp33_ASAP7_75t_SL g1214 ( 
.A1(n_993),
.A2(n_1159),
.B(n_1118),
.C(n_1126),
.Y(n_1214)
);

NOR3xp33_ASAP7_75t_SL g1215 ( 
.A(n_1005),
.B(n_13),
.C(n_15),
.Y(n_1215)
);

NAND3xp33_ASAP7_75t_L g1216 ( 
.A(n_1150),
.B(n_845),
.C(n_423),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_1026),
.Y(n_1217)
);

NOR2xp33_ASAP7_75t_L g1218 ( 
.A(n_1125),
.B(n_918),
.Y(n_1218)
);

BUFx2_ASAP7_75t_L g1219 ( 
.A(n_999),
.Y(n_1219)
);

OAI22xp33_ASAP7_75t_L g1220 ( 
.A1(n_985),
.A2(n_918),
.B1(n_423),
.B2(n_23),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_1042),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_SL g1222 ( 
.A(n_992),
.B(n_918),
.Y(n_1222)
);

BUFx6f_ASAP7_75t_L g1223 ( 
.A(n_1008),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1048),
.A2(n_423),
.B(n_172),
.Y(n_1224)
);

BUFx6f_ASAP7_75t_L g1225 ( 
.A(n_1008),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1048),
.A2(n_423),
.B(n_181),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1132),
.B(n_227),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1030),
.A2(n_168),
.B(n_106),
.Y(n_1228)
);

NOR2xp33_ASAP7_75t_L g1229 ( 
.A(n_988),
.B(n_15),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1121),
.B(n_21),
.Y(n_1230)
);

NOR2xp33_ASAP7_75t_SL g1231 ( 
.A(n_1099),
.B(n_309),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_SL g1232 ( 
.A(n_1054),
.B(n_309),
.Y(n_1232)
);

A2O1A1Ixp33_ASAP7_75t_L g1233 ( 
.A1(n_1080),
.A2(n_309),
.B(n_268),
.C(n_227),
.Y(n_1233)
);

NAND3xp33_ASAP7_75t_L g1234 ( 
.A(n_1148),
.B(n_21),
.C(n_27),
.Y(n_1234)
);

INVx3_ASAP7_75t_L g1235 ( 
.A(n_1008),
.Y(n_1235)
);

OAI22xp5_ASAP7_75t_L g1236 ( 
.A1(n_1130),
.A2(n_28),
.B1(n_30),
.B2(n_31),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1030),
.B(n_309),
.Y(n_1237)
);

INVx2_ASAP7_75t_SL g1238 ( 
.A(n_1054),
.Y(n_1238)
);

O2A1O1Ixp33_ASAP7_75t_SL g1239 ( 
.A1(n_1036),
.A2(n_30),
.B(n_31),
.C(n_32),
.Y(n_1239)
);

O2A1O1Ixp5_ASAP7_75t_L g1240 ( 
.A1(n_1122),
.A2(n_32),
.B(n_33),
.C(n_34),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1032),
.A2(n_182),
.B(n_108),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1032),
.A2(n_196),
.B(n_129),
.Y(n_1242)
);

INVx2_ASAP7_75t_L g1243 ( 
.A(n_1073),
.Y(n_1243)
);

NOR2xp33_ASAP7_75t_SL g1244 ( 
.A(n_1138),
.B(n_309),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1053),
.Y(n_1245)
);

HB1xp67_ASAP7_75t_L g1246 ( 
.A(n_1160),
.Y(n_1246)
);

NOR2xp33_ASAP7_75t_L g1247 ( 
.A(n_1079),
.B(n_33),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1084),
.Y(n_1248)
);

AND2x2_ASAP7_75t_L g1249 ( 
.A(n_1100),
.B(n_1124),
.Y(n_1249)
);

BUFx4f_ASAP7_75t_L g1250 ( 
.A(n_1168),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_SL g1251 ( 
.A(n_1043),
.B(n_309),
.Y(n_1251)
);

NOR2xp33_ASAP7_75t_L g1252 ( 
.A(n_1016),
.B(n_1131),
.Y(n_1252)
);

INVxp67_ASAP7_75t_L g1253 ( 
.A(n_1012),
.Y(n_1253)
);

A2O1A1Ixp33_ASAP7_75t_L g1254 ( 
.A1(n_1017),
.A2(n_309),
.B(n_268),
.C(n_227),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1090),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1129),
.B(n_1127),
.Y(n_1256)
);

AOI21x1_ASAP7_75t_L g1257 ( 
.A1(n_1078),
.A2(n_309),
.B(n_268),
.Y(n_1257)
);

AOI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1044),
.A2(n_166),
.B(n_132),
.Y(n_1258)
);

INVx3_ASAP7_75t_SL g1259 ( 
.A(n_1058),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1103),
.Y(n_1260)
);

NOR2xp33_ASAP7_75t_SL g1261 ( 
.A(n_1085),
.B(n_268),
.Y(n_1261)
);

O2A1O1Ixp5_ASAP7_75t_SL g1262 ( 
.A1(n_1166),
.A2(n_268),
.B(n_227),
.C(n_44),
.Y(n_1262)
);

INVx2_ASAP7_75t_L g1263 ( 
.A(n_1110),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1172),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1129),
.B(n_41),
.Y(n_1265)
);

AND2x2_ASAP7_75t_SL g1266 ( 
.A(n_1160),
.B(n_41),
.Y(n_1266)
);

AOI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_1028),
.A2(n_199),
.B(n_133),
.Y(n_1267)
);

BUFx6f_ASAP7_75t_L g1268 ( 
.A(n_1010),
.Y(n_1268)
);

OAI22xp5_ASAP7_75t_L g1269 ( 
.A1(n_1002),
.A2(n_43),
.B1(n_45),
.B2(n_46),
.Y(n_1269)
);

INVx5_ASAP7_75t_L g1270 ( 
.A(n_1010),
.Y(n_1270)
);

NAND2xp33_ASAP7_75t_SL g1271 ( 
.A(n_1010),
.B(n_45),
.Y(n_1271)
);

AOI22xp33_ASAP7_75t_L g1272 ( 
.A1(n_1152),
.A2(n_268),
.B1(n_227),
.B2(n_49),
.Y(n_1272)
);

HB1xp67_ASAP7_75t_L g1273 ( 
.A(n_1111),
.Y(n_1273)
);

NAND3xp33_ASAP7_75t_SL g1274 ( 
.A(n_1139),
.B(n_46),
.C(n_48),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1002),
.B(n_268),
.Y(n_1275)
);

OAI22xp5_ASAP7_75t_L g1276 ( 
.A1(n_1092),
.A2(n_48),
.B1(n_50),
.B2(n_52),
.Y(n_1276)
);

O2A1O1Ixp33_ASAP7_75t_L g1277 ( 
.A1(n_1119),
.A2(n_54),
.B(n_55),
.C(n_56),
.Y(n_1277)
);

INVx3_ASAP7_75t_SL g1278 ( 
.A(n_1162),
.Y(n_1278)
);

OAI22xp33_ASAP7_75t_L g1279 ( 
.A1(n_1146),
.A2(n_55),
.B1(n_57),
.B2(n_59),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_996),
.B(n_268),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_996),
.B(n_268),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_1174),
.Y(n_1282)
);

O2A1O1Ixp33_ASAP7_75t_L g1283 ( 
.A1(n_1094),
.A2(n_63),
.B(n_66),
.C(n_67),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1134),
.Y(n_1284)
);

O2A1O1Ixp33_ASAP7_75t_L g1285 ( 
.A1(n_1096),
.A2(n_69),
.B(n_70),
.C(n_71),
.Y(n_1285)
);

BUFx2_ASAP7_75t_L g1286 ( 
.A(n_1111),
.Y(n_1286)
);

AOI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1056),
.A2(n_147),
.B(n_220),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1165),
.B(n_1137),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1102),
.B(n_70),
.Y(n_1289)
);

BUFx2_ASAP7_75t_L g1290 ( 
.A(n_1023),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1023),
.B(n_72),
.Y(n_1291)
);

BUFx6f_ASAP7_75t_L g1292 ( 
.A(n_1018),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_SL g1293 ( 
.A(n_1145),
.B(n_227),
.Y(n_1293)
);

BUFx6f_ASAP7_75t_L g1294 ( 
.A(n_1018),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_1174),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1050),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1050),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_1068),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1091),
.B(n_75),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_1068),
.Y(n_1300)
);

NOR2xp33_ASAP7_75t_L g1301 ( 
.A(n_1098),
.B(n_75),
.Y(n_1301)
);

AOI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1128),
.A2(n_148),
.B(n_214),
.Y(n_1302)
);

OAI21xp33_ASAP7_75t_L g1303 ( 
.A1(n_1167),
.A2(n_76),
.B(n_77),
.Y(n_1303)
);

AOI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_986),
.A2(n_1060),
.B(n_1061),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1101),
.B(n_77),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1164),
.Y(n_1306)
);

AOI21xp5_ASAP7_75t_L g1307 ( 
.A1(n_986),
.A2(n_153),
.B(n_208),
.Y(n_1307)
);

NOR2xp33_ASAP7_75t_R g1308 ( 
.A(n_1018),
.B(n_145),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1086),
.B(n_79),
.Y(n_1309)
);

CKINVDCx20_ASAP7_75t_R g1310 ( 
.A(n_1027),
.Y(n_1310)
);

AOI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_1064),
.A2(n_155),
.B(n_206),
.Y(n_1311)
);

NOR2xp33_ASAP7_75t_L g1312 ( 
.A(n_1170),
.B(n_79),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_1164),
.Y(n_1313)
);

OAI22xp5_ASAP7_75t_L g1314 ( 
.A1(n_1070),
.A2(n_80),
.B1(n_81),
.B2(n_82),
.Y(n_1314)
);

OAI22xp5_ASAP7_75t_L g1315 ( 
.A1(n_1037),
.A2(n_1015),
.B1(n_1014),
.B2(n_1067),
.Y(n_1315)
);

AOI21xp5_ASAP7_75t_L g1316 ( 
.A1(n_1066),
.A2(n_90),
.B(n_161),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1029),
.Y(n_1317)
);

AOI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1074),
.A2(n_201),
.B(n_204),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1051),
.B(n_80),
.Y(n_1319)
);

NOR2xp33_ASAP7_75t_L g1320 ( 
.A(n_1135),
.B(n_84),
.Y(n_1320)
);

NOR2xp33_ASAP7_75t_L g1321 ( 
.A(n_1072),
.B(n_84),
.Y(n_1321)
);

AOI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_989),
.A2(n_216),
.B(n_1087),
.Y(n_1322)
);

INVx2_ASAP7_75t_SL g1323 ( 
.A(n_1027),
.Y(n_1323)
);

OAI22xp5_ASAP7_75t_L g1324 ( 
.A1(n_1025),
.A2(n_1109),
.B1(n_1113),
.B2(n_1107),
.Y(n_1324)
);

A2O1A1Ixp33_ASAP7_75t_L g1325 ( 
.A1(n_1077),
.A2(n_1049),
.B(n_1022),
.C(n_1115),
.Y(n_1325)
);

OAI22xp5_ASAP7_75t_L g1326 ( 
.A1(n_1107),
.A2(n_1109),
.B1(n_1113),
.B2(n_1071),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_1027),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_SL g1328 ( 
.A(n_1155),
.B(n_1038),
.Y(n_1328)
);

OAI22xp5_ASAP7_75t_L g1329 ( 
.A1(n_1055),
.A2(n_1175),
.B1(n_1088),
.B2(n_1095),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1063),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1033),
.Y(n_1331)
);

NOR2xp33_ASAP7_75t_R g1332 ( 
.A(n_1038),
.B(n_1097),
.Y(n_1332)
);

AO32x1_ASAP7_75t_L g1333 ( 
.A1(n_1059),
.A2(n_1040),
.A3(n_1081),
.B1(n_1065),
.B2(n_1021),
.Y(n_1333)
);

O2A1O1Ixp33_ASAP7_75t_L g1334 ( 
.A1(n_1076),
.A2(n_1154),
.B(n_1153),
.C(n_1151),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1069),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1163),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1149),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1149),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1097),
.B(n_1112),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1112),
.B(n_1106),
.Y(n_1340)
);

AOI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1093),
.A2(n_1105),
.B(n_1001),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1082),
.Y(n_1342)
);

INVx2_ASAP7_75t_SL g1343 ( 
.A(n_1031),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1256),
.B(n_1086),
.Y(n_1344)
);

AND2x4_ASAP7_75t_L g1345 ( 
.A(n_1206),
.B(n_1310),
.Y(n_1345)
);

OAI21x1_ASAP7_75t_SL g1346 ( 
.A1(n_1340),
.A2(n_1075),
.B(n_1011),
.Y(n_1346)
);

BUFx10_ASAP7_75t_L g1347 ( 
.A(n_1312),
.Y(n_1347)
);

INVxp67_ASAP7_75t_L g1348 ( 
.A(n_1203),
.Y(n_1348)
);

AOI22xp5_ASAP7_75t_L g1349 ( 
.A1(n_1266),
.A2(n_1106),
.B1(n_1095),
.B2(n_1088),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1249),
.B(n_1136),
.Y(n_1350)
);

OAI22xp5_ASAP7_75t_L g1351 ( 
.A1(n_1230),
.A2(n_1256),
.B1(n_1236),
.B2(n_1265),
.Y(n_1351)
);

NAND2xp33_ASAP7_75t_SL g1352 ( 
.A(n_1206),
.B(n_1083),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1190),
.Y(n_1353)
);

OAI21x1_ASAP7_75t_L g1354 ( 
.A1(n_1257),
.A2(n_1176),
.B(n_1020),
.Y(n_1354)
);

AOI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1324),
.A2(n_1003),
.B(n_1144),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1286),
.B(n_1031),
.Y(n_1356)
);

OAI21x1_ASAP7_75t_L g1357 ( 
.A1(n_1304),
.A2(n_1034),
.B(n_1041),
.Y(n_1357)
);

NAND3xp33_ASAP7_75t_L g1358 ( 
.A(n_1236),
.B(n_1173),
.C(n_1171),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1184),
.Y(n_1359)
);

AOI22xp33_ASAP7_75t_L g1360 ( 
.A1(n_1210),
.A2(n_1082),
.B1(n_1083),
.B2(n_1142),
.Y(n_1360)
);

OAI21x1_ASAP7_75t_L g1361 ( 
.A1(n_1341),
.A2(n_1114),
.B(n_1062),
.Y(n_1361)
);

AOI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1324),
.A2(n_1035),
.B(n_1045),
.Y(n_1362)
);

OAI22xp5_ASAP7_75t_SL g1363 ( 
.A1(n_1288),
.A2(n_1143),
.B1(n_1141),
.B2(n_1140),
.Y(n_1363)
);

NOR2xp33_ASAP7_75t_L g1364 ( 
.A(n_1252),
.B(n_1157),
.Y(n_1364)
);

AO31x2_ASAP7_75t_L g1365 ( 
.A1(n_1330),
.A2(n_1158),
.A3(n_1161),
.B(n_1169),
.Y(n_1365)
);

OR2x2_ASAP7_75t_L g1366 ( 
.A(n_1273),
.B(n_1117),
.Y(n_1366)
);

AO31x2_ASAP7_75t_L g1367 ( 
.A1(n_1233),
.A2(n_1331),
.A3(n_1315),
.B(n_1325),
.Y(n_1367)
);

O2A1O1Ixp33_ASAP7_75t_SL g1368 ( 
.A1(n_1214),
.A2(n_1116),
.B(n_1309),
.C(n_1222),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1296),
.B(n_1297),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1185),
.B(n_1282),
.Y(n_1370)
);

OAI21xp5_ASAP7_75t_L g1371 ( 
.A1(n_1329),
.A2(n_1202),
.B(n_1189),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1201),
.Y(n_1372)
);

OAI21x1_ASAP7_75t_L g1373 ( 
.A1(n_1192),
.A2(n_1322),
.B(n_1181),
.Y(n_1373)
);

AOI21x1_ASAP7_75t_L g1374 ( 
.A1(n_1329),
.A2(n_1336),
.B(n_1237),
.Y(n_1374)
);

OAI21xp5_ASAP7_75t_L g1375 ( 
.A1(n_1309),
.A2(n_1326),
.B(n_1315),
.Y(n_1375)
);

AOI31xp67_ASAP7_75t_L g1376 ( 
.A1(n_1237),
.A2(n_1275),
.A3(n_1281),
.B(n_1280),
.Y(n_1376)
);

AOI221xp5_ASAP7_75t_SL g1377 ( 
.A1(n_1279),
.A2(n_1276),
.B1(n_1283),
.B2(n_1285),
.C(n_1269),
.Y(n_1377)
);

NAND2x1p5_ASAP7_75t_L g1378 ( 
.A(n_1199),
.B(n_1270),
.Y(n_1378)
);

BUFx3_ASAP7_75t_L g1379 ( 
.A(n_1259),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1208),
.Y(n_1380)
);

AO31x2_ASAP7_75t_L g1381 ( 
.A1(n_1212),
.A2(n_1335),
.A3(n_1326),
.B(n_1204),
.Y(n_1381)
);

OAI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1178),
.A2(n_1188),
.B(n_1205),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1209),
.B(n_1284),
.Y(n_1383)
);

AOI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1188),
.A2(n_1333),
.B(n_1258),
.Y(n_1384)
);

AOI21xp5_ASAP7_75t_L g1385 ( 
.A1(n_1333),
.A2(n_1334),
.B(n_1342),
.Y(n_1385)
);

AOI21x1_ASAP7_75t_L g1386 ( 
.A1(n_1275),
.A2(n_1280),
.B(n_1281),
.Y(n_1386)
);

NAND2x1_ASAP7_75t_L g1387 ( 
.A(n_1235),
.B(n_1187),
.Y(n_1387)
);

O2A1O1Ixp33_ASAP7_75t_SL g1388 ( 
.A1(n_1328),
.A2(n_1291),
.B(n_1320),
.C(n_1289),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1211),
.B(n_1246),
.Y(n_1389)
);

AOI222xp33_ASAP7_75t_L g1390 ( 
.A1(n_1276),
.A2(n_1220),
.B1(n_1274),
.B2(n_1247),
.C1(n_1269),
.C2(n_1197),
.Y(n_1390)
);

BUFx2_ASAP7_75t_L g1391 ( 
.A(n_1327),
.Y(n_1391)
);

NOR2x1_ASAP7_75t_SL g1392 ( 
.A(n_1199),
.B(n_1270),
.Y(n_1392)
);

AOI21xp5_ASAP7_75t_L g1393 ( 
.A1(n_1333),
.A2(n_1226),
.B(n_1224),
.Y(n_1393)
);

NAND3x1_ASAP7_75t_L g1394 ( 
.A(n_1301),
.B(n_1229),
.C(n_1321),
.Y(n_1394)
);

AOI21xp5_ASAP7_75t_L g1395 ( 
.A1(n_1193),
.A2(n_1186),
.B(n_1191),
.Y(n_1395)
);

BUFx3_ASAP7_75t_L g1396 ( 
.A(n_1250),
.Y(n_1396)
);

AOI21xp5_ASAP7_75t_L g1397 ( 
.A1(n_1193),
.A2(n_1287),
.B(n_1267),
.Y(n_1397)
);

A2O1A1Ixp33_ASAP7_75t_L g1398 ( 
.A1(n_1303),
.A2(n_1182),
.B(n_1218),
.C(n_1200),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1213),
.B(n_1245),
.Y(n_1399)
);

OAI21xp5_ASAP7_75t_L g1400 ( 
.A1(n_1262),
.A2(n_1254),
.B(n_1197),
.Y(n_1400)
);

AND2x6_ASAP7_75t_L g1401 ( 
.A(n_1337),
.B(n_1338),
.Y(n_1401)
);

OA21x2_ASAP7_75t_L g1402 ( 
.A1(n_1227),
.A2(n_1216),
.B(n_1302),
.Y(n_1402)
);

OAI21x1_ASAP7_75t_L g1403 ( 
.A1(n_1311),
.A2(n_1316),
.B(n_1318),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1248),
.Y(n_1404)
);

AND2x4_ASAP7_75t_L g1405 ( 
.A(n_1196),
.B(n_1238),
.Y(n_1405)
);

OAI21x1_ASAP7_75t_L g1406 ( 
.A1(n_1227),
.A2(n_1242),
.B(n_1228),
.Y(n_1406)
);

OA21x2_ASAP7_75t_L g1407 ( 
.A1(n_1198),
.A2(n_1313),
.B(n_1306),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1278),
.B(n_1177),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1295),
.B(n_1298),
.Y(n_1409)
);

OAI22xp5_ASAP7_75t_L g1410 ( 
.A1(n_1319),
.A2(n_1215),
.B1(n_1234),
.B2(n_1255),
.Y(n_1410)
);

AOI21xp5_ASAP7_75t_L g1411 ( 
.A1(n_1241),
.A2(n_1307),
.B(n_1180),
.Y(n_1411)
);

A2O1A1Ixp33_ASAP7_75t_L g1412 ( 
.A1(n_1277),
.A2(n_1305),
.B(n_1272),
.C(n_1299),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1300),
.B(n_1207),
.Y(n_1413)
);

OAI21x1_ASAP7_75t_L g1414 ( 
.A1(n_1339),
.A2(n_1212),
.B(n_1183),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1196),
.B(n_1264),
.Y(n_1415)
);

OAI21x1_ASAP7_75t_L g1416 ( 
.A1(n_1317),
.A2(n_1235),
.B(n_1240),
.Y(n_1416)
);

AOI21xp5_ASAP7_75t_L g1417 ( 
.A1(n_1271),
.A2(n_1239),
.B(n_1270),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_SL g1418 ( 
.A(n_1199),
.B(n_1270),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1194),
.Y(n_1419)
);

OAI21x1_ASAP7_75t_L g1420 ( 
.A1(n_1251),
.A2(n_1232),
.B(n_1293),
.Y(n_1420)
);

CKINVDCx9p33_ASAP7_75t_R g1421 ( 
.A(n_1219),
.Y(n_1421)
);

AOI221x1_ASAP7_75t_L g1422 ( 
.A1(n_1314),
.A2(n_1243),
.B1(n_1260),
.B2(n_1263),
.C(n_1221),
.Y(n_1422)
);

O2A1O1Ixp33_ASAP7_75t_L g1423 ( 
.A1(n_1314),
.A2(n_1290),
.B(n_1253),
.C(n_1261),
.Y(n_1423)
);

BUFx3_ASAP7_75t_L g1424 ( 
.A(n_1250),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1196),
.B(n_1217),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1177),
.Y(n_1426)
);

O2A1O1Ixp33_ASAP7_75t_L g1427 ( 
.A1(n_1244),
.A2(n_1231),
.B(n_1179),
.C(n_1195),
.Y(n_1427)
);

NOR2xp67_ASAP7_75t_SL g1428 ( 
.A(n_1199),
.B(n_1187),
.Y(n_1428)
);

OAI21x1_ASAP7_75t_L g1429 ( 
.A1(n_1343),
.A2(n_1187),
.B(n_1223),
.Y(n_1429)
);

OA21x2_ASAP7_75t_L g1430 ( 
.A1(n_1323),
.A2(n_1308),
.B(n_1225),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1223),
.B(n_1225),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1223),
.Y(n_1432)
);

AOI21xp5_ASAP7_75t_L g1433 ( 
.A1(n_1225),
.A2(n_1268),
.B(n_1292),
.Y(n_1433)
);

BUFx2_ASAP7_75t_L g1434 ( 
.A(n_1332),
.Y(n_1434)
);

AO31x2_ASAP7_75t_L g1435 ( 
.A1(n_1268),
.A2(n_1330),
.A3(n_1233),
.B(n_1331),
.Y(n_1435)
);

NOR2xp33_ASAP7_75t_L g1436 ( 
.A(n_1294),
.B(n_1268),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1292),
.B(n_1294),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1292),
.B(n_1294),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1256),
.B(n_1296),
.Y(n_1439)
);

AOI21xp5_ASAP7_75t_L g1440 ( 
.A1(n_1324),
.A2(n_1326),
.B(n_1188),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1249),
.B(n_1133),
.Y(n_1441)
);

OAI21x1_ASAP7_75t_L g1442 ( 
.A1(n_1257),
.A2(n_1304),
.B(n_1341),
.Y(n_1442)
);

O2A1O1Ixp5_ASAP7_75t_L g1443 ( 
.A1(n_1230),
.A2(n_860),
.B(n_1089),
.C(n_990),
.Y(n_1443)
);

AOI22xp5_ASAP7_75t_L g1444 ( 
.A1(n_1266),
.A2(n_983),
.B1(n_1133),
.B2(n_713),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1256),
.B(n_1296),
.Y(n_1445)
);

AND2x4_ASAP7_75t_L g1446 ( 
.A(n_1206),
.B(n_1019),
.Y(n_1446)
);

AOI21xp5_ASAP7_75t_L g1447 ( 
.A1(n_1324),
.A2(n_1326),
.B(n_1188),
.Y(n_1447)
);

AOI221x1_ASAP7_75t_L g1448 ( 
.A1(n_1236),
.A2(n_1303),
.B1(n_1080),
.B2(n_1269),
.C(n_1089),
.Y(n_1448)
);

AOI21xp5_ASAP7_75t_L g1449 ( 
.A1(n_1324),
.A2(n_1326),
.B(n_1188),
.Y(n_1449)
);

AOI21xp5_ASAP7_75t_L g1450 ( 
.A1(n_1324),
.A2(n_1326),
.B(n_1188),
.Y(n_1450)
);

OAI21x1_ASAP7_75t_L g1451 ( 
.A1(n_1257),
.A2(n_1304),
.B(n_1341),
.Y(n_1451)
);

NAND3xp33_ASAP7_75t_SL g1452 ( 
.A(n_1230),
.B(n_674),
.C(n_592),
.Y(n_1452)
);

OA21x2_ASAP7_75t_L g1453 ( 
.A1(n_1304),
.A2(n_1257),
.B(n_1341),
.Y(n_1453)
);

OAI21xp5_ASAP7_75t_L g1454 ( 
.A1(n_1329),
.A2(n_1202),
.B(n_1189),
.Y(n_1454)
);

AOI21xp5_ASAP7_75t_L g1455 ( 
.A1(n_1324),
.A2(n_1326),
.B(n_1188),
.Y(n_1455)
);

O2A1O1Ixp5_ASAP7_75t_SL g1456 ( 
.A1(n_1236),
.A2(n_1080),
.B(n_1331),
.C(n_1269),
.Y(n_1456)
);

BUFx4f_ASAP7_75t_SL g1457 ( 
.A(n_1259),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1256),
.B(n_1296),
.Y(n_1458)
);

AOI21xp5_ASAP7_75t_L g1459 ( 
.A1(n_1324),
.A2(n_1326),
.B(n_1188),
.Y(n_1459)
);

AO31x2_ASAP7_75t_L g1460 ( 
.A1(n_1330),
.A2(n_1233),
.A3(n_1331),
.B(n_1315),
.Y(n_1460)
);

OA21x2_ASAP7_75t_L g1461 ( 
.A1(n_1304),
.A2(n_1257),
.B(n_1341),
.Y(n_1461)
);

AOI21xp5_ASAP7_75t_L g1462 ( 
.A1(n_1324),
.A2(n_1326),
.B(n_1188),
.Y(n_1462)
);

A2O1A1Ixp33_ASAP7_75t_L g1463 ( 
.A1(n_1320),
.A2(n_1230),
.B(n_1089),
.C(n_860),
.Y(n_1463)
);

INVx3_ASAP7_75t_SL g1464 ( 
.A(n_1259),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1256),
.B(n_1296),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1201),
.Y(n_1466)
);

AOI21xp5_ASAP7_75t_L g1467 ( 
.A1(n_1324),
.A2(n_1326),
.B(n_1188),
.Y(n_1467)
);

AO31x2_ASAP7_75t_L g1468 ( 
.A1(n_1330),
.A2(n_1233),
.A3(n_1331),
.B(n_1315),
.Y(n_1468)
);

CKINVDCx20_ASAP7_75t_R g1469 ( 
.A(n_1259),
.Y(n_1469)
);

AND2x4_ASAP7_75t_L g1470 ( 
.A(n_1206),
.B(n_1019),
.Y(n_1470)
);

OAI21xp5_ASAP7_75t_SL g1471 ( 
.A1(n_1236),
.A2(n_860),
.B(n_900),
.Y(n_1471)
);

INVx4_ASAP7_75t_L g1472 ( 
.A(n_1259),
.Y(n_1472)
);

CKINVDCx16_ASAP7_75t_R g1473 ( 
.A(n_1310),
.Y(n_1473)
);

OA21x2_ASAP7_75t_L g1474 ( 
.A1(n_1304),
.A2(n_1257),
.B(n_1341),
.Y(n_1474)
);

BUFx8_ASAP7_75t_L g1475 ( 
.A(n_1219),
.Y(n_1475)
);

OAI21x1_ASAP7_75t_L g1476 ( 
.A1(n_1257),
.A2(n_1304),
.B(n_1341),
.Y(n_1476)
);

AOI22xp33_ASAP7_75t_L g1477 ( 
.A1(n_1266),
.A2(n_900),
.B1(n_967),
.B2(n_631),
.Y(n_1477)
);

BUFx10_ASAP7_75t_L g1478 ( 
.A(n_1312),
.Y(n_1478)
);

BUFx2_ASAP7_75t_L g1479 ( 
.A(n_1310),
.Y(n_1479)
);

INVx1_ASAP7_75t_SL g1480 ( 
.A(n_1286),
.Y(n_1480)
);

AO21x2_ASAP7_75t_L g1481 ( 
.A1(n_1257),
.A2(n_1078),
.B(n_1331),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1190),
.Y(n_1482)
);

A2O1A1Ixp33_ASAP7_75t_L g1483 ( 
.A1(n_1320),
.A2(n_1230),
.B(n_1089),
.C(n_860),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1249),
.B(n_1133),
.Y(n_1484)
);

OAI21xp5_ASAP7_75t_L g1485 ( 
.A1(n_1329),
.A2(n_1202),
.B(n_1189),
.Y(n_1485)
);

A2O1A1Ixp33_ASAP7_75t_L g1486 ( 
.A1(n_1320),
.A2(n_1230),
.B(n_1089),
.C(n_860),
.Y(n_1486)
);

AOI21xp5_ASAP7_75t_L g1487 ( 
.A1(n_1324),
.A2(n_1326),
.B(n_1188),
.Y(n_1487)
);

AOI21xp5_ASAP7_75t_L g1488 ( 
.A1(n_1324),
.A2(n_1326),
.B(n_1188),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1249),
.B(n_1133),
.Y(n_1489)
);

OAI21x1_ASAP7_75t_L g1490 ( 
.A1(n_1257),
.A2(n_1304),
.B(n_1341),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1201),
.Y(n_1491)
);

INVx5_ASAP7_75t_L g1492 ( 
.A(n_1206),
.Y(n_1492)
);

NOR2xp33_ASAP7_75t_L g1493 ( 
.A(n_1288),
.B(n_983),
.Y(n_1493)
);

AOI21xp5_ASAP7_75t_L g1494 ( 
.A1(n_1324),
.A2(n_1326),
.B(n_1188),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1249),
.B(n_1133),
.Y(n_1495)
);

NOR2xp33_ASAP7_75t_SL g1496 ( 
.A(n_1266),
.B(n_1179),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_SL g1497 ( 
.A(n_1256),
.B(n_713),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1249),
.B(n_1133),
.Y(n_1498)
);

A2O1A1Ixp33_ASAP7_75t_L g1499 ( 
.A1(n_1320),
.A2(n_1230),
.B(n_1089),
.C(n_860),
.Y(n_1499)
);

A2O1A1Ixp33_ASAP7_75t_L g1500 ( 
.A1(n_1320),
.A2(n_1230),
.B(n_1089),
.C(n_860),
.Y(n_1500)
);

OAI21x1_ASAP7_75t_L g1501 ( 
.A1(n_1257),
.A2(n_1304),
.B(n_1341),
.Y(n_1501)
);

OAI21xp5_ASAP7_75t_L g1502 ( 
.A1(n_1329),
.A2(n_1202),
.B(n_1189),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1201),
.Y(n_1503)
);

AND2x6_ASAP7_75t_L g1504 ( 
.A(n_1182),
.B(n_1147),
.Y(n_1504)
);

CKINVDCx5p33_ASAP7_75t_R g1505 ( 
.A(n_1259),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1249),
.B(n_1133),
.Y(n_1506)
);

AO32x2_ASAP7_75t_L g1507 ( 
.A1(n_1236),
.A2(n_1269),
.A3(n_1329),
.B1(n_1197),
.B2(n_1276),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1249),
.B(n_1133),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1201),
.Y(n_1509)
);

AOI21xp5_ASAP7_75t_L g1510 ( 
.A1(n_1324),
.A2(n_1326),
.B(n_1188),
.Y(n_1510)
);

OAI21xp5_ASAP7_75t_L g1511 ( 
.A1(n_1329),
.A2(n_1202),
.B(n_1189),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1201),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1249),
.B(n_1133),
.Y(n_1513)
);

AOI21xp5_ASAP7_75t_L g1514 ( 
.A1(n_1324),
.A2(n_1326),
.B(n_1188),
.Y(n_1514)
);

CKINVDCx5p33_ASAP7_75t_R g1515 ( 
.A(n_1259),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1190),
.Y(n_1516)
);

AO31x2_ASAP7_75t_L g1517 ( 
.A1(n_1330),
.A2(n_1233),
.A3(n_1331),
.B(n_1315),
.Y(n_1517)
);

AOI21xp5_ASAP7_75t_L g1518 ( 
.A1(n_1324),
.A2(n_1326),
.B(n_1188),
.Y(n_1518)
);

AO31x2_ASAP7_75t_L g1519 ( 
.A1(n_1330),
.A2(n_1233),
.A3(n_1331),
.B(n_1315),
.Y(n_1519)
);

OAI22xp33_ASAP7_75t_L g1520 ( 
.A1(n_1471),
.A2(n_1496),
.B1(n_1444),
.B2(n_1448),
.Y(n_1520)
);

AOI22xp33_ASAP7_75t_L g1521 ( 
.A1(n_1390),
.A2(n_1477),
.B1(n_1493),
.B2(n_1351),
.Y(n_1521)
);

OAI22x1_ASAP7_75t_SL g1522 ( 
.A1(n_1469),
.A2(n_1515),
.B1(n_1505),
.B2(n_1472),
.Y(n_1522)
);

OAI21xp5_ASAP7_75t_L g1523 ( 
.A1(n_1463),
.A2(n_1486),
.B(n_1483),
.Y(n_1523)
);

BUFx8_ASAP7_75t_SL g1524 ( 
.A(n_1479),
.Y(n_1524)
);

BUFx3_ASAP7_75t_L g1525 ( 
.A(n_1457),
.Y(n_1525)
);

OAI21xp33_ASAP7_75t_L g1526 ( 
.A1(n_1499),
.A2(n_1500),
.B(n_1471),
.Y(n_1526)
);

BUFx3_ASAP7_75t_L g1527 ( 
.A(n_1379),
.Y(n_1527)
);

CKINVDCx20_ASAP7_75t_R g1528 ( 
.A(n_1464),
.Y(n_1528)
);

AOI22xp33_ASAP7_75t_L g1529 ( 
.A1(n_1390),
.A2(n_1351),
.B1(n_1504),
.B2(n_1496),
.Y(n_1529)
);

INVx3_ASAP7_75t_L g1530 ( 
.A(n_1378),
.Y(n_1530)
);

BUFx4f_ASAP7_75t_SL g1531 ( 
.A(n_1396),
.Y(n_1531)
);

BUFx6f_ASAP7_75t_L g1532 ( 
.A(n_1378),
.Y(n_1532)
);

AOI22xp33_ASAP7_75t_SL g1533 ( 
.A1(n_1504),
.A2(n_1375),
.B1(n_1410),
.B2(n_1394),
.Y(n_1533)
);

CKINVDCx6p67_ASAP7_75t_R g1534 ( 
.A(n_1421),
.Y(n_1534)
);

INVx1_ASAP7_75t_SL g1535 ( 
.A(n_1408),
.Y(n_1535)
);

AOI22xp33_ASAP7_75t_L g1536 ( 
.A1(n_1504),
.A2(n_1375),
.B1(n_1498),
.B2(n_1441),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1399),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1372),
.Y(n_1538)
);

OAI22xp5_ASAP7_75t_L g1539 ( 
.A1(n_1349),
.A2(n_1364),
.B1(n_1489),
.B2(n_1495),
.Y(n_1539)
);

INVx3_ASAP7_75t_L g1540 ( 
.A(n_1492),
.Y(n_1540)
);

AOI22xp33_ASAP7_75t_L g1541 ( 
.A1(n_1504),
.A2(n_1506),
.B1(n_1484),
.B2(n_1508),
.Y(n_1541)
);

AOI22xp33_ASAP7_75t_L g1542 ( 
.A1(n_1513),
.A2(n_1410),
.B1(n_1350),
.B2(n_1497),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1380),
.Y(n_1543)
);

BUFx8_ASAP7_75t_L g1544 ( 
.A(n_1391),
.Y(n_1544)
);

OAI22xp33_ASAP7_75t_L g1545 ( 
.A1(n_1439),
.A2(n_1458),
.B1(n_1465),
.B2(n_1445),
.Y(n_1545)
);

AOI22xp33_ASAP7_75t_L g1546 ( 
.A1(n_1383),
.A2(n_1347),
.B1(n_1478),
.B2(n_1465),
.Y(n_1546)
);

AOI22xp5_ASAP7_75t_L g1547 ( 
.A1(n_1348),
.A2(n_1377),
.B1(n_1452),
.B2(n_1478),
.Y(n_1547)
);

AOI22xp33_ASAP7_75t_SL g1548 ( 
.A1(n_1507),
.A2(n_1347),
.B1(n_1400),
.B2(n_1439),
.Y(n_1548)
);

BUFx8_ASAP7_75t_SL g1549 ( 
.A(n_1424),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1480),
.B(n_1473),
.Y(n_1550)
);

AOI22xp33_ASAP7_75t_L g1551 ( 
.A1(n_1445),
.A2(n_1458),
.B1(n_1344),
.B2(n_1389),
.Y(n_1551)
);

CKINVDCx6p67_ASAP7_75t_R g1552 ( 
.A(n_1472),
.Y(n_1552)
);

NAND2x1p5_ASAP7_75t_L g1553 ( 
.A(n_1428),
.B(n_1430),
.Y(n_1553)
);

BUFx12f_ASAP7_75t_L g1554 ( 
.A(n_1475),
.Y(n_1554)
);

OAI21xp5_ASAP7_75t_L g1555 ( 
.A1(n_1443),
.A2(n_1456),
.B(n_1388),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1404),
.Y(n_1556)
);

BUFx6f_ASAP7_75t_L g1557 ( 
.A(n_1430),
.Y(n_1557)
);

OAI22xp5_ASAP7_75t_L g1558 ( 
.A1(n_1440),
.A2(n_1467),
.B1(n_1518),
.B2(n_1514),
.Y(n_1558)
);

OAI21xp33_ASAP7_75t_L g1559 ( 
.A1(n_1371),
.A2(n_1485),
.B(n_1502),
.Y(n_1559)
);

AOI22xp33_ASAP7_75t_L g1560 ( 
.A1(n_1359),
.A2(n_1482),
.B1(n_1516),
.B2(n_1419),
.Y(n_1560)
);

BUFx3_ASAP7_75t_L g1561 ( 
.A(n_1475),
.Y(n_1561)
);

AO22x1_ASAP7_75t_L g1562 ( 
.A1(n_1401),
.A2(n_1434),
.B1(n_1405),
.B2(n_1492),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1466),
.Y(n_1563)
);

CKINVDCx11_ASAP7_75t_R g1564 ( 
.A(n_1426),
.Y(n_1564)
);

AOI22xp33_ASAP7_75t_L g1565 ( 
.A1(n_1344),
.A2(n_1425),
.B1(n_1409),
.B2(n_1401),
.Y(n_1565)
);

OAI21xp5_ASAP7_75t_L g1566 ( 
.A1(n_1398),
.A2(n_1412),
.B(n_1362),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1491),
.Y(n_1567)
);

AOI22xp33_ASAP7_75t_L g1568 ( 
.A1(n_1369),
.A2(n_1413),
.B1(n_1512),
.B2(n_1503),
.Y(n_1568)
);

AOI22xp33_ASAP7_75t_L g1569 ( 
.A1(n_1425),
.A2(n_1409),
.B1(n_1401),
.B2(n_1413),
.Y(n_1569)
);

BUFx12f_ASAP7_75t_L g1570 ( 
.A(n_1492),
.Y(n_1570)
);

AOI22xp33_ASAP7_75t_SL g1571 ( 
.A1(n_1507),
.A2(n_1400),
.B1(n_1449),
.B2(n_1510),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1509),
.Y(n_1572)
);

AOI22xp33_ASAP7_75t_L g1573 ( 
.A1(n_1401),
.A2(n_1415),
.B1(n_1366),
.B2(n_1358),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1370),
.Y(n_1574)
);

AOI22xp33_ASAP7_75t_SL g1575 ( 
.A1(n_1507),
.A2(n_1447),
.B1(n_1462),
.B2(n_1455),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1370),
.Y(n_1576)
);

CKINVDCx5p33_ASAP7_75t_R g1577 ( 
.A(n_1436),
.Y(n_1577)
);

AOI22xp33_ASAP7_75t_L g1578 ( 
.A1(n_1415),
.A2(n_1358),
.B1(n_1363),
.B2(n_1407),
.Y(n_1578)
);

AOI22xp33_ASAP7_75t_SL g1579 ( 
.A1(n_1450),
.A2(n_1487),
.B1(n_1459),
.B2(n_1488),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1432),
.Y(n_1580)
);

BUFx6f_ASAP7_75t_L g1581 ( 
.A(n_1446),
.Y(n_1581)
);

INVx6_ASAP7_75t_L g1582 ( 
.A(n_1446),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1356),
.B(n_1470),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1431),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1431),
.Y(n_1585)
);

OAI21xp5_ASAP7_75t_SL g1586 ( 
.A1(n_1423),
.A2(n_1427),
.B(n_1494),
.Y(n_1586)
);

BUFx4f_ASAP7_75t_L g1587 ( 
.A(n_1470),
.Y(n_1587)
);

OAI21xp5_ASAP7_75t_SL g1588 ( 
.A1(n_1371),
.A2(n_1511),
.B(n_1502),
.Y(n_1588)
);

INVx5_ASAP7_75t_L g1589 ( 
.A(n_1392),
.Y(n_1589)
);

AOI22xp33_ASAP7_75t_L g1590 ( 
.A1(n_1360),
.A2(n_1414),
.B1(n_1352),
.B2(n_1417),
.Y(n_1590)
);

AOI22xp33_ASAP7_75t_SL g1591 ( 
.A1(n_1377),
.A2(n_1454),
.B1(n_1511),
.B2(n_1485),
.Y(n_1591)
);

OAI22xp5_ASAP7_75t_L g1592 ( 
.A1(n_1454),
.A2(n_1355),
.B1(n_1382),
.B2(n_1397),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1437),
.Y(n_1593)
);

BUFx8_ASAP7_75t_L g1594 ( 
.A(n_1387),
.Y(n_1594)
);

OAI22xp5_ASAP7_75t_L g1595 ( 
.A1(n_1382),
.A2(n_1384),
.B1(n_1385),
.B2(n_1393),
.Y(n_1595)
);

CKINVDCx11_ASAP7_75t_R g1596 ( 
.A(n_1438),
.Y(n_1596)
);

AOI22xp33_ASAP7_75t_L g1597 ( 
.A1(n_1402),
.A2(n_1346),
.B1(n_1481),
.B2(n_1420),
.Y(n_1597)
);

INVx1_ASAP7_75t_SL g1598 ( 
.A(n_1437),
.Y(n_1598)
);

BUFx10_ASAP7_75t_L g1599 ( 
.A(n_1433),
.Y(n_1599)
);

INVx6_ASAP7_75t_L g1600 ( 
.A(n_1418),
.Y(n_1600)
);

BUFx4f_ASAP7_75t_SL g1601 ( 
.A(n_1429),
.Y(n_1601)
);

OAI21xp5_ASAP7_75t_SL g1602 ( 
.A1(n_1422),
.A2(n_1411),
.B(n_1395),
.Y(n_1602)
);

INVx8_ASAP7_75t_L g1603 ( 
.A(n_1416),
.Y(n_1603)
);

BUFx8_ASAP7_75t_L g1604 ( 
.A(n_1368),
.Y(n_1604)
);

AOI22xp5_ASAP7_75t_L g1605 ( 
.A1(n_1402),
.A2(n_1481),
.B1(n_1406),
.B2(n_1403),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1435),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1374),
.Y(n_1607)
);

OAI21xp5_ASAP7_75t_SL g1608 ( 
.A1(n_1386),
.A2(n_1367),
.B(n_1381),
.Y(n_1608)
);

INVx6_ASAP7_75t_L g1609 ( 
.A(n_1435),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1435),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1460),
.Y(n_1611)
);

BUFx3_ASAP7_75t_L g1612 ( 
.A(n_1367),
.Y(n_1612)
);

CKINVDCx5p33_ASAP7_75t_R g1613 ( 
.A(n_1376),
.Y(n_1613)
);

AOI22xp33_ASAP7_75t_L g1614 ( 
.A1(n_1354),
.A2(n_1474),
.B1(n_1461),
.B2(n_1453),
.Y(n_1614)
);

AOI22x1_ASAP7_75t_SL g1615 ( 
.A1(n_1367),
.A2(n_1381),
.B1(n_1365),
.B2(n_1519),
.Y(n_1615)
);

OAI21xp33_ASAP7_75t_SL g1616 ( 
.A1(n_1361),
.A2(n_1357),
.B(n_1373),
.Y(n_1616)
);

OAI22xp5_ASAP7_75t_SL g1617 ( 
.A1(n_1453),
.A2(n_1474),
.B1(n_1461),
.B2(n_1381),
.Y(n_1617)
);

AOI22xp33_ASAP7_75t_L g1618 ( 
.A1(n_1442),
.A2(n_1490),
.B1(n_1451),
.B2(n_1501),
.Y(n_1618)
);

AOI22xp33_ASAP7_75t_SL g1619 ( 
.A1(n_1468),
.A2(n_1517),
.B1(n_1519),
.B2(n_1476),
.Y(n_1619)
);

BUFx6f_ASAP7_75t_L g1620 ( 
.A(n_1468),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1517),
.B(n_1519),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1517),
.B(n_1365),
.Y(n_1622)
);

BUFx2_ASAP7_75t_L g1623 ( 
.A(n_1345),
.Y(n_1623)
);

CKINVDCx11_ASAP7_75t_R g1624 ( 
.A(n_1469),
.Y(n_1624)
);

CKINVDCx5p33_ASAP7_75t_R g1625 ( 
.A(n_1505),
.Y(n_1625)
);

OAI22xp33_ASAP7_75t_SL g1626 ( 
.A1(n_1496),
.A2(n_1150),
.B1(n_1230),
.B2(n_1288),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1399),
.Y(n_1627)
);

NAND2x1p5_ASAP7_75t_L g1628 ( 
.A(n_1428),
.B(n_1430),
.Y(n_1628)
);

AOI22xp33_ASAP7_75t_SL g1629 ( 
.A1(n_1496),
.A2(n_1266),
.B1(n_740),
.B2(n_1504),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1383),
.B(n_1493),
.Y(n_1630)
);

AOI22xp33_ASAP7_75t_L g1631 ( 
.A1(n_1477),
.A2(n_900),
.B1(n_1133),
.B2(n_1390),
.Y(n_1631)
);

AOI22xp33_ASAP7_75t_L g1632 ( 
.A1(n_1477),
.A2(n_900),
.B1(n_1133),
.B2(n_1390),
.Y(n_1632)
);

BUFx4f_ASAP7_75t_SL g1633 ( 
.A(n_1469),
.Y(n_1633)
);

BUFx6f_ASAP7_75t_L g1634 ( 
.A(n_1378),
.Y(n_1634)
);

INVx5_ASAP7_75t_L g1635 ( 
.A(n_1401),
.Y(n_1635)
);

BUFx10_ASAP7_75t_L g1636 ( 
.A(n_1505),
.Y(n_1636)
);

AOI22xp33_ASAP7_75t_SL g1637 ( 
.A1(n_1496),
.A2(n_1266),
.B1(n_740),
.B2(n_1504),
.Y(n_1637)
);

BUFx8_ASAP7_75t_SL g1638 ( 
.A(n_1469),
.Y(n_1638)
);

OAI22xp5_ASAP7_75t_L g1639 ( 
.A1(n_1463),
.A2(n_1486),
.B1(n_1499),
.B2(n_1483),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1441),
.B(n_1484),
.Y(n_1640)
);

AOI22xp33_ASAP7_75t_L g1641 ( 
.A1(n_1477),
.A2(n_900),
.B1(n_1133),
.B2(n_1390),
.Y(n_1641)
);

AOI22xp33_ASAP7_75t_SL g1642 ( 
.A1(n_1496),
.A2(n_1266),
.B1(n_740),
.B2(n_1504),
.Y(n_1642)
);

AOI22xp33_ASAP7_75t_SL g1643 ( 
.A1(n_1496),
.A2(n_1266),
.B1(n_740),
.B2(n_1504),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1383),
.B(n_1493),
.Y(n_1644)
);

AOI22xp33_ASAP7_75t_L g1645 ( 
.A1(n_1390),
.A2(n_900),
.B1(n_1477),
.B2(n_1266),
.Y(n_1645)
);

AOI22xp33_ASAP7_75t_SL g1646 ( 
.A1(n_1496),
.A2(n_1266),
.B1(n_740),
.B2(n_1504),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1383),
.B(n_1493),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1399),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1399),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1399),
.Y(n_1650)
);

AOI22xp33_ASAP7_75t_SL g1651 ( 
.A1(n_1496),
.A2(n_1266),
.B1(n_740),
.B2(n_1504),
.Y(n_1651)
);

CKINVDCx11_ASAP7_75t_R g1652 ( 
.A(n_1469),
.Y(n_1652)
);

BUFx6f_ASAP7_75t_SL g1653 ( 
.A(n_1396),
.Y(n_1653)
);

OAI22xp33_ASAP7_75t_L g1654 ( 
.A1(n_1471),
.A2(n_1496),
.B1(n_900),
.B2(n_1444),
.Y(n_1654)
);

BUFx12f_ASAP7_75t_L g1655 ( 
.A(n_1505),
.Y(n_1655)
);

AOI22xp33_ASAP7_75t_SL g1656 ( 
.A1(n_1496),
.A2(n_1266),
.B1(n_740),
.B2(n_1504),
.Y(n_1656)
);

BUFx4f_ASAP7_75t_SL g1657 ( 
.A(n_1469),
.Y(n_1657)
);

CKINVDCx11_ASAP7_75t_R g1658 ( 
.A(n_1469),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1399),
.Y(n_1659)
);

OAI22xp33_ASAP7_75t_L g1660 ( 
.A1(n_1471),
.A2(n_1496),
.B1(n_900),
.B2(n_1444),
.Y(n_1660)
);

BUFx2_ASAP7_75t_L g1661 ( 
.A(n_1345),
.Y(n_1661)
);

AOI22xp33_ASAP7_75t_L g1662 ( 
.A1(n_1477),
.A2(n_900),
.B1(n_1133),
.B2(n_1390),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1399),
.Y(n_1663)
);

AOI22xp33_ASAP7_75t_SL g1664 ( 
.A1(n_1496),
.A2(n_1266),
.B1(n_740),
.B2(n_1504),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1353),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1399),
.Y(n_1666)
);

AOI22xp33_ASAP7_75t_L g1667 ( 
.A1(n_1477),
.A2(n_900),
.B1(n_1133),
.B2(n_1390),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1399),
.Y(n_1668)
);

OAI22xp5_ASAP7_75t_L g1669 ( 
.A1(n_1463),
.A2(n_1486),
.B1(n_1499),
.B2(n_1483),
.Y(n_1669)
);

AOI22xp33_ASAP7_75t_L g1670 ( 
.A1(n_1477),
.A2(n_900),
.B1(n_1133),
.B2(n_1390),
.Y(n_1670)
);

CKINVDCx11_ASAP7_75t_R g1671 ( 
.A(n_1469),
.Y(n_1671)
);

OAI22xp5_ASAP7_75t_L g1672 ( 
.A1(n_1463),
.A2(n_1486),
.B1(n_1499),
.B2(n_1483),
.Y(n_1672)
);

OAI22xp33_ASAP7_75t_L g1673 ( 
.A1(n_1471),
.A2(n_1496),
.B1(n_900),
.B2(n_1444),
.Y(n_1673)
);

CKINVDCx11_ASAP7_75t_R g1674 ( 
.A(n_1469),
.Y(n_1674)
);

OAI22xp5_ASAP7_75t_L g1675 ( 
.A1(n_1463),
.A2(n_1486),
.B1(n_1499),
.B2(n_1483),
.Y(n_1675)
);

CKINVDCx5p33_ASAP7_75t_R g1676 ( 
.A(n_1505),
.Y(n_1676)
);

CKINVDCx20_ASAP7_75t_R g1677 ( 
.A(n_1457),
.Y(n_1677)
);

BUFx10_ASAP7_75t_L g1678 ( 
.A(n_1505),
.Y(n_1678)
);

OAI22xp33_ASAP7_75t_L g1679 ( 
.A1(n_1471),
.A2(n_1496),
.B1(n_900),
.B2(n_1444),
.Y(n_1679)
);

BUFx2_ASAP7_75t_L g1680 ( 
.A(n_1345),
.Y(n_1680)
);

AOI211xp5_ASAP7_75t_L g1681 ( 
.A1(n_1520),
.A2(n_1654),
.B(n_1673),
.C(n_1660),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1607),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1559),
.Y(n_1683)
);

INVx2_ASAP7_75t_SL g1684 ( 
.A(n_1603),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1588),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1611),
.Y(n_1686)
);

AOI21x1_ASAP7_75t_L g1687 ( 
.A1(n_1592),
.A2(n_1595),
.B(n_1639),
.Y(n_1687)
);

CKINVDCx6p67_ASAP7_75t_R g1688 ( 
.A(n_1534),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1591),
.B(n_1538),
.Y(n_1689)
);

OAI21x1_ASAP7_75t_L g1690 ( 
.A1(n_1558),
.A2(n_1614),
.B(n_1618),
.Y(n_1690)
);

BUFx3_ASAP7_75t_L g1691 ( 
.A(n_1635),
.Y(n_1691)
);

INVx1_ASAP7_75t_SL g1692 ( 
.A(n_1623),
.Y(n_1692)
);

INVx3_ASAP7_75t_L g1693 ( 
.A(n_1603),
.Y(n_1693)
);

NOR2xp33_ASAP7_75t_L g1694 ( 
.A(n_1630),
.B(n_1644),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1543),
.Y(n_1695)
);

INVx3_ASAP7_75t_L g1696 ( 
.A(n_1603),
.Y(n_1696)
);

HB1xp67_ASAP7_75t_L g1697 ( 
.A(n_1584),
.Y(n_1697)
);

BUFx2_ASAP7_75t_L g1698 ( 
.A(n_1613),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1591),
.B(n_1556),
.Y(n_1699)
);

OA21x2_ASAP7_75t_L g1700 ( 
.A1(n_1602),
.A2(n_1608),
.B(n_1605),
.Y(n_1700)
);

HB1xp67_ASAP7_75t_L g1701 ( 
.A(n_1622),
.Y(n_1701)
);

BUFx6f_ASAP7_75t_L g1702 ( 
.A(n_1635),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1545),
.B(n_1551),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1563),
.Y(n_1704)
);

OA21x2_ASAP7_75t_L g1705 ( 
.A1(n_1621),
.A2(n_1578),
.B(n_1555),
.Y(n_1705)
);

INVx3_ASAP7_75t_L g1706 ( 
.A(n_1604),
.Y(n_1706)
);

OA21x2_ASAP7_75t_L g1707 ( 
.A1(n_1597),
.A2(n_1566),
.B(n_1526),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1545),
.B(n_1551),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1567),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1572),
.Y(n_1710)
);

INVx3_ASAP7_75t_L g1711 ( 
.A(n_1604),
.Y(n_1711)
);

INVx3_ASAP7_75t_L g1712 ( 
.A(n_1612),
.Y(n_1712)
);

INVx1_ASAP7_75t_SL g1713 ( 
.A(n_1661),
.Y(n_1713)
);

OR2x2_ASAP7_75t_L g1714 ( 
.A(n_1529),
.B(n_1539),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1620),
.Y(n_1715)
);

HB1xp67_ASAP7_75t_L g1716 ( 
.A(n_1593),
.Y(n_1716)
);

AOI22xp33_ASAP7_75t_L g1717 ( 
.A1(n_1629),
.A2(n_1643),
.B1(n_1656),
.B2(n_1651),
.Y(n_1717)
);

BUFx3_ASAP7_75t_L g1718 ( 
.A(n_1635),
.Y(n_1718)
);

OA21x2_ASAP7_75t_L g1719 ( 
.A1(n_1597),
.A2(n_1610),
.B(n_1523),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1574),
.Y(n_1720)
);

HB1xp67_ASAP7_75t_L g1721 ( 
.A(n_1580),
.Y(n_1721)
);

OAI21x1_ASAP7_75t_L g1722 ( 
.A1(n_1590),
.A2(n_1606),
.B(n_1669),
.Y(n_1722)
);

HB1xp67_ASAP7_75t_L g1723 ( 
.A(n_1617),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1609),
.Y(n_1724)
);

AO21x2_ASAP7_75t_L g1725 ( 
.A1(n_1520),
.A2(n_1660),
.B(n_1654),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1576),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1615),
.Y(n_1727)
);

CKINVDCx11_ASAP7_75t_R g1728 ( 
.A(n_1677),
.Y(n_1728)
);

OR2x2_ASAP7_75t_L g1729 ( 
.A(n_1529),
.B(n_1536),
.Y(n_1729)
);

NOR2xp33_ASAP7_75t_L g1730 ( 
.A(n_1647),
.B(n_1633),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1548),
.B(n_1536),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1609),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1575),
.Y(n_1733)
);

OR2x2_ASAP7_75t_L g1734 ( 
.A(n_1568),
.B(n_1537),
.Y(n_1734)
);

HB1xp67_ASAP7_75t_L g1735 ( 
.A(n_1616),
.Y(n_1735)
);

INVx2_ASAP7_75t_L g1736 ( 
.A(n_1557),
.Y(n_1736)
);

NOR2xp33_ASAP7_75t_L g1737 ( 
.A(n_1633),
.B(n_1657),
.Y(n_1737)
);

AOI21xp5_ASAP7_75t_SL g1738 ( 
.A1(n_1672),
.A2(n_1675),
.B(n_1679),
.Y(n_1738)
);

OAI21x1_ASAP7_75t_L g1739 ( 
.A1(n_1573),
.A2(n_1628),
.B(n_1553),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1575),
.Y(n_1740)
);

OA21x2_ASAP7_75t_L g1741 ( 
.A1(n_1586),
.A2(n_1565),
.B(n_1569),
.Y(n_1741)
);

AO21x1_ASAP7_75t_L g1742 ( 
.A1(n_1673),
.A2(n_1679),
.B(n_1626),
.Y(n_1742)
);

INVx1_ASAP7_75t_SL g1743 ( 
.A(n_1680),
.Y(n_1743)
);

BUFx2_ASAP7_75t_L g1744 ( 
.A(n_1557),
.Y(n_1744)
);

HB1xp67_ASAP7_75t_L g1745 ( 
.A(n_1557),
.Y(n_1745)
);

BUFx12f_ASAP7_75t_L g1746 ( 
.A(n_1624),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1571),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1548),
.B(n_1571),
.Y(n_1748)
);

OAI21x1_ASAP7_75t_L g1749 ( 
.A1(n_1628),
.A2(n_1540),
.B(n_1568),
.Y(n_1749)
);

BUFx2_ASAP7_75t_L g1750 ( 
.A(n_1601),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1533),
.B(n_1640),
.Y(n_1751)
);

HB1xp67_ASAP7_75t_L g1752 ( 
.A(n_1585),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1579),
.B(n_1627),
.Y(n_1753)
);

INVx3_ASAP7_75t_L g1754 ( 
.A(n_1601),
.Y(n_1754)
);

AOI22xp33_ASAP7_75t_SL g1755 ( 
.A1(n_1629),
.A2(n_1656),
.B1(n_1646),
.B2(n_1651),
.Y(n_1755)
);

AO21x1_ASAP7_75t_L g1756 ( 
.A1(n_1533),
.A2(n_1666),
.B(n_1663),
.Y(n_1756)
);

INVx3_ASAP7_75t_L g1757 ( 
.A(n_1599),
.Y(n_1757)
);

BUFx3_ASAP7_75t_L g1758 ( 
.A(n_1570),
.Y(n_1758)
);

OA21x2_ASAP7_75t_L g1759 ( 
.A1(n_1542),
.A2(n_1649),
.B(n_1659),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1579),
.Y(n_1760)
);

INVx2_ASAP7_75t_SL g1761 ( 
.A(n_1599),
.Y(n_1761)
);

OAI22xp33_ASAP7_75t_L g1762 ( 
.A1(n_1547),
.A2(n_1645),
.B1(n_1637),
.B2(n_1642),
.Y(n_1762)
);

INVx3_ASAP7_75t_L g1763 ( 
.A(n_1589),
.Y(n_1763)
);

AOI22xp33_ASAP7_75t_SL g1764 ( 
.A1(n_1637),
.A2(n_1664),
.B1(n_1646),
.B2(n_1643),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1648),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1650),
.Y(n_1766)
);

BUFx4f_ASAP7_75t_SL g1767 ( 
.A(n_1554),
.Y(n_1767)
);

BUFx2_ASAP7_75t_L g1768 ( 
.A(n_1550),
.Y(n_1768)
);

INVx4_ASAP7_75t_L g1769 ( 
.A(n_1589),
.Y(n_1769)
);

INVx1_ASAP7_75t_SL g1770 ( 
.A(n_1535),
.Y(n_1770)
);

HB1xp67_ASAP7_75t_L g1771 ( 
.A(n_1668),
.Y(n_1771)
);

AO21x1_ASAP7_75t_L g1772 ( 
.A1(n_1521),
.A2(n_1645),
.B(n_1642),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1619),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1541),
.B(n_1546),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1521),
.B(n_1598),
.Y(n_1775)
);

OAI21x1_ASAP7_75t_L g1776 ( 
.A1(n_1530),
.A2(n_1546),
.B(n_1665),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1583),
.B(n_1664),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1560),
.Y(n_1778)
);

HB1xp67_ASAP7_75t_L g1779 ( 
.A(n_1600),
.Y(n_1779)
);

OAI21x1_ASAP7_75t_L g1780 ( 
.A1(n_1631),
.A2(n_1670),
.B(n_1632),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1562),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1600),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1577),
.B(n_1596),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1641),
.B(n_1662),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1532),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1634),
.Y(n_1786)
);

AOI22xp33_ASAP7_75t_L g1787 ( 
.A1(n_1667),
.A2(n_1564),
.B1(n_1587),
.B2(n_1653),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1634),
.Y(n_1788)
);

INVx11_ASAP7_75t_L g1789 ( 
.A(n_1655),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1581),
.Y(n_1790)
);

INVx2_ASAP7_75t_L g1791 ( 
.A(n_1582),
.Y(n_1791)
);

BUFx3_ASAP7_75t_L g1792 ( 
.A(n_1594),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1594),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1587),
.Y(n_1794)
);

INVx1_ASAP7_75t_SL g1795 ( 
.A(n_1527),
.Y(n_1795)
);

AO21x1_ASAP7_75t_SL g1796 ( 
.A1(n_1552),
.A2(n_1522),
.B(n_1544),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1544),
.Y(n_1797)
);

HB1xp67_ASAP7_75t_L g1798 ( 
.A(n_1524),
.Y(n_1798)
);

OA21x2_ASAP7_75t_L g1799 ( 
.A1(n_1756),
.A2(n_1676),
.B(n_1625),
.Y(n_1799)
);

NOR2x1_ASAP7_75t_SL g1800 ( 
.A(n_1796),
.B(n_1561),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1768),
.B(n_1678),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1683),
.B(n_1657),
.Y(n_1802)
);

OAI21xp5_ASAP7_75t_L g1803 ( 
.A1(n_1738),
.A2(n_1528),
.B(n_1525),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1771),
.Y(n_1804)
);

OAI21xp5_ASAP7_75t_L g1805 ( 
.A1(n_1738),
.A2(n_1531),
.B(n_1549),
.Y(n_1805)
);

OR2x2_ASAP7_75t_L g1806 ( 
.A(n_1768),
.B(n_1658),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1698),
.B(n_1636),
.Y(n_1807)
);

AOI22xp5_ASAP7_75t_L g1808 ( 
.A1(n_1762),
.A2(n_1531),
.B1(n_1652),
.B2(n_1671),
.Y(n_1808)
);

OAI21xp33_ASAP7_75t_L g1809 ( 
.A1(n_1748),
.A2(n_1674),
.B(n_1638),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1698),
.B(n_1636),
.Y(n_1810)
);

OR2x2_ASAP7_75t_L g1811 ( 
.A(n_1721),
.B(n_1678),
.Y(n_1811)
);

A2O1A1Ixp33_ASAP7_75t_L g1812 ( 
.A1(n_1681),
.A2(n_1714),
.B(n_1748),
.C(n_1708),
.Y(n_1812)
);

AOI21xp5_ASAP7_75t_L g1813 ( 
.A1(n_1681),
.A2(n_1735),
.B(n_1725),
.Y(n_1813)
);

A2O1A1Ixp33_ASAP7_75t_L g1814 ( 
.A1(n_1714),
.A2(n_1703),
.B(n_1708),
.C(n_1731),
.Y(n_1814)
);

OA21x2_ASAP7_75t_L g1815 ( 
.A1(n_1756),
.A2(n_1749),
.B(n_1690),
.Y(n_1815)
);

OAI22xp5_ASAP7_75t_L g1816 ( 
.A1(n_1729),
.A2(n_1755),
.B1(n_1764),
.B2(n_1717),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1695),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1683),
.B(n_1685),
.Y(n_1818)
);

AND2x4_ASAP7_75t_L g1819 ( 
.A(n_1750),
.B(n_1754),
.Y(n_1819)
);

INVx3_ASAP7_75t_L g1820 ( 
.A(n_1754),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1692),
.B(n_1713),
.Y(n_1821)
);

INVxp67_ASAP7_75t_L g1822 ( 
.A(n_1730),
.Y(n_1822)
);

AOI31xp33_ASAP7_75t_L g1823 ( 
.A1(n_1742),
.A2(n_1703),
.A3(n_1772),
.B(n_1764),
.Y(n_1823)
);

OR3x1_ASAP7_75t_L g1824 ( 
.A(n_1685),
.B(n_1760),
.C(n_1740),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1695),
.Y(n_1825)
);

INVx4_ASAP7_75t_L g1826 ( 
.A(n_1706),
.Y(n_1826)
);

OAI22xp5_ASAP7_75t_L g1827 ( 
.A1(n_1729),
.A2(n_1755),
.B1(n_1784),
.B2(n_1733),
.Y(n_1827)
);

CKINVDCx5p33_ASAP7_75t_R g1828 ( 
.A(n_1728),
.Y(n_1828)
);

CKINVDCx5p33_ASAP7_75t_R g1829 ( 
.A(n_1746),
.Y(n_1829)
);

OAI21xp5_ASAP7_75t_L g1830 ( 
.A1(n_1687),
.A2(n_1707),
.B(n_1780),
.Y(n_1830)
);

AOI221xp5_ASAP7_75t_L g1831 ( 
.A1(n_1742),
.A2(n_1772),
.B1(n_1747),
.B2(n_1740),
.C(n_1733),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1689),
.B(n_1699),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1692),
.B(n_1713),
.Y(n_1833)
);

AOI22xp5_ASAP7_75t_L g1834 ( 
.A1(n_1725),
.A2(n_1784),
.B1(n_1731),
.B2(n_1741),
.Y(n_1834)
);

OAI21xp5_ASAP7_75t_L g1835 ( 
.A1(n_1707),
.A2(n_1780),
.B(n_1753),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1743),
.B(n_1751),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1743),
.B(n_1751),
.Y(n_1837)
);

NOR2xp33_ASAP7_75t_L g1838 ( 
.A(n_1694),
.B(n_1795),
.Y(n_1838)
);

NOR2xp33_ASAP7_75t_L g1839 ( 
.A(n_1795),
.B(n_1783),
.Y(n_1839)
);

A2O1A1Ixp33_ASAP7_75t_L g1840 ( 
.A1(n_1780),
.A2(n_1723),
.B(n_1747),
.C(n_1787),
.Y(n_1840)
);

BUFx2_ASAP7_75t_L g1841 ( 
.A(n_1779),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1704),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1723),
.B(n_1770),
.Y(n_1843)
);

OAI211xp5_ASAP7_75t_L g1844 ( 
.A1(n_1753),
.A2(n_1741),
.B(n_1707),
.C(n_1700),
.Y(n_1844)
);

NOR2xp33_ASAP7_75t_L g1845 ( 
.A(n_1783),
.B(n_1737),
.Y(n_1845)
);

OR2x2_ASAP7_75t_L g1846 ( 
.A(n_1697),
.B(n_1716),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1770),
.B(n_1779),
.Y(n_1847)
);

AOI221xp5_ASAP7_75t_L g1848 ( 
.A1(n_1725),
.A2(n_1773),
.B1(n_1775),
.B2(n_1774),
.C(n_1727),
.Y(n_1848)
);

AO32x2_ASAP7_75t_L g1849 ( 
.A1(n_1761),
.A2(n_1684),
.A3(n_1769),
.B1(n_1734),
.B2(n_1759),
.Y(n_1849)
);

AOI221xp5_ASAP7_75t_L g1850 ( 
.A1(n_1725),
.A2(n_1773),
.B1(n_1775),
.B2(n_1774),
.C(n_1727),
.Y(n_1850)
);

OA21x2_ASAP7_75t_L g1851 ( 
.A1(n_1749),
.A2(n_1690),
.B(n_1739),
.Y(n_1851)
);

AO21x1_ASAP7_75t_L g1852 ( 
.A1(n_1709),
.A2(n_1710),
.B(n_1766),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_L g1853 ( 
.A(n_1720),
.B(n_1726),
.Y(n_1853)
);

O2A1O1Ixp33_ASAP7_75t_L g1854 ( 
.A1(n_1707),
.A2(n_1741),
.B(n_1793),
.C(n_1761),
.Y(n_1854)
);

OAI211xp5_ASAP7_75t_L g1855 ( 
.A1(n_1741),
.A2(n_1700),
.B(n_1735),
.C(n_1705),
.Y(n_1855)
);

BUFx3_ASAP7_75t_L g1856 ( 
.A(n_1746),
.Y(n_1856)
);

NOR2xp33_ASAP7_75t_L g1857 ( 
.A(n_1798),
.B(n_1746),
.Y(n_1857)
);

A2O1A1Ixp33_ASAP7_75t_L g1858 ( 
.A1(n_1722),
.A2(n_1739),
.B(n_1734),
.C(n_1792),
.Y(n_1858)
);

A2O1A1Ixp33_ASAP7_75t_L g1859 ( 
.A1(n_1722),
.A2(n_1739),
.B(n_1792),
.C(n_1781),
.Y(n_1859)
);

AOI221xp5_ASAP7_75t_SL g1860 ( 
.A1(n_1782),
.A2(n_1682),
.B1(n_1720),
.B2(n_1726),
.C(n_1706),
.Y(n_1860)
);

O2A1O1Ixp33_ASAP7_75t_L g1861 ( 
.A1(n_1793),
.A2(n_1705),
.B(n_1711),
.C(n_1706),
.Y(n_1861)
);

A2O1A1Ixp33_ASAP7_75t_L g1862 ( 
.A1(n_1792),
.A2(n_1781),
.B(n_1777),
.C(n_1691),
.Y(n_1862)
);

NOR2xp33_ASAP7_75t_L g1863 ( 
.A(n_1798),
.B(n_1797),
.Y(n_1863)
);

A2O1A1Ixp33_ASAP7_75t_L g1864 ( 
.A1(n_1777),
.A2(n_1691),
.B(n_1718),
.C(n_1690),
.Y(n_1864)
);

AO32x2_ASAP7_75t_L g1865 ( 
.A1(n_1684),
.A2(n_1769),
.A3(n_1759),
.B1(n_1752),
.B2(n_1701),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1700),
.B(n_1790),
.Y(n_1866)
);

INVx1_ASAP7_75t_SL g1867 ( 
.A(n_1744),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1765),
.B(n_1766),
.Y(n_1868)
);

NOR2xp33_ASAP7_75t_L g1869 ( 
.A(n_1688),
.B(n_1767),
.Y(n_1869)
);

OA21x2_ASAP7_75t_L g1870 ( 
.A1(n_1749),
.A2(n_1776),
.B(n_1736),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1700),
.B(n_1790),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1682),
.Y(n_1872)
);

OR2x2_ASAP7_75t_L g1873 ( 
.A(n_1759),
.B(n_1705),
.Y(n_1873)
);

AND2x4_ASAP7_75t_L g1874 ( 
.A(n_1693),
.B(n_1696),
.Y(n_1874)
);

NOR2xp33_ASAP7_75t_L g1875 ( 
.A(n_1688),
.B(n_1789),
.Y(n_1875)
);

AOI22xp33_ASAP7_75t_L g1876 ( 
.A1(n_1778),
.A2(n_1759),
.B1(n_1705),
.B2(n_1700),
.Y(n_1876)
);

INVx1_ASAP7_75t_SL g1877 ( 
.A(n_1744),
.Y(n_1877)
);

AO21x1_ASAP7_75t_L g1878 ( 
.A1(n_1785),
.A2(n_1786),
.B(n_1788),
.Y(n_1878)
);

INVx3_ASAP7_75t_L g1879 ( 
.A(n_1763),
.Y(n_1879)
);

INVx3_ASAP7_75t_L g1880 ( 
.A(n_1879),
.Y(n_1880)
);

OR2x2_ASAP7_75t_L g1881 ( 
.A(n_1818),
.B(n_1719),
.Y(n_1881)
);

AND2x2_ASAP7_75t_L g1882 ( 
.A(n_1866),
.B(n_1719),
.Y(n_1882)
);

AND2x4_ASAP7_75t_L g1883 ( 
.A(n_1871),
.B(n_1693),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1852),
.Y(n_1884)
);

INVx1_ASAP7_75t_SL g1885 ( 
.A(n_1841),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1872),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1817),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1849),
.B(n_1719),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1825),
.Y(n_1889)
);

AND2x2_ASAP7_75t_L g1890 ( 
.A(n_1849),
.B(n_1719),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1842),
.Y(n_1891)
);

INVxp67_ASAP7_75t_SL g1892 ( 
.A(n_1854),
.Y(n_1892)
);

AND2x2_ASAP7_75t_L g1893 ( 
.A(n_1849),
.B(n_1719),
.Y(n_1893)
);

HB1xp67_ASAP7_75t_L g1894 ( 
.A(n_1846),
.Y(n_1894)
);

INVx2_ASAP7_75t_SL g1895 ( 
.A(n_1819),
.Y(n_1895)
);

BUFx3_ASAP7_75t_L g1896 ( 
.A(n_1856),
.Y(n_1896)
);

INVxp67_ASAP7_75t_SL g1897 ( 
.A(n_1860),
.Y(n_1897)
);

AOI22xp33_ASAP7_75t_L g1898 ( 
.A1(n_1831),
.A2(n_1778),
.B1(n_1686),
.B2(n_1794),
.Y(n_1898)
);

AND2x2_ASAP7_75t_SL g1899 ( 
.A(n_1799),
.B(n_1702),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1813),
.B(n_1757),
.Y(n_1900)
);

OR2x2_ASAP7_75t_L g1901 ( 
.A(n_1832),
.B(n_1745),
.Y(n_1901)
);

INVxp67_ASAP7_75t_SL g1902 ( 
.A(n_1860),
.Y(n_1902)
);

INVx1_ASAP7_75t_SL g1903 ( 
.A(n_1811),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1868),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1813),
.B(n_1757),
.Y(n_1905)
);

INVxp67_ASAP7_75t_SL g1906 ( 
.A(n_1861),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1868),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1853),
.Y(n_1908)
);

AND2x4_ASAP7_75t_L g1909 ( 
.A(n_1874),
.B(n_1757),
.Y(n_1909)
);

AND2x2_ASAP7_75t_L g1910 ( 
.A(n_1855),
.B(n_1865),
.Y(n_1910)
);

AND2x2_ASAP7_75t_L g1911 ( 
.A(n_1855),
.B(n_1715),
.Y(n_1911)
);

AND2x4_ASAP7_75t_L g1912 ( 
.A(n_1874),
.B(n_1712),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1804),
.B(n_1834),
.Y(n_1913)
);

CKINVDCx11_ASAP7_75t_R g1914 ( 
.A(n_1826),
.Y(n_1914)
);

BUFx2_ASAP7_75t_L g1915 ( 
.A(n_1867),
.Y(n_1915)
);

AND2x2_ASAP7_75t_L g1916 ( 
.A(n_1865),
.B(n_1851),
.Y(n_1916)
);

AOI22xp33_ASAP7_75t_L g1917 ( 
.A1(n_1831),
.A2(n_1724),
.B1(n_1732),
.B2(n_1791),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_SL g1918 ( 
.A(n_1803),
.B(n_1711),
.Y(n_1918)
);

INVx2_ASAP7_75t_L g1919 ( 
.A(n_1870),
.Y(n_1919)
);

BUFx3_ASAP7_75t_L g1920 ( 
.A(n_1878),
.Y(n_1920)
);

AOI22xp33_ASAP7_75t_L g1921 ( 
.A1(n_1898),
.A2(n_1827),
.B1(n_1816),
.B2(n_1850),
.Y(n_1921)
);

AND2x2_ASAP7_75t_L g1922 ( 
.A(n_1882),
.B(n_1821),
.Y(n_1922)
);

INVxp67_ASAP7_75t_SL g1923 ( 
.A(n_1920),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1886),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1886),
.Y(n_1925)
);

OAI221xp5_ASAP7_75t_L g1926 ( 
.A1(n_1898),
.A2(n_1812),
.B1(n_1808),
.B2(n_1823),
.C(n_1814),
.Y(n_1926)
);

BUFx3_ASAP7_75t_L g1927 ( 
.A(n_1914),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1897),
.B(n_1861),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1897),
.B(n_1844),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1887),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1889),
.Y(n_1931)
);

OAI22xp5_ASAP7_75t_L g1932 ( 
.A1(n_1902),
.A2(n_1823),
.B1(n_1827),
.B2(n_1824),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1889),
.Y(n_1933)
);

AOI211xp5_ASAP7_75t_L g1934 ( 
.A1(n_1906),
.A2(n_1803),
.B(n_1844),
.C(n_1816),
.Y(n_1934)
);

OR2x2_ASAP7_75t_L g1935 ( 
.A(n_1881),
.B(n_1873),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1902),
.B(n_1830),
.Y(n_1936)
);

AND2x2_ASAP7_75t_L g1937 ( 
.A(n_1882),
.B(n_1833),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1891),
.Y(n_1938)
);

AND2x2_ASAP7_75t_L g1939 ( 
.A(n_1882),
.B(n_1864),
.Y(n_1939)
);

BUFx3_ASAP7_75t_L g1940 ( 
.A(n_1915),
.Y(n_1940)
);

AND2x2_ASAP7_75t_L g1941 ( 
.A(n_1888),
.B(n_1815),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_L g1942 ( 
.A(n_1892),
.B(n_1830),
.Y(n_1942)
);

AND2x2_ASAP7_75t_L g1943 ( 
.A(n_1888),
.B(n_1815),
.Y(n_1943)
);

OAI33xp33_ASAP7_75t_L g1944 ( 
.A1(n_1884),
.A2(n_1802),
.A3(n_1809),
.B1(n_1822),
.B2(n_1806),
.B3(n_1829),
.Y(n_1944)
);

OAI31xp33_ASAP7_75t_L g1945 ( 
.A1(n_1917),
.A2(n_1840),
.A3(n_1858),
.B(n_1862),
.Y(n_1945)
);

INVx4_ASAP7_75t_L g1946 ( 
.A(n_1920),
.Y(n_1946)
);

AND2x2_ASAP7_75t_L g1947 ( 
.A(n_1888),
.B(n_1847),
.Y(n_1947)
);

INVx2_ASAP7_75t_L g1948 ( 
.A(n_1919),
.Y(n_1948)
);

NOR2xp33_ASAP7_75t_L g1949 ( 
.A(n_1903),
.B(n_1802),
.Y(n_1949)
);

OAI21xp5_ASAP7_75t_L g1950 ( 
.A1(n_1906),
.A2(n_1799),
.B(n_1850),
.Y(n_1950)
);

NAND3xp33_ASAP7_75t_L g1951 ( 
.A(n_1892),
.B(n_1848),
.C(n_1835),
.Y(n_1951)
);

AOI31xp33_ASAP7_75t_L g1952 ( 
.A1(n_1910),
.A2(n_1805),
.A3(n_1848),
.B(n_1857),
.Y(n_1952)
);

BUFx2_ASAP7_75t_L g1953 ( 
.A(n_1915),
.Y(n_1953)
);

NOR2xp33_ASAP7_75t_L g1954 ( 
.A(n_1903),
.B(n_1838),
.Y(n_1954)
);

INVx3_ASAP7_75t_L g1955 ( 
.A(n_1883),
.Y(n_1955)
);

AOI22xp33_ASAP7_75t_L g1956 ( 
.A1(n_1910),
.A2(n_1835),
.B1(n_1876),
.B2(n_1843),
.Y(n_1956)
);

AO21x2_ASAP7_75t_L g1957 ( 
.A1(n_1910),
.A2(n_1859),
.B(n_1776),
.Y(n_1957)
);

AND2x2_ASAP7_75t_L g1958 ( 
.A(n_1890),
.B(n_1867),
.Y(n_1958)
);

INVx2_ASAP7_75t_L g1959 ( 
.A(n_1919),
.Y(n_1959)
);

BUFx3_ASAP7_75t_L g1960 ( 
.A(n_1896),
.Y(n_1960)
);

AOI221xp5_ASAP7_75t_L g1961 ( 
.A1(n_1884),
.A2(n_1805),
.B1(n_1837),
.B2(n_1836),
.C(n_1863),
.Y(n_1961)
);

AND2x2_ASAP7_75t_L g1962 ( 
.A(n_1890),
.B(n_1877),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_L g1963 ( 
.A(n_1904),
.B(n_1877),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_SL g1964 ( 
.A(n_1920),
.B(n_1826),
.Y(n_1964)
);

INVx1_ASAP7_75t_SL g1965 ( 
.A(n_1885),
.Y(n_1965)
);

INVx5_ASAP7_75t_L g1966 ( 
.A(n_1890),
.Y(n_1966)
);

BUFx3_ASAP7_75t_L g1967 ( 
.A(n_1896),
.Y(n_1967)
);

INVx3_ASAP7_75t_L g1968 ( 
.A(n_1883),
.Y(n_1968)
);

INVx4_ASAP7_75t_L g1969 ( 
.A(n_1896),
.Y(n_1969)
);

AND2x4_ASAP7_75t_L g1970 ( 
.A(n_1883),
.B(n_1820),
.Y(n_1970)
);

NAND2x1_ASAP7_75t_L g1971 ( 
.A(n_1946),
.B(n_1895),
.Y(n_1971)
);

OR2x2_ASAP7_75t_L g1972 ( 
.A(n_1929),
.B(n_1913),
.Y(n_1972)
);

BUFx3_ASAP7_75t_L g1973 ( 
.A(n_1927),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_L g1974 ( 
.A(n_1929),
.B(n_1904),
.Y(n_1974)
);

AND2x4_ASAP7_75t_L g1975 ( 
.A(n_1966),
.B(n_1946),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1924),
.Y(n_1976)
);

HB1xp67_ASAP7_75t_L g1977 ( 
.A(n_1936),
.Y(n_1977)
);

INVx2_ASAP7_75t_SL g1978 ( 
.A(n_1966),
.Y(n_1978)
);

INVx2_ASAP7_75t_L g1979 ( 
.A(n_1948),
.Y(n_1979)
);

AND2x4_ASAP7_75t_L g1980 ( 
.A(n_1966),
.B(n_1893),
.Y(n_1980)
);

AOI22xp5_ASAP7_75t_L g1981 ( 
.A1(n_1921),
.A2(n_1893),
.B1(n_1918),
.B2(n_1913),
.Y(n_1981)
);

OR2x2_ASAP7_75t_L g1982 ( 
.A(n_1936),
.B(n_1894),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1924),
.Y(n_1983)
);

AND2x2_ASAP7_75t_L g1984 ( 
.A(n_1939),
.B(n_1922),
.Y(n_1984)
);

AND2x2_ASAP7_75t_L g1985 ( 
.A(n_1939),
.B(n_1883),
.Y(n_1985)
);

NAND2x1_ASAP7_75t_L g1986 ( 
.A(n_1946),
.B(n_1880),
.Y(n_1986)
);

BUFx2_ASAP7_75t_L g1987 ( 
.A(n_1946),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1925),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_L g1989 ( 
.A(n_1942),
.B(n_1907),
.Y(n_1989)
);

AND2x2_ASAP7_75t_L g1990 ( 
.A(n_1939),
.B(n_1909),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_L g1991 ( 
.A(n_1942),
.B(n_1907),
.Y(n_1991)
);

NAND2xp33_ASAP7_75t_R g1992 ( 
.A(n_1953),
.B(n_1828),
.Y(n_1992)
);

AND2x2_ASAP7_75t_L g1993 ( 
.A(n_1922),
.B(n_1909),
.Y(n_1993)
);

AND2x2_ASAP7_75t_L g1994 ( 
.A(n_1922),
.B(n_1909),
.Y(n_1994)
);

HB1xp67_ASAP7_75t_L g1995 ( 
.A(n_1928),
.Y(n_1995)
);

AND2x4_ASAP7_75t_L g1996 ( 
.A(n_1946),
.B(n_1893),
.Y(n_1996)
);

INVx1_ASAP7_75t_SL g1997 ( 
.A(n_1965),
.Y(n_1997)
);

INVx2_ASAP7_75t_L g1998 ( 
.A(n_1948),
.Y(n_1998)
);

OR2x2_ASAP7_75t_L g1999 ( 
.A(n_1928),
.B(n_1901),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1925),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_L g2001 ( 
.A(n_1923),
.B(n_1935),
.Y(n_2001)
);

BUFx3_ASAP7_75t_L g2002 ( 
.A(n_1927),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_L g2003 ( 
.A(n_1923),
.B(n_1908),
.Y(n_2003)
);

OR2x2_ASAP7_75t_L g2004 ( 
.A(n_1935),
.B(n_1901),
.Y(n_2004)
);

AOI21xp5_ASAP7_75t_L g2005 ( 
.A1(n_1950),
.A2(n_1900),
.B(n_1905),
.Y(n_2005)
);

INVx2_ASAP7_75t_L g2006 ( 
.A(n_1948),
.Y(n_2006)
);

OAI31xp33_ASAP7_75t_L g2007 ( 
.A1(n_1932),
.A2(n_1926),
.A3(n_1921),
.B(n_1951),
.Y(n_2007)
);

AND2x2_ASAP7_75t_L g2008 ( 
.A(n_1937),
.B(n_1912),
.Y(n_2008)
);

AND2x4_ASAP7_75t_L g2009 ( 
.A(n_1955),
.B(n_1916),
.Y(n_2009)
);

AND2x4_ASAP7_75t_L g2010 ( 
.A(n_1955),
.B(n_1916),
.Y(n_2010)
);

OR2x2_ASAP7_75t_L g2011 ( 
.A(n_1953),
.B(n_1881),
.Y(n_2011)
);

INVx2_ASAP7_75t_L g2012 ( 
.A(n_1959),
.Y(n_2012)
);

INVx2_ASAP7_75t_L g2013 ( 
.A(n_1979),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1976),
.Y(n_2014)
);

NOR2xp33_ASAP7_75t_L g2015 ( 
.A(n_1973),
.B(n_1927),
.Y(n_2015)
);

OAI21xp5_ASAP7_75t_L g2016 ( 
.A1(n_2007),
.A2(n_1926),
.B(n_1952),
.Y(n_2016)
);

AND2x2_ASAP7_75t_L g2017 ( 
.A(n_1984),
.B(n_1955),
.Y(n_2017)
);

INVx2_ASAP7_75t_L g2018 ( 
.A(n_1979),
.Y(n_2018)
);

AND2x2_ASAP7_75t_L g2019 ( 
.A(n_1984),
.B(n_1955),
.Y(n_2019)
);

OAI21xp5_ASAP7_75t_SL g2020 ( 
.A1(n_2007),
.A2(n_1952),
.B(n_1950),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1976),
.Y(n_2021)
);

INVx1_ASAP7_75t_SL g2022 ( 
.A(n_1973),
.Y(n_2022)
);

INVxp33_ASAP7_75t_L g2023 ( 
.A(n_1973),
.Y(n_2023)
);

INVx3_ASAP7_75t_L g2024 ( 
.A(n_1980),
.Y(n_2024)
);

AOI21xp5_ASAP7_75t_L g2025 ( 
.A1(n_2005),
.A2(n_1934),
.B(n_1951),
.Y(n_2025)
);

INVx2_ASAP7_75t_L g2026 ( 
.A(n_1979),
.Y(n_2026)
);

NAND2xp5_ASAP7_75t_L g2027 ( 
.A(n_1995),
.B(n_1930),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1983),
.Y(n_2028)
);

OR2x2_ASAP7_75t_L g2029 ( 
.A(n_1995),
.B(n_1963),
.Y(n_2029)
);

AND2x2_ASAP7_75t_L g2030 ( 
.A(n_1990),
.B(n_1968),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_1977),
.B(n_1931),
.Y(n_2031)
);

INVx2_ASAP7_75t_L g2032 ( 
.A(n_1998),
.Y(n_2032)
);

HB1xp67_ASAP7_75t_L g2033 ( 
.A(n_2003),
.Y(n_2033)
);

INVxp67_ASAP7_75t_L g2034 ( 
.A(n_2002),
.Y(n_2034)
);

INVx2_ASAP7_75t_L g2035 ( 
.A(n_1998),
.Y(n_2035)
);

OR2x2_ASAP7_75t_L g2036 ( 
.A(n_1972),
.B(n_1963),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_1983),
.Y(n_2037)
);

OR2x2_ASAP7_75t_L g2038 ( 
.A(n_1972),
.B(n_1965),
.Y(n_2038)
);

INVx2_ASAP7_75t_L g2039 ( 
.A(n_1998),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1988),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1988),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_SL g2042 ( 
.A(n_1997),
.B(n_1961),
.Y(n_2042)
);

AND2x2_ASAP7_75t_L g2043 ( 
.A(n_1985),
.B(n_1968),
.Y(n_2043)
);

OR2x2_ASAP7_75t_L g2044 ( 
.A(n_1974),
.B(n_1931),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_L g2045 ( 
.A(n_1977),
.B(n_1933),
.Y(n_2045)
);

INVx2_ASAP7_75t_L g2046 ( 
.A(n_2006),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_L g2047 ( 
.A(n_1974),
.B(n_1933),
.Y(n_2047)
);

AND2x2_ASAP7_75t_L g2048 ( 
.A(n_2008),
.B(n_1969),
.Y(n_2048)
);

NAND2xp5_ASAP7_75t_L g2049 ( 
.A(n_1999),
.B(n_1938),
.Y(n_2049)
);

AND2x2_ASAP7_75t_L g2050 ( 
.A(n_1993),
.B(n_1969),
.Y(n_2050)
);

OR2x2_ASAP7_75t_L g2051 ( 
.A(n_1999),
.B(n_1938),
.Y(n_2051)
);

AND2x2_ASAP7_75t_L g2052 ( 
.A(n_1993),
.B(n_1969),
.Y(n_2052)
);

NAND2x1p5_ASAP7_75t_L g2053 ( 
.A(n_1971),
.B(n_1969),
.Y(n_2053)
);

CKINVDCx16_ASAP7_75t_R g2054 ( 
.A(n_1992),
.Y(n_2054)
);

AND2x4_ASAP7_75t_SL g2055 ( 
.A(n_1975),
.B(n_1970),
.Y(n_2055)
);

INVx1_ASAP7_75t_SL g2056 ( 
.A(n_2002),
.Y(n_2056)
);

AND2x2_ASAP7_75t_L g2057 ( 
.A(n_1980),
.B(n_1940),
.Y(n_2057)
);

A2O1A1Ixp33_ASAP7_75t_L g2058 ( 
.A1(n_1981),
.A2(n_1934),
.B(n_1945),
.C(n_1956),
.Y(n_2058)
);

OAI21xp33_ASAP7_75t_L g2059 ( 
.A1(n_2005),
.A2(n_1956),
.B(n_1932),
.Y(n_2059)
);

AND2x2_ASAP7_75t_L g2060 ( 
.A(n_1994),
.B(n_1960),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_2000),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_2000),
.Y(n_2062)
);

NAND2xp5_ASAP7_75t_L g2063 ( 
.A(n_2025),
.B(n_1997),
.Y(n_2063)
);

OR2x2_ASAP7_75t_L g2064 ( 
.A(n_2038),
.B(n_1982),
.Y(n_2064)
);

INVx5_ASAP7_75t_L g2065 ( 
.A(n_2054),
.Y(n_2065)
);

INVx2_ASAP7_75t_L g2066 ( 
.A(n_2019),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_2014),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_2014),
.Y(n_2068)
);

INVx2_ASAP7_75t_L g2069 ( 
.A(n_2019),
.Y(n_2069)
);

AND2x2_ASAP7_75t_L g2070 ( 
.A(n_2060),
.B(n_2054),
.Y(n_2070)
);

NAND2xp5_ASAP7_75t_L g2071 ( 
.A(n_2025),
.B(n_2020),
.Y(n_2071)
);

OR2x2_ASAP7_75t_L g2072 ( 
.A(n_2038),
.B(n_1982),
.Y(n_2072)
);

NOR2xp33_ASAP7_75t_L g2073 ( 
.A(n_2020),
.B(n_2002),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_2021),
.Y(n_2074)
);

INVx2_ASAP7_75t_R g2075 ( 
.A(n_2021),
.Y(n_2075)
);

INVx1_ASAP7_75t_SL g2076 ( 
.A(n_2022),
.Y(n_2076)
);

AOI21xp5_ASAP7_75t_L g2077 ( 
.A1(n_2016),
.A2(n_1944),
.B(n_1981),
.Y(n_2077)
);

NOR2xp33_ASAP7_75t_L g2078 ( 
.A(n_2016),
.B(n_1944),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_2028),
.Y(n_2079)
);

INVxp67_ASAP7_75t_L g2080 ( 
.A(n_2015),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_2028),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_2037),
.Y(n_2082)
);

INVxp67_ASAP7_75t_L g2083 ( 
.A(n_2022),
.Y(n_2083)
);

NAND2xp33_ASAP7_75t_SL g2084 ( 
.A(n_2023),
.B(n_1971),
.Y(n_2084)
);

INVxp67_ASAP7_75t_L g2085 ( 
.A(n_2056),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_2037),
.Y(n_2086)
);

OR2x2_ASAP7_75t_L g2087 ( 
.A(n_2036),
.B(n_1989),
.Y(n_2087)
);

NAND2xp5_ASAP7_75t_L g2088 ( 
.A(n_2058),
.B(n_1989),
.Y(n_2088)
);

AOI21xp5_ASAP7_75t_L g2089 ( 
.A1(n_2042),
.A2(n_1945),
.B(n_1991),
.Y(n_2089)
);

OR2x2_ASAP7_75t_L g2090 ( 
.A(n_2036),
.B(n_1991),
.Y(n_2090)
);

NAND2xp5_ASAP7_75t_L g2091 ( 
.A(n_2056),
.B(n_2001),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_2040),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_L g2093 ( 
.A(n_2034),
.B(n_2001),
.Y(n_2093)
);

AND2x2_ASAP7_75t_L g2094 ( 
.A(n_2060),
.B(n_2055),
.Y(n_2094)
);

AND2x2_ASAP7_75t_L g2095 ( 
.A(n_2055),
.B(n_1975),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_2040),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_2041),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_L g2098 ( 
.A(n_2034),
.B(n_1954),
.Y(n_2098)
);

INVx2_ASAP7_75t_L g2099 ( 
.A(n_2019),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_L g2100 ( 
.A(n_2033),
.B(n_1954),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_L g2101 ( 
.A(n_2033),
.B(n_2003),
.Y(n_2101)
);

AND2x2_ASAP7_75t_L g2102 ( 
.A(n_2055),
.B(n_1975),
.Y(n_2102)
);

NAND2xp5_ASAP7_75t_L g2103 ( 
.A(n_2071),
.B(n_2089),
.Y(n_2103)
);

AOI22xp33_ASAP7_75t_L g2104 ( 
.A1(n_2078),
.A2(n_2059),
.B1(n_1957),
.B2(n_1943),
.Y(n_2104)
);

NAND2xp5_ASAP7_75t_L g2105 ( 
.A(n_2078),
.B(n_2059),
.Y(n_2105)
);

OR2x2_ASAP7_75t_L g2106 ( 
.A(n_2063),
.B(n_2029),
.Y(n_2106)
);

OAI21xp5_ASAP7_75t_L g2107 ( 
.A1(n_2077),
.A2(n_2027),
.B(n_2029),
.Y(n_2107)
);

AOI21xp5_ASAP7_75t_L g2108 ( 
.A1(n_2088),
.A2(n_2027),
.B(n_2031),
.Y(n_2108)
);

NOR2xp67_ASAP7_75t_L g2109 ( 
.A(n_2065),
.B(n_2024),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_2067),
.Y(n_2110)
);

NOR2xp33_ASAP7_75t_L g2111 ( 
.A(n_2065),
.B(n_1869),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_2068),
.Y(n_2112)
);

OR2x2_ASAP7_75t_L g2113 ( 
.A(n_2087),
.B(n_2051),
.Y(n_2113)
);

NAND2xp5_ASAP7_75t_SL g2114 ( 
.A(n_2065),
.B(n_1987),
.Y(n_2114)
);

AOI32xp33_ASAP7_75t_L g2115 ( 
.A1(n_2073),
.A2(n_1996),
.A3(n_1943),
.B1(n_1941),
.B2(n_1980),
.Y(n_2115)
);

INVx2_ASAP7_75t_L g2116 ( 
.A(n_2066),
.Y(n_2116)
);

NAND2xp5_ASAP7_75t_L g2117 ( 
.A(n_2076),
.B(n_2049),
.Y(n_2117)
);

INVx2_ASAP7_75t_L g2118 ( 
.A(n_2066),
.Y(n_2118)
);

AOI22xp33_ASAP7_75t_SL g2119 ( 
.A1(n_2065),
.A2(n_1941),
.B1(n_1943),
.B2(n_1957),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_2074),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_2079),
.Y(n_2121)
);

INVxp67_ASAP7_75t_SL g2122 ( 
.A(n_2073),
.Y(n_2122)
);

OAI31xp33_ASAP7_75t_L g2123 ( 
.A1(n_2070),
.A2(n_1941),
.A3(n_1996),
.B(n_1980),
.Y(n_2123)
);

AOI211x1_ASAP7_75t_L g2124 ( 
.A1(n_2070),
.A2(n_2017),
.B(n_2049),
.C(n_2043),
.Y(n_2124)
);

HB1xp67_ASAP7_75t_L g2125 ( 
.A(n_2083),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_2081),
.Y(n_2126)
);

AOI222xp33_ASAP7_75t_L g2127 ( 
.A1(n_2065),
.A2(n_1961),
.B1(n_1996),
.B2(n_2013),
.C1(n_2026),
.C2(n_2039),
.Y(n_2127)
);

INVx2_ASAP7_75t_L g2128 ( 
.A(n_2069),
.Y(n_2128)
);

AOI221xp5_ASAP7_75t_L g2129 ( 
.A1(n_2100),
.A2(n_2101),
.B1(n_2085),
.B2(n_2093),
.C(n_2091),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_2082),
.Y(n_2130)
);

AOI211xp5_ASAP7_75t_SL g2131 ( 
.A1(n_2080),
.A2(n_2024),
.B(n_1975),
.C(n_2057),
.Y(n_2131)
);

NAND2xp5_ASAP7_75t_L g2132 ( 
.A(n_2103),
.B(n_2098),
.Y(n_2132)
);

AOI221xp5_ASAP7_75t_L g2133 ( 
.A1(n_2105),
.A2(n_2092),
.B1(n_2086),
.B2(n_2097),
.C(n_2096),
.Y(n_2133)
);

OR2x2_ASAP7_75t_L g2134 ( 
.A(n_2106),
.B(n_2064),
.Y(n_2134)
);

NAND2xp5_ASAP7_75t_L g2135 ( 
.A(n_2108),
.B(n_2072),
.Y(n_2135)
);

AOI22xp5_ASAP7_75t_L g2136 ( 
.A1(n_2104),
.A2(n_1957),
.B1(n_1996),
.B2(n_2094),
.Y(n_2136)
);

OAI322xp33_ASAP7_75t_L g2137 ( 
.A1(n_2106),
.A2(n_2090),
.A3(n_2087),
.B1(n_2069),
.B2(n_2099),
.C1(n_2045),
.C2(n_2031),
.Y(n_2137)
);

AND2x2_ASAP7_75t_L g2138 ( 
.A(n_2111),
.B(n_2094),
.Y(n_2138)
);

OAI22xp33_ASAP7_75t_L g2139 ( 
.A1(n_2107),
.A2(n_1978),
.B1(n_1881),
.B2(n_2090),
.Y(n_2139)
);

O2A1O1Ixp5_ASAP7_75t_L g2140 ( 
.A1(n_2131),
.A2(n_2084),
.B(n_2099),
.C(n_2095),
.Y(n_2140)
);

OAI221xp5_ASAP7_75t_L g2141 ( 
.A1(n_2119),
.A2(n_2084),
.B1(n_2075),
.B2(n_1987),
.C(n_2045),
.Y(n_2141)
);

INVx2_ASAP7_75t_L g2142 ( 
.A(n_2116),
.Y(n_2142)
);

INVxp67_ASAP7_75t_SL g2143 ( 
.A(n_2109),
.Y(n_2143)
);

OR2x2_ASAP7_75t_L g2144 ( 
.A(n_2125),
.B(n_2051),
.Y(n_2144)
);

INVx1_ASAP7_75t_SL g2145 ( 
.A(n_2117),
.Y(n_2145)
);

OAI22xp33_ASAP7_75t_L g2146 ( 
.A1(n_2122),
.A2(n_1978),
.B1(n_2011),
.B2(n_2024),
.Y(n_2146)
);

AOI22xp5_ASAP7_75t_L g2147 ( 
.A1(n_2127),
.A2(n_1957),
.B1(n_1899),
.B2(n_2013),
.Y(n_2147)
);

INVx1_ASAP7_75t_SL g2148 ( 
.A(n_2113),
.Y(n_2148)
);

OAI32xp33_ASAP7_75t_L g2149 ( 
.A1(n_2113),
.A2(n_2024),
.A3(n_2095),
.B1(n_2102),
.B2(n_2075),
.Y(n_2149)
);

NOR2xp33_ASAP7_75t_SL g2150 ( 
.A(n_2123),
.B(n_1875),
.Y(n_2150)
);

NOR3xp33_ASAP7_75t_SL g2151 ( 
.A(n_2114),
.B(n_1964),
.C(n_1845),
.Y(n_2151)
);

AOI321xp33_ASAP7_75t_L g2152 ( 
.A1(n_2129),
.A2(n_2102),
.A3(n_1911),
.B1(n_2013),
.B2(n_2018),
.C(n_2026),
.Y(n_2152)
);

OAI211xp5_ASAP7_75t_L g2153 ( 
.A1(n_2124),
.A2(n_2114),
.B(n_2115),
.C(n_2121),
.Y(n_2153)
);

INVx2_ASAP7_75t_L g2154 ( 
.A(n_2116),
.Y(n_2154)
);

NOR2xp33_ASAP7_75t_L g2155 ( 
.A(n_2132),
.B(n_2118),
.Y(n_2155)
);

NAND3xp33_ASAP7_75t_L g2156 ( 
.A(n_2152),
.B(n_2128),
.C(n_2118),
.Y(n_2156)
);

NAND2xp33_ASAP7_75t_SL g2157 ( 
.A(n_2151),
.B(n_2128),
.Y(n_2157)
);

AO22x1_ASAP7_75t_L g2158 ( 
.A1(n_2143),
.A2(n_2126),
.B1(n_2130),
.B2(n_2121),
.Y(n_2158)
);

OAI21xp33_ASAP7_75t_L g2159 ( 
.A1(n_2150),
.A2(n_2112),
.B(n_2110),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_2134),
.Y(n_2160)
);

INVx1_ASAP7_75t_SL g2161 ( 
.A(n_2148),
.Y(n_2161)
);

OAI21xp33_ASAP7_75t_L g2162 ( 
.A1(n_2138),
.A2(n_2120),
.B(n_2126),
.Y(n_2162)
);

INVxp67_ASAP7_75t_L g2163 ( 
.A(n_2135),
.Y(n_2163)
);

NAND2xp5_ASAP7_75t_L g2164 ( 
.A(n_2145),
.B(n_2144),
.Y(n_2164)
);

AND2x4_ASAP7_75t_L g2165 ( 
.A(n_2142),
.B(n_2130),
.Y(n_2165)
);

OAI22xp5_ASAP7_75t_L g2166 ( 
.A1(n_2141),
.A2(n_1978),
.B1(n_2010),
.B2(n_2009),
.Y(n_2166)
);

NOR2xp33_ASAP7_75t_L g2167 ( 
.A(n_2137),
.B(n_1789),
.Y(n_2167)
);

AOI22xp5_ASAP7_75t_L g2168 ( 
.A1(n_2147),
.A2(n_2039),
.B1(n_2018),
.B2(n_2026),
.Y(n_2168)
);

INVxp67_ASAP7_75t_L g2169 ( 
.A(n_2154),
.Y(n_2169)
);

INVxp67_ASAP7_75t_SL g2170 ( 
.A(n_2133),
.Y(n_2170)
);

NOR2x1_ASAP7_75t_L g2171 ( 
.A(n_2161),
.B(n_2153),
.Y(n_2171)
);

NOR5xp2_ASAP7_75t_L g2172 ( 
.A(n_2170),
.B(n_2141),
.C(n_2149),
.D(n_2153),
.E(n_2140),
.Y(n_2172)
);

NAND3xp33_ASAP7_75t_L g2173 ( 
.A(n_2163),
.B(n_2133),
.C(n_2155),
.Y(n_2173)
);

NAND4xp75_ASAP7_75t_L g2174 ( 
.A(n_2164),
.B(n_2136),
.C(n_2057),
.D(n_2146),
.Y(n_2174)
);

NAND4xp25_ASAP7_75t_L g2175 ( 
.A(n_2167),
.B(n_2057),
.C(n_2017),
.D(n_2043),
.Y(n_2175)
);

O2A1O1Ixp33_ASAP7_75t_L g2176 ( 
.A1(n_2169),
.A2(n_2139),
.B(n_2047),
.C(n_2044),
.Y(n_2176)
);

OR2x2_ASAP7_75t_L g2177 ( 
.A(n_2160),
.B(n_2044),
.Y(n_2177)
);

OAI21xp5_ASAP7_75t_L g2178 ( 
.A1(n_2156),
.A2(n_2061),
.B(n_2041),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_2165),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_2165),
.Y(n_2180)
);

HB1xp67_ASAP7_75t_L g2181 ( 
.A(n_2158),
.Y(n_2181)
);

NOR2xp33_ASAP7_75t_L g2182 ( 
.A(n_2162),
.B(n_2053),
.Y(n_2182)
);

NOR4xp25_ASAP7_75t_L g2183 ( 
.A(n_2159),
.B(n_2061),
.C(n_2062),
.D(n_2035),
.Y(n_2183)
);

OAI22xp5_ASAP7_75t_L g2184 ( 
.A1(n_2171),
.A2(n_2166),
.B1(n_2168),
.B2(n_2047),
.Y(n_2184)
);

OAI21xp5_ASAP7_75t_L g2185 ( 
.A1(n_2173),
.A2(n_2157),
.B(n_2062),
.Y(n_2185)
);

AOI221xp5_ASAP7_75t_L g2186 ( 
.A1(n_2181),
.A2(n_2035),
.B1(n_2032),
.B2(n_2046),
.C(n_2018),
.Y(n_2186)
);

OAI211xp5_ASAP7_75t_L g2187 ( 
.A1(n_2183),
.A2(n_1986),
.B(n_1964),
.C(n_2043),
.Y(n_2187)
);

NAND2xp5_ASAP7_75t_SL g2188 ( 
.A(n_2179),
.B(n_2053),
.Y(n_2188)
);

AOI221xp5_ASAP7_75t_L g2189 ( 
.A1(n_2178),
.A2(n_2032),
.B1(n_2035),
.B2(n_2039),
.C(n_2046),
.Y(n_2189)
);

NAND2xp5_ASAP7_75t_L g2190 ( 
.A(n_2180),
.B(n_2030),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_2190),
.Y(n_2191)
);

AOI22xp5_ASAP7_75t_L g2192 ( 
.A1(n_2184),
.A2(n_2174),
.B1(n_2182),
.B2(n_2177),
.Y(n_2192)
);

NAND3xp33_ASAP7_75t_SL g2193 ( 
.A(n_2185),
.B(n_2172),
.C(n_2176),
.Y(n_2193)
);

AOI22xp5_ASAP7_75t_L g2194 ( 
.A1(n_2186),
.A2(n_2175),
.B1(n_2032),
.B2(n_2046),
.Y(n_2194)
);

NOR2x1_ASAP7_75t_L g2195 ( 
.A(n_2188),
.B(n_1960),
.Y(n_2195)
);

AOI322xp5_ASAP7_75t_L g2196 ( 
.A1(n_2189),
.A2(n_1899),
.A3(n_1958),
.B1(n_1962),
.B2(n_2006),
.C1(n_2012),
.C2(n_1947),
.Y(n_2196)
);

AOI21xp5_ASAP7_75t_L g2197 ( 
.A1(n_2187),
.A2(n_1800),
.B(n_2053),
.Y(n_2197)
);

OAI211xp5_ASAP7_75t_SL g2198 ( 
.A1(n_2185),
.A2(n_2011),
.B(n_1839),
.C(n_2004),
.Y(n_2198)
);

XNOR2xp5_ASAP7_75t_L g2199 ( 
.A(n_2193),
.B(n_1796),
.Y(n_2199)
);

NAND2xp5_ASAP7_75t_L g2200 ( 
.A(n_2191),
.B(n_1940),
.Y(n_2200)
);

NOR2x1_ASAP7_75t_L g2201 ( 
.A(n_2195),
.B(n_1960),
.Y(n_2201)
);

NOR2x1_ASAP7_75t_L g2202 ( 
.A(n_2198),
.B(n_1967),
.Y(n_2202)
);

INVx2_ASAP7_75t_L g2203 ( 
.A(n_2194),
.Y(n_2203)
);

XNOR2x1_ASAP7_75t_L g2204 ( 
.A(n_2192),
.B(n_1807),
.Y(n_2204)
);

OAI22xp33_ASAP7_75t_L g2205 ( 
.A1(n_2203),
.A2(n_2197),
.B1(n_2196),
.B2(n_2053),
.Y(n_2205)
);

NOR3xp33_ASAP7_75t_L g2206 ( 
.A(n_2200),
.B(n_1810),
.C(n_1758),
.Y(n_2206)
);

OA22x2_ASAP7_75t_L g2207 ( 
.A1(n_2199),
.A2(n_1986),
.B1(n_2052),
.B2(n_2050),
.Y(n_2207)
);

OAI221xp5_ASAP7_75t_L g2208 ( 
.A1(n_2201),
.A2(n_1967),
.B1(n_2006),
.B2(n_2012),
.C(n_1949),
.Y(n_2208)
);

HB1xp67_ASAP7_75t_L g2209 ( 
.A(n_2207),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_2208),
.Y(n_2210)
);

CKINVDCx20_ASAP7_75t_R g2211 ( 
.A(n_2209),
.Y(n_2211)
);

NAND2xp5_ASAP7_75t_L g2212 ( 
.A(n_2211),
.B(n_2204),
.Y(n_2212)
);

INVx4_ASAP7_75t_L g2213 ( 
.A(n_2211),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_2213),
.Y(n_2214)
);

OAI22xp5_ASAP7_75t_L g2215 ( 
.A1(n_2212),
.A2(n_2205),
.B1(n_2210),
.B2(n_2202),
.Y(n_2215)
);

AOI221xp5_ASAP7_75t_L g2216 ( 
.A1(n_2215),
.A2(n_2206),
.B1(n_2012),
.B2(n_2009),
.C(n_2010),
.Y(n_2216)
);

AOI21xp5_ASAP7_75t_L g2217 ( 
.A1(n_2214),
.A2(n_2010),
.B(n_2009),
.Y(n_2217)
);

OAI21xp5_ASAP7_75t_L g2218 ( 
.A1(n_2217),
.A2(n_2050),
.B(n_2048),
.Y(n_2218)
);

NAND2xp5_ASAP7_75t_SL g2219 ( 
.A(n_2218),
.B(n_2216),
.Y(n_2219)
);

INVx2_ASAP7_75t_L g2220 ( 
.A(n_2219),
.Y(n_2220)
);

AOI221xp5_ASAP7_75t_L g2221 ( 
.A1(n_2220),
.A2(n_1949),
.B1(n_2009),
.B2(n_2010),
.C(n_1967),
.Y(n_2221)
);

AOI211xp5_ASAP7_75t_L g2222 ( 
.A1(n_2221),
.A2(n_1688),
.B(n_1758),
.C(n_1801),
.Y(n_2222)
);


endmodule