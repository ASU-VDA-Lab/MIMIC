module fake_jpeg_13996_n_179 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_179);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_179;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_122;
wire n_75;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

INVx11_ASAP7_75t_SL g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_35),
.Y(n_51)
);

INVx4_ASAP7_75t_SL g36 ( 
.A(n_29),
.Y(n_36)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_30),
.B(n_1),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_37),
.B(n_40),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_29),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_42),
.Y(n_60)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_15),
.B(n_5),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_15),
.B(n_5),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_46),
.B(n_19),
.Y(n_70)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_49),
.B(n_31),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_47),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_50),
.B(n_65),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_18),
.C(n_27),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_53),
.B(n_1),
.C(n_2),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_41),
.A2(n_18),
.B1(n_27),
.B2(n_24),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_57),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_48),
.A2(n_23),
.B1(n_21),
.B2(n_24),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_61),
.A2(n_25),
.B1(n_17),
.B2(n_23),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_21),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_16),
.Y(n_77)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_64),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_47),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_41),
.B(n_33),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_70),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_73),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_49),
.A2(n_16),
.B1(n_23),
.B2(n_32),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_16),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_44),
.B(n_33),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_35),
.B(n_25),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_16),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_77),
.B(n_85),
.Y(n_105)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

O2A1O1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_62),
.A2(n_36),
.B(n_32),
.C(n_20),
.Y(n_81)
);

O2A1O1Ixp33_ASAP7_75t_SL g108 ( 
.A1(n_81),
.A2(n_55),
.B(n_56),
.C(n_54),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_82),
.A2(n_56),
.B1(n_63),
.B2(n_59),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_86),
.Y(n_100)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_84),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_52),
.B(n_17),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_60),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_L g106 ( 
.A1(n_87),
.A2(n_54),
.B1(n_64),
.B2(n_58),
.Y(n_106)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_55),
.C(n_66),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_50),
.B(n_6),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_93),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_53),
.B(n_1),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_2),
.Y(n_104)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_92),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_51),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_59),
.Y(n_94)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_51),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_3),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_65),
.B(n_6),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_97),
.Y(n_114)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_96),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_103),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_89),
.C(n_79),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_104),
.B(n_115),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_106),
.A2(n_76),
.B(n_92),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_108),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_80),
.A2(n_63),
.B1(n_58),
.B2(n_66),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_109),
.A2(n_110),
.B1(n_95),
.B2(n_88),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_80),
.A2(n_2),
.B1(n_3),
.B2(n_8),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_76),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_113),
.B(n_93),
.Y(n_119)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_111),
.Y(n_117)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_117),
.Y(n_137)
);

A2O1A1Ixp33_ASAP7_75t_SL g118 ( 
.A1(n_108),
.A2(n_106),
.B(n_87),
.C(n_81),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_118),
.A2(n_127),
.B(n_128),
.Y(n_136)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_119),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_91),
.Y(n_120)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_120),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_77),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_121),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_122),
.B(n_101),
.C(n_115),
.Y(n_134)
);

NOR3xp33_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_85),
.C(n_75),
.Y(n_123)
);

CKINVDCx12_ASAP7_75t_R g133 ( 
.A(n_123),
.Y(n_133)
);

AO22x1_ASAP7_75t_SL g126 ( 
.A1(n_108),
.A2(n_87),
.B1(n_78),
.B2(n_84),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_126),
.A2(n_129),
.B1(n_109),
.B2(n_103),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_100),
.B(n_86),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_112),
.Y(n_130)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_130),
.Y(n_143)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_112),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_131),
.A2(n_98),
.B(n_107),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_134),
.B(n_144),
.C(n_120),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_135),
.A2(n_140),
.B1(n_8),
.B2(n_11),
.Y(n_153)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_138),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_132),
.A2(n_82),
.B1(n_98),
.B2(n_107),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_132),
.A2(n_116),
.B(n_94),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_142),
.A2(n_118),
.B(n_96),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_122),
.B(n_116),
.C(n_114),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_139),
.B(n_121),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_146),
.B(n_149),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_147),
.B(n_134),
.C(n_136),
.Y(n_156)
);

AOI322xp5_ASAP7_75t_L g149 ( 
.A1(n_145),
.A2(n_125),
.A3(n_126),
.B1(n_118),
.B2(n_129),
.C1(n_127),
.C2(n_124),
.Y(n_149)
);

NOR2x1_ASAP7_75t_L g150 ( 
.A(n_141),
.B(n_126),
.Y(n_150)
);

OAI21x1_ASAP7_75t_L g161 ( 
.A1(n_150),
.A2(n_152),
.B(n_155),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_136),
.A2(n_118),
.B(n_99),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_151),
.B(n_142),
.Y(n_159)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_153),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g154 ( 
.A(n_133),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_154),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_144),
.B(n_11),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_156),
.B(n_152),
.C(n_135),
.Y(n_167)
);

NOR2xp67_ASAP7_75t_L g158 ( 
.A(n_147),
.B(n_140),
.Y(n_158)
);

NOR3xp33_ASAP7_75t_L g166 ( 
.A(n_158),
.B(n_150),
.C(n_148),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_159),
.B(n_148),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_156),
.B(n_151),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_163),
.B(n_166),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_164),
.B(n_165),
.Y(n_170)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_160),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_167),
.B(n_159),
.C(n_153),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_164),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_168),
.Y(n_172)
);

OAI21x1_ASAP7_75t_L g174 ( 
.A1(n_171),
.A2(n_162),
.B(n_138),
.Y(n_174)
);

OA21x2_ASAP7_75t_SL g173 ( 
.A1(n_169),
.A2(n_157),
.B(n_161),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_173),
.A2(n_174),
.B(n_171),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_172),
.B(n_170),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_175),
.A2(n_176),
.B(n_162),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_177),
.A2(n_143),
.B(n_137),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_143),
.Y(n_179)
);


endmodule