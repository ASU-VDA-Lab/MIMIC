module fake_ariane_885_n_1712 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1712);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1712;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_1083;
wire n_967;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_600;
wire n_481;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_727;
wire n_590;
wire n_699;
wire n_301;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_166;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_683;
wire n_236;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_679;
wire n_244;
wire n_1630;
wire n_220;
wire n_663;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_1067;
wire n_968;
wire n_1323;
wire n_1235;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1684;
wire n_1148;
wire n_1588;
wire n_1409;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1670;
wire n_1707;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_156;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_1102;
wire n_719;
wire n_263;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_484;
wire n_411;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_0),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_55),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_28),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_127),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_40),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_100),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_149),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_141),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_116),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_119),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_56),
.Y(n_166)
);

BUFx10_ASAP7_75t_L g167 ( 
.A(n_39),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_140),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_28),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_57),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_44),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_61),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_152),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_155),
.Y(n_174)
);

INVx2_ASAP7_75t_SL g175 ( 
.A(n_93),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_37),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_129),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_13),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_107),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_83),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_21),
.Y(n_181)
);

BUFx10_ASAP7_75t_L g182 ( 
.A(n_45),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_118),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_128),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_145),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_130),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_80),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_13),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_38),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_1),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_9),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_85),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_49),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_78),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_19),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_94),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_122),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_143),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_105),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_66),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_30),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_48),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_79),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_44),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_69),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_142),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_62),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_137),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_121),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_6),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_2),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_4),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_111),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_18),
.Y(n_214)
);

INVx2_ASAP7_75t_SL g215 ( 
.A(n_47),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_16),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_0),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_108),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_16),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_15),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_148),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_1),
.Y(n_222)
);

BUFx10_ASAP7_75t_L g223 ( 
.A(n_102),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_19),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_17),
.Y(n_225)
);

BUFx2_ASAP7_75t_L g226 ( 
.A(n_35),
.Y(n_226)
);

INVxp33_ASAP7_75t_SL g227 ( 
.A(n_77),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_2),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_64),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_97),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_4),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_50),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_114),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_9),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_150),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_131),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_76),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_136),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g239 ( 
.A(n_95),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_135),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_74),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_7),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_75),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_65),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_86),
.Y(n_245)
);

CKINVDCx14_ASAP7_75t_R g246 ( 
.A(n_146),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_104),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_60),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_33),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_117),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_49),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_24),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_144),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_91),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_151),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_53),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_6),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_17),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_40),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_46),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_31),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_98),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_20),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_92),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_22),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_125),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_8),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_31),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_153),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_14),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_20),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_18),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_37),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_81),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_22),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_132),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_7),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_126),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_89),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_133),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_52),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_106),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_134),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_21),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_139),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_147),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_27),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_10),
.Y(n_288)
);

BUFx3_ASAP7_75t_L g289 ( 
.A(n_42),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_42),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_14),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_8),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_59),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_99),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_10),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_109),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_36),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_27),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_110),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_124),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_96),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_84),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_51),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_120),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g305 ( 
.A(n_90),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_3),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_73),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_23),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_113),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_24),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_163),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_230),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_253),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_189),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_158),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_158),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_158),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_246),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_190),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_220),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_158),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_158),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_193),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_201),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_195),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_195),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_195),
.Y(n_327)
);

NOR2xp67_ASAP7_75t_L g328 ( 
.A(n_215),
.B(n_3),
.Y(n_328)
);

BUFx2_ASAP7_75t_L g329 ( 
.A(n_226),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_195),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_195),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_222),
.Y(n_332)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_191),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_204),
.Y(n_334)
);

NOR2xp67_ASAP7_75t_L g335 ( 
.A(n_215),
.B(n_5),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_222),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_210),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_306),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_224),
.Y(n_339)
);

CKINVDCx16_ASAP7_75t_R g340 ( 
.A(n_223),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_306),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_251),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_164),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_211),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_183),
.B(n_157),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_164),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_166),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_166),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_212),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_219),
.Y(n_350)
);

INVxp67_ASAP7_75t_SL g351 ( 
.A(n_217),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_238),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_238),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_176),
.Y(n_354)
);

INVxp67_ASAP7_75t_SL g355 ( 
.A(n_217),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_288),
.Y(n_356)
);

INVxp67_ASAP7_75t_SL g357 ( 
.A(n_289),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_223),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_225),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_180),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_181),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_223),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_188),
.Y(n_363)
);

CKINVDCx16_ASAP7_75t_R g364 ( 
.A(n_180),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_231),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_202),
.Y(n_366)
);

INVxp67_ASAP7_75t_SL g367 ( 
.A(n_289),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_214),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_232),
.Y(n_369)
);

INVxp67_ASAP7_75t_SL g370 ( 
.A(n_216),
.Y(n_370)
);

BUFx2_ASAP7_75t_SL g371 ( 
.A(n_175),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_228),
.Y(n_372)
);

INVxp67_ASAP7_75t_SL g373 ( 
.A(n_252),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_234),
.Y(n_374)
);

CKINVDCx16_ASAP7_75t_R g375 ( 
.A(n_167),
.Y(n_375)
);

CKINVDCx16_ASAP7_75t_R g376 ( 
.A(n_167),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_257),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_258),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_159),
.B(n_5),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_165),
.B(n_11),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_242),
.Y(n_381)
);

AND2x4_ASAP7_75t_L g382 ( 
.A(n_175),
.B(n_11),
.Y(n_382)
);

OA21x2_ASAP7_75t_L g383 ( 
.A1(n_315),
.A2(n_173),
.B(n_170),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_382),
.B(n_318),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_321),
.Y(n_385)
);

INVx3_ASAP7_75t_L g386 ( 
.A(n_321),
.Y(n_386)
);

INVx3_ASAP7_75t_L g387 ( 
.A(n_315),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_382),
.B(n_318),
.Y(n_388)
);

OA21x2_ASAP7_75t_L g389 ( 
.A1(n_316),
.A2(n_186),
.B(n_179),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_316),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_360),
.B(n_192),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_317),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_317),
.Y(n_393)
);

AND2x4_ASAP7_75t_L g394 ( 
.A(n_382),
.B(n_263),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_322),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_322),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_325),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_325),
.Y(n_398)
);

NAND2x1_ASAP7_75t_L g399 ( 
.A(n_382),
.B(n_161),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_326),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_326),
.Y(n_401)
);

AND2x6_ASAP7_75t_L g402 ( 
.A(n_343),
.B(n_161),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_327),
.Y(n_403)
);

NAND2xp33_ASAP7_75t_L g404 ( 
.A(n_380),
.B(n_161),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_327),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_330),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_351),
.B(n_265),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_330),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_331),
.Y(n_409)
);

AND2x4_ASAP7_75t_L g410 ( 
.A(n_360),
.B(n_277),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_331),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_343),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_329),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_346),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_346),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_347),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_329),
.A2(n_333),
.B1(n_340),
.B2(n_345),
.Y(n_417)
);

AND2x4_ASAP7_75t_L g418 ( 
.A(n_347),
.B(n_281),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_364),
.B(n_227),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_311),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_348),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_348),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_355),
.B(n_291),
.Y(n_423)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_352),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_352),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_353),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_353),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_332),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_357),
.B(n_367),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_332),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_312),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_336),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_336),
.Y(n_433)
);

BUFx2_ASAP7_75t_L g434 ( 
.A(n_314),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_338),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_338),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_371),
.B(n_194),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_341),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_341),
.Y(n_439)
);

AND2x4_ASAP7_75t_L g440 ( 
.A(n_370),
.B(n_297),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_364),
.B(n_310),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_354),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_354),
.Y(n_443)
);

INVx3_ASAP7_75t_L g444 ( 
.A(n_361),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_361),
.Y(n_445)
);

NAND2xp33_ASAP7_75t_SL g446 ( 
.A(n_358),
.B(n_156),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_313),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_387),
.Y(n_448)
);

BUFx3_ASAP7_75t_L g449 ( 
.A(n_444),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_387),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_429),
.B(n_371),
.Y(n_451)
);

NAND3xp33_ASAP7_75t_L g452 ( 
.A(n_444),
.B(n_379),
.C(n_335),
.Y(n_452)
);

AOI22xp33_ASAP7_75t_L g453 ( 
.A1(n_440),
.A2(n_328),
.B1(n_373),
.B2(n_362),
.Y(n_453)
);

BUFx4f_ASAP7_75t_L g454 ( 
.A(n_383),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_390),
.Y(n_455)
);

AND2x4_ASAP7_75t_L g456 ( 
.A(n_440),
.B(n_363),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_390),
.Y(n_457)
);

AOI22xp33_ASAP7_75t_L g458 ( 
.A1(n_440),
.A2(n_340),
.B1(n_284),
.B2(n_167),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_390),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_387),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g461 ( 
.A(n_442),
.B(n_363),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_392),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_387),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_434),
.B(n_319),
.Y(n_464)
);

OAI22xp33_ASAP7_75t_SL g465 ( 
.A1(n_417),
.A2(n_375),
.B1(n_376),
.B2(n_298),
.Y(n_465)
);

INVx2_ASAP7_75t_SL g466 ( 
.A(n_399),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_417),
.B(n_320),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_384),
.B(n_388),
.Y(n_468)
);

AND2x6_ASAP7_75t_L g469 ( 
.A(n_394),
.B(n_441),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_441),
.A2(n_156),
.B1(n_160),
.B2(n_169),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_392),
.Y(n_471)
);

BUFx10_ASAP7_75t_L g472 ( 
.A(n_394),
.Y(n_472)
);

BUFx3_ASAP7_75t_L g473 ( 
.A(n_444),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_392),
.Y(n_474)
);

INVx4_ASAP7_75t_SL g475 ( 
.A(n_402),
.Y(n_475)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_415),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_387),
.Y(n_477)
);

INVx3_ASAP7_75t_L g478 ( 
.A(n_415),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_429),
.B(n_437),
.Y(n_479)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_415),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_393),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_393),
.Y(n_482)
);

BUFx10_ASAP7_75t_L g483 ( 
.A(n_394),
.Y(n_483)
);

BUFx4f_ASAP7_75t_L g484 ( 
.A(n_383),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_384),
.B(n_388),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_393),
.Y(n_486)
);

AOI22xp33_ASAP7_75t_L g487 ( 
.A1(n_440),
.A2(n_182),
.B1(n_381),
.B2(n_350),
.Y(n_487)
);

AO21x2_ASAP7_75t_L g488 ( 
.A1(n_419),
.A2(n_199),
.B(n_197),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_387),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_400),
.Y(n_490)
);

BUFx10_ASAP7_75t_L g491 ( 
.A(n_394),
.Y(n_491)
);

BUFx4f_ASAP7_75t_L g492 ( 
.A(n_383),
.Y(n_492)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_415),
.Y(n_493)
);

BUFx3_ASAP7_75t_L g494 ( 
.A(n_444),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_400),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_437),
.B(n_323),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_434),
.B(n_324),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_395),
.Y(n_498)
);

BUFx6f_ASAP7_75t_L g499 ( 
.A(n_415),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_419),
.B(n_334),
.Y(n_500)
);

AND2x6_ASAP7_75t_L g501 ( 
.A(n_394),
.B(n_161),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_SL g502 ( 
.A(n_420),
.B(n_337),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_395),
.Y(n_503)
);

BUFx3_ASAP7_75t_L g504 ( 
.A(n_444),
.Y(n_504)
);

NAND3xp33_ASAP7_75t_L g505 ( 
.A(n_444),
.B(n_349),
.C(n_344),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_400),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_405),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_394),
.B(n_359),
.Y(n_508)
);

AOI22xp33_ASAP7_75t_L g509 ( 
.A1(n_440),
.A2(n_182),
.B1(n_369),
.B2(n_374),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_405),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_440),
.B(n_365),
.Y(n_511)
);

INVx3_ASAP7_75t_L g512 ( 
.A(n_415),
.Y(n_512)
);

AOI22xp33_ASAP7_75t_L g513 ( 
.A1(n_410),
.A2(n_182),
.B1(n_377),
.B2(n_372),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_441),
.A2(n_275),
.B1(n_171),
.B2(n_160),
.Y(n_514)
);

OR2x6_ASAP7_75t_L g515 ( 
.A(n_399),
.B(n_366),
.Y(n_515)
);

INVx3_ASAP7_75t_L g516 ( 
.A(n_415),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_395),
.Y(n_517)
);

BUFx10_ASAP7_75t_L g518 ( 
.A(n_420),
.Y(n_518)
);

INVx2_ASAP7_75t_SL g519 ( 
.A(n_399),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_415),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_442),
.B(n_366),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_434),
.B(n_368),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_413),
.B(n_368),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_442),
.B(n_372),
.Y(n_524)
);

INVx3_ASAP7_75t_L g525 ( 
.A(n_415),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_413),
.B(n_377),
.Y(n_526)
);

OR2x6_ASAP7_75t_L g527 ( 
.A(n_407),
.B(n_378),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_407),
.B(n_162),
.Y(n_528)
);

INVx4_ASAP7_75t_L g529 ( 
.A(n_389),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_395),
.Y(n_530)
);

INVx3_ASAP7_75t_L g531 ( 
.A(n_424),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_397),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_397),
.Y(n_533)
);

AOI22xp33_ASAP7_75t_L g534 ( 
.A1(n_410),
.A2(n_378),
.B1(n_239),
.B2(n_305),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_424),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_405),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_418),
.B(n_169),
.Y(n_537)
);

OR2x2_ASAP7_75t_L g538 ( 
.A(n_407),
.B(n_171),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_397),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_397),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_424),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_424),
.Y(n_542)
);

INVx4_ASAP7_75t_L g543 ( 
.A(n_389),
.Y(n_543)
);

INVx1_ASAP7_75t_SL g544 ( 
.A(n_431),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_398),
.Y(n_545)
);

AOI22xp33_ASAP7_75t_L g546 ( 
.A1(n_410),
.A2(n_247),
.B1(n_259),
.B2(n_261),
.Y(n_546)
);

INVx1_ASAP7_75t_SL g547 ( 
.A(n_431),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_423),
.B(n_162),
.Y(n_548)
);

INVx5_ASAP7_75t_L g549 ( 
.A(n_402),
.Y(n_549)
);

BUFx4f_ASAP7_75t_L g550 ( 
.A(n_383),
.Y(n_550)
);

BUFx3_ASAP7_75t_L g551 ( 
.A(n_410),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_424),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_423),
.B(n_168),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_424),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_414),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_414),
.Y(n_556)
);

INVx3_ASAP7_75t_L g557 ( 
.A(n_428),
.Y(n_557)
);

BUFx3_ASAP7_75t_L g558 ( 
.A(n_410),
.Y(n_558)
);

INVx5_ASAP7_75t_L g559 ( 
.A(n_402),
.Y(n_559)
);

XOR2x2_ASAP7_75t_SL g560 ( 
.A(n_446),
.B(n_339),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_398),
.Y(n_561)
);

BUFx3_ASAP7_75t_L g562 ( 
.A(n_443),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_447),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_414),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_398),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g566 ( 
.A(n_418),
.B(n_178),
.Y(n_566)
);

AO22x2_ASAP7_75t_L g567 ( 
.A1(n_423),
.A2(n_296),
.B1(n_285),
.B2(n_309),
.Y(n_567)
);

BUFx4f_ASAP7_75t_L g568 ( 
.A(n_383),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_414),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_398),
.Y(n_570)
);

XOR2xp5_ASAP7_75t_L g571 ( 
.A(n_447),
.B(n_342),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_418),
.B(n_443),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_401),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_401),
.Y(n_574)
);

BUFx8_ASAP7_75t_SL g575 ( 
.A(n_410),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_412),
.B(n_168),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_412),
.B(n_172),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_416),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_401),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_446),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_416),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_401),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_391),
.B(n_209),
.Y(n_583)
);

OR2x6_ASAP7_75t_L g584 ( 
.A(n_418),
.B(n_221),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_403),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_412),
.B(n_172),
.Y(n_586)
);

INVx2_ASAP7_75t_SL g587 ( 
.A(n_389),
.Y(n_587)
);

INVx4_ASAP7_75t_L g588 ( 
.A(n_389),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_416),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_403),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_418),
.Y(n_591)
);

AOI22xp33_ASAP7_75t_L g592 ( 
.A1(n_418),
.A2(n_271),
.B1(n_270),
.B2(n_249),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_416),
.Y(n_593)
);

AOI22xp33_ASAP7_75t_L g594 ( 
.A1(n_383),
.A2(n_272),
.B1(n_268),
.B2(n_260),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_425),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_496),
.B(n_391),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_562),
.Y(n_597)
);

AOI22xp33_ASAP7_75t_L g598 ( 
.A1(n_567),
.A2(n_389),
.B1(n_383),
.B2(n_445),
.Y(n_598)
);

OR2x2_ASAP7_75t_L g599 ( 
.A(n_544),
.B(n_443),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_479),
.B(n_443),
.Y(n_600)
);

BUFx3_ASAP7_75t_L g601 ( 
.A(n_449),
.Y(n_601)
);

INVx2_ASAP7_75t_SL g602 ( 
.A(n_518),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_562),
.Y(n_603)
);

OR2x6_ASAP7_75t_L g604 ( 
.A(n_527),
.B(n_456),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_451),
.B(n_445),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_522),
.B(n_445),
.Y(n_606)
);

INVx3_ASAP7_75t_L g607 ( 
.A(n_472),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_472),
.B(n_445),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_541),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_SL g610 ( 
.A(n_502),
.B(n_356),
.Y(n_610)
);

AOI22xp5_ASAP7_75t_L g611 ( 
.A1(n_469),
.A2(n_404),
.B1(n_421),
.B2(n_422),
.Y(n_611)
);

AOI22xp5_ASAP7_75t_L g612 ( 
.A1(n_469),
.A2(n_404),
.B1(n_421),
.B2(n_422),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_468),
.B(n_421),
.Y(n_613)
);

INVx2_ASAP7_75t_SL g614 ( 
.A(n_518),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_541),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_485),
.B(n_456),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_456),
.B(n_422),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_456),
.B(n_426),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_542),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_498),
.Y(n_620)
);

INVx3_ASAP7_75t_L g621 ( 
.A(n_472),
.Y(n_621)
);

AOI22xp33_ASAP7_75t_L g622 ( 
.A1(n_567),
.A2(n_389),
.B1(n_425),
.B2(n_426),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_542),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_523),
.B(n_426),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_500),
.B(n_427),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_498),
.Y(n_626)
);

NAND2xp33_ASAP7_75t_L g627 ( 
.A(n_469),
.B(n_174),
.Y(n_627)
);

NOR3xp33_ASAP7_75t_L g628 ( 
.A(n_464),
.B(n_292),
.C(n_303),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_472),
.B(n_428),
.Y(n_629)
);

NAND2xp33_ASAP7_75t_SL g630 ( 
.A(n_511),
.B(n_178),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_552),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_526),
.B(n_427),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_503),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_508),
.B(n_427),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_503),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_591),
.B(n_433),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_466),
.B(n_433),
.Y(n_637)
);

NOR2xp67_ASAP7_75t_L g638 ( 
.A(n_505),
.B(n_433),
.Y(n_638)
);

INVx2_ASAP7_75t_SL g639 ( 
.A(n_518),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_552),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_591),
.B(n_438),
.Y(n_641)
);

INVxp67_ASAP7_75t_L g642 ( 
.A(n_571),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_517),
.Y(n_643)
);

NAND2xp33_ASAP7_75t_L g644 ( 
.A(n_469),
.B(n_174),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_466),
.B(n_438),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_483),
.B(n_428),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_505),
.B(n_438),
.Y(n_647)
);

NOR2xp67_ASAP7_75t_L g648 ( 
.A(n_497),
.B(n_425),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_519),
.B(n_425),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_528),
.B(n_267),
.Y(n_650)
);

OAI22xp5_ASAP7_75t_L g651 ( 
.A1(n_452),
.A2(n_290),
.B1(n_273),
.B2(n_275),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_519),
.B(n_430),
.Y(n_652)
);

AND2x2_ASAP7_75t_SL g653 ( 
.A(n_594),
.B(n_229),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_469),
.B(n_430),
.Y(n_654)
);

INVxp67_ASAP7_75t_L g655 ( 
.A(n_571),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_517),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_527),
.B(n_439),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_554),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_554),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_572),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_483),
.B(n_428),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_469),
.B(n_430),
.Y(n_662)
);

NAND2xp33_ASAP7_75t_L g663 ( 
.A(n_469),
.B(n_177),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_483),
.B(n_428),
.Y(n_664)
);

OAI22xp5_ASAP7_75t_L g665 ( 
.A1(n_452),
.A2(n_292),
.B1(n_273),
.B2(n_287),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_572),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_483),
.B(n_428),
.Y(n_667)
);

BUFx6f_ASAP7_75t_SL g668 ( 
.A(n_518),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_530),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_461),
.B(n_430),
.Y(n_670)
);

NAND2x1p5_ASAP7_75t_L g671 ( 
.A(n_551),
.B(n_428),
.Y(n_671)
);

OAI221xp5_ASAP7_75t_L g672 ( 
.A1(n_487),
.A2(n_295),
.B1(n_287),
.B2(n_290),
.C(n_298),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_530),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_532),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_461),
.B(n_436),
.Y(n_675)
);

AOI21xp5_ASAP7_75t_L g676 ( 
.A1(n_454),
.A2(n_439),
.B(n_436),
.Y(n_676)
);

NAND3xp33_ASAP7_75t_L g677 ( 
.A(n_509),
.B(n_295),
.C(n_303),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_583),
.B(n_436),
.Y(n_678)
);

AND2x6_ASAP7_75t_SL g679 ( 
.A(n_563),
.B(n_308),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_527),
.B(n_436),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_527),
.B(n_439),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_532),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_491),
.B(n_428),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_533),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_455),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_527),
.B(n_439),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_548),
.B(n_553),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_531),
.B(n_428),
.Y(n_688)
);

NAND2xp33_ASAP7_75t_L g689 ( 
.A(n_501),
.B(n_499),
.Y(n_689)
);

O2A1O1Ixp33_ASAP7_75t_L g690 ( 
.A1(n_521),
.A2(n_409),
.B(n_408),
.C(n_403),
.Y(n_690)
);

AOI22xp5_ASAP7_75t_L g691 ( 
.A1(n_515),
.A2(n_185),
.B1(n_307),
.B2(n_304),
.Y(n_691)
);

NOR3xp33_ASAP7_75t_L g692 ( 
.A(n_563),
.B(n_308),
.C(n_250),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_470),
.B(n_432),
.Y(n_693)
);

AND2x4_ASAP7_75t_L g694 ( 
.A(n_551),
.B(n_432),
.Y(n_694)
);

AOI22xp5_ASAP7_75t_L g695 ( 
.A1(n_515),
.A2(n_184),
.B1(n_307),
.B2(n_304),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_491),
.B(n_432),
.Y(n_696)
);

INVxp67_ASAP7_75t_L g697 ( 
.A(n_547),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_531),
.B(n_535),
.Y(n_698)
);

AOI22xp5_ASAP7_75t_L g699 ( 
.A1(n_515),
.A2(n_187),
.B1(n_185),
.B2(n_184),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_470),
.B(n_432),
.Y(n_700)
);

INVx2_ASAP7_75t_SL g701 ( 
.A(n_538),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_531),
.B(n_432),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_535),
.B(n_432),
.Y(n_703)
);

NOR2xp67_ASAP7_75t_L g704 ( 
.A(n_514),
.B(n_386),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_535),
.B(n_432),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_491),
.B(n_432),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_488),
.B(n_432),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_533),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_514),
.B(n_435),
.Y(n_709)
);

A2O1A1Ixp33_ASAP7_75t_L g710 ( 
.A1(n_454),
.A2(n_568),
.B(n_550),
.C(n_484),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_491),
.B(n_435),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_488),
.B(n_435),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_539),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_454),
.B(n_435),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_488),
.B(n_435),
.Y(n_715)
);

OAI22xp5_ASAP7_75t_L g716 ( 
.A1(n_584),
.A2(n_280),
.B1(n_187),
.B2(n_177),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_539),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_551),
.B(n_435),
.Y(n_718)
);

INVxp67_ASAP7_75t_L g719 ( 
.A(n_538),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_558),
.B(n_576),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_540),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_558),
.B(n_435),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_455),
.Y(n_723)
);

AOI22xp33_ASAP7_75t_L g724 ( 
.A1(n_567),
.A2(n_435),
.B1(n_409),
.B2(n_408),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_540),
.Y(n_725)
);

NAND2xp33_ASAP7_75t_L g726 ( 
.A(n_501),
.B(n_276),
.Y(n_726)
);

BUFx6f_ASAP7_75t_L g727 ( 
.A(n_499),
.Y(n_727)
);

AOI221xp5_ASAP7_75t_L g728 ( 
.A1(n_465),
.A2(n_283),
.B1(n_302),
.B2(n_276),
.C(n_300),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_558),
.B(n_435),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_545),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_545),
.Y(n_731)
);

CKINVDCx20_ASAP7_75t_R g732 ( 
.A(n_560),
.Y(n_732)
);

BUFx6f_ASAP7_75t_L g733 ( 
.A(n_499),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_484),
.B(n_279),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_577),
.B(n_279),
.Y(n_735)
);

NAND2x1_ASAP7_75t_L g736 ( 
.A(n_515),
.B(n_402),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_586),
.B(n_280),
.Y(n_737)
);

INVxp67_ASAP7_75t_SL g738 ( 
.A(n_587),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_515),
.B(n_283),
.Y(n_739)
);

INVx3_ASAP7_75t_L g740 ( 
.A(n_449),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_561),
.Y(n_741)
);

BUFx6f_ASAP7_75t_L g742 ( 
.A(n_499),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_453),
.B(n_403),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_537),
.B(n_286),
.Y(n_744)
);

INVxp67_ASAP7_75t_L g745 ( 
.A(n_575),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_561),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_537),
.B(n_286),
.Y(n_747)
);

INVxp67_ASAP7_75t_L g748 ( 
.A(n_467),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_565),
.Y(n_749)
);

AOI22xp5_ASAP7_75t_L g750 ( 
.A1(n_567),
.A2(n_302),
.B1(n_299),
.B2(n_300),
.Y(n_750)
);

OAI22xp33_ASAP7_75t_L g751 ( 
.A1(n_580),
.A2(n_299),
.B1(n_294),
.B2(n_256),
.Y(n_751)
);

OR2x2_ASAP7_75t_L g752 ( 
.A(n_467),
.B(n_386),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_565),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_457),
.Y(n_754)
);

AOI22xp5_ASAP7_75t_L g755 ( 
.A1(n_584),
.A2(n_294),
.B1(n_274),
.B2(n_282),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_473),
.B(n_266),
.Y(n_756)
);

INVx1_ASAP7_75t_SL g757 ( 
.A(n_580),
.Y(n_757)
);

OAI22xp5_ASAP7_75t_L g758 ( 
.A1(n_584),
.A2(n_293),
.B1(n_301),
.B2(n_254),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_473),
.B(n_494),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_566),
.B(n_386),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_566),
.B(n_386),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_494),
.B(n_386),
.Y(n_762)
);

AOI221xp5_ASAP7_75t_L g763 ( 
.A1(n_465),
.A2(n_241),
.B1(n_208),
.B2(n_213),
.C(n_196),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_459),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_504),
.B(n_524),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_504),
.B(n_386),
.Y(n_766)
);

A2O1A1Ixp33_ASAP7_75t_L g767 ( 
.A1(n_625),
.A2(n_484),
.B(n_550),
.C(n_492),
.Y(n_767)
);

BUFx6f_ASAP7_75t_L g768 ( 
.A(n_727),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_685),
.Y(n_769)
);

OAI22xp5_ASAP7_75t_L g770 ( 
.A1(n_625),
.A2(n_584),
.B1(n_550),
.B2(n_568),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_596),
.B(n_534),
.Y(n_771)
);

INVx2_ASAP7_75t_SL g772 ( 
.A(n_599),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_687),
.B(n_458),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_719),
.B(n_513),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_668),
.Y(n_775)
);

BUFx6f_ASAP7_75t_L g776 ( 
.A(n_727),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_723),
.Y(n_777)
);

OAI22xp33_ASAP7_75t_L g778 ( 
.A1(n_616),
.A2(n_584),
.B1(n_560),
.B2(n_471),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_SL g779 ( 
.A(n_610),
.B(n_529),
.Y(n_779)
);

AOI21xp5_ASAP7_75t_L g780 ( 
.A1(n_714),
.A2(n_492),
.B(n_568),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_607),
.B(n_492),
.Y(n_781)
);

BUFx24_ASAP7_75t_L g782 ( 
.A(n_668),
.Y(n_782)
);

AOI21x1_ASAP7_75t_L g783 ( 
.A1(n_714),
.A2(n_506),
.B(n_459),
.Y(n_783)
);

AOI21xp5_ASAP7_75t_L g784 ( 
.A1(n_600),
.A2(n_587),
.B(n_460),
.Y(n_784)
);

OAI22xp5_ASAP7_75t_L g785 ( 
.A1(n_636),
.A2(n_641),
.B1(n_687),
.B2(n_604),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_607),
.B(n_499),
.Y(n_786)
);

AO21x1_ASAP7_75t_L g787 ( 
.A1(n_647),
.A2(n_543),
.B(n_529),
.Y(n_787)
);

AND2x4_ASAP7_75t_L g788 ( 
.A(n_604),
.B(n_475),
.Y(n_788)
);

AOI21xp5_ASAP7_75t_L g789 ( 
.A1(n_738),
.A2(n_448),
.B(n_450),
.Y(n_789)
);

OAI22xp5_ASAP7_75t_L g790 ( 
.A1(n_636),
.A2(n_592),
.B1(n_495),
.B2(n_490),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_596),
.B(n_529),
.Y(n_791)
);

BUFx2_ASAP7_75t_L g792 ( 
.A(n_697),
.Y(n_792)
);

INVx4_ASAP7_75t_L g793 ( 
.A(n_604),
.Y(n_793)
);

OAI21xp5_ASAP7_75t_L g794 ( 
.A1(n_676),
.A2(n_543),
.B(n_529),
.Y(n_794)
);

AOI21xp5_ASAP7_75t_L g795 ( 
.A1(n_698),
.A2(n_448),
.B(n_450),
.Y(n_795)
);

OAI21xp33_ASAP7_75t_L g796 ( 
.A1(n_641),
.A2(n_546),
.B(n_462),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_621),
.B(n_460),
.Y(n_797)
);

AO21x1_ASAP7_75t_L g798 ( 
.A1(n_647),
.A2(n_715),
.B(n_734),
.Y(n_798)
);

INVxp67_ASAP7_75t_L g799 ( 
.A(n_657),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_634),
.B(n_555),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_634),
.B(n_555),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_621),
.B(n_463),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_754),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_757),
.B(n_543),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_624),
.B(n_556),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_632),
.B(n_556),
.Y(n_806)
);

INVxp67_ASAP7_75t_L g807 ( 
.A(n_657),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_679),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_606),
.B(n_564),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_701),
.B(n_543),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_613),
.B(n_564),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_764),
.Y(n_812)
);

OAI21xp5_ASAP7_75t_L g813 ( 
.A1(n_688),
.A2(n_588),
.B(n_462),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_702),
.A2(n_489),
.B(n_463),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_703),
.A2(n_489),
.B(n_477),
.Y(n_815)
);

OAI21xp5_ASAP7_75t_L g816 ( 
.A1(n_705),
.A2(n_615),
.B(n_609),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_660),
.B(n_569),
.Y(n_817)
);

AOI21xp5_ASAP7_75t_L g818 ( 
.A1(n_678),
.A2(n_477),
.B(n_476),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_666),
.B(n_569),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_765),
.A2(n_520),
.B(n_476),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_619),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_623),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_686),
.B(n_617),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_734),
.A2(n_520),
.B(n_476),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_710),
.A2(n_520),
.B(n_478),
.Y(n_825)
);

OAI21xp5_ASAP7_75t_L g826 ( 
.A1(n_631),
.A2(n_588),
.B(n_536),
.Y(n_826)
);

AOI21x1_ASAP7_75t_L g827 ( 
.A1(n_707),
.A2(n_495),
.B(n_471),
.Y(n_827)
);

INVx2_ASAP7_75t_SL g828 ( 
.A(n_752),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_710),
.A2(n_478),
.B(n_480),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_686),
.B(n_578),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_626),
.Y(n_831)
);

AO21x1_ASAP7_75t_L g832 ( 
.A1(n_715),
.A2(n_588),
.B(n_490),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_608),
.A2(n_605),
.B(n_720),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_618),
.B(n_578),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_640),
.Y(n_835)
);

INVx11_ASAP7_75t_L g836 ( 
.A(n_745),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_743),
.B(n_581),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_739),
.B(n_581),
.Y(n_838)
);

NOR3xp33_ASAP7_75t_L g839 ( 
.A(n_672),
.B(n_482),
.C(n_510),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_602),
.B(n_614),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_608),
.A2(n_525),
.B(n_478),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_650),
.B(n_744),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_762),
.A2(n_480),
.B(n_493),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_766),
.A2(n_480),
.B(n_493),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_650),
.B(n_588),
.Y(n_845)
);

AOI33xp33_ASAP7_75t_L g846 ( 
.A1(n_728),
.A2(n_536),
.A3(n_474),
.B1(n_481),
.B2(n_482),
.B3(n_486),
.Y(n_846)
);

INVx4_ASAP7_75t_L g847 ( 
.A(n_694),
.Y(n_847)
);

INVx3_ASAP7_75t_L g848 ( 
.A(n_601),
.Y(n_848)
);

O2A1O1Ixp33_ASAP7_75t_L g849 ( 
.A1(n_651),
.A2(n_595),
.B(n_593),
.C(n_589),
.Y(n_849)
);

AOI21xp33_ASAP7_75t_L g850 ( 
.A1(n_653),
.A2(n_507),
.B(n_510),
.Y(n_850)
);

O2A1O1Ixp33_ASAP7_75t_L g851 ( 
.A1(n_665),
.A2(n_595),
.B(n_593),
.C(n_589),
.Y(n_851)
);

AOI21x1_ASAP7_75t_L g852 ( 
.A1(n_712),
.A2(n_486),
.B(n_474),
.Y(n_852)
);

OAI21xp5_ASAP7_75t_L g853 ( 
.A1(n_658),
.A2(n_507),
.B(n_481),
.Y(n_853)
);

NAND3xp33_ASAP7_75t_SL g854 ( 
.A(n_692),
.B(n_506),
.C(n_200),
.Y(n_854)
);

INVx3_ASAP7_75t_L g855 ( 
.A(n_601),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_629),
.A2(n_493),
.B(n_512),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_747),
.B(n_512),
.Y(n_857)
);

A2O1A1Ixp33_ASAP7_75t_L g858 ( 
.A1(n_739),
.A2(n_750),
.B(n_756),
.C(n_654),
.Y(n_858)
);

AO21x1_ASAP7_75t_L g859 ( 
.A1(n_690),
.A2(n_590),
.B(n_585),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_639),
.B(n_501),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_629),
.A2(n_512),
.B(n_516),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_637),
.B(n_501),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_645),
.B(n_501),
.Y(n_863)
);

A2O1A1Ixp33_ASAP7_75t_L g864 ( 
.A1(n_756),
.A2(n_590),
.B(n_585),
.C(n_582),
.Y(n_864)
);

OAI21xp5_ASAP7_75t_L g865 ( 
.A1(n_659),
.A2(n_525),
.B(n_516),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_693),
.B(n_501),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_748),
.B(n_642),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_700),
.B(n_501),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_670),
.Y(n_869)
);

OAI21xp5_ASAP7_75t_L g870 ( 
.A1(n_662),
.A2(n_525),
.B(n_557),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_755),
.B(n_516),
.Y(n_871)
);

AOI22xp5_ASAP7_75t_L g872 ( 
.A1(n_653),
.A2(n_557),
.B1(n_579),
.B2(n_574),
.Y(n_872)
);

NAND2x1p5_ASAP7_75t_L g873 ( 
.A(n_694),
.B(n_557),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_709),
.B(n_570),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_633),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_646),
.A2(n_582),
.B(n_579),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_677),
.B(n_570),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_655),
.B(n_573),
.Y(n_878)
);

BUFx6f_ASAP7_75t_L g879 ( 
.A(n_727),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_646),
.A2(n_574),
.B(n_573),
.Y(n_880)
);

INVx3_ASAP7_75t_L g881 ( 
.A(n_671),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_661),
.A2(n_248),
.B(n_198),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_635),
.Y(n_883)
);

INVx5_ASAP7_75t_L g884 ( 
.A(n_727),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_661),
.A2(n_255),
.B(n_205),
.Y(n_885)
);

AOI21x1_ASAP7_75t_L g886 ( 
.A1(n_649),
.A2(n_409),
.B(n_408),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_735),
.B(n_408),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_675),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_680),
.Y(n_889)
);

AO21x1_ASAP7_75t_L g890 ( 
.A1(n_758),
.A2(n_409),
.B(n_385),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_635),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_664),
.A2(n_245),
.B(n_206),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_682),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_664),
.A2(n_262),
.B(n_207),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_681),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_667),
.A2(n_264),
.B(n_218),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_733),
.B(n_411),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_667),
.A2(n_269),
.B(n_233),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_733),
.B(n_411),
.Y(n_899)
);

AND2x4_ASAP7_75t_L g900 ( 
.A(n_704),
.B(n_475),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_737),
.B(n_385),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_759),
.B(n_597),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_759),
.B(n_385),
.Y(n_903)
);

AOI21x1_ASAP7_75t_L g904 ( 
.A1(n_652),
.A2(n_385),
.B(n_396),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_683),
.A2(n_236),
.B(n_240),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_597),
.B(n_235),
.Y(n_906)
);

O2A1O1Ixp33_ASAP7_75t_L g907 ( 
.A1(n_760),
.A2(n_12),
.B(n_15),
.C(n_23),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_683),
.A2(n_237),
.B(n_243),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_603),
.B(n_12),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_L g910 ( 
.A(n_691),
.B(n_25),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_603),
.B(n_25),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_696),
.A2(n_559),
.B(n_549),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_682),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_628),
.B(n_475),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_706),
.A2(n_711),
.B(n_718),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_684),
.Y(n_916)
);

INVx11_ASAP7_75t_L g917 ( 
.A(n_648),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_706),
.A2(n_559),
.B(n_549),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_711),
.A2(n_729),
.B(n_722),
.Y(n_919)
);

OAI21xp5_ASAP7_75t_L g920 ( 
.A1(n_638),
.A2(n_402),
.B(n_549),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_L g921 ( 
.A(n_695),
.B(n_26),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_761),
.A2(n_559),
.B(n_549),
.Y(n_922)
);

OAI21xp5_ASAP7_75t_L g923 ( 
.A1(n_611),
.A2(n_402),
.B(n_549),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_740),
.B(n_26),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_684),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_627),
.A2(n_663),
.B(n_644),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_733),
.B(n_396),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_708),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_708),
.A2(n_559),
.B(n_396),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_717),
.A2(n_559),
.B(n_396),
.Y(n_930)
);

OAI21xp5_ASAP7_75t_L g931 ( 
.A1(n_612),
.A2(n_402),
.B(n_475),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_SL g932 ( 
.A(n_733),
.B(n_411),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_740),
.B(n_29),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_732),
.B(n_29),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_724),
.B(n_30),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_724),
.B(n_32),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_751),
.B(n_32),
.Y(n_937)
);

OR2x6_ASAP7_75t_SL g938 ( 
.A(n_716),
.B(n_33),
.Y(n_938)
);

OAI22xp5_ASAP7_75t_L g939 ( 
.A1(n_671),
.A2(n_411),
.B1(n_406),
.B2(n_396),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_699),
.B(n_34),
.Y(n_940)
);

AND2x4_ASAP7_75t_L g941 ( 
.A(n_742),
.B(n_402),
.Y(n_941)
);

AND2x4_ASAP7_75t_L g942 ( 
.A(n_742),
.B(n_402),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_622),
.B(n_721),
.Y(n_943)
);

OAI22xp5_ASAP7_75t_L g944 ( 
.A1(n_742),
.A2(n_411),
.B1(n_406),
.B2(n_396),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_717),
.A2(n_411),
.B(n_406),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_SL g946 ( 
.A(n_742),
.B(n_411),
.Y(n_946)
);

OAI21xp5_ASAP7_75t_L g947 ( 
.A1(n_721),
.A2(n_402),
.B(n_406),
.Y(n_947)
);

AO21x1_ASAP7_75t_L g948 ( 
.A1(n_630),
.A2(n_411),
.B(n_406),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_622),
.B(n_34),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_725),
.B(n_35),
.Y(n_950)
);

INVx3_ASAP7_75t_L g951 ( 
.A(n_736),
.Y(n_951)
);

INVx3_ASAP7_75t_L g952 ( 
.A(n_788),
.Y(n_952)
);

INVxp67_ASAP7_75t_L g953 ( 
.A(n_792),
.Y(n_953)
);

HB1xp67_ASAP7_75t_L g954 ( 
.A(n_772),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_869),
.B(n_725),
.Y(n_955)
);

A2O1A1Ixp33_ASAP7_75t_L g956 ( 
.A1(n_842),
.A2(n_763),
.B(n_730),
.C(n_731),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_769),
.Y(n_957)
);

OA21x2_ASAP7_75t_L g958 ( 
.A1(n_832),
.A2(n_598),
.B(n_730),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_777),
.Y(n_959)
);

O2A1O1Ixp33_ASAP7_75t_L g960 ( 
.A1(n_785),
.A2(n_842),
.B(n_921),
.C(n_910),
.Y(n_960)
);

NOR2x1_ASAP7_75t_L g961 ( 
.A(n_848),
.B(n_689),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_774),
.B(n_598),
.Y(n_962)
);

INVx4_ASAP7_75t_L g963 ( 
.A(n_788),
.Y(n_963)
);

NAND2x1p5_ASAP7_75t_L g964 ( 
.A(n_793),
.B(n_731),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_800),
.A2(n_741),
.B(n_749),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_782),
.Y(n_966)
);

NAND3xp33_ASAP7_75t_SL g967 ( 
.A(n_773),
.B(n_673),
.C(n_746),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_888),
.B(n_741),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_L g969 ( 
.A(n_773),
.B(n_771),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_R g970 ( 
.A(n_775),
.B(n_726),
.Y(n_970)
);

AOI21x1_ASAP7_75t_L g971 ( 
.A1(n_827),
.A2(n_852),
.B(n_886),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_803),
.Y(n_972)
);

OAI22xp5_ASAP7_75t_L g973 ( 
.A1(n_823),
.A2(n_753),
.B1(n_713),
.B2(n_674),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_799),
.B(n_669),
.Y(n_974)
);

A2O1A1Ixp33_ASAP7_75t_L g975 ( 
.A1(n_910),
.A2(n_643),
.B(n_620),
.C(n_656),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_799),
.B(n_36),
.Y(n_976)
);

BUFx2_ASAP7_75t_L g977 ( 
.A(n_867),
.Y(n_977)
);

INVx3_ASAP7_75t_L g978 ( 
.A(n_793),
.Y(n_978)
);

BUFx2_ASAP7_75t_L g979 ( 
.A(n_878),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_801),
.A2(n_278),
.B(n_244),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_807),
.B(n_38),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_SL g982 ( 
.A(n_807),
.B(n_411),
.Y(n_982)
);

AOI221xp5_ASAP7_75t_L g983 ( 
.A1(n_921),
.A2(n_396),
.B1(n_406),
.B2(n_278),
.C(n_244),
.Y(n_983)
);

INVx3_ASAP7_75t_L g984 ( 
.A(n_847),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_L g985 ( 
.A(n_778),
.B(n_39),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_791),
.A2(n_278),
.B(n_244),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_812),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_889),
.B(n_41),
.Y(n_988)
);

OAI22xp5_ASAP7_75t_L g989 ( 
.A1(n_791),
.A2(n_406),
.B1(n_396),
.B2(n_278),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_767),
.A2(n_278),
.B(n_244),
.Y(n_990)
);

AO21x1_ASAP7_75t_L g991 ( 
.A1(n_845),
.A2(n_244),
.B(n_203),
.Y(n_991)
);

BUFx3_ASAP7_75t_L g992 ( 
.A(n_934),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_SL g993 ( 
.A(n_847),
.B(n_406),
.Y(n_993)
);

BUFx2_ASAP7_75t_L g994 ( 
.A(n_828),
.Y(n_994)
);

HB1xp67_ASAP7_75t_L g995 ( 
.A(n_873),
.Y(n_995)
);

AO21x1_ASAP7_75t_L g996 ( 
.A1(n_845),
.A2(n_203),
.B(n_161),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_895),
.B(n_830),
.Y(n_997)
);

CKINVDCx11_ASAP7_75t_R g998 ( 
.A(n_938),
.Y(n_998)
);

BUFx8_ASAP7_75t_L g999 ( 
.A(n_914),
.Y(n_999)
);

BUFx3_ASAP7_75t_L g1000 ( 
.A(n_848),
.Y(n_1000)
);

AND2x2_ASAP7_75t_L g1001 ( 
.A(n_808),
.B(n_41),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_770),
.A2(n_203),
.B(n_406),
.Y(n_1002)
);

A2O1A1Ixp33_ASAP7_75t_L g1003 ( 
.A1(n_858),
.A2(n_396),
.B(n_203),
.C(n_402),
.Y(n_1003)
);

BUFx6f_ASAP7_75t_L g1004 ( 
.A(n_768),
.Y(n_1004)
);

O2A1O1Ixp33_ASAP7_75t_L g1005 ( 
.A1(n_937),
.A2(n_43),
.B(n_45),
.C(n_46),
.Y(n_1005)
);

BUFx12f_ASAP7_75t_L g1006 ( 
.A(n_941),
.Y(n_1006)
);

OAI22xp5_ASAP7_75t_L g1007 ( 
.A1(n_778),
.A2(n_203),
.B1(n_51),
.B2(n_52),
.Y(n_1007)
);

NOR3xp33_ASAP7_75t_L g1008 ( 
.A(n_854),
.B(n_50),
.C(n_402),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_SL g1009 ( 
.A(n_804),
.B(n_54),
.Y(n_1009)
);

BUFx6f_ASAP7_75t_L g1010 ( 
.A(n_768),
.Y(n_1010)
);

O2A1O1Ixp33_ASAP7_75t_L g1011 ( 
.A1(n_940),
.A2(n_796),
.B(n_854),
.C(n_790),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_926),
.A2(n_58),
.B(n_63),
.Y(n_1012)
);

OR2x6_ASAP7_75t_SL g1013 ( 
.A(n_949),
.B(n_67),
.Y(n_1013)
);

AND2x4_ASAP7_75t_L g1014 ( 
.A(n_900),
.B(n_68),
.Y(n_1014)
);

HB1xp67_ASAP7_75t_L g1015 ( 
.A(n_873),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_SL g1016 ( 
.A(n_804),
.B(n_70),
.Y(n_1016)
);

INVx3_ASAP7_75t_L g1017 ( 
.A(n_941),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_836),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_831),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_805),
.A2(n_71),
.B(n_72),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_SL g1021 ( 
.A(n_810),
.B(n_82),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_821),
.B(n_87),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_810),
.B(n_855),
.Y(n_1023)
);

BUFx6f_ASAP7_75t_L g1024 ( 
.A(n_768),
.Y(n_1024)
);

O2A1O1Ixp33_ASAP7_75t_L g1025 ( 
.A1(n_907),
.A2(n_88),
.B(n_101),
.C(n_103),
.Y(n_1025)
);

BUFx2_ASAP7_75t_L g1026 ( 
.A(n_855),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_SL g1027 ( 
.A(n_779),
.B(n_112),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_SL g1028 ( 
.A(n_884),
.B(n_115),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_SL g1029 ( 
.A(n_935),
.B(n_154),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_884),
.B(n_123),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_806),
.B(n_138),
.Y(n_1031)
);

HB1xp67_ASAP7_75t_L g1032 ( 
.A(n_950),
.Y(n_1032)
);

INVxp67_ASAP7_75t_L g1033 ( 
.A(n_822),
.Y(n_1033)
);

A2O1A1Ixp33_ASAP7_75t_L g1034 ( 
.A1(n_850),
.A2(n_846),
.B(n_950),
.C(n_838),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_811),
.A2(n_809),
.B(n_784),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_835),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_R g1037 ( 
.A(n_884),
.B(n_776),
.Y(n_1037)
);

BUFx6f_ASAP7_75t_L g1038 ( 
.A(n_776),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_925),
.Y(n_1039)
);

AND2x4_ASAP7_75t_L g1040 ( 
.A(n_900),
.B(n_884),
.Y(n_1040)
);

INVx4_ASAP7_75t_L g1041 ( 
.A(n_776),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_837),
.B(n_834),
.Y(n_1042)
);

NAND2x1p5_ASAP7_75t_L g1043 ( 
.A(n_881),
.B(n_951),
.Y(n_1043)
);

BUFx3_ASAP7_75t_L g1044 ( 
.A(n_942),
.Y(n_1044)
);

AND2x2_ASAP7_75t_L g1045 ( 
.A(n_839),
.B(n_936),
.Y(n_1045)
);

HB1xp67_ASAP7_75t_L g1046 ( 
.A(n_909),
.Y(n_1046)
);

INVx6_ASAP7_75t_L g1047 ( 
.A(n_776),
.Y(n_1047)
);

OAI22x1_ASAP7_75t_L g1048 ( 
.A1(n_840),
.A2(n_877),
.B1(n_872),
.B2(n_871),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_875),
.Y(n_1049)
);

OAI22xp5_ASAP7_75t_L g1050 ( 
.A1(n_817),
.A2(n_819),
.B1(n_853),
.B2(n_839),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_833),
.A2(n_813),
.B(n_794),
.Y(n_1051)
);

NAND3xp33_ASAP7_75t_L g1052 ( 
.A(n_877),
.B(n_857),
.C(n_933),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_943),
.B(n_857),
.Y(n_1053)
);

INVx4_ASAP7_75t_L g1054 ( 
.A(n_879),
.Y(n_1054)
);

O2A1O1Ixp33_ASAP7_75t_L g1055 ( 
.A1(n_924),
.A2(n_887),
.B(n_851),
.C(n_849),
.Y(n_1055)
);

INVx1_ASAP7_75t_SL g1056 ( 
.A(n_942),
.Y(n_1056)
);

NOR3xp33_ASAP7_75t_L g1057 ( 
.A(n_781),
.B(n_911),
.C(n_816),
.Y(n_1057)
);

AO32x2_ASAP7_75t_L g1058 ( 
.A1(n_798),
.A2(n_944),
.A3(n_787),
.B1(n_939),
.B2(n_890),
.Y(n_1058)
);

OAI22x1_ASAP7_75t_L g1059 ( 
.A1(n_883),
.A2(n_891),
.B1(n_928),
.B2(n_893),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_902),
.B(n_913),
.Y(n_1060)
);

INVx3_ASAP7_75t_L g1061 ( 
.A(n_879),
.Y(n_1061)
);

A2O1A1Ixp33_ASAP7_75t_L g1062 ( 
.A1(n_915),
.A2(n_826),
.B(n_863),
.C(n_862),
.Y(n_1062)
);

AOI222xp33_ASAP7_75t_L g1063 ( 
.A1(n_931),
.A2(n_923),
.B1(n_866),
.B2(n_868),
.C1(n_916),
.C2(n_802),
.Y(n_1063)
);

OR2x2_ASAP7_75t_L g1064 ( 
.A(n_906),
.B(n_874),
.Y(n_1064)
);

BUFx6f_ASAP7_75t_L g1065 ( 
.A(n_879),
.Y(n_1065)
);

AND2x2_ASAP7_75t_L g1066 ( 
.A(n_881),
.B(n_879),
.Y(n_1066)
);

O2A1O1Ixp33_ASAP7_75t_L g1067 ( 
.A1(n_797),
.A2(n_802),
.B(n_864),
.C(n_786),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_919),
.B(n_951),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_882),
.B(n_892),
.Y(n_1069)
);

A2O1A1Ixp33_ASAP7_75t_SL g1070 ( 
.A1(n_865),
.A2(n_829),
.B(n_825),
.C(n_824),
.Y(n_1070)
);

AND2x2_ASAP7_75t_L g1071 ( 
.A(n_885),
.B(n_908),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_901),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_780),
.B(n_903),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_820),
.A2(n_818),
.B(n_843),
.Y(n_1074)
);

BUFx6f_ASAP7_75t_L g1075 ( 
.A(n_897),
.Y(n_1075)
);

A2O1A1Ixp33_ASAP7_75t_L g1076 ( 
.A1(n_876),
.A2(n_880),
.B(n_795),
.C(n_789),
.Y(n_1076)
);

AND2x4_ASAP7_75t_L g1077 ( 
.A(n_786),
.B(n_860),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_797),
.B(n_814),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_815),
.B(n_870),
.Y(n_1079)
);

BUFx3_ASAP7_75t_L g1080 ( 
.A(n_948),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_856),
.B(n_861),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_R g1082 ( 
.A(n_783),
.B(n_904),
.Y(n_1082)
);

AOI21x1_ASAP7_75t_L g1083 ( 
.A1(n_859),
.A2(n_927),
.B(n_946),
.Y(n_1083)
);

BUFx2_ASAP7_75t_L g1084 ( 
.A(n_920),
.Y(n_1084)
);

BUFx2_ASAP7_75t_L g1085 ( 
.A(n_947),
.Y(n_1085)
);

CKINVDCx14_ASAP7_75t_R g1086 ( 
.A(n_917),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_841),
.B(n_844),
.Y(n_1087)
);

BUFx2_ASAP7_75t_L g1088 ( 
.A(n_897),
.Y(n_1088)
);

O2A1O1Ixp33_ASAP7_75t_L g1089 ( 
.A1(n_899),
.A2(n_946),
.B(n_932),
.C(n_927),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_899),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_932),
.A2(n_922),
.B(n_930),
.Y(n_1091)
);

INVx1_ASAP7_75t_SL g1092 ( 
.A(n_945),
.Y(n_1092)
);

A2O1A1Ixp33_ASAP7_75t_L g1093 ( 
.A1(n_894),
.A2(n_896),
.B(n_898),
.C(n_905),
.Y(n_1093)
);

OAI21x1_ASAP7_75t_L g1094 ( 
.A1(n_1074),
.A2(n_929),
.B(n_912),
.Y(n_1094)
);

AOI22xp33_ASAP7_75t_L g1095 ( 
.A1(n_985),
.A2(n_918),
.B1(n_969),
.B2(n_1007),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_979),
.B(n_997),
.Y(n_1096)
);

BUFx10_ASAP7_75t_L g1097 ( 
.A(n_1018),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_1035),
.A2(n_1051),
.B(n_960),
.Y(n_1098)
);

OAI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_1011),
.A2(n_1034),
.B(n_1062),
.Y(n_1099)
);

BUFx2_ASAP7_75t_L g1100 ( 
.A(n_953),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_1031),
.A2(n_1073),
.B(n_1079),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_1031),
.A2(n_1073),
.B(n_1079),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_1050),
.A2(n_1087),
.B(n_1042),
.Y(n_1103)
);

BUFx8_ASAP7_75t_L g1104 ( 
.A(n_1001),
.Y(n_1104)
);

OAI21x1_ASAP7_75t_SL g1105 ( 
.A1(n_1007),
.A2(n_1067),
.B(n_1042),
.Y(n_1105)
);

OAI21x1_ASAP7_75t_L g1106 ( 
.A1(n_1091),
.A2(n_971),
.B(n_1087),
.Y(n_1106)
);

OAI21x1_ASAP7_75t_L g1107 ( 
.A1(n_1081),
.A2(n_990),
.B(n_1068),
.Y(n_1107)
);

NAND3xp33_ASAP7_75t_L g1108 ( 
.A(n_1005),
.B(n_1032),
.C(n_1045),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_1050),
.A2(n_989),
.B(n_1053),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_L g1110 ( 
.A(n_977),
.B(n_994),
.Y(n_1110)
);

O2A1O1Ixp5_ASAP7_75t_L g1111 ( 
.A1(n_1009),
.A2(n_1016),
.B(n_1021),
.C(n_1002),
.Y(n_1111)
);

AO31x2_ASAP7_75t_L g1112 ( 
.A1(n_991),
.A2(n_996),
.A3(n_1059),
.B(n_1076),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_997),
.B(n_962),
.Y(n_1113)
);

AND2x2_ASAP7_75t_L g1114 ( 
.A(n_992),
.B(n_954),
.Y(n_1114)
);

AND2x4_ASAP7_75t_L g1115 ( 
.A(n_963),
.B(n_1044),
.Y(n_1115)
);

AND2x2_ASAP7_75t_L g1116 ( 
.A(n_1033),
.B(n_959),
.Y(n_1116)
);

CKINVDCx9p33_ASAP7_75t_R g1117 ( 
.A(n_1026),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_966),
.Y(n_1118)
);

AOI31xp67_ASAP7_75t_L g1119 ( 
.A1(n_1078),
.A2(n_1090),
.A3(n_1053),
.B(n_1023),
.Y(n_1119)
);

A2O1A1Ixp33_ASAP7_75t_L g1120 ( 
.A1(n_1052),
.A2(n_983),
.B(n_1055),
.C(n_981),
.Y(n_1120)
);

AOI22xp5_ASAP7_75t_L g1121 ( 
.A1(n_1029),
.A2(n_976),
.B1(n_1027),
.B2(n_1063),
.Y(n_1121)
);

BUFx6f_ASAP7_75t_L g1122 ( 
.A(n_1006),
.Y(n_1122)
);

OAI22xp5_ASAP7_75t_L g1123 ( 
.A1(n_989),
.A2(n_988),
.B1(n_984),
.B2(n_1013),
.Y(n_1123)
);

INVx5_ASAP7_75t_L g1124 ( 
.A(n_1040),
.Y(n_1124)
);

AOI22xp5_ASAP7_75t_L g1125 ( 
.A1(n_1029),
.A2(n_1027),
.B1(n_1063),
.B2(n_1008),
.Y(n_1125)
);

OAI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_956),
.A2(n_1003),
.B(n_986),
.Y(n_1126)
);

OA21x2_ASAP7_75t_L g1127 ( 
.A1(n_980),
.A2(n_1083),
.B(n_1057),
.Y(n_1127)
);

BUFx10_ASAP7_75t_L g1128 ( 
.A(n_1047),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_1070),
.A2(n_1012),
.B(n_1093),
.Y(n_1129)
);

OAI21x1_ASAP7_75t_L g1130 ( 
.A1(n_965),
.A2(n_1089),
.B(n_973),
.Y(n_1130)
);

NOR2xp67_ASAP7_75t_L g1131 ( 
.A(n_1041),
.B(n_1054),
.Y(n_1131)
);

CKINVDCx12_ASAP7_75t_R g1132 ( 
.A(n_1086),
.Y(n_1132)
);

NAND3xp33_ASAP7_75t_SL g1133 ( 
.A(n_970),
.B(n_1025),
.C(n_1046),
.Y(n_1133)
);

AND2x2_ASAP7_75t_L g1134 ( 
.A(n_972),
.B(n_987),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1036),
.Y(n_1135)
);

OAI21x1_ASAP7_75t_L g1136 ( 
.A1(n_973),
.A2(n_1071),
.B(n_1069),
.Y(n_1136)
);

AO31x2_ASAP7_75t_L g1137 ( 
.A1(n_1048),
.A2(n_975),
.A3(n_1072),
.B(n_1084),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1092),
.A2(n_1020),
.B(n_1022),
.Y(n_1138)
);

AO31x2_ASAP7_75t_L g1139 ( 
.A1(n_1060),
.A2(n_955),
.A3(n_968),
.B(n_1039),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_1092),
.A2(n_955),
.B(n_968),
.Y(n_1140)
);

BUFx2_ASAP7_75t_L g1141 ( 
.A(n_1000),
.Y(n_1141)
);

OAI22x1_ASAP7_75t_L g1142 ( 
.A1(n_998),
.A2(n_1014),
.B1(n_995),
.B2(n_1015),
.Y(n_1142)
);

BUFx3_ASAP7_75t_L g1143 ( 
.A(n_999),
.Y(n_1143)
);

AO21x2_ASAP7_75t_L g1144 ( 
.A1(n_1082),
.A2(n_967),
.B(n_982),
.Y(n_1144)
);

AOI22xp5_ASAP7_75t_L g1145 ( 
.A1(n_1056),
.A2(n_1064),
.B1(n_1017),
.B2(n_1014),
.Y(n_1145)
);

A2O1A1Ixp33_ASAP7_75t_L g1146 ( 
.A1(n_974),
.A2(n_1077),
.B(n_1080),
.C(n_1017),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1049),
.Y(n_1147)
);

HB1xp67_ASAP7_75t_L g1148 ( 
.A(n_1088),
.Y(n_1148)
);

CKINVDCx20_ASAP7_75t_R g1149 ( 
.A(n_999),
.Y(n_1149)
);

A2O1A1Ixp33_ASAP7_75t_L g1150 ( 
.A1(n_1077),
.A2(n_961),
.B(n_1085),
.C(n_984),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_993),
.A2(n_1030),
.B(n_1028),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1047),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_1061),
.A2(n_1075),
.B(n_958),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1047),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_1061),
.A2(n_1075),
.B(n_958),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_952),
.B(n_978),
.Y(n_1156)
);

BUFx2_ASAP7_75t_L g1157 ( 
.A(n_1037),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_SL g1158 ( 
.A(n_978),
.B(n_1075),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1040),
.B(n_1066),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1004),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1010),
.Y(n_1161)
);

O2A1O1Ixp33_ASAP7_75t_SL g1162 ( 
.A1(n_1041),
.A2(n_1054),
.B(n_1010),
.C(n_1024),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_964),
.Y(n_1163)
);

BUFx10_ASAP7_75t_L g1164 ( 
.A(n_1024),
.Y(n_1164)
);

AO32x2_ASAP7_75t_L g1165 ( 
.A1(n_1058),
.A2(n_1007),
.A3(n_1050),
.B1(n_785),
.B2(n_989),
.Y(n_1165)
);

OAI21x1_ASAP7_75t_L g1166 ( 
.A1(n_1043),
.A2(n_1058),
.B(n_1038),
.Y(n_1166)
);

OAI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_1058),
.A2(n_960),
.B(n_791),
.Y(n_1167)
);

OAI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1065),
.A2(n_960),
.B(n_785),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_SL g1169 ( 
.A(n_1065),
.B(n_960),
.Y(n_1169)
);

OAI21x1_ASAP7_75t_L g1170 ( 
.A1(n_1065),
.A2(n_1074),
.B(n_1091),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_SL g1171 ( 
.A(n_960),
.B(n_785),
.Y(n_1171)
);

NAND3xp33_ASAP7_75t_L g1172 ( 
.A(n_960),
.B(n_842),
.C(n_785),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_1035),
.A2(n_785),
.B(n_1051),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_969),
.B(n_773),
.Y(n_1174)
);

INVxp67_ASAP7_75t_L g1175 ( 
.A(n_954),
.Y(n_1175)
);

AO31x2_ASAP7_75t_L g1176 ( 
.A1(n_991),
.A2(n_996),
.A3(n_832),
.B(n_798),
.Y(n_1176)
);

AO31x2_ASAP7_75t_L g1177 ( 
.A1(n_991),
.A2(n_996),
.A3(n_832),
.B(n_798),
.Y(n_1177)
);

OR2x2_ASAP7_75t_L g1178 ( 
.A(n_979),
.B(n_977),
.Y(n_1178)
);

BUFx10_ASAP7_75t_L g1179 ( 
.A(n_1018),
.Y(n_1179)
);

A2O1A1Ixp33_ASAP7_75t_L g1180 ( 
.A1(n_960),
.A2(n_842),
.B(n_969),
.C(n_773),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_969),
.B(n_773),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1035),
.A2(n_785),
.B(n_1051),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_957),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_957),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_1019),
.Y(n_1185)
);

BUFx2_ASAP7_75t_L g1186 ( 
.A(n_953),
.Y(n_1186)
);

OAI22xp5_ASAP7_75t_L g1187 ( 
.A1(n_960),
.A2(n_785),
.B1(n_842),
.B2(n_773),
.Y(n_1187)
);

INVx3_ASAP7_75t_SL g1188 ( 
.A(n_1018),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_969),
.B(n_773),
.Y(n_1189)
);

AND2x4_ASAP7_75t_L g1190 ( 
.A(n_963),
.B(n_1044),
.Y(n_1190)
);

OAI21x1_ASAP7_75t_L g1191 ( 
.A1(n_1074),
.A2(n_1091),
.B(n_971),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1035),
.A2(n_785),
.B(n_1051),
.Y(n_1192)
);

O2A1O1Ixp33_ASAP7_75t_L g1193 ( 
.A1(n_960),
.A2(n_842),
.B(n_785),
.C(n_773),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_957),
.Y(n_1194)
);

BUFx10_ASAP7_75t_L g1195 ( 
.A(n_1018),
.Y(n_1195)
);

AOI221xp5_ASAP7_75t_SL g1196 ( 
.A1(n_960),
.A2(n_1007),
.B1(n_785),
.B2(n_921),
.C(n_910),
.Y(n_1196)
);

AO31x2_ASAP7_75t_L g1197 ( 
.A1(n_991),
.A2(n_996),
.A3(n_832),
.B(n_798),
.Y(n_1197)
);

AOI221xp5_ASAP7_75t_SL g1198 ( 
.A1(n_960),
.A2(n_1007),
.B1(n_785),
.B2(n_921),
.C(n_910),
.Y(n_1198)
);

OAI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_960),
.A2(n_791),
.B(n_845),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_957),
.Y(n_1200)
);

A2O1A1Ixp33_ASAP7_75t_L g1201 ( 
.A1(n_960),
.A2(n_842),
.B(n_969),
.C(n_773),
.Y(n_1201)
);

AOI221x1_ASAP7_75t_L g1202 ( 
.A1(n_1007),
.A2(n_985),
.B1(n_1008),
.B2(n_785),
.C(n_1048),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1035),
.A2(n_785),
.B(n_1051),
.Y(n_1203)
);

OAI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_960),
.A2(n_791),
.B(n_845),
.Y(n_1204)
);

BUFx2_ASAP7_75t_L g1205 ( 
.A(n_953),
.Y(n_1205)
);

INVx8_ASAP7_75t_L g1206 ( 
.A(n_1006),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_969),
.B(n_773),
.Y(n_1207)
);

AO31x2_ASAP7_75t_L g1208 ( 
.A1(n_991),
.A2(n_996),
.A3(n_832),
.B(n_798),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1035),
.A2(n_785),
.B(n_1051),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1035),
.A2(n_785),
.B(n_1051),
.Y(n_1210)
);

AO32x2_ASAP7_75t_L g1211 ( 
.A1(n_1007),
.A2(n_1050),
.A3(n_785),
.B1(n_989),
.B2(n_973),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1019),
.Y(n_1212)
);

O2A1O1Ixp33_ASAP7_75t_L g1213 ( 
.A1(n_960),
.A2(n_842),
.B(n_785),
.C(n_773),
.Y(n_1213)
);

AOI221xp5_ASAP7_75t_L g1214 ( 
.A1(n_960),
.A2(n_773),
.B1(n_417),
.B2(n_1007),
.C(n_969),
.Y(n_1214)
);

O2A1O1Ixp33_ASAP7_75t_SL g1215 ( 
.A1(n_960),
.A2(n_785),
.B(n_791),
.C(n_1034),
.Y(n_1215)
);

OA21x2_ASAP7_75t_L g1216 ( 
.A1(n_1074),
.A2(n_1051),
.B(n_1087),
.Y(n_1216)
);

AOI221xp5_ASAP7_75t_L g1217 ( 
.A1(n_960),
.A2(n_773),
.B1(n_417),
.B2(n_1007),
.C(n_969),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1035),
.A2(n_785),
.B(n_1051),
.Y(n_1218)
);

AND2x2_ASAP7_75t_L g1219 ( 
.A(n_979),
.B(n_934),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_969),
.B(n_773),
.Y(n_1220)
);

OAI21x1_ASAP7_75t_L g1221 ( 
.A1(n_1074),
.A2(n_1091),
.B(n_971),
.Y(n_1221)
);

OAI21x1_ASAP7_75t_L g1222 ( 
.A1(n_1074),
.A2(n_1091),
.B(n_971),
.Y(n_1222)
);

OA21x2_ASAP7_75t_L g1223 ( 
.A1(n_1074),
.A2(n_1051),
.B(n_1087),
.Y(n_1223)
);

INVxp67_ASAP7_75t_L g1224 ( 
.A(n_954),
.Y(n_1224)
);

AOI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1035),
.A2(n_785),
.B(n_1051),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1113),
.B(n_1174),
.Y(n_1226)
);

INVx4_ASAP7_75t_L g1227 ( 
.A(n_1188),
.Y(n_1227)
);

INVx3_ASAP7_75t_L g1228 ( 
.A(n_1164),
.Y(n_1228)
);

INVx2_ASAP7_75t_SL g1229 ( 
.A(n_1206),
.Y(n_1229)
);

AOI22xp33_ASAP7_75t_L g1230 ( 
.A1(n_1214),
.A2(n_1217),
.B1(n_1187),
.B2(n_1207),
.Y(n_1230)
);

HB1xp67_ASAP7_75t_L g1231 ( 
.A(n_1148),
.Y(n_1231)
);

AOI22xp33_ASAP7_75t_L g1232 ( 
.A1(n_1181),
.A2(n_1220),
.B1(n_1189),
.B2(n_1172),
.Y(n_1232)
);

OAI22xp5_ASAP7_75t_L g1233 ( 
.A1(n_1180),
.A2(n_1201),
.B1(n_1172),
.B2(n_1213),
.Y(n_1233)
);

AOI22xp33_ASAP7_75t_L g1234 ( 
.A1(n_1121),
.A2(n_1171),
.B1(n_1219),
.B2(n_1125),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1103),
.B(n_1193),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1134),
.Y(n_1236)
);

AOI22xp33_ASAP7_75t_SL g1237 ( 
.A1(n_1105),
.A2(n_1204),
.B1(n_1199),
.B2(n_1167),
.Y(n_1237)
);

INVx3_ASAP7_75t_L g1238 ( 
.A(n_1164),
.Y(n_1238)
);

INVx6_ASAP7_75t_L g1239 ( 
.A(n_1097),
.Y(n_1239)
);

OAI22xp5_ASAP7_75t_SL g1240 ( 
.A1(n_1149),
.A2(n_1132),
.B1(n_1121),
.B2(n_1142),
.Y(n_1240)
);

OAI22x1_ASAP7_75t_L g1241 ( 
.A1(n_1125),
.A2(n_1145),
.B1(n_1108),
.B2(n_1200),
.Y(n_1241)
);

INVx1_ASAP7_75t_SL g1242 ( 
.A(n_1117),
.Y(n_1242)
);

AOI22xp5_ASAP7_75t_L g1243 ( 
.A1(n_1196),
.A2(n_1198),
.B1(n_1123),
.B2(n_1108),
.Y(n_1243)
);

INVx6_ASAP7_75t_L g1244 ( 
.A(n_1179),
.Y(n_1244)
);

AOI22xp33_ASAP7_75t_SL g1245 ( 
.A1(n_1199),
.A2(n_1204),
.B1(n_1167),
.B2(n_1198),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1135),
.Y(n_1246)
);

AOI22xp33_ASAP7_75t_L g1247 ( 
.A1(n_1095),
.A2(n_1185),
.B1(n_1212),
.B2(n_1133),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1183),
.Y(n_1248)
);

INVx6_ASAP7_75t_L g1249 ( 
.A(n_1179),
.Y(n_1249)
);

AOI22xp33_ASAP7_75t_SL g1250 ( 
.A1(n_1196),
.A2(n_1168),
.B1(n_1099),
.B2(n_1104),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1184),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_1118),
.Y(n_1252)
);

INVx6_ASAP7_75t_L g1253 ( 
.A(n_1195),
.Y(n_1253)
);

INVx2_ASAP7_75t_SL g1254 ( 
.A(n_1206),
.Y(n_1254)
);

CKINVDCx11_ASAP7_75t_R g1255 ( 
.A(n_1195),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_1143),
.Y(n_1256)
);

BUFx2_ASAP7_75t_L g1257 ( 
.A(n_1178),
.Y(n_1257)
);

AOI22xp33_ASAP7_75t_L g1258 ( 
.A1(n_1147),
.A2(n_1116),
.B1(n_1096),
.B2(n_1114),
.Y(n_1258)
);

INVx3_ASAP7_75t_L g1259 ( 
.A(n_1128),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1109),
.B(n_1139),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_1194),
.Y(n_1261)
);

BUFx3_ASAP7_75t_L g1262 ( 
.A(n_1141),
.Y(n_1262)
);

BUFx3_ASAP7_75t_L g1263 ( 
.A(n_1100),
.Y(n_1263)
);

INVx6_ASAP7_75t_L g1264 ( 
.A(n_1122),
.Y(n_1264)
);

INVx5_ASAP7_75t_L g1265 ( 
.A(n_1157),
.Y(n_1265)
);

AOI22xp33_ASAP7_75t_L g1266 ( 
.A1(n_1099),
.A2(n_1110),
.B1(n_1169),
.B2(n_1122),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1139),
.Y(n_1267)
);

CKINVDCx11_ASAP7_75t_R g1268 ( 
.A(n_1122),
.Y(n_1268)
);

OAI22xp5_ASAP7_75t_L g1269 ( 
.A1(n_1120),
.A2(n_1098),
.B1(n_1210),
.B2(n_1225),
.Y(n_1269)
);

OAI22xp33_ASAP7_75t_L g1270 ( 
.A1(n_1202),
.A2(n_1175),
.B1(n_1224),
.B2(n_1186),
.Y(n_1270)
);

AOI22xp33_ASAP7_75t_SL g1271 ( 
.A1(n_1104),
.A2(n_1126),
.B1(n_1124),
.B2(n_1211),
.Y(n_1271)
);

CKINVDCx11_ASAP7_75t_R g1272 ( 
.A(n_1205),
.Y(n_1272)
);

CKINVDCx11_ASAP7_75t_R g1273 ( 
.A(n_1128),
.Y(n_1273)
);

BUFx3_ASAP7_75t_L g1274 ( 
.A(n_1115),
.Y(n_1274)
);

OAI21xp5_ASAP7_75t_SL g1275 ( 
.A1(n_1173),
.A2(n_1209),
.B(n_1192),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1139),
.Y(n_1276)
);

BUFx12f_ASAP7_75t_L g1277 ( 
.A(n_1115),
.Y(n_1277)
);

BUFx10_ASAP7_75t_L g1278 ( 
.A(n_1190),
.Y(n_1278)
);

CKINVDCx5p33_ASAP7_75t_R g1279 ( 
.A(n_1190),
.Y(n_1279)
);

AOI22xp33_ASAP7_75t_SL g1280 ( 
.A1(n_1126),
.A2(n_1124),
.B1(n_1211),
.B2(n_1165),
.Y(n_1280)
);

AOI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1144),
.A2(n_1159),
.B1(n_1140),
.B2(n_1163),
.Y(n_1281)
);

INVx8_ASAP7_75t_L g1282 ( 
.A(n_1124),
.Y(n_1282)
);

OAI221xp5_ASAP7_75t_L g1283 ( 
.A1(n_1215),
.A2(n_1111),
.B1(n_1182),
.B2(n_1218),
.C(n_1203),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_L g1284 ( 
.A1(n_1144),
.A2(n_1158),
.B1(n_1152),
.B2(n_1154),
.Y(n_1284)
);

BUFx4f_ASAP7_75t_SL g1285 ( 
.A(n_1160),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1119),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_1161),
.Y(n_1287)
);

OAI21xp5_ASAP7_75t_SL g1288 ( 
.A1(n_1211),
.A2(n_1151),
.B(n_1129),
.Y(n_1288)
);

AOI22xp33_ASAP7_75t_SL g1289 ( 
.A1(n_1165),
.A2(n_1136),
.B1(n_1101),
.B2(n_1102),
.Y(n_1289)
);

INVx3_ASAP7_75t_L g1290 ( 
.A(n_1166),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1138),
.A2(n_1216),
.B(n_1223),
.Y(n_1291)
);

OAI22xp5_ASAP7_75t_L g1292 ( 
.A1(n_1150),
.A2(n_1165),
.B1(n_1146),
.B2(n_1156),
.Y(n_1292)
);

AOI22xp33_ASAP7_75t_SL g1293 ( 
.A1(n_1130),
.A2(n_1127),
.B1(n_1153),
.B2(n_1155),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_SL g1294 ( 
.A1(n_1216),
.A2(n_1223),
.B1(n_1137),
.B2(n_1107),
.Y(n_1294)
);

INVx5_ASAP7_75t_L g1295 ( 
.A(n_1162),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1137),
.Y(n_1296)
);

INVx6_ASAP7_75t_L g1297 ( 
.A(n_1131),
.Y(n_1297)
);

AOI22xp33_ASAP7_75t_L g1298 ( 
.A1(n_1094),
.A2(n_1106),
.B1(n_1170),
.B2(n_1222),
.Y(n_1298)
);

CKINVDCx10_ASAP7_75t_R g1299 ( 
.A(n_1176),
.Y(n_1299)
);

BUFx2_ASAP7_75t_SL g1300 ( 
.A(n_1112),
.Y(n_1300)
);

AOI22xp5_ASAP7_75t_L g1301 ( 
.A1(n_1191),
.A2(n_1221),
.B1(n_1112),
.B2(n_1197),
.Y(n_1301)
);

AOI22xp33_ASAP7_75t_SL g1302 ( 
.A1(n_1177),
.A2(n_985),
.B1(n_1007),
.B2(n_773),
.Y(n_1302)
);

AOI22xp33_ASAP7_75t_SL g1303 ( 
.A1(n_1197),
.A2(n_985),
.B1(n_1007),
.B2(n_773),
.Y(n_1303)
);

AOI22xp33_ASAP7_75t_L g1304 ( 
.A1(n_1197),
.A2(n_778),
.B1(n_467),
.B2(n_985),
.Y(n_1304)
);

OAI22xp5_ASAP7_75t_L g1305 ( 
.A1(n_1208),
.A2(n_1201),
.B1(n_1180),
.B2(n_960),
.Y(n_1305)
);

AOI22xp33_ASAP7_75t_SL g1306 ( 
.A1(n_1187),
.A2(n_985),
.B1(n_1007),
.B2(n_732),
.Y(n_1306)
);

AOI22xp33_ASAP7_75t_SL g1307 ( 
.A1(n_1187),
.A2(n_985),
.B1(n_1007),
.B2(n_732),
.Y(n_1307)
);

OAI22xp5_ASAP7_75t_L g1308 ( 
.A1(n_1180),
.A2(n_1201),
.B1(n_960),
.B2(n_1187),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1134),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_1188),
.Y(n_1310)
);

INVx1_ASAP7_75t_SL g1311 ( 
.A(n_1117),
.Y(n_1311)
);

CKINVDCx6p67_ASAP7_75t_R g1312 ( 
.A(n_1132),
.Y(n_1312)
);

AOI22xp33_ASAP7_75t_L g1313 ( 
.A1(n_1214),
.A2(n_778),
.B1(n_467),
.B2(n_985),
.Y(n_1313)
);

OAI21xp5_ASAP7_75t_L g1314 ( 
.A1(n_1180),
.A2(n_960),
.B(n_1201),
.Y(n_1314)
);

INVx6_ASAP7_75t_L g1315 ( 
.A(n_1097),
.Y(n_1315)
);

OAI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_1180),
.A2(n_1201),
.B1(n_960),
.B2(n_1187),
.Y(n_1316)
);

CKINVDCx8_ASAP7_75t_R g1317 ( 
.A(n_1118),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1134),
.Y(n_1318)
);

AOI22xp33_ASAP7_75t_L g1319 ( 
.A1(n_1214),
.A2(n_778),
.B1(n_467),
.B2(n_985),
.Y(n_1319)
);

CKINVDCx20_ASAP7_75t_R g1320 ( 
.A(n_1132),
.Y(n_1320)
);

INVx6_ASAP7_75t_L g1321 ( 
.A(n_1097),
.Y(n_1321)
);

CKINVDCx20_ASAP7_75t_R g1322 ( 
.A(n_1132),
.Y(n_1322)
);

BUFx6f_ASAP7_75t_L g1323 ( 
.A(n_1157),
.Y(n_1323)
);

INVx8_ASAP7_75t_L g1324 ( 
.A(n_1206),
.Y(n_1324)
);

CKINVDCx11_ASAP7_75t_R g1325 ( 
.A(n_1149),
.Y(n_1325)
);

BUFx6f_ASAP7_75t_L g1326 ( 
.A(n_1157),
.Y(n_1326)
);

AOI22xp33_ASAP7_75t_L g1327 ( 
.A1(n_1214),
.A2(n_778),
.B1(n_467),
.B2(n_985),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_SL g1328 ( 
.A1(n_1187),
.A2(n_985),
.B1(n_1007),
.B2(n_732),
.Y(n_1328)
);

AOI21xp5_ASAP7_75t_L g1329 ( 
.A1(n_1173),
.A2(n_1192),
.B(n_1182),
.Y(n_1329)
);

AOI22xp5_ASAP7_75t_L g1330 ( 
.A1(n_1214),
.A2(n_1217),
.B1(n_773),
.B2(n_985),
.Y(n_1330)
);

OAI21xp5_ASAP7_75t_SL g1331 ( 
.A1(n_1214),
.A2(n_960),
.B(n_1217),
.Y(n_1331)
);

CKINVDCx20_ASAP7_75t_R g1332 ( 
.A(n_1132),
.Y(n_1332)
);

BUFx10_ASAP7_75t_L g1333 ( 
.A(n_1118),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_1267),
.Y(n_1334)
);

INVx2_ASAP7_75t_SL g1335 ( 
.A(n_1265),
.Y(n_1335)
);

AND2x4_ASAP7_75t_L g1336 ( 
.A(n_1265),
.B(n_1261),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1280),
.B(n_1236),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1276),
.Y(n_1338)
);

OR2x6_ASAP7_75t_L g1339 ( 
.A(n_1282),
.B(n_1300),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1226),
.B(n_1232),
.Y(n_1340)
);

BUFx3_ASAP7_75t_L g1341 ( 
.A(n_1277),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1260),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1260),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_1325),
.Y(n_1344)
);

INVx2_ASAP7_75t_SL g1345 ( 
.A(n_1265),
.Y(n_1345)
);

INVx3_ASAP7_75t_L g1346 ( 
.A(n_1290),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1296),
.Y(n_1347)
);

HB1xp67_ASAP7_75t_L g1348 ( 
.A(n_1231),
.Y(n_1348)
);

OAI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1331),
.A2(n_1330),
.B(n_1230),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1286),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1309),
.B(n_1318),
.Y(n_1351)
);

INVx1_ASAP7_75t_SL g1352 ( 
.A(n_1272),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1246),
.Y(n_1353)
);

AND2x4_ASAP7_75t_L g1354 ( 
.A(n_1248),
.B(n_1251),
.Y(n_1354)
);

AO21x2_ASAP7_75t_L g1355 ( 
.A1(n_1291),
.A2(n_1301),
.B(n_1329),
.Y(n_1355)
);

INVx3_ASAP7_75t_L g1356 ( 
.A(n_1290),
.Y(n_1356)
);

BUFx3_ASAP7_75t_L g1357 ( 
.A(n_1323),
.Y(n_1357)
);

NOR2xp33_ASAP7_75t_L g1358 ( 
.A(n_1242),
.B(n_1311),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1235),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1235),
.Y(n_1360)
);

INVx3_ASAP7_75t_L g1361 ( 
.A(n_1295),
.Y(n_1361)
);

HB1xp67_ASAP7_75t_L g1362 ( 
.A(n_1257),
.Y(n_1362)
);

NOR2xp33_ASAP7_75t_L g1363 ( 
.A(n_1242),
.B(n_1311),
.Y(n_1363)
);

OR2x2_ASAP7_75t_L g1364 ( 
.A(n_1234),
.B(n_1258),
.Y(n_1364)
);

A2O1A1Ixp33_ASAP7_75t_L g1365 ( 
.A1(n_1331),
.A2(n_1319),
.B(n_1313),
.C(n_1327),
.Y(n_1365)
);

INVxp67_ASAP7_75t_L g1366 ( 
.A(n_1263),
.Y(n_1366)
);

OAI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1291),
.A2(n_1329),
.B(n_1269),
.Y(n_1367)
);

NAND2xp33_ASAP7_75t_R g1368 ( 
.A(n_1256),
.B(n_1279),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1241),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1292),
.Y(n_1370)
);

AOI22xp33_ASAP7_75t_L g1371 ( 
.A1(n_1304),
.A2(n_1307),
.B1(n_1328),
.B2(n_1306),
.Y(n_1371)
);

HB1xp67_ASAP7_75t_L g1372 ( 
.A(n_1262),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1292),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1243),
.Y(n_1374)
);

OA21x2_ASAP7_75t_L g1375 ( 
.A1(n_1275),
.A2(n_1288),
.B(n_1298),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1305),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1305),
.Y(n_1377)
);

OAI21x1_ASAP7_75t_L g1378 ( 
.A1(n_1269),
.A2(n_1275),
.B(n_1314),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1270),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1283),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1281),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1283),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1288),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1226),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1289),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1289),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1245),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1308),
.B(n_1316),
.Y(n_1388)
);

OAI21x1_ASAP7_75t_L g1389 ( 
.A1(n_1314),
.A2(n_1233),
.B(n_1316),
.Y(n_1389)
);

OAI21x1_ASAP7_75t_L g1390 ( 
.A1(n_1233),
.A2(n_1308),
.B(n_1284),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1294),
.Y(n_1391)
);

OAI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1247),
.A2(n_1266),
.B(n_1228),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1294),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1237),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1271),
.B(n_1250),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1293),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1299),
.Y(n_1397)
);

BUFx2_ASAP7_75t_R g1398 ( 
.A(n_1317),
.Y(n_1398)
);

AOI21xp5_ASAP7_75t_SL g1399 ( 
.A1(n_1274),
.A2(n_1287),
.B(n_1282),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1302),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1302),
.Y(n_1401)
);

BUFx2_ASAP7_75t_L g1402 ( 
.A(n_1326),
.Y(n_1402)
);

AOI222xp33_ASAP7_75t_L g1403 ( 
.A1(n_1240),
.A2(n_1303),
.B1(n_1268),
.B2(n_1285),
.C1(n_1322),
.C2(n_1320),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1303),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1259),
.Y(n_1405)
);

AOI22xp5_ASAP7_75t_L g1406 ( 
.A1(n_1332),
.A2(n_1312),
.B1(n_1264),
.B2(n_1229),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1383),
.B(n_1259),
.Y(n_1407)
);

AOI22xp5_ASAP7_75t_L g1408 ( 
.A1(n_1349),
.A2(n_1264),
.B1(n_1254),
.B2(n_1297),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1362),
.B(n_1227),
.Y(n_1409)
);

NOR2xp33_ASAP7_75t_L g1410 ( 
.A(n_1388),
.B(n_1227),
.Y(n_1410)
);

OAI21xp5_ASAP7_75t_L g1411 ( 
.A1(n_1389),
.A2(n_1228),
.B(n_1238),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1402),
.B(n_1333),
.Y(n_1412)
);

OR2x6_ASAP7_75t_L g1413 ( 
.A(n_1399),
.B(n_1282),
.Y(n_1413)
);

INVxp67_ASAP7_75t_L g1414 ( 
.A(n_1342),
.Y(n_1414)
);

OAI21xp5_ASAP7_75t_L g1415 ( 
.A1(n_1389),
.A2(n_1238),
.B(n_1310),
.Y(n_1415)
);

AO21x2_ASAP7_75t_L g1416 ( 
.A1(n_1396),
.A2(n_1381),
.B(n_1385),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1372),
.B(n_1273),
.Y(n_1417)
);

OAI22xp5_ASAP7_75t_L g1418 ( 
.A1(n_1371),
.A2(n_1239),
.B1(n_1244),
.B2(n_1249),
.Y(n_1418)
);

HB1xp67_ASAP7_75t_L g1419 ( 
.A(n_1342),
.Y(n_1419)
);

AND2x4_ASAP7_75t_L g1420 ( 
.A(n_1336),
.B(n_1252),
.Y(n_1420)
);

OR2x2_ASAP7_75t_L g1421 ( 
.A(n_1348),
.B(n_1354),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1384),
.B(n_1244),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1384),
.B(n_1249),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1351),
.B(n_1354),
.Y(n_1424)
);

OR2x2_ASAP7_75t_L g1425 ( 
.A(n_1354),
.B(n_1324),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1351),
.B(n_1357),
.Y(n_1426)
);

AO32x2_ASAP7_75t_L g1427 ( 
.A1(n_1335),
.A2(n_1278),
.A3(n_1253),
.B1(n_1315),
.B2(n_1321),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1353),
.Y(n_1428)
);

OAI22xp5_ASAP7_75t_SL g1429 ( 
.A1(n_1394),
.A2(n_1315),
.B1(n_1321),
.B2(n_1255),
.Y(n_1429)
);

OAI21xp5_ASAP7_75t_L g1430 ( 
.A1(n_1390),
.A2(n_1387),
.B(n_1378),
.Y(n_1430)
);

NOR2xp33_ASAP7_75t_L g1431 ( 
.A(n_1340),
.B(n_1297),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1366),
.B(n_1324),
.Y(n_1432)
);

O2A1O1Ixp33_ASAP7_75t_L g1433 ( 
.A1(n_1365),
.A2(n_1387),
.B(n_1394),
.C(n_1374),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1358),
.B(n_1363),
.Y(n_1434)
);

NAND2xp33_ASAP7_75t_L g1435 ( 
.A(n_1380),
.B(n_1382),
.Y(n_1435)
);

OR2x6_ASAP7_75t_L g1436 ( 
.A(n_1399),
.B(n_1339),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1359),
.B(n_1360),
.Y(n_1437)
);

AO32x2_ASAP7_75t_L g1438 ( 
.A1(n_1335),
.A2(n_1345),
.A3(n_1400),
.B1(n_1401),
.B2(n_1370),
.Y(n_1438)
);

OAI22xp5_ASAP7_75t_L g1439 ( 
.A1(n_1376),
.A2(n_1377),
.B1(n_1382),
.B2(n_1380),
.Y(n_1439)
);

OAI21x1_ASAP7_75t_L g1440 ( 
.A1(n_1367),
.A2(n_1378),
.B(n_1390),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1385),
.B(n_1386),
.Y(n_1441)
);

AO32x2_ASAP7_75t_L g1442 ( 
.A1(n_1345),
.A2(n_1401),
.A3(n_1400),
.B1(n_1404),
.B2(n_1386),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1347),
.Y(n_1443)
);

NAND3xp33_ASAP7_75t_L g1444 ( 
.A(n_1379),
.B(n_1369),
.C(n_1396),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1391),
.B(n_1393),
.Y(n_1445)
);

NAND2xp33_ASAP7_75t_SL g1446 ( 
.A(n_1395),
.B(n_1344),
.Y(n_1446)
);

O2A1O1Ixp33_ASAP7_75t_SL g1447 ( 
.A1(n_1352),
.A2(n_1405),
.B(n_1406),
.C(n_1361),
.Y(n_1447)
);

AOI211xp5_ASAP7_75t_L g1448 ( 
.A1(n_1395),
.A2(n_1391),
.B(n_1393),
.C(n_1373),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1419),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1443),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1424),
.B(n_1375),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1426),
.B(n_1375),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1407),
.B(n_1375),
.Y(n_1453)
);

OR2x2_ASAP7_75t_SL g1454 ( 
.A(n_1425),
.B(n_1375),
.Y(n_1454)
);

INVx4_ASAP7_75t_L g1455 ( 
.A(n_1436),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1419),
.B(n_1343),
.Y(n_1456)
);

NOR3xp33_ASAP7_75t_L g1457 ( 
.A(n_1433),
.B(n_1392),
.C(n_1367),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1440),
.B(n_1355),
.Y(n_1458)
);

INVx5_ASAP7_75t_L g1459 ( 
.A(n_1436),
.Y(n_1459)
);

BUFx2_ASAP7_75t_L g1460 ( 
.A(n_1427),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1414),
.B(n_1343),
.Y(n_1461)
);

HB1xp67_ASAP7_75t_L g1462 ( 
.A(n_1414),
.Y(n_1462)
);

BUFx2_ASAP7_75t_L g1463 ( 
.A(n_1427),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1440),
.B(n_1355),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1430),
.B(n_1355),
.Y(n_1465)
);

INVxp67_ASAP7_75t_SL g1466 ( 
.A(n_1437),
.Y(n_1466)
);

INVx1_ASAP7_75t_SL g1467 ( 
.A(n_1421),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1438),
.B(n_1350),
.Y(n_1468)
);

INVxp67_ASAP7_75t_L g1469 ( 
.A(n_1431),
.Y(n_1469)
);

HB1xp67_ASAP7_75t_L g1470 ( 
.A(n_1428),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1438),
.B(n_1346),
.Y(n_1471)
);

INVx2_ASAP7_75t_SL g1472 ( 
.A(n_1420),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1438),
.B(n_1346),
.Y(n_1473)
);

AOI22xp33_ASAP7_75t_L g1474 ( 
.A1(n_1444),
.A2(n_1364),
.B1(n_1337),
.B2(n_1403),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1438),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1470),
.Y(n_1476)
);

BUFx3_ASAP7_75t_L g1477 ( 
.A(n_1460),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1451),
.B(n_1453),
.Y(n_1478)
);

INVx5_ASAP7_75t_L g1479 ( 
.A(n_1459),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1449),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1449),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1451),
.B(n_1453),
.Y(n_1482)
);

INVx2_ASAP7_75t_SL g1483 ( 
.A(n_1471),
.Y(n_1483)
);

INVx2_ASAP7_75t_SL g1484 ( 
.A(n_1471),
.Y(n_1484)
);

AOI31xp33_ASAP7_75t_L g1485 ( 
.A1(n_1474),
.A2(n_1446),
.A3(n_1448),
.B(n_1447),
.Y(n_1485)
);

OAI33xp33_ASAP7_75t_L g1486 ( 
.A1(n_1475),
.A2(n_1439),
.A3(n_1429),
.B1(n_1418),
.B2(n_1422),
.B3(n_1423),
.Y(n_1486)
);

INVx3_ASAP7_75t_L g1487 ( 
.A(n_1458),
.Y(n_1487)
);

OA21x2_ASAP7_75t_L g1488 ( 
.A1(n_1458),
.A2(n_1411),
.B(n_1415),
.Y(n_1488)
);

INVx3_ASAP7_75t_L g1489 ( 
.A(n_1458),
.Y(n_1489)
);

NOR3xp33_ASAP7_75t_L g1490 ( 
.A(n_1457),
.B(n_1465),
.C(n_1446),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1473),
.B(n_1356),
.Y(n_1491)
);

INVx2_ASAP7_75t_SL g1492 ( 
.A(n_1473),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1468),
.Y(n_1493)
);

HB1xp67_ASAP7_75t_L g1494 ( 
.A(n_1462),
.Y(n_1494)
);

NAND3xp33_ASAP7_75t_L g1495 ( 
.A(n_1457),
.B(n_1410),
.C(n_1435),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1468),
.Y(n_1496)
);

INVx3_ASAP7_75t_L g1497 ( 
.A(n_1464),
.Y(n_1497)
);

AOI31xp67_ASAP7_75t_L g1498 ( 
.A1(n_1450),
.A2(n_1408),
.A3(n_1334),
.B(n_1338),
.Y(n_1498)
);

AOI22xp33_ASAP7_75t_SL g1499 ( 
.A1(n_1475),
.A2(n_1435),
.B1(n_1416),
.B2(n_1441),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1452),
.B(n_1445),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1452),
.B(n_1442),
.Y(n_1501)
);

INVx3_ASAP7_75t_L g1502 ( 
.A(n_1464),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1468),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1464),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1460),
.B(n_1442),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1466),
.B(n_1416),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1463),
.B(n_1442),
.Y(n_1507)
);

NOR2xp33_ASAP7_75t_L g1508 ( 
.A(n_1486),
.B(n_1469),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1478),
.B(n_1482),
.Y(n_1509)
);

OR2x2_ASAP7_75t_L g1510 ( 
.A(n_1501),
.B(n_1493),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1498),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1478),
.B(n_1463),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1498),
.Y(n_1513)
);

OR2x2_ASAP7_75t_L g1514 ( 
.A(n_1501),
.B(n_1466),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1478),
.B(n_1462),
.Y(n_1515)
);

AND2x4_ASAP7_75t_L g1516 ( 
.A(n_1483),
.B(n_1459),
.Y(n_1516)
);

OR2x2_ASAP7_75t_L g1517 ( 
.A(n_1501),
.B(n_1456),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1480),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1480),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1498),
.Y(n_1520)
);

INVx2_ASAP7_75t_SL g1521 ( 
.A(n_1491),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1483),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_SL g1523 ( 
.A(n_1490),
.B(n_1472),
.Y(n_1523)
);

NOR2x1_ASAP7_75t_L g1524 ( 
.A(n_1495),
.B(n_1417),
.Y(n_1524)
);

AND2x2_ASAP7_75t_SL g1525 ( 
.A(n_1490),
.B(n_1455),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1480),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1482),
.B(n_1469),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1476),
.B(n_1461),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1483),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1481),
.Y(n_1530)
);

BUFx3_ASAP7_75t_L g1531 ( 
.A(n_1479),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1481),
.Y(n_1532)
);

AOI22xp5_ASAP7_75t_L g1533 ( 
.A1(n_1486),
.A2(n_1441),
.B1(n_1397),
.B2(n_1410),
.Y(n_1533)
);

NAND2x1p5_ASAP7_75t_L g1534 ( 
.A(n_1479),
.B(n_1459),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1481),
.Y(n_1535)
);

INVxp67_ASAP7_75t_L g1536 ( 
.A(n_1495),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1476),
.B(n_1461),
.Y(n_1537)
);

BUFx2_ASAP7_75t_L g1538 ( 
.A(n_1477),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1476),
.B(n_1456),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1484),
.B(n_1467),
.Y(n_1540)
);

HB1xp67_ASAP7_75t_L g1541 ( 
.A(n_1477),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1509),
.B(n_1477),
.Y(n_1542)
);

NAND2x1p5_ASAP7_75t_L g1543 ( 
.A(n_1525),
.B(n_1479),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1509),
.B(n_1477),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1509),
.B(n_1484),
.Y(n_1545)
);

INVx2_ASAP7_75t_SL g1546 ( 
.A(n_1538),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1518),
.Y(n_1547)
);

HB1xp67_ASAP7_75t_L g1548 ( 
.A(n_1541),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1518),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1519),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1524),
.B(n_1484),
.Y(n_1551)
);

INVx6_ASAP7_75t_L g1552 ( 
.A(n_1531),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1510),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1519),
.Y(n_1554)
);

INVxp67_ASAP7_75t_SL g1555 ( 
.A(n_1536),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1524),
.B(n_1484),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1510),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1536),
.B(n_1501),
.Y(n_1558)
);

INVx4_ASAP7_75t_L g1559 ( 
.A(n_1525),
.Y(n_1559)
);

A2O1A1Ixp33_ASAP7_75t_L g1560 ( 
.A1(n_1508),
.A2(n_1485),
.B(n_1507),
.C(n_1505),
.Y(n_1560)
);

NAND2x2_ASAP7_75t_L g1561 ( 
.A(n_1531),
.B(n_1341),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1510),
.Y(n_1562)
);

OR2x6_ASAP7_75t_L g1563 ( 
.A(n_1534),
.B(n_1413),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1526),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1526),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1530),
.Y(n_1566)
);

HB1xp67_ASAP7_75t_L g1567 ( 
.A(n_1541),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1508),
.B(n_1500),
.Y(n_1568)
);

INVxp67_ASAP7_75t_L g1569 ( 
.A(n_1533),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1530),
.Y(n_1570)
);

OR2x2_ASAP7_75t_L g1571 ( 
.A(n_1514),
.B(n_1517),
.Y(n_1571)
);

INVx2_ASAP7_75t_SL g1572 ( 
.A(n_1538),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1532),
.Y(n_1573)
);

OAI21xp33_ASAP7_75t_L g1574 ( 
.A1(n_1523),
.A2(n_1487),
.B(n_1489),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1532),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1527),
.B(n_1492),
.Y(n_1576)
);

OA21x2_ASAP7_75t_SL g1577 ( 
.A1(n_1523),
.A2(n_1467),
.B(n_1485),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1533),
.B(n_1527),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1522),
.Y(n_1579)
);

NOR2xp33_ASAP7_75t_L g1580 ( 
.A(n_1527),
.B(n_1344),
.Y(n_1580)
);

AND2x4_ASAP7_75t_L g1581 ( 
.A(n_1516),
.B(n_1492),
.Y(n_1581)
);

OR2x2_ASAP7_75t_L g1582 ( 
.A(n_1514),
.B(n_1493),
.Y(n_1582)
);

OR2x2_ASAP7_75t_L g1583 ( 
.A(n_1514),
.B(n_1493),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1555),
.B(n_1568),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1559),
.B(n_1525),
.Y(n_1585)
);

AND2x4_ASAP7_75t_L g1586 ( 
.A(n_1559),
.B(n_1516),
.Y(n_1586)
);

NAND2x1p5_ASAP7_75t_L g1587 ( 
.A(n_1559),
.B(n_1479),
.Y(n_1587)
);

OAI21xp5_ASAP7_75t_SL g1588 ( 
.A1(n_1560),
.A2(n_1489),
.B(n_1487),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1549),
.Y(n_1589)
);

AOI221xp5_ASAP7_75t_L g1590 ( 
.A1(n_1569),
.A2(n_1520),
.B1(n_1513),
.B2(n_1511),
.C(n_1505),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1542),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1546),
.B(n_1500),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1546),
.B(n_1500),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1572),
.B(n_1500),
.Y(n_1594)
);

OAI211xp5_ASAP7_75t_L g1595 ( 
.A1(n_1578),
.A2(n_1531),
.B(n_1487),
.C(n_1489),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1549),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1554),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1543),
.B(n_1525),
.Y(n_1598)
);

NAND2x1_ASAP7_75t_L g1599 ( 
.A(n_1552),
.B(n_1551),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1543),
.B(n_1551),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1543),
.B(n_1556),
.Y(n_1601)
);

INVxp67_ASAP7_75t_L g1602 ( 
.A(n_1580),
.Y(n_1602)
);

OAI21xp33_ASAP7_75t_L g1603 ( 
.A1(n_1558),
.A2(n_1489),
.B(n_1487),
.Y(n_1603)
);

OR2x2_ASAP7_75t_L g1604 ( 
.A(n_1571),
.B(n_1517),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1572),
.B(n_1515),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1548),
.B(n_1515),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1542),
.Y(n_1607)
);

NOR2x1_ASAP7_75t_L g1608 ( 
.A(n_1556),
.B(n_1516),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1544),
.B(n_1576),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1544),
.B(n_1512),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1567),
.B(n_1515),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1554),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1576),
.B(n_1505),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1564),
.Y(n_1614)
);

OR2x2_ASAP7_75t_L g1615 ( 
.A(n_1571),
.B(n_1517),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1564),
.Y(n_1616)
);

OAI22xp5_ASAP7_75t_L g1617 ( 
.A1(n_1577),
.A2(n_1454),
.B1(n_1492),
.B2(n_1488),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1575),
.Y(n_1618)
);

OAI32xp33_ASAP7_75t_L g1619 ( 
.A1(n_1617),
.A2(n_1574),
.A3(n_1561),
.B1(n_1562),
.B2(n_1557),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1609),
.B(n_1545),
.Y(n_1620)
);

AOI21xp5_ASAP7_75t_L g1621 ( 
.A1(n_1584),
.A2(n_1507),
.B(n_1505),
.Y(n_1621)
);

A2O1A1Ixp33_ASAP7_75t_L g1622 ( 
.A1(n_1590),
.A2(n_1507),
.B(n_1513),
.C(n_1511),
.Y(n_1622)
);

INVx1_ASAP7_75t_SL g1623 ( 
.A(n_1585),
.Y(n_1623)
);

AOI22xp5_ASAP7_75t_L g1624 ( 
.A1(n_1588),
.A2(n_1507),
.B1(n_1499),
.B2(n_1488),
.Y(n_1624)
);

INVx1_ASAP7_75t_SL g1625 ( 
.A(n_1585),
.Y(n_1625)
);

NAND3xp33_ASAP7_75t_L g1626 ( 
.A(n_1599),
.B(n_1513),
.C(n_1511),
.Y(n_1626)
);

AOI21xp33_ASAP7_75t_L g1627 ( 
.A1(n_1599),
.A2(n_1579),
.B(n_1557),
.Y(n_1627)
);

AOI21xp33_ASAP7_75t_L g1628 ( 
.A1(n_1597),
.A2(n_1579),
.B(n_1562),
.Y(n_1628)
);

HB1xp67_ASAP7_75t_L g1629 ( 
.A(n_1591),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1597),
.Y(n_1630)
);

OAI21xp5_ASAP7_75t_L g1631 ( 
.A1(n_1595),
.A2(n_1520),
.B(n_1581),
.Y(n_1631)
);

HB1xp67_ASAP7_75t_L g1632 ( 
.A(n_1591),
.Y(n_1632)
);

OAI21xp5_ASAP7_75t_L g1633 ( 
.A1(n_1602),
.A2(n_1520),
.B(n_1581),
.Y(n_1633)
);

NOR3xp33_ASAP7_75t_SL g1634 ( 
.A(n_1603),
.B(n_1605),
.C(n_1606),
.Y(n_1634)
);

INVxp67_ASAP7_75t_SL g1635 ( 
.A(n_1587),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_SL g1636 ( 
.A(n_1586),
.B(n_1581),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1589),
.Y(n_1637)
);

O2A1O1Ixp33_ASAP7_75t_L g1638 ( 
.A1(n_1618),
.A2(n_1502),
.B(n_1487),
.C(n_1489),
.Y(n_1638)
);

NOR2xp33_ASAP7_75t_L g1639 ( 
.A(n_1607),
.B(n_1609),
.Y(n_1639)
);

AOI32xp33_ASAP7_75t_L g1640 ( 
.A1(n_1598),
.A2(n_1553),
.A3(n_1487),
.B1(n_1489),
.B2(n_1497),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1596),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1612),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1607),
.B(n_1553),
.Y(n_1643)
);

OR2x2_ASAP7_75t_L g1644 ( 
.A(n_1623),
.B(n_1625),
.Y(n_1644)
);

OAI221xp5_ASAP7_75t_L g1645 ( 
.A1(n_1622),
.A2(n_1608),
.B1(n_1587),
.B2(n_1604),
.C(n_1615),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1639),
.B(n_1610),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1620),
.B(n_1610),
.Y(n_1647)
);

INVxp67_ASAP7_75t_L g1648 ( 
.A(n_1629),
.Y(n_1648)
);

INVxp67_ASAP7_75t_L g1649 ( 
.A(n_1632),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1630),
.Y(n_1650)
);

AOI221xp5_ASAP7_75t_L g1651 ( 
.A1(n_1622),
.A2(n_1616),
.B1(n_1614),
.B2(n_1613),
.C(n_1604),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1637),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1641),
.Y(n_1653)
);

AOI22xp5_ASAP7_75t_L g1654 ( 
.A1(n_1624),
.A2(n_1488),
.B1(n_1601),
.B2(n_1600),
.Y(n_1654)
);

INVxp67_ASAP7_75t_SL g1655 ( 
.A(n_1626),
.Y(n_1655)
);

A2O1A1Ixp33_ASAP7_75t_L g1656 ( 
.A1(n_1621),
.A2(n_1598),
.B(n_1601),
.C(n_1600),
.Y(n_1656)
);

OAI32xp33_ASAP7_75t_L g1657 ( 
.A1(n_1627),
.A2(n_1615),
.A3(n_1587),
.B1(n_1611),
.B2(n_1561),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1620),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1639),
.B(n_1586),
.Y(n_1659)
);

OAI221xp5_ASAP7_75t_L g1660 ( 
.A1(n_1633),
.A2(n_1499),
.B1(n_1552),
.B2(n_1582),
.C(n_1583),
.Y(n_1660)
);

AND2x2_ASAP7_75t_SL g1661 ( 
.A(n_1643),
.B(n_1586),
.Y(n_1661)
);

OR2x2_ASAP7_75t_L g1662 ( 
.A(n_1636),
.B(n_1592),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1647),
.B(n_1642),
.Y(n_1663)
);

A2O1A1Ixp33_ASAP7_75t_L g1664 ( 
.A1(n_1655),
.A2(n_1619),
.B(n_1634),
.C(n_1628),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1644),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1658),
.Y(n_1666)
);

AOI222xp33_ASAP7_75t_L g1667 ( 
.A1(n_1655),
.A2(n_1631),
.B1(n_1635),
.B2(n_1636),
.C1(n_1506),
.C2(n_1397),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1648),
.Y(n_1668)
);

AOI221xp5_ASAP7_75t_L g1669 ( 
.A1(n_1651),
.A2(n_1640),
.B1(n_1638),
.B2(n_1575),
.C(n_1506),
.Y(n_1669)
);

AOI221xp5_ASAP7_75t_L g1670 ( 
.A1(n_1651),
.A2(n_1504),
.B1(n_1547),
.B2(n_1565),
.C(n_1550),
.Y(n_1670)
);

AOI21xp33_ASAP7_75t_L g1671 ( 
.A1(n_1648),
.A2(n_1570),
.B(n_1566),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_SL g1672 ( 
.A(n_1661),
.B(n_1516),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1646),
.B(n_1649),
.Y(n_1673)
);

OAI221xp5_ASAP7_75t_L g1674 ( 
.A1(n_1654),
.A2(n_1552),
.B1(n_1582),
.B2(n_1583),
.C(n_1563),
.Y(n_1674)
);

HB1xp67_ASAP7_75t_L g1675 ( 
.A(n_1665),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1663),
.Y(n_1676)
);

NAND3xp33_ASAP7_75t_L g1677 ( 
.A(n_1664),
.B(n_1649),
.C(n_1645),
.Y(n_1677)
);

NOR2x1_ASAP7_75t_L g1678 ( 
.A(n_1668),
.B(n_1650),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1666),
.Y(n_1679)
);

NAND3xp33_ASAP7_75t_L g1680 ( 
.A(n_1667),
.B(n_1653),
.C(n_1652),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1673),
.Y(n_1681)
);

OAI21xp33_ASAP7_75t_SL g1682 ( 
.A1(n_1670),
.A2(n_1659),
.B(n_1662),
.Y(n_1682)
);

INVxp67_ASAP7_75t_L g1683 ( 
.A(n_1672),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1675),
.B(n_1656),
.Y(n_1684)
);

OAI221xp5_ASAP7_75t_L g1685 ( 
.A1(n_1677),
.A2(n_1660),
.B1(n_1674),
.B2(n_1669),
.C(n_1671),
.Y(n_1685)
);

NOR2xp33_ASAP7_75t_R g1686 ( 
.A(n_1681),
.B(n_1368),
.Y(n_1686)
);

NAND4xp75_ASAP7_75t_L g1687 ( 
.A(n_1678),
.B(n_1657),
.C(n_1594),
.D(n_1593),
.Y(n_1687)
);

NAND4xp25_ASAP7_75t_L g1688 ( 
.A(n_1680),
.B(n_1545),
.C(n_1341),
.D(n_1398),
.Y(n_1688)
);

AOI211xp5_ASAP7_75t_L g1689 ( 
.A1(n_1685),
.A2(n_1682),
.B(n_1679),
.C(n_1676),
.Y(n_1689)
);

OAI21xp5_ASAP7_75t_L g1690 ( 
.A1(n_1687),
.A2(n_1683),
.B(n_1522),
.Y(n_1690)
);

INVx2_ASAP7_75t_SL g1691 ( 
.A(n_1686),
.Y(n_1691)
);

OAI22xp5_ASAP7_75t_L g1692 ( 
.A1(n_1684),
.A2(n_1552),
.B1(n_1529),
.B2(n_1522),
.Y(n_1692)
);

XNOR2x1_ASAP7_75t_L g1693 ( 
.A(n_1688),
.B(n_1563),
.Y(n_1693)
);

AOI211xp5_ASAP7_75t_SL g1694 ( 
.A1(n_1684),
.A2(n_1447),
.B(n_1573),
.C(n_1529),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1693),
.Y(n_1695)
);

AOI22xp33_ASAP7_75t_L g1696 ( 
.A1(n_1691),
.A2(n_1488),
.B1(n_1563),
.B2(n_1516),
.Y(n_1696)
);

AOI22xp5_ASAP7_75t_L g1697 ( 
.A1(n_1689),
.A2(n_1563),
.B1(n_1512),
.B2(n_1529),
.Y(n_1697)
);

NOR2x1_ASAP7_75t_L g1698 ( 
.A(n_1690),
.B(n_1540),
.Y(n_1698)
);

NOR2x1_ASAP7_75t_L g1699 ( 
.A(n_1692),
.B(n_1540),
.Y(n_1699)
);

OAI221xp5_ASAP7_75t_L g1700 ( 
.A1(n_1698),
.A2(n_1694),
.B1(n_1492),
.B2(n_1534),
.C(n_1496),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1699),
.Y(n_1701)
);

OR2x2_ASAP7_75t_L g1702 ( 
.A(n_1697),
.B(n_1528),
.Y(n_1702)
);

CKINVDCx20_ASAP7_75t_R g1703 ( 
.A(n_1701),
.Y(n_1703)
);

AOI22xp5_ASAP7_75t_SL g1704 ( 
.A1(n_1703),
.A2(n_1695),
.B1(n_1700),
.B2(n_1702),
.Y(n_1704)
);

XNOR2xp5_ASAP7_75t_L g1705 ( 
.A(n_1704),
.B(n_1696),
.Y(n_1705)
);

OAI22x1_ASAP7_75t_SL g1706 ( 
.A1(n_1705),
.A2(n_1521),
.B1(n_1503),
.B2(n_1496),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1706),
.Y(n_1707)
);

OAI221xp5_ASAP7_75t_L g1708 ( 
.A1(n_1707),
.A2(n_1534),
.B1(n_1535),
.B2(n_1537),
.C(n_1497),
.Y(n_1708)
);

AOI21xp33_ASAP7_75t_SL g1709 ( 
.A1(n_1708),
.A2(n_1534),
.B(n_1434),
.Y(n_1709)
);

INVxp67_ASAP7_75t_L g1710 ( 
.A(n_1709),
.Y(n_1710)
);

OAI221xp5_ASAP7_75t_R g1711 ( 
.A1(n_1710),
.A2(n_1494),
.B1(n_1521),
.B2(n_1512),
.C(n_1539),
.Y(n_1711)
);

AOI211xp5_ASAP7_75t_L g1712 ( 
.A1(n_1711),
.A2(n_1409),
.B(n_1432),
.C(n_1412),
.Y(n_1712)
);


endmodule