module fake_jpeg_3485_n_493 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_493);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_493;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx8_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx8_ASAP7_75t_SL g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx24_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_15),
.B(n_13),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx8_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

INVx6_ASAP7_75t_SL g37 ( 
.A(n_14),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_17),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_13),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_11),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_13),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

INVx11_ASAP7_75t_SL g46 ( 
.A(n_12),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_4),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_13),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_7),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_34),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_55),
.B(n_65),
.Y(n_131)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_56),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_57),
.Y(n_122)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_58),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_59),
.Y(n_125)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_60),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

INVx5_ASAP7_75t_L g203 ( 
.A(n_61),
.Y(n_203)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_62),
.Y(n_147)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_63),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_64),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_34),
.B(n_16),
.C(n_1),
.Y(n_65)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

BUFx4f_ASAP7_75t_SL g152 ( 
.A(n_66),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_22),
.B(n_16),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_67),
.B(n_84),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_32),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_68),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_69),
.Y(n_136)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_20),
.Y(n_70)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_70),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_71),
.Y(n_167)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_72),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_32),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_73),
.Y(n_168)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_20),
.Y(n_74)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_74),
.Y(n_194)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_19),
.Y(n_75)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_75),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_30),
.B(n_0),
.Y(n_76)
);

OAI21xp33_ASAP7_75t_L g179 ( 
.A1(n_76),
.A2(n_83),
.B(n_90),
.Y(n_179)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_77),
.Y(n_196)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_19),
.Y(n_78)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_78),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_79),
.Y(n_202)
);

BUFx8_ASAP7_75t_L g80 ( 
.A(n_26),
.Y(n_80)
);

BUFx5_ASAP7_75t_L g182 ( 
.A(n_80),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_26),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_81),
.Y(n_172)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_82),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_30),
.B(n_0),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_38),
.B(n_14),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_85),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_38),
.B(n_0),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_86),
.B(n_87),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_18),
.B(n_12),
.Y(n_87)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_19),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g146 ( 
.A(n_88),
.Y(n_146)
);

BUFx24_ASAP7_75t_L g89 ( 
.A(n_26),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g158 ( 
.A(n_89),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_28),
.B(n_1),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_41),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_91),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_28),
.B(n_1),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_92),
.B(n_94),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_41),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_93),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_33),
.B(n_39),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

INVx6_ASAP7_75t_L g178 ( 
.A(n_95),
.Y(n_178)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_96),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_47),
.Y(n_97)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_97),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_27),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_98),
.B(n_103),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_47),
.Y(n_99)
);

INVx8_ASAP7_75t_L g137 ( 
.A(n_99),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_36),
.Y(n_100)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_100),
.Y(n_171)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_50),
.Y(n_101)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_101),
.Y(n_132)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_102),
.Y(n_195)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_36),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_36),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_104),
.B(n_109),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_33),
.B(n_2),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_105),
.B(n_24),
.Y(n_155)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_52),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_106),
.B(n_112),
.Y(n_164)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_23),
.Y(n_107)
);

INVx2_ASAP7_75t_R g199 ( 
.A(n_107),
.Y(n_199)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_54),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_108),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_36),
.Y(n_109)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_52),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_110),
.B(n_113),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_54),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_111),
.Y(n_141)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_52),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g113 ( 
.A(n_27),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_18),
.B(n_2),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_114),
.B(n_115),
.Y(n_170)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_52),
.Y(n_115)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_52),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_116),
.B(n_118),
.Y(n_166)
);

INVx11_ASAP7_75t_L g117 ( 
.A(n_31),
.Y(n_117)
);

AOI21xp33_ASAP7_75t_L g126 ( 
.A1(n_117),
.A2(n_31),
.B(n_45),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_54),
.Y(n_118)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_35),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_119),
.B(n_120),
.Y(n_173)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_31),
.Y(n_120)
);

AOI21xp33_ASAP7_75t_L g257 ( 
.A1(n_126),
.A2(n_182),
.B(n_199),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_63),
.A2(n_29),
.B1(n_51),
.B2(n_49),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_128),
.A2(n_129),
.B1(n_180),
.B2(n_179),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_108),
.A2(n_29),
.B1(n_51),
.B2(n_49),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_90),
.A2(n_24),
.B1(n_48),
.B2(n_44),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_130),
.A2(n_145),
.B1(n_151),
.B2(n_157),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_92),
.A2(n_53),
.B(n_45),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_134),
.B(n_191),
.C(n_138),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_105),
.B(n_53),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_139),
.B(n_143),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_80),
.A2(n_35),
.B1(n_43),
.B2(n_44),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_140),
.A2(n_162),
.B1(n_190),
.B2(n_192),
.Y(n_211)
);

NOR2x1_ASAP7_75t_L g142 ( 
.A(n_94),
.B(n_83),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g225 ( 
.A(n_142),
.B(n_135),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_76),
.B(n_43),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_57),
.A2(n_42),
.B1(n_40),
.B2(n_39),
.Y(n_145)
);

OA22x2_ASAP7_75t_L g148 ( 
.A1(n_59),
.A2(n_31),
.B1(n_23),
.B2(n_4),
.Y(n_148)
);

AO22x2_ASAP7_75t_L g256 ( 
.A1(n_148),
.A2(n_171),
.B1(n_127),
.B2(n_121),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_68),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_149),
.B(n_153),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_71),
.A2(n_48),
.B1(n_42),
.B2(n_40),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_73),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_155),
.B(n_179),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_85),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_91),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_161),
.A2(n_165),
.B1(n_180),
.B2(n_183),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_104),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_93),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_61),
.B(n_9),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_169),
.B(n_175),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_60),
.B(n_9),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_104),
.B(n_10),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_177),
.B(n_181),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_95),
.A2(n_11),
.B1(n_12),
.B2(n_99),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_62),
.B(n_11),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_97),
.A2(n_111),
.B1(n_118),
.B2(n_89),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_88),
.A2(n_102),
.B1(n_120),
.B2(n_113),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_187),
.A2(n_158),
.B1(n_152),
.B2(n_161),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_113),
.B(n_66),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_189),
.B(n_200),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_80),
.A2(n_36),
.B1(n_26),
.B2(n_46),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_90),
.B(n_92),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_191),
.B(n_142),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_80),
.A2(n_36),
.B1(n_26),
.B2(n_46),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_55),
.B(n_94),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_94),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_201),
.B(n_200),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_204),
.B(n_207),
.Y(n_274)
);

INVx13_ASAP7_75t_L g205 ( 
.A(n_152),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_205),
.Y(n_278)
);

CKINVDCx14_ASAP7_75t_R g207 ( 
.A(n_160),
.Y(n_207)
);

OAI22xp33_ASAP7_75t_SL g299 ( 
.A1(n_209),
.A2(n_225),
.B1(n_244),
.B2(n_211),
.Y(n_299)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_150),
.Y(n_210)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_210),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_164),
.B(n_170),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_212),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_152),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_213),
.B(n_216),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_128),
.A2(n_129),
.B1(n_148),
.B2(n_158),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_214),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_176),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_186),
.Y(n_217)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_217),
.Y(n_277)
);

BUFx2_ASAP7_75t_L g218 ( 
.A(n_172),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g303 ( 
.A(n_218),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_219),
.B(n_221),
.Y(n_289)
);

OAI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_139),
.A2(n_143),
.B1(n_148),
.B2(n_124),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_222),
.A2(n_264),
.B1(n_272),
.B2(n_220),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_L g287 ( 
.A1(n_223),
.A2(n_208),
.B1(n_233),
.B2(n_258),
.Y(n_287)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_158),
.Y(n_224)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_224),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_225),
.B(n_233),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_131),
.A2(n_173),
.B1(n_148),
.B2(n_134),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_226),
.A2(n_257),
.B(n_221),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_123),
.B(n_159),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_227),
.B(n_260),
.Y(n_318)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_147),
.Y(n_228)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_228),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_176),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_229),
.B(n_241),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_122),
.Y(n_230)
);

INVx5_ASAP7_75t_L g288 ( 
.A(n_230),
.Y(n_288)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_150),
.Y(n_231)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_231),
.Y(n_291)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_196),
.Y(n_232)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_232),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_166),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_186),
.Y(n_234)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_234),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_132),
.B(n_198),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_235),
.B(n_255),
.Y(n_273)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_195),
.Y(n_238)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_238),
.Y(n_310)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_195),
.Y(n_239)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_239),
.Y(n_311)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_196),
.Y(n_240)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_240),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_163),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_141),
.A2(n_178),
.B1(n_122),
.B2(n_125),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_242),
.A2(n_252),
.B1(n_256),
.B2(n_265),
.Y(n_319)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_197),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_243),
.B(n_248),
.Y(n_301)
);

OR2x2_ASAP7_75t_L g244 ( 
.A(n_121),
.B(n_199),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_244),
.B(n_245),
.Y(n_316)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_197),
.Y(n_245)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_147),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_246),
.Y(n_276)
);

INVx5_ASAP7_75t_L g247 ( 
.A(n_172),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_247),
.Y(n_280)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_198),
.Y(n_248)
);

INVx4_ASAP7_75t_L g249 ( 
.A(n_203),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_249),
.Y(n_283)
);

INVx5_ASAP7_75t_L g250 ( 
.A(n_146),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_250),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_178),
.A2(n_168),
.B1(n_125),
.B2(n_188),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_154),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_253),
.B(n_261),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_171),
.A2(n_127),
.B1(n_194),
.B2(n_154),
.Y(n_254)
);

OAI22xp33_ASAP7_75t_L g322 ( 
.A1(n_254),
.A2(n_262),
.B1(n_267),
.B2(n_224),
.Y(n_322)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_203),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_194),
.B(n_144),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_258),
.B(n_259),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_144),
.B(n_167),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_156),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_174),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_202),
.A2(n_136),
.B1(n_184),
.B2(n_174),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_156),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_263),
.B(n_268),
.Y(n_309)
);

BUFx2_ASAP7_75t_L g264 ( 
.A(n_136),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_167),
.A2(n_193),
.B1(n_168),
.B2(n_188),
.Y(n_265)
);

A2O1A1Ixp33_ASAP7_75t_L g266 ( 
.A1(n_182),
.A2(n_184),
.B(n_202),
.C(n_146),
.Y(n_266)
);

A2O1A1Ixp33_ASAP7_75t_L g306 ( 
.A1(n_266),
.A2(n_256),
.B(n_216),
.C(n_270),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_146),
.A2(n_133),
.B1(n_137),
.B2(n_185),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_133),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_137),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_269),
.B(n_270),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_185),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_193),
.B(n_191),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_271),
.B(n_259),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_226),
.A2(n_209),
.B1(n_271),
.B2(n_212),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_275),
.A2(n_281),
.B1(n_292),
.B2(n_297),
.Y(n_337)
);

MAJx2_ASAP7_75t_L g279 ( 
.A(n_212),
.B(n_219),
.C(n_220),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_279),
.B(n_302),
.C(n_293),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_282),
.B(n_299),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_287),
.A2(n_320),
.B1(n_253),
.B2(n_261),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_292),
.A2(n_293),
.B(n_304),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_215),
.A2(n_206),
.B1(n_241),
.B2(n_251),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_296),
.B(n_312),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_235),
.B(n_236),
.C(n_248),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_266),
.A2(n_237),
.B(n_256),
.Y(n_304)
);

O2A1O1Ixp33_ASAP7_75t_L g341 ( 
.A1(n_306),
.A2(n_273),
.B(n_285),
.C(n_289),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_238),
.B(n_239),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_240),
.B(n_243),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_313),
.B(n_314),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_210),
.B(n_231),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_217),
.B(n_234),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_317),
.B(n_269),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_256),
.A2(n_245),
.B1(n_232),
.B2(n_268),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_SL g355 ( 
.A1(n_322),
.A2(n_280),
.B1(n_283),
.B2(n_284),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_323),
.A2(n_335),
.B1(n_346),
.B2(n_276),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_318),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_325),
.B(n_329),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_312),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_286),
.Y(n_329)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_303),
.Y(n_330)
);

INVx4_ASAP7_75t_L g366 ( 
.A(n_330),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_318),
.B(n_298),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g386 ( 
.A(n_331),
.B(n_332),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_298),
.B(n_228),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_334),
.B(n_336),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_282),
.A2(n_230),
.B1(n_246),
.B2(n_218),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_296),
.B(n_255),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_337),
.B(n_347),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_275),
.A2(n_316),
.B1(n_274),
.B2(n_273),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_SL g376 ( 
.A1(n_338),
.A2(n_340),
.B(n_284),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_306),
.A2(n_264),
.B1(n_247),
.B2(n_249),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_339),
.A2(n_353),
.B1(n_276),
.B2(n_283),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_304),
.A2(n_205),
.B(n_250),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_341),
.B(n_345),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_302),
.B(n_295),
.Y(n_342)
);

CKINVDCx14_ASAP7_75t_R g368 ( 
.A(n_342),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_343),
.B(n_359),
.C(n_360),
.Y(n_388)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_286),
.Y(n_344)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_344),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_285),
.B(n_289),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_319),
.A2(n_320),
.B1(n_279),
.B2(n_274),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_SL g347 ( 
.A(n_290),
.B(n_279),
.Y(n_347)
);

BUFx12f_ASAP7_75t_L g348 ( 
.A(n_294),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_310),
.Y(n_349)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_349),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_313),
.B(n_317),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_350),
.B(n_351),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_301),
.B(n_309),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_310),
.Y(n_352)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_352),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_319),
.A2(n_309),
.B1(n_301),
.B2(n_311),
.Y(n_353)
);

CKINVDCx16_ASAP7_75t_R g354 ( 
.A(n_290),
.Y(n_354)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_354),
.Y(n_372)
);

OAI21xp33_ASAP7_75t_SL g385 ( 
.A1(n_355),
.A2(n_294),
.B(n_303),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_311),
.B(n_314),
.Y(n_356)
);

OR2x2_ASAP7_75t_L g381 ( 
.A(n_356),
.B(n_357),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_305),
.B(n_321),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_305),
.Y(n_358)
);

CKINVDCx16_ASAP7_75t_R g389 ( 
.A(n_358),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_277),
.B(n_321),
.C(n_308),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_277),
.B(n_308),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_362),
.A2(n_367),
.B1(n_373),
.B2(n_378),
.Y(n_395)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_349),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_353),
.A2(n_338),
.B1(n_337),
.B2(n_326),
.Y(n_367)
);

INVx1_ASAP7_75t_SL g369 ( 
.A(n_340),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_369),
.B(n_371),
.Y(n_396)
);

OAI32xp33_ASAP7_75t_L g371 ( 
.A1(n_347),
.A2(n_315),
.A3(n_291),
.B1(n_300),
.B2(n_307),
.Y(n_371)
);

NOR2x1_ASAP7_75t_L g375 ( 
.A(n_327),
.B(n_315),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_375),
.B(n_379),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_376),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_346),
.A2(n_280),
.B1(n_288),
.B2(n_291),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_377),
.A2(n_387),
.B1(n_358),
.B2(n_334),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_329),
.A2(n_288),
.B1(n_300),
.B2(n_307),
.Y(n_378)
);

AND2x6_ASAP7_75t_L g379 ( 
.A(n_343),
.B(n_278),
.Y(n_379)
);

AND2x6_ASAP7_75t_L g380 ( 
.A(n_333),
.B(n_278),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_380),
.B(n_341),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_385),
.A2(n_335),
.B1(n_354),
.B2(n_352),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_323),
.A2(n_344),
.B1(n_339),
.B2(n_336),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_390),
.A2(n_402),
.B1(n_407),
.B2(n_409),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_388),
.B(n_345),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_391),
.B(n_397),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_389),
.B(n_359),
.Y(n_392)
);

INVxp33_ASAP7_75t_L g424 ( 
.A(n_392),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_388),
.B(n_342),
.C(n_333),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_393),
.B(n_413),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_389),
.B(n_332),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_394),
.B(n_370),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_383),
.B(n_324),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_376),
.A2(n_341),
.B(n_327),
.Y(n_398)
);

AOI21xp33_ASAP7_75t_L g415 ( 
.A1(n_398),
.A2(n_382),
.B(n_369),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g421 ( 
.A(n_399),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_374),
.Y(n_401)
);

NOR3xp33_ASAP7_75t_L g432 ( 
.A(n_401),
.B(n_361),
.C(n_363),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_362),
.A2(n_324),
.B1(n_350),
.B2(n_328),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_364),
.Y(n_403)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_403),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_404),
.B(n_375),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g405 ( 
.A(n_366),
.Y(n_405)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_405),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g407 ( 
.A1(n_387),
.A2(n_328),
.B1(n_327),
.B2(n_356),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_365),
.Y(n_408)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_408),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_367),
.A2(n_351),
.B1(n_331),
.B2(n_357),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_373),
.A2(n_360),
.B1(n_330),
.B2(n_348),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_410),
.B(n_377),
.Y(n_414)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_386),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_411),
.B(n_386),
.Y(n_417)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_365),
.Y(n_412)
);

INVx1_ASAP7_75t_SL g423 ( 
.A(n_412),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_383),
.B(n_348),
.C(n_368),
.Y(n_413)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_414),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_L g444 ( 
.A1(n_415),
.A2(n_400),
.B(n_396),
.Y(n_444)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_417),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_401),
.B(n_382),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_418),
.B(n_419),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_413),
.B(n_372),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_SL g422 ( 
.A(n_397),
.B(n_384),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_SL g442 ( 
.A(n_422),
.B(n_363),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_391),
.B(n_384),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_426),
.B(n_371),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_409),
.B(n_381),
.Y(n_427)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_427),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_392),
.B(n_372),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_429),
.B(n_432),
.Y(n_445)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_430),
.Y(n_440)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_433),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_434),
.B(n_393),
.C(n_406),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_435),
.B(n_434),
.C(n_426),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_431),
.A2(n_395),
.B1(n_399),
.B2(n_398),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_437),
.A2(n_430),
.B1(n_396),
.B2(n_427),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_L g438 ( 
.A1(n_431),
.A2(n_395),
.B1(n_402),
.B2(n_404),
.Y(n_438)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_438),
.Y(n_462)
);

AOI321xp33_ASAP7_75t_L g441 ( 
.A1(n_424),
.A2(n_379),
.A3(n_407),
.B1(n_394),
.B2(n_361),
.C(n_380),
.Y(n_441)
);

OAI21xp33_ASAP7_75t_L g457 ( 
.A1(n_441),
.A2(n_381),
.B(n_375),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_442),
.B(n_443),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_L g451 ( 
.A1(n_444),
.A2(n_415),
.B(n_430),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_416),
.B(n_406),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_447),
.B(n_414),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_416),
.B(n_390),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_448),
.B(n_435),
.Y(n_454)
);

OR2x2_ASAP7_75t_L g472 ( 
.A(n_451),
.B(n_443),
.Y(n_472)
);

HB1xp67_ASAP7_75t_L g464 ( 
.A(n_453),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_454),
.B(n_456),
.C(n_460),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_L g467 ( 
.A1(n_455),
.A2(n_457),
.B1(n_461),
.B2(n_440),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_447),
.B(n_421),
.C(n_422),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_436),
.B(n_425),
.Y(n_458)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_458),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_SL g459 ( 
.A(n_449),
.B(n_425),
.Y(n_459)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_459),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_439),
.A2(n_410),
.B1(n_381),
.B2(n_423),
.Y(n_461)
);

AOI221xp5_ASAP7_75t_L g463 ( 
.A1(n_451),
.A2(n_446),
.B1(n_440),
.B2(n_455),
.C(n_444),
.Y(n_463)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_463),
.Y(n_475)
);

OAI221xp5_ASAP7_75t_L g466 ( 
.A1(n_453),
.A2(n_450),
.B1(n_445),
.B2(n_441),
.C(n_442),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_466),
.B(n_456),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_467),
.B(n_448),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_462),
.A2(n_450),
.B1(n_437),
.B2(n_439),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_468),
.B(n_423),
.Y(n_476)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_461),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_470),
.B(n_460),
.Y(n_473)
);

INVxp67_ASAP7_75t_SL g477 ( 
.A(n_472),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_473),
.B(n_476),
.Y(n_484)
);

OAI21x1_ASAP7_75t_SL g480 ( 
.A1(n_474),
.A2(n_465),
.B(n_464),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_472),
.A2(n_420),
.B1(n_428),
.B2(n_452),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_478),
.B(n_477),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_479),
.B(n_454),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_480),
.B(n_481),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_475),
.B(n_469),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_482),
.B(n_471),
.C(n_479),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_483),
.A2(n_474),
.B1(n_481),
.B2(n_484),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_485),
.B(n_487),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_485),
.B(n_471),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_489),
.B(n_486),
.C(n_487),
.Y(n_490)
);

AOI21xp5_ASAP7_75t_L g491 ( 
.A1(n_490),
.A2(n_488),
.B(n_478),
.Y(n_491)
);

AOI21xp5_ASAP7_75t_L g492 ( 
.A1(n_491),
.A2(n_452),
.B(n_420),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g493 ( 
.A(n_492),
.Y(n_493)
);


endmodule