module fake_ariane_2457_n_2110 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_213, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_208, n_96, n_156, n_209, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_200, n_51, n_166, n_76, n_218, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_217, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_214, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_211, n_194, n_97, n_154, n_215, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_216, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_2110);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_96;
input n_156;
input n_209;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_200;
input n_51;
input n_166;
input n_76;
input n_218;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_217;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_214;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_211;
input n_194;
input n_97;
input n_154;
input n_215;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_216;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_2110;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_2084;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_1985;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_238;
wire n_365;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_2098;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_2043;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2072;
wire n_306;
wire n_436;
wire n_324;
wire n_2087;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_2100;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2041;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_2099;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_2059;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_2075;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_2057;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_342;
wire n_2035;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_2032;
wire n_2090;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1429;
wire n_1324;
wire n_2064;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_2022;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1288;
wire n_1201;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_2070;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_689;
wire n_400;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_1978;
wire n_571;
wire n_414;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_1986;
wire n_540;
wire n_692;
wire n_2054;
wire n_1857;
wire n_984;
wire n_1687;
wire n_2073;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_2093;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_2014;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_2065;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_2096;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_2012;
wire n_1937;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_2103;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_2062;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_2101;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_2088;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2108;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_2085;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_954;
wire n_596;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_252;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1967;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_2081;
wire n_265;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_718;
wire n_329;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_484;
wire n_411;
wire n_849;
wire n_2095;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_198),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_58),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_201),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_43),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_103),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_189),
.Y(n_224)
);

BUFx5_ASAP7_75t_L g225 ( 
.A(n_116),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_94),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_6),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_187),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_31),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_10),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_7),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_119),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_54),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_216),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_8),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_1),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_72),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_109),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_97),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_126),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_73),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_218),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_70),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_73),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_35),
.Y(n_245)
);

BUFx2_ASAP7_75t_L g246 ( 
.A(n_102),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_174),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_161),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_158),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_48),
.Y(n_250)
);

BUFx10_ASAP7_75t_L g251 ( 
.A(n_47),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_111),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_210),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_98),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_136),
.Y(n_255)
);

BUFx2_ASAP7_75t_L g256 ( 
.A(n_72),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_213),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_184),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_168),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_129),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_8),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_208),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_74),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_107),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_55),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_177),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_90),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_133),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_71),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_214),
.Y(n_270)
);

INVx1_ASAP7_75t_SL g271 ( 
.A(n_197),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_188),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_128),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_143),
.Y(n_274)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_91),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_104),
.Y(n_276)
);

CKINVDCx14_ASAP7_75t_R g277 ( 
.A(n_67),
.Y(n_277)
);

INVx2_ASAP7_75t_SL g278 ( 
.A(n_93),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_130),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_18),
.Y(n_280)
);

BUFx5_ASAP7_75t_L g281 ( 
.A(n_170),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_150),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_167),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_186),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g285 ( 
.A(n_30),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_217),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_125),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_171),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_20),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_16),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_86),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_176),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_191),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_28),
.Y(n_294)
);

INVx2_ASAP7_75t_SL g295 ( 
.A(n_215),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_211),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_9),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_30),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_70),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_75),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_137),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_2),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_2),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_34),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_47),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_132),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_0),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_100),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_175),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_204),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_96),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_141),
.Y(n_312)
);

BUFx3_ASAP7_75t_L g313 ( 
.A(n_71),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_75),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_38),
.Y(n_315)
);

BUFx2_ASAP7_75t_SL g316 ( 
.A(n_76),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_25),
.Y(n_317)
);

BUFx10_ASAP7_75t_L g318 ( 
.A(n_62),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_85),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_81),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_36),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_163),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_1),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_156),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_46),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_16),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_95),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_87),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_206),
.Y(n_329)
);

BUFx5_ASAP7_75t_L g330 ( 
.A(n_27),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_140),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_0),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_142),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_38),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_45),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_118),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_44),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_33),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_67),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_5),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_21),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_18),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_32),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_127),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_82),
.Y(n_345)
);

INVx1_ASAP7_75t_SL g346 ( 
.A(n_112),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_196),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_11),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_181),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_115),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_145),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_124),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_122),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_66),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_48),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_83),
.Y(n_356)
);

BUFx3_ASAP7_75t_L g357 ( 
.A(n_23),
.Y(n_357)
);

HB1xp67_ASAP7_75t_L g358 ( 
.A(n_54),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_66),
.Y(n_359)
);

BUFx10_ASAP7_75t_L g360 ( 
.A(n_44),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_22),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_178),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_110),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_105),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_92),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_80),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_113),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_165),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_11),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_63),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_51),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_13),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_52),
.Y(n_373)
);

BUFx2_ASAP7_75t_SL g374 ( 
.A(n_154),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_6),
.Y(n_375)
);

BUFx2_ASAP7_75t_L g376 ( 
.A(n_41),
.Y(n_376)
);

CKINVDCx16_ASAP7_75t_R g377 ( 
.A(n_37),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_56),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_65),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_27),
.Y(n_380)
);

INVx2_ASAP7_75t_SL g381 ( 
.A(n_50),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_146),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_37),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_159),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_147),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_121),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_68),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_15),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_40),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_24),
.Y(n_390)
);

BUFx2_ASAP7_75t_L g391 ( 
.A(n_185),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_42),
.Y(n_392)
);

INVx1_ASAP7_75t_SL g393 ( 
.A(n_144),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_202),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_78),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_209),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_43),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_56),
.Y(n_398)
);

INVx2_ASAP7_75t_SL g399 ( 
.A(n_160),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_12),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_152),
.Y(n_401)
);

BUFx2_ASAP7_75t_L g402 ( 
.A(n_23),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_212),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_99),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_24),
.Y(n_405)
);

INVx1_ASAP7_75t_SL g406 ( 
.A(n_183),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_106),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_123),
.Y(n_408)
);

INVx2_ASAP7_75t_SL g409 ( 
.A(n_5),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_200),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_17),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_108),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g413 ( 
.A(n_149),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_63),
.Y(n_414)
);

BUFx2_ASAP7_75t_L g415 ( 
.A(n_9),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_120),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_68),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_157),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_69),
.Y(n_419)
);

INVx2_ASAP7_75t_SL g420 ( 
.A(n_20),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_52),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_169),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_4),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_114),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_34),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_7),
.Y(n_426)
);

BUFx3_ASAP7_75t_L g427 ( 
.A(n_194),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_117),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_207),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_36),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g431 ( 
.A(n_58),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_148),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_297),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_377),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_330),
.Y(n_435)
);

CKINVDCx16_ASAP7_75t_R g436 ( 
.A(n_277),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_330),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_330),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_330),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_223),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_330),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_330),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_242),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_330),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_330),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_230),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_287),
.Y(n_447)
);

CKINVDCx16_ASAP7_75t_R g448 ( 
.A(n_270),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_230),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_256),
.B(n_3),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_319),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_230),
.Y(n_452)
);

HB1xp67_ASAP7_75t_L g453 ( 
.A(n_358),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_230),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_320),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_230),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_250),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_327),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_250),
.Y(n_459)
);

HB1xp67_ASAP7_75t_L g460 ( 
.A(n_375),
.Y(n_460)
);

INVxp67_ASAP7_75t_SL g461 ( 
.A(n_313),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_250),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_347),
.Y(n_463)
);

BUFx6f_ASAP7_75t_SL g464 ( 
.A(n_275),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_250),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_250),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_418),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_361),
.Y(n_468)
);

NOR2xp67_ASAP7_75t_L g469 ( 
.A(n_381),
.B(n_3),
.Y(n_469)
);

INVxp67_ASAP7_75t_L g470 ( 
.A(n_376),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_289),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_361),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_417),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_294),
.Y(n_474)
);

BUFx2_ASAP7_75t_SL g475 ( 
.A(n_278),
.Y(n_475)
);

HB1xp67_ASAP7_75t_L g476 ( 
.A(n_431),
.Y(n_476)
);

BUFx2_ASAP7_75t_L g477 ( 
.A(n_402),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_299),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_231),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_417),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_300),
.Y(n_481)
);

INVxp67_ASAP7_75t_SL g482 ( 
.A(n_313),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_357),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_357),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_220),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_229),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_236),
.Y(n_487)
);

CKINVDCx16_ASAP7_75t_R g488 ( 
.A(n_251),
.Y(n_488)
);

INVxp67_ASAP7_75t_L g489 ( 
.A(n_415),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_238),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_275),
.Y(n_491)
);

INVxp33_ASAP7_75t_L g492 ( 
.A(n_244),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_238),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_255),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_255),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_279),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_279),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_283),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_283),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_246),
.B(n_4),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_328),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_328),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_302),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_298),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_303),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_391),
.B(n_10),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_304),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_317),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_345),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_323),
.Y(n_510)
);

HB1xp67_ASAP7_75t_L g511 ( 
.A(n_222),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_325),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_413),
.B(n_12),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_326),
.Y(n_514)
);

BUFx6f_ASAP7_75t_SL g515 ( 
.A(n_427),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_345),
.Y(n_516)
);

BUFx3_ASAP7_75t_L g517 ( 
.A(n_427),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_334),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_410),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_337),
.Y(n_520)
);

INVxp33_ASAP7_75t_L g521 ( 
.A(n_265),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_355),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_381),
.B(n_13),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_410),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_338),
.Y(n_525)
);

CKINVDCx16_ASAP7_75t_R g526 ( 
.A(n_251),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_390),
.Y(n_527)
);

CKINVDCx16_ASAP7_75t_R g528 ( 
.A(n_251),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_340),
.Y(n_529)
);

HB1xp67_ASAP7_75t_L g530 ( 
.A(n_222),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_428),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_409),
.B(n_14),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_428),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_341),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_269),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_280),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_290),
.Y(n_537)
);

OR2x2_ASAP7_75t_L g538 ( 
.A(n_409),
.B(n_14),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_305),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_307),
.Y(n_540)
);

BUFx2_ASAP7_75t_L g541 ( 
.A(n_227),
.Y(n_541)
);

NOR2xp67_ASAP7_75t_L g542 ( 
.A(n_420),
.B(n_15),
.Y(n_542)
);

INVxp67_ASAP7_75t_SL g543 ( 
.A(n_314),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_315),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_321),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_342),
.Y(n_546)
);

BUFx2_ASAP7_75t_L g547 ( 
.A(n_227),
.Y(n_547)
);

BUFx3_ASAP7_75t_L g548 ( 
.A(n_491),
.Y(n_548)
);

HB1xp67_ASAP7_75t_L g549 ( 
.A(n_541),
.Y(n_549)
);

AND2x4_ASAP7_75t_L g550 ( 
.A(n_517),
.B(n_420),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_435),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_492),
.B(n_332),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_435),
.Y(n_553)
);

HB1xp67_ASAP7_75t_L g554 ( 
.A(n_541),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_437),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_437),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_438),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_438),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_440),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_521),
.B(n_335),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_439),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g562 ( 
.A(n_439),
.Y(n_562)
);

BUFx3_ASAP7_75t_L g563 ( 
.A(n_491),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_461),
.B(n_482),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_441),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_441),
.B(n_224),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_442),
.Y(n_567)
);

INVx3_ASAP7_75t_L g568 ( 
.A(n_442),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_444),
.B(n_445),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_444),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_443),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_445),
.B(n_228),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_446),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_490),
.B(n_232),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_446),
.Y(n_575)
);

INVx2_ASAP7_75t_SL g576 ( 
.A(n_517),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_447),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_449),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_449),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_452),
.Y(n_580)
);

BUFx2_ASAP7_75t_L g581 ( 
.A(n_433),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_452),
.Y(n_582)
);

BUFx2_ASAP7_75t_L g583 ( 
.A(n_434),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_490),
.B(n_247),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_454),
.Y(n_585)
);

HB1xp67_ASAP7_75t_L g586 ( 
.A(n_547),
.Y(n_586)
);

NAND2xp33_ASAP7_75t_SL g587 ( 
.A(n_450),
.B(n_233),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_454),
.Y(n_588)
);

NOR2x1_ASAP7_75t_L g589 ( 
.A(n_475),
.B(n_374),
.Y(n_589)
);

AND2x2_ASAP7_75t_L g590 ( 
.A(n_483),
.B(n_339),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_456),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_456),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_457),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_457),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_459),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_459),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_462),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_462),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_465),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_493),
.B(n_248),
.Y(n_600)
);

BUFx2_ASAP7_75t_L g601 ( 
.A(n_547),
.Y(n_601)
);

OAI22xp5_ASAP7_75t_SL g602 ( 
.A1(n_479),
.A2(n_425),
.B1(n_430),
.B2(n_237),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_465),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_466),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_466),
.Y(n_605)
);

INVx3_ASAP7_75t_L g606 ( 
.A(n_493),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_451),
.Y(n_607)
);

OAI21x1_ASAP7_75t_L g608 ( 
.A1(n_494),
.A2(n_257),
.B(n_254),
.Y(n_608)
);

INVxp67_ASAP7_75t_L g609 ( 
.A(n_511),
.Y(n_609)
);

BUFx6f_ASAP7_75t_L g610 ( 
.A(n_494),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_475),
.B(n_278),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_495),
.Y(n_612)
);

INVx3_ASAP7_75t_L g613 ( 
.A(n_495),
.Y(n_613)
);

INVx3_ASAP7_75t_L g614 ( 
.A(n_496),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_496),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_497),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_497),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_498),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_498),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_499),
.Y(n_620)
);

AND2x2_ASAP7_75t_SL g621 ( 
.A(n_538),
.B(n_234),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_499),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_501),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_484),
.B(n_359),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_501),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_502),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_455),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_502),
.Y(n_628)
);

BUFx2_ASAP7_75t_L g629 ( 
.A(n_471),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_509),
.Y(n_630)
);

INVx3_ASAP7_75t_L g631 ( 
.A(n_509),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_516),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_516),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_519),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_SL g635 ( 
.A(n_436),
.B(n_318),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_519),
.Y(n_636)
);

HB1xp67_ASAP7_75t_L g637 ( 
.A(n_470),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_555),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_621),
.B(n_448),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_637),
.B(n_488),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_548),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_576),
.B(n_611),
.Y(n_642)
);

NOR2x1p5_ASAP7_75t_L g643 ( 
.A(n_571),
.B(n_474),
.Y(n_643)
);

AND2x6_ASAP7_75t_L g644 ( 
.A(n_589),
.B(n_450),
.Y(n_644)
);

INVx3_ASAP7_75t_L g645 ( 
.A(n_568),
.Y(n_645)
);

INVx2_ASAP7_75t_SL g646 ( 
.A(n_621),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_571),
.Y(n_647)
);

INVx2_ASAP7_75t_SL g648 ( 
.A(n_621),
.Y(n_648)
);

OAI22xp5_ASAP7_75t_L g649 ( 
.A1(n_621),
.A2(n_513),
.B1(n_538),
.B2(n_500),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_637),
.B(n_526),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_548),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_548),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_548),
.Y(n_653)
);

INVx3_ASAP7_75t_L g654 ( 
.A(n_568),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_576),
.B(n_464),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_563),
.Y(n_656)
);

INVx2_ASAP7_75t_SL g657 ( 
.A(n_576),
.Y(n_657)
);

AO22x2_ASAP7_75t_L g658 ( 
.A1(n_552),
.A2(n_489),
.B1(n_543),
.B2(n_531),
.Y(n_658)
);

INVx1_ASAP7_75t_SL g659 ( 
.A(n_581),
.Y(n_659)
);

BUFx2_ASAP7_75t_L g660 ( 
.A(n_581),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_563),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_610),
.Y(n_662)
);

AND2x6_ASAP7_75t_L g663 ( 
.A(n_589),
.B(n_234),
.Y(n_663)
);

INVx6_ASAP7_75t_L g664 ( 
.A(n_550),
.Y(n_664)
);

INVx1_ASAP7_75t_SL g665 ( 
.A(n_581),
.Y(n_665)
);

INVx1_ASAP7_75t_SL g666 ( 
.A(n_583),
.Y(n_666)
);

AOI22xp33_ASAP7_75t_L g667 ( 
.A1(n_587),
.A2(n_532),
.B1(n_523),
.B2(n_506),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_611),
.B(n_478),
.Y(n_668)
);

INVx5_ASAP7_75t_L g669 ( 
.A(n_557),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_569),
.B(n_481),
.Y(n_670)
);

BUFx3_ASAP7_75t_L g671 ( 
.A(n_563),
.Y(n_671)
);

AOI22xp33_ASAP7_75t_L g672 ( 
.A1(n_587),
.A2(n_542),
.B1(n_469),
.B2(n_531),
.Y(n_672)
);

INVx2_ASAP7_75t_SL g673 ( 
.A(n_629),
.Y(n_673)
);

INVxp67_ASAP7_75t_L g674 ( 
.A(n_583),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_555),
.Y(n_675)
);

BUFx2_ASAP7_75t_L g676 ( 
.A(n_583),
.Y(n_676)
);

AOI22xp5_ASAP7_75t_L g677 ( 
.A1(n_564),
.A2(n_505),
.B1(n_508),
.B2(n_503),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_555),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_565),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_563),
.Y(n_680)
);

BUFx10_ASAP7_75t_L g681 ( 
.A(n_559),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_601),
.B(n_549),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_569),
.Y(n_683)
);

INVx2_ASAP7_75t_SL g684 ( 
.A(n_564),
.Y(n_684)
);

BUFx10_ASAP7_75t_L g685 ( 
.A(n_607),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_565),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_565),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_612),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_612),
.Y(n_689)
);

NAND2xp33_ASAP7_75t_R g690 ( 
.A(n_629),
.B(n_463),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_564),
.B(n_510),
.Y(n_691)
);

OAI22xp5_ASAP7_75t_L g692 ( 
.A1(n_609),
.A2(n_235),
.B1(n_237),
.B2(n_233),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_570),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_570),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_551),
.B(n_512),
.Y(n_695)
);

OR2x2_ASAP7_75t_L g696 ( 
.A(n_601),
.B(n_528),
.Y(n_696)
);

OAI21xp5_ASAP7_75t_L g697 ( 
.A1(n_608),
.A2(n_259),
.B(n_258),
.Y(n_697)
);

BUFx6f_ASAP7_75t_L g698 ( 
.A(n_610),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_551),
.B(n_514),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_568),
.B(n_518),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_553),
.B(n_520),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_615),
.Y(n_702)
);

AND2x6_ASAP7_75t_L g703 ( 
.A(n_570),
.B(n_234),
.Y(n_703)
);

CKINVDCx16_ASAP7_75t_R g704 ( 
.A(n_635),
.Y(n_704)
);

BUFx10_ASAP7_75t_L g705 ( 
.A(n_627),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_553),
.B(n_464),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_556),
.B(n_464),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_597),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_597),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_615),
.Y(n_710)
);

NAND2xp33_ASAP7_75t_L g711 ( 
.A(n_557),
.B(n_225),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_601),
.B(n_530),
.Y(n_712)
);

BUFx8_ASAP7_75t_SL g713 ( 
.A(n_577),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_617),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_568),
.B(n_525),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_617),
.Y(n_716)
);

OR2x6_ASAP7_75t_L g717 ( 
.A(n_602),
.B(n_477),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_618),
.Y(n_718)
);

BUFx10_ASAP7_75t_L g719 ( 
.A(n_577),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_618),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_619),
.Y(n_721)
);

INVxp67_ASAP7_75t_L g722 ( 
.A(n_629),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_619),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_620),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_597),
.Y(n_725)
);

INVx4_ASAP7_75t_L g726 ( 
.A(n_557),
.Y(n_726)
);

INVx5_ASAP7_75t_L g727 ( 
.A(n_557),
.Y(n_727)
);

AND2x2_ASAP7_75t_L g728 ( 
.A(n_549),
.B(n_529),
.Y(n_728)
);

INVx3_ASAP7_75t_L g729 ( 
.A(n_568),
.Y(n_729)
);

BUFx6f_ASAP7_75t_SL g730 ( 
.A(n_550),
.Y(n_730)
);

OR2x2_ASAP7_75t_L g731 ( 
.A(n_554),
.B(n_477),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_620),
.Y(n_732)
);

INVx4_ASAP7_75t_L g733 ( 
.A(n_557),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_556),
.B(n_534),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_622),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_622),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_558),
.B(n_546),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_597),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_623),
.Y(n_739)
);

BUFx6f_ASAP7_75t_L g740 ( 
.A(n_610),
.Y(n_740)
);

AOI22xp5_ASAP7_75t_L g741 ( 
.A1(n_609),
.A2(n_285),
.B1(n_245),
.B2(n_343),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_558),
.B(n_561),
.Y(n_742)
);

INVx6_ASAP7_75t_L g743 ( 
.A(n_550),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_623),
.Y(n_744)
);

NAND2xp33_ASAP7_75t_L g745 ( 
.A(n_557),
.B(n_225),
.Y(n_745)
);

AND2x6_ASAP7_75t_L g746 ( 
.A(n_561),
.B(n_234),
.Y(n_746)
);

INVxp33_ASAP7_75t_L g747 ( 
.A(n_554),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_597),
.Y(n_748)
);

BUFx8_ASAP7_75t_SL g749 ( 
.A(n_552),
.Y(n_749)
);

AND2x4_ASAP7_75t_L g750 ( 
.A(n_550),
.B(n_545),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_603),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_603),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_603),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_567),
.B(n_524),
.Y(n_754)
);

INVx4_ASAP7_75t_L g755 ( 
.A(n_557),
.Y(n_755)
);

AOI22xp5_ASAP7_75t_L g756 ( 
.A1(n_635),
.A2(n_354),
.B1(n_348),
.B2(n_241),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_625),
.Y(n_757)
);

AND2x6_ASAP7_75t_L g758 ( 
.A(n_567),
.B(n_234),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_603),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_625),
.Y(n_760)
);

BUFx6f_ASAP7_75t_L g761 ( 
.A(n_610),
.Y(n_761)
);

INVx3_ASAP7_75t_L g762 ( 
.A(n_557),
.Y(n_762)
);

INVx2_ASAP7_75t_SL g763 ( 
.A(n_586),
.Y(n_763)
);

AND2x4_ASAP7_75t_L g764 ( 
.A(n_550),
.B(n_590),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_626),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_606),
.B(n_524),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_566),
.B(n_515),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_566),
.B(n_572),
.Y(n_768)
);

INVx4_ASAP7_75t_L g769 ( 
.A(n_562),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_603),
.Y(n_770)
);

BUFx6f_ASAP7_75t_L g771 ( 
.A(n_610),
.Y(n_771)
);

BUFx6f_ASAP7_75t_L g772 ( 
.A(n_610),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_626),
.Y(n_773)
);

NOR3xp33_ASAP7_75t_L g774 ( 
.A(n_602),
.B(n_241),
.C(n_235),
.Y(n_774)
);

INVx2_ASAP7_75t_SL g775 ( 
.A(n_552),
.Y(n_775)
);

AND3x2_ASAP7_75t_L g776 ( 
.A(n_586),
.B(n_460),
.C(n_453),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_562),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_630),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_562),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_562),
.Y(n_780)
);

BUFx10_ASAP7_75t_L g781 ( 
.A(n_630),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_606),
.B(n_533),
.Y(n_782)
);

BUFx2_ASAP7_75t_L g783 ( 
.A(n_560),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_634),
.Y(n_784)
);

INVx2_ASAP7_75t_SL g785 ( 
.A(n_560),
.Y(n_785)
);

BUFx10_ASAP7_75t_L g786 ( 
.A(n_634),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_572),
.B(n_262),
.Y(n_787)
);

INVx3_ASAP7_75t_L g788 ( 
.A(n_562),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_560),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_636),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_636),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_562),
.Y(n_792)
);

OR2x2_ASAP7_75t_L g793 ( 
.A(n_590),
.B(n_467),
.Y(n_793)
);

BUFx2_ASAP7_75t_L g794 ( 
.A(n_590),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_688),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_646),
.B(n_562),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_646),
.B(n_562),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_689),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_642),
.B(n_606),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_677),
.B(n_219),
.Y(n_800)
);

BUFx6f_ASAP7_75t_L g801 ( 
.A(n_671),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_668),
.B(n_219),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_659),
.B(n_476),
.Y(n_803)
);

NAND3xp33_ASAP7_75t_L g804 ( 
.A(n_667),
.B(n_261),
.C(n_243),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_642),
.B(n_606),
.Y(n_805)
);

OR2x2_ASAP7_75t_L g806 ( 
.A(n_665),
.B(n_624),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_673),
.B(n_221),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_683),
.B(n_606),
.Y(n_808)
);

AND2x6_ASAP7_75t_SL g809 ( 
.A(n_717),
.B(n_369),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_638),
.Y(n_810)
);

NAND2xp33_ASAP7_75t_L g811 ( 
.A(n_695),
.B(n_221),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_691),
.B(n_613),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_638),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_684),
.B(n_767),
.Y(n_814)
);

OAI22xp33_ASAP7_75t_L g815 ( 
.A1(n_649),
.A2(n_614),
.B1(n_631),
.B2(n_613),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_675),
.Y(n_816)
);

AND2x6_ASAP7_75t_SL g817 ( 
.A(n_717),
.B(n_370),
.Y(n_817)
);

NOR3xp33_ASAP7_75t_L g818 ( 
.A(n_722),
.B(n_378),
.C(n_372),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_684),
.B(n_613),
.Y(n_819)
);

AOI22xp5_ASAP7_75t_L g820 ( 
.A1(n_648),
.A2(n_614),
.B1(n_631),
.B2(n_613),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_670),
.B(n_639),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_702),
.Y(n_822)
);

INVx2_ASAP7_75t_SL g823 ( 
.A(n_666),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_767),
.B(n_613),
.Y(n_824)
);

OAI22xp5_ASAP7_75t_L g825 ( 
.A1(n_667),
.A2(n_261),
.B1(n_263),
.B2(n_243),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_670),
.B(n_639),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_781),
.B(n_226),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_648),
.B(n_614),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_675),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_699),
.B(n_614),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_781),
.B(n_226),
.Y(n_831)
);

BUFx6f_ASAP7_75t_L g832 ( 
.A(n_662),
.Y(n_832)
);

BUFx6f_ASAP7_75t_SL g833 ( 
.A(n_681),
.Y(n_833)
);

BUFx5_ASAP7_75t_L g834 ( 
.A(n_703),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_728),
.B(n_458),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_781),
.B(n_239),
.Y(n_836)
);

NOR3xp33_ASAP7_75t_L g837 ( 
.A(n_674),
.B(n_395),
.C(n_389),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_768),
.B(n_614),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_786),
.B(n_239),
.Y(n_839)
);

AOI221xp5_ASAP7_75t_L g840 ( 
.A1(n_692),
.A2(n_426),
.B1(n_423),
.B2(n_430),
.C(n_371),
.Y(n_840)
);

AOI22xp33_ASAP7_75t_L g841 ( 
.A1(n_658),
.A2(n_631),
.B1(n_632),
.B2(n_616),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_786),
.B(n_240),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_701),
.B(n_631),
.Y(n_843)
);

AND2x6_ASAP7_75t_SL g844 ( 
.A(n_717),
.B(n_535),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_786),
.B(n_240),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_710),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_768),
.B(n_631),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_775),
.B(n_616),
.Y(n_848)
);

INVx2_ASAP7_75t_SL g849 ( 
.A(n_660),
.Y(n_849)
);

OAI22xp5_ASAP7_75t_L g850 ( 
.A1(n_789),
.A2(n_371),
.B1(n_373),
.B2(n_263),
.Y(n_850)
);

OAI21xp5_ASAP7_75t_L g851 ( 
.A1(n_697),
.A2(n_608),
.B(n_584),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_775),
.B(n_249),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_SL g853 ( 
.A(n_645),
.B(n_610),
.Y(n_853)
);

AND2x2_ASAP7_75t_L g854 ( 
.A(n_682),
.B(n_624),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_785),
.B(n_616),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_734),
.B(n_624),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_712),
.B(n_504),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_785),
.B(n_632),
.Y(n_858)
);

AND2x6_ASAP7_75t_L g859 ( 
.A(n_764),
.B(n_632),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_644),
.B(n_633),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_644),
.B(n_750),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_644),
.B(n_633),
.Y(n_862)
);

AOI22xp33_ASAP7_75t_L g863 ( 
.A1(n_658),
.A2(n_633),
.B1(n_610),
.B2(n_628),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_714),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_644),
.B(n_574),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_644),
.B(n_574),
.Y(n_866)
);

AND2x6_ASAP7_75t_L g867 ( 
.A(n_764),
.B(n_268),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_750),
.B(n_584),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_750),
.B(n_600),
.Y(n_869)
);

BUFx12f_ASAP7_75t_L g870 ( 
.A(n_681),
.Y(n_870)
);

INVx3_ASAP7_75t_L g871 ( 
.A(n_645),
.Y(n_871)
);

NAND2x1_ASAP7_75t_L g872 ( 
.A(n_645),
.B(n_573),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_657),
.B(n_764),
.Y(n_873)
);

NOR2xp67_ASAP7_75t_L g874 ( 
.A(n_647),
.B(n_600),
.Y(n_874)
);

OAI22x1_ASAP7_75t_SL g875 ( 
.A1(n_647),
.A2(n_522),
.B1(n_527),
.B2(n_507),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_678),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_657),
.B(n_628),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_734),
.B(n_515),
.Y(n_878)
);

NAND2x1p5_ASAP7_75t_L g879 ( 
.A(n_700),
.B(n_715),
.Y(n_879)
);

O2A1O1Ixp33_ASAP7_75t_L g880 ( 
.A1(n_742),
.A2(n_536),
.B(n_537),
.C(n_535),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_716),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_706),
.B(n_628),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_678),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_706),
.B(n_628),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_789),
.B(n_249),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_L g886 ( 
.A(n_737),
.B(n_515),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_679),
.Y(n_887)
);

OAI22xp5_ASAP7_75t_L g888 ( 
.A1(n_664),
.A2(n_387),
.B1(n_373),
.B2(n_379),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_707),
.B(n_628),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_718),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_756),
.B(n_252),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_679),
.Y(n_892)
);

BUFx6f_ASAP7_75t_L g893 ( 
.A(n_662),
.Y(n_893)
);

NOR2xp67_ASAP7_75t_L g894 ( 
.A(n_696),
.B(n_533),
.Y(n_894)
);

NOR2xp67_ASAP7_75t_L g895 ( 
.A(n_763),
.B(n_485),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_720),
.Y(n_896)
);

INVxp67_ASAP7_75t_L g897 ( 
.A(n_676),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_783),
.B(n_252),
.Y(n_898)
);

AOI22xp33_ASAP7_75t_L g899 ( 
.A1(n_658),
.A2(n_628),
.B1(n_593),
.B2(n_605),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_707),
.B(n_628),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_654),
.B(n_628),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_721),
.B(n_573),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_777),
.A2(n_608),
.B(n_579),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_723),
.B(n_578),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_640),
.B(n_486),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_724),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_L g907 ( 
.A(n_737),
.B(n_379),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_732),
.B(n_578),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_735),
.Y(n_909)
);

AOI22xp5_ASAP7_75t_L g910 ( 
.A1(n_664),
.A2(n_295),
.B1(n_399),
.B2(n_429),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_654),
.B(n_260),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_736),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_SL g913 ( 
.A(n_704),
.B(n_318),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_739),
.B(n_579),
.Y(n_914)
);

INVx2_ASAP7_75t_SL g915 ( 
.A(n_650),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_744),
.B(n_580),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_SL g917 ( 
.A(n_654),
.B(n_260),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_686),
.Y(n_918)
);

OAI22xp5_ASAP7_75t_SL g919 ( 
.A1(n_741),
.A2(n_414),
.B1(n_411),
.B2(n_405),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_747),
.B(n_794),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_L g921 ( 
.A(n_700),
.B(n_380),
.Y(n_921)
);

BUFx6f_ASAP7_75t_L g922 ( 
.A(n_662),
.Y(n_922)
);

BUFx6f_ASAP7_75t_L g923 ( 
.A(n_662),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_SL g924 ( 
.A(n_672),
.B(n_366),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_715),
.B(n_380),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_757),
.B(n_580),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_760),
.B(n_582),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_747),
.B(n_719),
.Y(n_928)
);

O2A1O1Ixp33_ASAP7_75t_L g929 ( 
.A1(n_765),
.A2(n_545),
.B(n_536),
.C(n_537),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_773),
.B(n_582),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_778),
.Y(n_931)
);

AND2x6_ASAP7_75t_L g932 ( 
.A(n_729),
.B(n_268),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_664),
.B(n_383),
.Y(n_933)
);

CKINVDCx20_ASAP7_75t_R g934 ( 
.A(n_713),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_719),
.B(n_487),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_672),
.B(n_366),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_784),
.B(n_585),
.Y(n_937)
);

OAI22xp33_ASAP7_75t_SL g938 ( 
.A1(n_743),
.A2(n_414),
.B1(n_419),
.B2(n_421),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_681),
.B(n_367),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_687),
.Y(n_940)
);

AND2x2_ASAP7_75t_L g941 ( 
.A(n_719),
.B(n_793),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_790),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_SL g943 ( 
.A(n_729),
.B(n_367),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_791),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_L g945 ( 
.A(n_743),
.B(n_383),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_SL g946 ( 
.A(n_729),
.B(n_368),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_655),
.B(n_585),
.Y(n_947)
);

AOI22xp5_ASAP7_75t_L g948 ( 
.A1(n_743),
.A2(n_295),
.B1(n_399),
.B2(n_429),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_754),
.Y(n_949)
);

INVxp67_ASAP7_75t_L g950 ( 
.A(n_690),
.Y(n_950)
);

AOI22xp33_ASAP7_75t_L g951 ( 
.A1(n_774),
.A2(n_605),
.B1(n_604),
.B2(n_591),
.Y(n_951)
);

INVx4_ASAP7_75t_L g952 ( 
.A(n_730),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_698),
.B(n_368),
.Y(n_953)
);

A2O1A1Ixp33_ASAP7_75t_L g954 ( 
.A1(n_708),
.A2(n_604),
.B(n_598),
.C(n_595),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_698),
.B(n_382),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_687),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_655),
.B(n_591),
.Y(n_957)
);

CKINVDCx20_ASAP7_75t_R g958 ( 
.A(n_713),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_787),
.B(n_592),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_698),
.B(n_382),
.Y(n_960)
);

OAI22xp5_ASAP7_75t_SL g961 ( 
.A1(n_731),
.A2(n_426),
.B1(n_405),
.B2(n_398),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_698),
.B(n_384),
.Y(n_962)
);

AOI22xp5_ASAP7_75t_L g963 ( 
.A1(n_730),
.A2(n_408),
.B1(n_386),
.B2(n_396),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_787),
.B(n_592),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_693),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_799),
.A2(n_779),
.B(n_777),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_805),
.A2(n_780),
.B(n_779),
.Y(n_967)
);

NOR2xp33_ASAP7_75t_L g968 ( 
.A(n_950),
.B(n_749),
.Y(n_968)
);

INVx3_ASAP7_75t_L g969 ( 
.A(n_801),
.Y(n_969)
);

O2A1O1Ixp33_ASAP7_75t_L g970 ( 
.A1(n_825),
.A2(n_782),
.B(n_766),
.C(n_709),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_868),
.B(n_663),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_L g972 ( 
.A(n_821),
.B(n_749),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_869),
.B(n_663),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_824),
.A2(n_792),
.B(n_780),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_838),
.A2(n_792),
.B(n_733),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_795),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_821),
.B(n_826),
.Y(n_977)
);

O2A1O1Ixp33_ASAP7_75t_L g978 ( 
.A1(n_907),
.A2(n_709),
.B(n_725),
.C(n_708),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_847),
.A2(n_733),
.B(n_726),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_810),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_813),
.Y(n_981)
);

BUFx3_ASAP7_75t_L g982 ( 
.A(n_870),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_947),
.A2(n_733),
.B(n_726),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_812),
.B(n_663),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_798),
.Y(n_985)
);

BUFx2_ASAP7_75t_L g986 ( 
.A(n_823),
.Y(n_986)
);

INVxp67_ASAP7_75t_L g987 ( 
.A(n_849),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_812),
.B(n_663),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_826),
.B(n_685),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_957),
.A2(n_755),
.B(n_726),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_L g991 ( 
.A(n_814),
.B(n_685),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_856),
.B(n_663),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_856),
.B(n_693),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_803),
.B(n_685),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_949),
.B(n_830),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_830),
.B(n_694),
.Y(n_996)
);

INVx3_ASAP7_75t_L g997 ( 
.A(n_801),
.Y(n_997)
);

AOI22xp5_ASAP7_75t_L g998 ( 
.A1(n_921),
.A2(n_690),
.B1(n_705),
.B2(n_643),
.Y(n_998)
);

OAI21xp5_ASAP7_75t_L g999 ( 
.A1(n_851),
.A2(n_694),
.B(n_725),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_843),
.B(n_738),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_843),
.B(n_738),
.Y(n_1001)
);

A2O1A1Ixp33_ASAP7_75t_L g1002 ( 
.A1(n_921),
.A2(n_751),
.B(n_770),
.C(n_748),
.Y(n_1002)
);

O2A1O1Ixp33_ASAP7_75t_L g1003 ( 
.A1(n_907),
.A2(n_751),
.B(n_770),
.C(n_748),
.Y(n_1003)
);

AND2x2_ASAP7_75t_L g1004 ( 
.A(n_920),
.B(n_705),
.Y(n_1004)
);

HB1xp67_ASAP7_75t_L g1005 ( 
.A(n_897),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_L g1006 ( 
.A(n_915),
.B(n_705),
.Y(n_1006)
);

OAI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_903),
.A2(n_753),
.B(n_752),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_877),
.A2(n_769),
.B(n_755),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_816),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_874),
.B(n_752),
.Y(n_1010)
);

O2A1O1Ixp33_ASAP7_75t_L g1011 ( 
.A1(n_925),
.A2(n_753),
.B(n_759),
.C(n_641),
.Y(n_1011)
);

INVx3_ASAP7_75t_L g1012 ( 
.A(n_801),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_822),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_808),
.A2(n_769),
.B(n_755),
.Y(n_1014)
);

BUFx12f_ASAP7_75t_L g1015 ( 
.A(n_844),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_905),
.B(n_759),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_925),
.B(n_854),
.Y(n_1017)
);

BUFx6f_ASAP7_75t_L g1018 ( 
.A(n_801),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_882),
.A2(n_889),
.B(n_884),
.Y(n_1019)
);

OAI22xp5_ASAP7_75t_L g1020 ( 
.A1(n_873),
.A2(n_769),
.B1(n_788),
.B2(n_762),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_933),
.B(n_651),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_829),
.Y(n_1022)
);

OAI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_820),
.A2(n_788),
.B(n_762),
.Y(n_1023)
);

HB1xp67_ASAP7_75t_L g1024 ( 
.A(n_857),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_876),
.Y(n_1025)
);

OAI21x1_ASAP7_75t_L g1026 ( 
.A1(n_860),
.A2(n_788),
.B(n_762),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_933),
.B(n_945),
.Y(n_1027)
);

AOI21x1_ASAP7_75t_L g1028 ( 
.A1(n_796),
.A2(n_653),
.B(n_652),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_900),
.A2(n_661),
.B(n_656),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_853),
.A2(n_680),
.B(n_669),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_853),
.A2(n_727),
.B(n_669),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_878),
.B(n_740),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_833),
.Y(n_1033)
);

AND2x2_ASAP7_75t_L g1034 ( 
.A(n_806),
.B(n_776),
.Y(n_1034)
);

OAI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_828),
.A2(n_745),
.B(n_711),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_L g1036 ( 
.A(n_804),
.B(n_740),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_901),
.A2(n_727),
.B(n_669),
.Y(n_1037)
);

HB1xp67_ASAP7_75t_L g1038 ( 
.A(n_835),
.Y(n_1038)
);

INVx11_ASAP7_75t_L g1039 ( 
.A(n_867),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_SL g1040 ( 
.A(n_861),
.B(n_740),
.Y(n_1040)
);

OAI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_879),
.A2(n_771),
.B1(n_761),
.B2(n_772),
.Y(n_1041)
);

NOR3xp33_ASAP7_75t_L g1042 ( 
.A(n_941),
.B(n_388),
.C(n_387),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_878),
.B(n_761),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_901),
.A2(n_727),
.B(n_669),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_886),
.B(n_761),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_872),
.A2(n_727),
.B(n_711),
.Y(n_1046)
);

AND2x2_ASAP7_75t_L g1047 ( 
.A(n_928),
.B(n_539),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_935),
.B(n_539),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_886),
.B(n_761),
.Y(n_1049)
);

BUFx4f_ASAP7_75t_L g1050 ( 
.A(n_859),
.Y(n_1050)
);

BUFx6f_ASAP7_75t_L g1051 ( 
.A(n_832),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_SL g1052 ( 
.A(n_879),
.B(n_815),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_841),
.B(n_771),
.Y(n_1053)
);

BUFx2_ASAP7_75t_SL g1054 ( 
.A(n_833),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_846),
.Y(n_1055)
);

AOI22xp5_ASAP7_75t_L g1056 ( 
.A1(n_859),
.A2(n_745),
.B1(n_772),
.B2(n_771),
.Y(n_1056)
);

NOR2x2_ASAP7_75t_L g1057 ( 
.A(n_961),
.B(n_318),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_864),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_819),
.A2(n_772),
.B(n_771),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_796),
.A2(n_772),
.B(n_386),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_797),
.A2(n_396),
.B(n_384),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_815),
.B(n_401),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_841),
.B(n_388),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_797),
.A2(n_407),
.B(n_401),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_881),
.B(n_392),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_848),
.A2(n_408),
.B(n_407),
.Y(n_1066)
);

OAI22x1_ASAP7_75t_L g1067 ( 
.A1(n_924),
.A2(n_411),
.B1(n_400),
.B2(n_419),
.Y(n_1067)
);

INVxp67_ASAP7_75t_L g1068 ( 
.A(n_895),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_855),
.A2(n_424),
.B(n_416),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_858),
.A2(n_424),
.B(n_416),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_902),
.A2(n_274),
.B(n_273),
.Y(n_1071)
);

OAI22xp5_ASAP7_75t_L g1072 ( 
.A1(n_871),
.A2(n_392),
.B1(n_397),
.B2(n_398),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_904),
.A2(n_914),
.B(n_908),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_L g1074 ( 
.A(n_871),
.B(n_397),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_916),
.A2(n_286),
.B(n_276),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_890),
.B(n_400),
.Y(n_1076)
);

OAI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_954),
.A2(n_594),
.B(n_593),
.Y(n_1077)
);

HB1xp67_ASAP7_75t_L g1078 ( 
.A(n_894),
.Y(n_1078)
);

AND2x2_ASAP7_75t_L g1079 ( 
.A(n_913),
.B(n_540),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_896),
.B(n_421),
.Y(n_1080)
);

INVxp67_ASAP7_75t_L g1081 ( 
.A(n_875),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_926),
.A2(n_296),
.B(n_291),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_927),
.A2(n_306),
.B(n_301),
.Y(n_1083)
);

AOI21x1_ASAP7_75t_L g1084 ( 
.A1(n_862),
.A2(n_595),
.B(n_594),
.Y(n_1084)
);

AND2x4_ASAP7_75t_L g1085 ( 
.A(n_952),
.B(n_540),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_883),
.Y(n_1086)
);

CKINVDCx20_ASAP7_75t_R g1087 ( 
.A(n_934),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_930),
.A2(n_937),
.B(n_917),
.Y(n_1088)
);

NAND2x1p5_ASAP7_75t_L g1089 ( 
.A(n_952),
.B(n_598),
.Y(n_1089)
);

OAI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_865),
.A2(n_404),
.B(n_349),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_906),
.B(n_423),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_909),
.B(n_544),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_912),
.B(n_544),
.Y(n_1093)
);

AND2x2_ASAP7_75t_L g1094 ( 
.A(n_850),
.B(n_468),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_931),
.B(n_316),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_911),
.A2(n_352),
.B(n_308),
.Y(n_1096)
);

NOR2x1_ASAP7_75t_R g1097 ( 
.A(n_939),
.B(n_309),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_911),
.A2(n_356),
.B(n_311),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_942),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_917),
.A2(n_362),
.B(n_324),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_SL g1101 ( 
.A(n_832),
.B(n_575),
.Y(n_1101)
);

NOR2xp33_ASAP7_75t_L g1102 ( 
.A(n_885),
.B(n_360),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_SL g1103 ( 
.A(n_832),
.B(n_575),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_887),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_SL g1105 ( 
.A(n_832),
.B(n_575),
.Y(n_1105)
);

OR2x6_ASAP7_75t_SL g1106 ( 
.A(n_888),
.B(n_329),
.Y(n_1106)
);

INVx3_ASAP7_75t_L g1107 ( 
.A(n_859),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_943),
.A2(n_351),
.B(n_331),
.Y(n_1108)
);

A2O1A1Ixp33_ASAP7_75t_L g1109 ( 
.A1(n_944),
.A2(n_292),
.B(n_288),
.C(n_284),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_L g1110 ( 
.A(n_936),
.B(n_360),
.Y(n_1110)
);

NOR2xp33_ASAP7_75t_L g1111 ( 
.A(n_866),
.B(n_360),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_899),
.B(n_253),
.Y(n_1112)
);

NOR2xp67_ASAP7_75t_L g1113 ( 
.A(n_963),
.B(n_468),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_899),
.B(n_266),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_859),
.B(n_271),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_943),
.A2(n_364),
.B(n_336),
.Y(n_1116)
);

AND2x2_ASAP7_75t_L g1117 ( 
.A(n_818),
.B(n_472),
.Y(n_1117)
);

INVx1_ASAP7_75t_SL g1118 ( 
.A(n_958),
.Y(n_1118)
);

O2A1O1Ixp33_ASAP7_75t_L g1119 ( 
.A1(n_946),
.A2(n_264),
.B(n_267),
.C(n_272),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_859),
.B(n_346),
.Y(n_1120)
);

AOI22xp5_ASAP7_75t_L g1121 ( 
.A1(n_827),
.A2(n_365),
.B1(n_282),
.B2(n_293),
.Y(n_1121)
);

NOR2xp33_ASAP7_75t_L g1122 ( 
.A(n_898),
.B(n_393),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_946),
.A2(n_802),
.B(n_953),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_892),
.Y(n_1124)
);

NOR2xp33_ASAP7_75t_L g1125 ( 
.A(n_831),
.B(n_406),
.Y(n_1125)
);

O2A1O1Ixp5_ASAP7_75t_L g1126 ( 
.A1(n_953),
.A2(n_596),
.B(n_599),
.C(n_310),
.Y(n_1126)
);

NOR2xp33_ASAP7_75t_L g1127 ( 
.A(n_836),
.B(n_839),
.Y(n_1127)
);

NOR2x1p5_ASAP7_75t_SL g1128 ( 
.A(n_834),
.B(n_225),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_863),
.B(n_472),
.Y(n_1129)
);

AND2x2_ASAP7_75t_L g1130 ( 
.A(n_837),
.B(n_473),
.Y(n_1130)
);

BUFx2_ASAP7_75t_L g1131 ( 
.A(n_809),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_863),
.B(n_473),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_955),
.A2(n_344),
.B(n_353),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_SL g1134 ( 
.A(n_893),
.B(n_575),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_918),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_955),
.A2(n_962),
.B(n_960),
.Y(n_1136)
);

INVx3_ASAP7_75t_L g1137 ( 
.A(n_893),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_960),
.A2(n_363),
.B(n_432),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_940),
.Y(n_1139)
);

NOR2xp33_ASAP7_75t_R g1140 ( 
.A(n_817),
.B(n_746),
.Y(n_1140)
);

O2A1O1Ixp33_ASAP7_75t_L g1141 ( 
.A1(n_842),
.A2(n_312),
.B(n_322),
.C(n_333),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_956),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_962),
.A2(n_422),
.B(n_403),
.Y(n_1143)
);

INVxp67_ASAP7_75t_L g1144 ( 
.A(n_852),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_951),
.B(n_480),
.Y(n_1145)
);

OAI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_959),
.A2(n_412),
.B(n_394),
.Y(n_1146)
);

A2O1A1Ixp33_ASAP7_75t_L g1147 ( 
.A1(n_929),
.A2(n_350),
.B(n_385),
.C(n_599),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_951),
.B(n_480),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_965),
.Y(n_1149)
);

OAI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_964),
.A2(n_599),
.B(n_596),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_845),
.B(n_596),
.Y(n_1151)
);

NOR2xp33_ASAP7_75t_L g1152 ( 
.A(n_800),
.B(n_17),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_SL g1153 ( 
.A(n_893),
.B(n_575),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_867),
.B(n_746),
.Y(n_1154)
);

BUFx6f_ASAP7_75t_L g1155 ( 
.A(n_893),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_867),
.B(n_746),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_SL g1157 ( 
.A(n_994),
.B(n_938),
.Y(n_1157)
);

BUFx2_ASAP7_75t_L g1158 ( 
.A(n_987),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_980),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_980),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_976),
.Y(n_1161)
);

BUFx3_ASAP7_75t_L g1162 ( 
.A(n_986),
.Y(n_1162)
);

NAND2x1p5_ASAP7_75t_L g1163 ( 
.A(n_1050),
.B(n_922),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_977),
.B(n_910),
.Y(n_1164)
);

NOR2xp33_ASAP7_75t_L g1165 ( 
.A(n_989),
.B(n_807),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_995),
.A2(n_923),
.B(n_922),
.Y(n_1166)
);

NOR2xp33_ASAP7_75t_SL g1167 ( 
.A(n_1050),
.B(n_867),
.Y(n_1167)
);

NOR2xp33_ASAP7_75t_L g1168 ( 
.A(n_989),
.B(n_891),
.Y(n_1168)
);

HB1xp67_ASAP7_75t_L g1169 ( 
.A(n_1005),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_977),
.B(n_948),
.Y(n_1170)
);

OR2x6_ASAP7_75t_SL g1171 ( 
.A(n_1033),
.B(n_1106),
.Y(n_1171)
);

INVx5_ASAP7_75t_L g1172 ( 
.A(n_1107),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_981),
.Y(n_1173)
);

OR2x2_ASAP7_75t_L g1174 ( 
.A(n_1024),
.B(n_919),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_SL g1175 ( 
.A(n_1027),
.B(n_922),
.Y(n_1175)
);

AND2x2_ASAP7_75t_L g1176 ( 
.A(n_1048),
.B(n_840),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_981),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1019),
.A2(n_923),
.B(n_922),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1017),
.B(n_867),
.Y(n_1179)
);

OAI22xp5_ASAP7_75t_L g1180 ( 
.A1(n_1062),
.A2(n_880),
.B1(n_923),
.B2(n_811),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_1073),
.A2(n_996),
.B(n_1000),
.Y(n_1181)
);

INVx3_ASAP7_75t_SL g1182 ( 
.A(n_1087),
.Y(n_1182)
);

BUFx6f_ASAP7_75t_L g1183 ( 
.A(n_1051),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_1009),
.Y(n_1184)
);

BUFx2_ASAP7_75t_L g1185 ( 
.A(n_1038),
.Y(n_1185)
);

AND2x4_ASAP7_75t_L g1186 ( 
.A(n_1107),
.B(n_923),
.Y(n_1186)
);

NOR2xp33_ASAP7_75t_L g1187 ( 
.A(n_991),
.B(n_932),
.Y(n_1187)
);

INVx3_ASAP7_75t_L g1188 ( 
.A(n_1018),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_991),
.B(n_932),
.Y(n_1189)
);

OAI22xp5_ASAP7_75t_SL g1190 ( 
.A1(n_972),
.A2(n_268),
.B1(n_21),
.B2(n_22),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_SL g1191 ( 
.A(n_998),
.B(n_834),
.Y(n_1191)
);

OAI21x1_ASAP7_75t_L g1192 ( 
.A1(n_1007),
.A2(n_834),
.B(n_932),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_985),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1047),
.B(n_932),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_SL g1195 ( 
.A(n_1004),
.B(n_834),
.Y(n_1195)
);

NOR3xp33_ASAP7_75t_SL g1196 ( 
.A(n_972),
.B(n_19),
.C(n_25),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1094),
.B(n_932),
.Y(n_1197)
);

O2A1O1Ixp33_ASAP7_75t_L g1198 ( 
.A1(n_1062),
.A2(n_19),
.B(n_26),
.C(n_28),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1001),
.A2(n_268),
.B(n_588),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1052),
.A2(n_268),
.B(n_588),
.Y(n_1200)
);

NOR2xp33_ASAP7_75t_L g1201 ( 
.A(n_1144),
.B(n_26),
.Y(n_1201)
);

OAI22xp5_ASAP7_75t_L g1202 ( 
.A1(n_1052),
.A2(n_575),
.B1(n_588),
.B2(n_32),
.Y(n_1202)
);

NOR2xp33_ASAP7_75t_L g1203 ( 
.A(n_1122),
.B(n_29),
.Y(n_1203)
);

NOR3xp33_ASAP7_75t_SL g1204 ( 
.A(n_968),
.B(n_29),
.C(n_31),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1013),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1111),
.B(n_834),
.Y(n_1206)
);

O2A1O1Ixp33_ASAP7_75t_L g1207 ( 
.A1(n_1152),
.A2(n_33),
.B(n_35),
.C(n_39),
.Y(n_1207)
);

O2A1O1Ixp33_ASAP7_75t_SL g1208 ( 
.A1(n_1002),
.A2(n_834),
.B(n_40),
.C(n_41),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_SL g1209 ( 
.A(n_1006),
.B(n_588),
.Y(n_1209)
);

AOI21x1_ASAP7_75t_L g1210 ( 
.A1(n_1136),
.A2(n_758),
.B(n_746),
.Y(n_1210)
);

OAI22xp5_ASAP7_75t_L g1211 ( 
.A1(n_1016),
.A2(n_575),
.B1(n_588),
.B2(n_45),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1111),
.B(n_758),
.Y(n_1212)
);

AOI22xp33_ASAP7_75t_L g1213 ( 
.A1(n_1034),
.A2(n_758),
.B1(n_746),
.B2(n_703),
.Y(n_1213)
);

NOR3xp33_ASAP7_75t_SL g1214 ( 
.A(n_968),
.B(n_39),
.C(n_42),
.Y(n_1214)
);

BUFx6f_ASAP7_75t_L g1215 ( 
.A(n_1051),
.Y(n_1215)
);

O2A1O1Ixp33_ASAP7_75t_SL g1216 ( 
.A1(n_1002),
.A2(n_46),
.B(n_49),
.C(n_50),
.Y(n_1216)
);

AND2x4_ASAP7_75t_L g1217 ( 
.A(n_1085),
.B(n_1055),
.Y(n_1217)
);

BUFx6f_ASAP7_75t_L g1218 ( 
.A(n_1051),
.Y(n_1218)
);

AND2x2_ASAP7_75t_L g1219 ( 
.A(n_1079),
.B(n_49),
.Y(n_1219)
);

INVx5_ASAP7_75t_L g1220 ( 
.A(n_1051),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_1009),
.Y(n_1221)
);

INVxp67_ASAP7_75t_L g1222 ( 
.A(n_1085),
.Y(n_1222)
);

AND2x4_ASAP7_75t_L g1223 ( 
.A(n_1058),
.B(n_703),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1099),
.Y(n_1224)
);

NOR2xp33_ASAP7_75t_L g1225 ( 
.A(n_1122),
.B(n_1125),
.Y(n_1225)
);

NOR3xp33_ASAP7_75t_L g1226 ( 
.A(n_1152),
.B(n_1127),
.C(n_1102),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_1022),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1135),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1026),
.A2(n_703),
.B(n_758),
.Y(n_1229)
);

O2A1O1Ixp33_ASAP7_75t_L g1230 ( 
.A1(n_1102),
.A2(n_51),
.B(n_53),
.C(n_55),
.Y(n_1230)
);

A2O1A1Ixp33_ASAP7_75t_L g1231 ( 
.A1(n_1146),
.A2(n_588),
.B(n_575),
.C(n_758),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1125),
.B(n_53),
.Y(n_1232)
);

AND2x4_ASAP7_75t_L g1233 ( 
.A(n_982),
.B(n_703),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_966),
.A2(n_588),
.B(n_138),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_SL g1235 ( 
.A(n_1006),
.B(n_588),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1139),
.Y(n_1236)
);

OR2x2_ASAP7_75t_L g1237 ( 
.A(n_1065),
.B(n_57),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1142),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1117),
.B(n_57),
.Y(n_1239)
);

OAI22xp5_ASAP7_75t_L g1240 ( 
.A1(n_1092),
.A2(n_59),
.B1(n_60),
.B2(n_61),
.Y(n_1240)
);

O2A1O1Ixp33_ASAP7_75t_L g1241 ( 
.A1(n_1109),
.A2(n_59),
.B(n_60),
.C(n_61),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1130),
.B(n_62),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_967),
.A2(n_153),
.B(n_205),
.Y(n_1243)
);

NOR2xp33_ASAP7_75t_R g1244 ( 
.A(n_982),
.B(n_151),
.Y(n_1244)
);

OAI22xp5_ASAP7_75t_L g1245 ( 
.A1(n_1093),
.A2(n_1127),
.B1(n_1090),
.B2(n_1021),
.Y(n_1245)
);

NAND2x1p5_ASAP7_75t_L g1246 ( 
.A(n_969),
.B(n_139),
.Y(n_1246)
);

INVx5_ASAP7_75t_L g1247 ( 
.A(n_1155),
.Y(n_1247)
);

A2O1A1Ixp33_ASAP7_75t_L g1248 ( 
.A1(n_1088),
.A2(n_281),
.B(n_225),
.C(n_69),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1149),
.Y(n_1249)
);

NOR2xp67_ASAP7_75t_L g1250 ( 
.A(n_1068),
.B(n_155),
.Y(n_1250)
);

O2A1O1Ixp33_ASAP7_75t_L g1251 ( 
.A1(n_1109),
.A2(n_64),
.B(n_65),
.C(n_74),
.Y(n_1251)
);

NOR2xp33_ASAP7_75t_L g1252 ( 
.A(n_1078),
.B(n_1110),
.Y(n_1252)
);

AOI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_983),
.A2(n_164),
.B(n_203),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_990),
.A2(n_162),
.B(n_199),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1074),
.B(n_64),
.Y(n_1255)
);

NAND2xp33_ASAP7_75t_L g1256 ( 
.A(n_1155),
.B(n_1018),
.Y(n_1256)
);

NOR3xp33_ASAP7_75t_SL g1257 ( 
.A(n_1072),
.B(n_76),
.C(n_77),
.Y(n_1257)
);

O2A1O1Ixp33_ASAP7_75t_L g1258 ( 
.A1(n_1095),
.A2(n_77),
.B(n_78),
.C(n_281),
.Y(n_1258)
);

INVx2_ASAP7_75t_L g1259 ( 
.A(n_1022),
.Y(n_1259)
);

NOR2xp33_ASAP7_75t_L g1260 ( 
.A(n_1110),
.B(n_79),
.Y(n_1260)
);

NOR2xp67_ASAP7_75t_SL g1261 ( 
.A(n_1054),
.B(n_84),
.Y(n_1261)
);

O2A1O1Ixp33_ASAP7_75t_L g1262 ( 
.A1(n_1074),
.A2(n_281),
.B(n_225),
.C(n_101),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_974),
.A2(n_88),
.B(n_89),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_984),
.A2(n_131),
.B(n_134),
.Y(n_1264)
);

OAI22xp5_ASAP7_75t_L g1265 ( 
.A1(n_1145),
.A2(n_281),
.B1(n_225),
.B2(n_172),
.Y(n_1265)
);

INVx3_ASAP7_75t_L g1266 ( 
.A(n_1018),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1025),
.Y(n_1267)
);

AND2x4_ASAP7_75t_L g1268 ( 
.A(n_969),
.B(n_135),
.Y(n_1268)
);

NOR2xp33_ASAP7_75t_L g1269 ( 
.A(n_1097),
.B(n_166),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1063),
.B(n_281),
.Y(n_1270)
);

BUFx6f_ASAP7_75t_L g1271 ( 
.A(n_1155),
.Y(n_1271)
);

INVx2_ASAP7_75t_SL g1272 ( 
.A(n_1118),
.Y(n_1272)
);

O2A1O1Ixp33_ASAP7_75t_L g1273 ( 
.A1(n_1042),
.A2(n_281),
.B(n_225),
.C(n_180),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1148),
.B(n_281),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1112),
.B(n_281),
.Y(n_1275)
);

OAI22xp33_ASAP7_75t_L g1276 ( 
.A1(n_1121),
.A2(n_225),
.B1(n_179),
.B2(n_182),
.Y(n_1276)
);

AOI21x1_ASAP7_75t_L g1277 ( 
.A1(n_1084),
.A2(n_173),
.B(n_190),
.Y(n_1277)
);

INVx4_ASAP7_75t_L g1278 ( 
.A(n_1039),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1114),
.B(n_192),
.Y(n_1279)
);

AOI21x1_ASAP7_75t_L g1280 ( 
.A1(n_1032),
.A2(n_193),
.B(n_195),
.Y(n_1280)
);

OA21x2_ASAP7_75t_L g1281 ( 
.A1(n_999),
.A2(n_1029),
.B(n_1077),
.Y(n_1281)
);

BUFx6f_ASAP7_75t_L g1282 ( 
.A(n_1155),
.Y(n_1282)
);

OAI22xp5_ASAP7_75t_L g1283 ( 
.A1(n_993),
.A2(n_1053),
.B1(n_1091),
.B2(n_1080),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_988),
.A2(n_975),
.B(n_1014),
.Y(n_1284)
);

OAI22xp5_ASAP7_75t_L g1285 ( 
.A1(n_1076),
.A2(n_1010),
.B1(n_1147),
.B2(n_1056),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1113),
.B(n_1129),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_SL g1287 ( 
.A(n_1018),
.B(n_1043),
.Y(n_1287)
);

O2A1O1Ixp33_ASAP7_75t_L g1288 ( 
.A1(n_1119),
.A2(n_1141),
.B(n_1011),
.C(n_1147),
.Y(n_1288)
);

AOI221xp5_ASAP7_75t_L g1289 ( 
.A1(n_1067),
.A2(n_1143),
.B1(n_1138),
.B2(n_1081),
.C(n_1131),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1025),
.Y(n_1290)
);

AOI22xp5_ASAP7_75t_L g1291 ( 
.A1(n_1036),
.A2(n_1115),
.B1(n_1120),
.B2(n_992),
.Y(n_1291)
);

NOR2xp33_ASAP7_75t_L g1292 ( 
.A(n_1089),
.B(n_1012),
.Y(n_1292)
);

OAI22xp5_ASAP7_75t_L g1293 ( 
.A1(n_1132),
.A2(n_1123),
.B1(n_1036),
.B2(n_1023),
.Y(n_1293)
);

AOI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_979),
.A2(n_1008),
.B(n_1049),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1086),
.Y(n_1295)
);

OAI22xp5_ASAP7_75t_L g1296 ( 
.A1(n_1045),
.A2(n_971),
.B1(n_973),
.B2(n_970),
.Y(n_1296)
);

OAI22xp5_ASAP7_75t_L g1297 ( 
.A1(n_1151),
.A2(n_978),
.B1(n_1003),
.B2(n_1041),
.Y(n_1297)
);

NOR2x1_ASAP7_75t_SL g1298 ( 
.A(n_1040),
.B(n_1134),
.Y(n_1298)
);

NOR2xp33_ASAP7_75t_L g1299 ( 
.A(n_997),
.B(n_1012),
.Y(n_1299)
);

NAND2x1p5_ASAP7_75t_L g1300 ( 
.A(n_997),
.B(n_1137),
.Y(n_1300)
);

AO221x2_ASAP7_75t_L g1301 ( 
.A1(n_1057),
.A2(n_1020),
.B1(n_1035),
.B2(n_1150),
.C(n_1140),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1104),
.Y(n_1302)
);

BUFx2_ASAP7_75t_L g1303 ( 
.A(n_1140),
.Y(n_1303)
);

BUFx8_ASAP7_75t_SL g1304 ( 
.A(n_1015),
.Y(n_1304)
);

A2O1A1Ixp33_ASAP7_75t_L g1305 ( 
.A1(n_1066),
.A2(n_1070),
.B(n_1069),
.C(n_1126),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1104),
.B(n_1124),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1124),
.B(n_1137),
.Y(n_1307)
);

AOI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1059),
.A2(n_1030),
.B(n_1134),
.Y(n_1308)
);

NOR3xp33_ASAP7_75t_SL g1309 ( 
.A(n_1096),
.B(n_1116),
.C(n_1108),
.Y(n_1309)
);

NOR2xp33_ASAP7_75t_L g1310 ( 
.A(n_1040),
.B(n_1064),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_1028),
.Y(n_1311)
);

NOR2xp33_ASAP7_75t_L g1312 ( 
.A(n_1061),
.B(n_1101),
.Y(n_1312)
);

AOI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1101),
.A2(n_1105),
.B(n_1103),
.Y(n_1313)
);

AOI21xp5_ASAP7_75t_L g1314 ( 
.A1(n_1103),
.A2(n_1153),
.B(n_1105),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1098),
.B(n_1100),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_SL g1316 ( 
.A(n_1071),
.B(n_1082),
.Y(n_1316)
);

BUFx2_ASAP7_75t_L g1317 ( 
.A(n_1154),
.Y(n_1317)
);

NAND2x1_ASAP7_75t_L g1318 ( 
.A(n_1046),
.B(n_1031),
.Y(n_1318)
);

BUFx2_ASAP7_75t_SL g1319 ( 
.A(n_1153),
.Y(n_1319)
);

O2A1O1Ixp33_ASAP7_75t_L g1320 ( 
.A1(n_1075),
.A2(n_1083),
.B(n_1133),
.C(n_1060),
.Y(n_1320)
);

INVx2_ASAP7_75t_L g1321 ( 
.A(n_1159),
.Y(n_1321)
);

NOR2xp33_ASAP7_75t_L g1322 ( 
.A(n_1225),
.B(n_1156),
.Y(n_1322)
);

AOI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1181),
.A2(n_1037),
.B(n_1044),
.Y(n_1323)
);

OAI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1164),
.A2(n_1128),
.B(n_1170),
.Y(n_1324)
);

AOI21xp5_ASAP7_75t_L g1325 ( 
.A1(n_1294),
.A2(n_1284),
.B(n_1178),
.Y(n_1325)
);

OAI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1293),
.A2(n_1296),
.B(n_1245),
.Y(n_1326)
);

AOI21xp5_ASAP7_75t_L g1327 ( 
.A1(n_1318),
.A2(n_1206),
.B(n_1308),
.Y(n_1327)
);

AOI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1245),
.A2(n_1316),
.B(n_1166),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1161),
.Y(n_1329)
);

AOI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1281),
.A2(n_1293),
.B(n_1296),
.Y(n_1330)
);

OAI22x1_ASAP7_75t_L g1331 ( 
.A1(n_1203),
.A2(n_1252),
.B1(n_1165),
.B2(n_1260),
.Y(n_1331)
);

AOI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1281),
.A2(n_1315),
.B(n_1187),
.Y(n_1332)
);

BUFx12f_ASAP7_75t_L g1333 ( 
.A(n_1272),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1193),
.Y(n_1334)
);

O2A1O1Ixp33_ASAP7_75t_L g1335 ( 
.A1(n_1226),
.A2(n_1232),
.B(n_1168),
.C(n_1230),
.Y(n_1335)
);

INVx1_ASAP7_75t_SL g1336 ( 
.A(n_1162),
.Y(n_1336)
);

INVxp67_ASAP7_75t_SL g1337 ( 
.A(n_1169),
.Y(n_1337)
);

OA21x2_ASAP7_75t_L g1338 ( 
.A1(n_1311),
.A2(n_1200),
.B(n_1199),
.Y(n_1338)
);

AOI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1320),
.A2(n_1234),
.B(n_1189),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1205),
.Y(n_1340)
);

OAI22xp5_ASAP7_75t_L g1341 ( 
.A1(n_1255),
.A2(n_1202),
.B1(n_1242),
.B2(n_1239),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1283),
.B(n_1286),
.Y(n_1342)
);

CKINVDCx20_ASAP7_75t_R g1343 ( 
.A(n_1182),
.Y(n_1343)
);

OR2x2_ASAP7_75t_L g1344 ( 
.A(n_1185),
.B(n_1174),
.Y(n_1344)
);

AO31x2_ASAP7_75t_L g1345 ( 
.A1(n_1265),
.A2(n_1283),
.A3(n_1275),
.B(n_1248),
.Y(n_1345)
);

A2O1A1Ixp33_ASAP7_75t_L g1346 ( 
.A1(n_1288),
.A2(n_1273),
.B(n_1262),
.C(n_1207),
.Y(n_1346)
);

AOI22xp5_ASAP7_75t_L g1347 ( 
.A1(n_1301),
.A2(n_1190),
.B1(n_1217),
.B2(n_1222),
.Y(n_1347)
);

INVx2_ASAP7_75t_SL g1348 ( 
.A(n_1303),
.Y(n_1348)
);

INVx4_ASAP7_75t_L g1349 ( 
.A(n_1220),
.Y(n_1349)
);

AND2x4_ASAP7_75t_L g1350 ( 
.A(n_1278),
.B(n_1220),
.Y(n_1350)
);

OAI21x1_ASAP7_75t_L g1351 ( 
.A1(n_1192),
.A2(n_1314),
.B(n_1313),
.Y(n_1351)
);

AOI21xp5_ASAP7_75t_L g1352 ( 
.A1(n_1256),
.A2(n_1254),
.B(n_1253),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1224),
.B(n_1291),
.Y(n_1353)
);

AO31x2_ASAP7_75t_L g1354 ( 
.A1(n_1265),
.A2(n_1285),
.A3(n_1310),
.B(n_1297),
.Y(n_1354)
);

AOI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1180),
.A2(n_1297),
.B(n_1175),
.Y(n_1355)
);

AOI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1180),
.A2(n_1285),
.B(n_1167),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1301),
.B(n_1267),
.Y(n_1357)
);

AO31x2_ASAP7_75t_L g1358 ( 
.A1(n_1279),
.A2(n_1270),
.A3(n_1298),
.B(n_1274),
.Y(n_1358)
);

OAI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1229),
.A2(n_1277),
.B(n_1280),
.Y(n_1359)
);

AOI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1167),
.A2(n_1305),
.B(n_1212),
.Y(n_1360)
);

BUFx4_ASAP7_75t_SL g1361 ( 
.A(n_1304),
.Y(n_1361)
);

NOR2x1_ASAP7_75t_L g1362 ( 
.A(n_1278),
.B(n_1269),
.Y(n_1362)
);

O2A1O1Ixp33_ASAP7_75t_SL g1363 ( 
.A1(n_1209),
.A2(n_1235),
.B(n_1179),
.C(n_1202),
.Y(n_1363)
);

O2A1O1Ixp33_ASAP7_75t_SL g1364 ( 
.A1(n_1195),
.A2(n_1191),
.B(n_1198),
.C(n_1276),
.Y(n_1364)
);

AOI21xp5_ASAP7_75t_L g1365 ( 
.A1(n_1243),
.A2(n_1263),
.B(n_1312),
.Y(n_1365)
);

INVx3_ASAP7_75t_L g1366 ( 
.A(n_1163),
.Y(n_1366)
);

O2A1O1Ixp33_ASAP7_75t_SL g1367 ( 
.A1(n_1240),
.A2(n_1237),
.B(n_1194),
.C(n_1197),
.Y(n_1367)
);

NOR4xp25_ASAP7_75t_L g1368 ( 
.A(n_1241),
.B(n_1251),
.C(n_1240),
.D(n_1258),
.Y(n_1368)
);

AND2x4_ASAP7_75t_L g1369 ( 
.A(n_1220),
.B(n_1247),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1290),
.B(n_1295),
.Y(n_1370)
);

INVx3_ASAP7_75t_L g1371 ( 
.A(n_1163),
.Y(n_1371)
);

OAI21x1_ASAP7_75t_L g1372 ( 
.A1(n_1210),
.A2(n_1287),
.B(n_1264),
.Y(n_1372)
);

AND2x4_ASAP7_75t_L g1373 ( 
.A(n_1220),
.B(n_1247),
.Y(n_1373)
);

OAI22xp5_ASAP7_75t_L g1374 ( 
.A1(n_1257),
.A2(n_1196),
.B1(n_1211),
.B2(n_1219),
.Y(n_1374)
);

BUFx12f_ASAP7_75t_L g1375 ( 
.A(n_1183),
.Y(n_1375)
);

BUFx10_ASAP7_75t_L g1376 ( 
.A(n_1201),
.Y(n_1376)
);

AOI22xp33_ASAP7_75t_L g1377 ( 
.A1(n_1157),
.A2(n_1236),
.B1(n_1249),
.B2(n_1238),
.Y(n_1377)
);

INVx3_ASAP7_75t_L g1378 ( 
.A(n_1247),
.Y(n_1378)
);

AND2x4_ASAP7_75t_L g1379 ( 
.A(n_1247),
.B(n_1186),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1160),
.Y(n_1380)
);

CKINVDCx5p33_ASAP7_75t_R g1381 ( 
.A(n_1171),
.Y(n_1381)
);

OAI21x1_ASAP7_75t_L g1382 ( 
.A1(n_1246),
.A2(n_1307),
.B(n_1266),
.Y(n_1382)
);

NOR2xp33_ASAP7_75t_L g1383 ( 
.A(n_1292),
.B(n_1299),
.Y(n_1383)
);

CKINVDCx5p33_ASAP7_75t_R g1384 ( 
.A(n_1244),
.Y(n_1384)
);

AOI21xp5_ASAP7_75t_L g1385 ( 
.A1(n_1208),
.A2(n_1211),
.B(n_1231),
.Y(n_1385)
);

A2O1A1Ixp33_ASAP7_75t_L g1386 ( 
.A1(n_1289),
.A2(n_1250),
.B(n_1204),
.C(n_1214),
.Y(n_1386)
);

OR2x2_ASAP7_75t_L g1387 ( 
.A(n_1228),
.B(n_1302),
.Y(n_1387)
);

OAI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1309),
.A2(n_1216),
.B(n_1186),
.Y(n_1388)
);

AOI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1268),
.A2(n_1172),
.B(n_1266),
.Y(n_1389)
);

INVx1_ASAP7_75t_SL g1390 ( 
.A(n_1319),
.Y(n_1390)
);

AOI21xp5_ASAP7_75t_L g1391 ( 
.A1(n_1268),
.A2(n_1172),
.B(n_1188),
.Y(n_1391)
);

INVx2_ASAP7_75t_L g1392 ( 
.A(n_1173),
.Y(n_1392)
);

AOI221x1_ASAP7_75t_L g1393 ( 
.A1(n_1306),
.A2(n_1177),
.B1(n_1184),
.B2(n_1259),
.C(n_1227),
.Y(n_1393)
);

INVx6_ASAP7_75t_L g1394 ( 
.A(n_1215),
.Y(n_1394)
);

O2A1O1Ixp33_ASAP7_75t_L g1395 ( 
.A1(n_1300),
.A2(n_1188),
.B(n_1223),
.C(n_1317),
.Y(n_1395)
);

AO21x1_ASAP7_75t_L g1396 ( 
.A1(n_1300),
.A2(n_1223),
.B(n_1221),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1172),
.B(n_1282),
.Y(n_1397)
);

INVx4_ASAP7_75t_L g1398 ( 
.A(n_1215),
.Y(n_1398)
);

BUFx12f_ASAP7_75t_L g1399 ( 
.A(n_1215),
.Y(n_1399)
);

O2A1O1Ixp33_ASAP7_75t_L g1400 ( 
.A1(n_1233),
.A2(n_1213),
.B(n_1261),
.C(n_1172),
.Y(n_1400)
);

O2A1O1Ixp5_ASAP7_75t_L g1401 ( 
.A1(n_1233),
.A2(n_1218),
.B(n_1271),
.C(n_1282),
.Y(n_1401)
);

CKINVDCx5p33_ASAP7_75t_R g1402 ( 
.A(n_1218),
.Y(n_1402)
);

OAI21xp5_ASAP7_75t_SL g1403 ( 
.A1(n_1271),
.A2(n_1203),
.B(n_1225),
.Y(n_1403)
);

INVx1_ASAP7_75t_SL g1404 ( 
.A(n_1162),
.Y(n_1404)
);

AO31x2_ASAP7_75t_L g1405 ( 
.A1(n_1311),
.A2(n_1296),
.A3(n_1265),
.B(n_1293),
.Y(n_1405)
);

BUFx3_ASAP7_75t_L g1406 ( 
.A(n_1162),
.Y(n_1406)
);

BUFx6f_ASAP7_75t_L g1407 ( 
.A(n_1220),
.Y(n_1407)
);

OAI22xp5_ASAP7_75t_L g1408 ( 
.A1(n_1164),
.A2(n_1170),
.B1(n_977),
.B2(n_1062),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1176),
.B(n_994),
.Y(n_1409)
);

AO31x2_ASAP7_75t_L g1410 ( 
.A1(n_1311),
.A2(n_1296),
.A3(n_1265),
.B(n_1293),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1176),
.B(n_994),
.Y(n_1411)
);

AOI22xp5_ASAP7_75t_L g1412 ( 
.A1(n_1225),
.A2(n_1203),
.B1(n_647),
.B2(n_1226),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1176),
.B(n_994),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_SL g1414 ( 
.A(n_1225),
.B(n_989),
.Y(n_1414)
);

AOI21xp5_ASAP7_75t_L g1415 ( 
.A1(n_1181),
.A2(n_995),
.B(n_1019),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1164),
.B(n_977),
.Y(n_1416)
);

AND2x4_ASAP7_75t_L g1417 ( 
.A(n_1278),
.B(n_1217),
.Y(n_1417)
);

A2O1A1Ixp33_ASAP7_75t_L g1418 ( 
.A1(n_1225),
.A2(n_1203),
.B(n_977),
.C(n_1260),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_SL g1419 ( 
.A1(n_1225),
.A2(n_458),
.B1(n_504),
.B2(n_479),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1164),
.B(n_977),
.Y(n_1420)
);

A2O1A1Ixp33_ASAP7_75t_L g1421 ( 
.A1(n_1225),
.A2(n_1203),
.B(n_977),
.C(n_1260),
.Y(n_1421)
);

OAI21x1_ASAP7_75t_L g1422 ( 
.A1(n_1284),
.A2(n_1294),
.B(n_1308),
.Y(n_1422)
);

BUFx12f_ASAP7_75t_L g1423 ( 
.A(n_1272),
.Y(n_1423)
);

AO31x2_ASAP7_75t_L g1424 ( 
.A1(n_1311),
.A2(n_1296),
.A3(n_1265),
.B(n_1293),
.Y(n_1424)
);

OAI21x1_ASAP7_75t_L g1425 ( 
.A1(n_1284),
.A2(n_1294),
.B(n_1308),
.Y(n_1425)
);

AO31x2_ASAP7_75t_L g1426 ( 
.A1(n_1311),
.A2(n_1296),
.A3(n_1265),
.B(n_1293),
.Y(n_1426)
);

BUFx8_ASAP7_75t_L g1427 ( 
.A(n_1158),
.Y(n_1427)
);

AOI21xp5_ASAP7_75t_L g1428 ( 
.A1(n_1181),
.A2(n_995),
.B(n_1019),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1164),
.B(n_977),
.Y(n_1429)
);

OAI21x1_ASAP7_75t_L g1430 ( 
.A1(n_1284),
.A2(n_1294),
.B(n_1308),
.Y(n_1430)
);

A2O1A1Ixp33_ASAP7_75t_L g1431 ( 
.A1(n_1225),
.A2(n_1203),
.B(n_977),
.C(n_1260),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1176),
.B(n_994),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1164),
.B(n_977),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1159),
.Y(n_1434)
);

AOI21xp5_ASAP7_75t_L g1435 ( 
.A1(n_1181),
.A2(n_995),
.B(n_1019),
.Y(n_1435)
);

OAI21x1_ASAP7_75t_L g1436 ( 
.A1(n_1284),
.A2(n_1294),
.B(n_1308),
.Y(n_1436)
);

AOI22xp5_ASAP7_75t_L g1437 ( 
.A1(n_1225),
.A2(n_1203),
.B1(n_647),
.B2(n_1226),
.Y(n_1437)
);

INVx3_ASAP7_75t_L g1438 ( 
.A(n_1163),
.Y(n_1438)
);

OAI22x1_ASAP7_75t_L g1439 ( 
.A1(n_1225),
.A2(n_1203),
.B1(n_998),
.B2(n_647),
.Y(n_1439)
);

OAI21xp5_ASAP7_75t_L g1440 ( 
.A1(n_1164),
.A2(n_977),
.B(n_1052),
.Y(n_1440)
);

INVx1_ASAP7_75t_SL g1441 ( 
.A(n_1162),
.Y(n_1441)
);

NOR4xp25_ASAP7_75t_L g1442 ( 
.A(n_1207),
.B(n_1230),
.C(n_1251),
.D(n_1241),
.Y(n_1442)
);

NOR2xp67_ASAP7_75t_L g1443 ( 
.A(n_1278),
.B(n_823),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1164),
.B(n_977),
.Y(n_1444)
);

O2A1O1Ixp33_ASAP7_75t_SL g1445 ( 
.A1(n_1164),
.A2(n_1170),
.B(n_1062),
.C(n_995),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1176),
.B(n_994),
.Y(n_1446)
);

NOR2xp33_ASAP7_75t_L g1447 ( 
.A(n_1225),
.B(n_647),
.Y(n_1447)
);

CKINVDCx20_ASAP7_75t_R g1448 ( 
.A(n_1182),
.Y(n_1448)
);

BUFx6f_ASAP7_75t_L g1449 ( 
.A(n_1220),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1225),
.B(n_789),
.Y(n_1450)
);

BUFx6f_ASAP7_75t_L g1451 ( 
.A(n_1220),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1225),
.B(n_789),
.Y(n_1452)
);

BUFx8_ASAP7_75t_SL g1453 ( 
.A(n_1304),
.Y(n_1453)
);

AOI21xp5_ASAP7_75t_L g1454 ( 
.A1(n_1181),
.A2(n_995),
.B(n_1019),
.Y(n_1454)
);

BUFx12f_ASAP7_75t_L g1455 ( 
.A(n_1272),
.Y(n_1455)
);

AO31x2_ASAP7_75t_L g1456 ( 
.A1(n_1311),
.A2(n_1296),
.A3(n_1265),
.B(n_1293),
.Y(n_1456)
);

AOI221x1_ASAP7_75t_L g1457 ( 
.A1(n_1225),
.A2(n_1226),
.B1(n_1202),
.B2(n_1265),
.C(n_1203),
.Y(n_1457)
);

OAI21x1_ASAP7_75t_L g1458 ( 
.A1(n_1284),
.A2(n_1294),
.B(n_1308),
.Y(n_1458)
);

AO31x2_ASAP7_75t_L g1459 ( 
.A1(n_1311),
.A2(n_1296),
.A3(n_1265),
.B(n_1293),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1159),
.Y(n_1460)
);

OAI21x1_ASAP7_75t_L g1461 ( 
.A1(n_1284),
.A2(n_1294),
.B(n_1308),
.Y(n_1461)
);

OAI22xp5_ASAP7_75t_L g1462 ( 
.A1(n_1164),
.A2(n_1170),
.B1(n_977),
.B2(n_1062),
.Y(n_1462)
);

AOI21xp5_ASAP7_75t_L g1463 ( 
.A1(n_1181),
.A2(n_995),
.B(n_1019),
.Y(n_1463)
);

OAI21x1_ASAP7_75t_L g1464 ( 
.A1(n_1284),
.A2(n_1294),
.B(n_1308),
.Y(n_1464)
);

BUFx2_ASAP7_75t_L g1465 ( 
.A(n_1162),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1164),
.B(n_977),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1159),
.Y(n_1467)
);

AO22x2_ASAP7_75t_L g1468 ( 
.A1(n_1226),
.A2(n_1202),
.B1(n_1245),
.B2(n_1283),
.Y(n_1468)
);

OAI21x1_ASAP7_75t_L g1469 ( 
.A1(n_1284),
.A2(n_1294),
.B(n_1308),
.Y(n_1469)
);

OAI21x1_ASAP7_75t_L g1470 ( 
.A1(n_1284),
.A2(n_1294),
.B(n_1308),
.Y(n_1470)
);

AOI21xp5_ASAP7_75t_L g1471 ( 
.A1(n_1181),
.A2(n_995),
.B(n_1019),
.Y(n_1471)
);

INVxp67_ASAP7_75t_L g1472 ( 
.A(n_1169),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1164),
.B(n_977),
.Y(n_1473)
);

AOI21xp5_ASAP7_75t_L g1474 ( 
.A1(n_1181),
.A2(n_995),
.B(n_1019),
.Y(n_1474)
);

AND3x2_ASAP7_75t_L g1475 ( 
.A(n_1225),
.B(n_1081),
.C(n_635),
.Y(n_1475)
);

AOI221xp5_ASAP7_75t_L g1476 ( 
.A1(n_1176),
.A2(n_1225),
.B1(n_1203),
.B2(n_774),
.C(n_919),
.Y(n_1476)
);

AO31x2_ASAP7_75t_L g1477 ( 
.A1(n_1311),
.A2(n_1296),
.A3(n_1265),
.B(n_1293),
.Y(n_1477)
);

AOI21xp5_ASAP7_75t_L g1478 ( 
.A1(n_1181),
.A2(n_995),
.B(n_1019),
.Y(n_1478)
);

OAI21x1_ASAP7_75t_L g1479 ( 
.A1(n_1284),
.A2(n_1294),
.B(n_1308),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1161),
.Y(n_1480)
);

AOI21x1_ASAP7_75t_L g1481 ( 
.A1(n_1318),
.A2(n_1284),
.B(n_1181),
.Y(n_1481)
);

INVx4_ASAP7_75t_L g1482 ( 
.A(n_1220),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1225),
.B(n_789),
.Y(n_1483)
);

AOI21xp5_ASAP7_75t_L g1484 ( 
.A1(n_1181),
.A2(n_995),
.B(n_1019),
.Y(n_1484)
);

BUFx4_ASAP7_75t_SL g1485 ( 
.A(n_1162),
.Y(n_1485)
);

AOI22xp5_ASAP7_75t_L g1486 ( 
.A1(n_1476),
.A2(n_1331),
.B1(n_1421),
.B2(n_1418),
.Y(n_1486)
);

BUFx3_ASAP7_75t_L g1487 ( 
.A(n_1406),
.Y(n_1487)
);

BUFx2_ASAP7_75t_L g1488 ( 
.A(n_1402),
.Y(n_1488)
);

AOI22xp5_ASAP7_75t_L g1489 ( 
.A1(n_1431),
.A2(n_1447),
.B1(n_1412),
.B2(n_1437),
.Y(n_1489)
);

AOI22xp33_ASAP7_75t_SL g1490 ( 
.A1(n_1341),
.A2(n_1468),
.B1(n_1462),
.B2(n_1408),
.Y(n_1490)
);

BUFx8_ASAP7_75t_L g1491 ( 
.A(n_1361),
.Y(n_1491)
);

INVx6_ASAP7_75t_L g1492 ( 
.A(n_1417),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1387),
.Y(n_1493)
);

CKINVDCx20_ASAP7_75t_R g1494 ( 
.A(n_1453),
.Y(n_1494)
);

INVx4_ASAP7_75t_L g1495 ( 
.A(n_1375),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1329),
.Y(n_1496)
);

AOI22xp33_ASAP7_75t_L g1497 ( 
.A1(n_1341),
.A2(n_1462),
.B1(n_1408),
.B2(n_1446),
.Y(n_1497)
);

OAI22xp5_ASAP7_75t_SL g1498 ( 
.A1(n_1439),
.A2(n_1381),
.B1(n_1450),
.B2(n_1483),
.Y(n_1498)
);

AOI22xp33_ASAP7_75t_SL g1499 ( 
.A1(n_1468),
.A2(n_1473),
.B1(n_1433),
.B2(n_1429),
.Y(n_1499)
);

AOI22xp33_ASAP7_75t_L g1500 ( 
.A1(n_1409),
.A2(n_1411),
.B1(n_1432),
.B2(n_1413),
.Y(n_1500)
);

CKINVDCx11_ASAP7_75t_R g1501 ( 
.A(n_1333),
.Y(n_1501)
);

BUFx6f_ASAP7_75t_L g1502 ( 
.A(n_1407),
.Y(n_1502)
);

OAI22xp33_ASAP7_75t_L g1503 ( 
.A1(n_1457),
.A2(n_1473),
.B1(n_1420),
.B2(n_1466),
.Y(n_1503)
);

CKINVDCx11_ASAP7_75t_R g1504 ( 
.A(n_1423),
.Y(n_1504)
);

AOI22xp33_ASAP7_75t_L g1505 ( 
.A1(n_1416),
.A2(n_1466),
.B1(n_1433),
.B2(n_1429),
.Y(n_1505)
);

INVx6_ASAP7_75t_L g1506 ( 
.A(n_1399),
.Y(n_1506)
);

INVxp67_ASAP7_75t_SL g1507 ( 
.A(n_1326),
.Y(n_1507)
);

AOI21xp5_ASAP7_75t_L g1508 ( 
.A1(n_1365),
.A2(n_1352),
.B(n_1326),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1334),
.Y(n_1509)
);

AOI22xp33_ASAP7_75t_L g1510 ( 
.A1(n_1416),
.A2(n_1420),
.B1(n_1444),
.B2(n_1452),
.Y(n_1510)
);

OAI21xp33_ASAP7_75t_SL g1511 ( 
.A1(n_1444),
.A2(n_1440),
.B(n_1414),
.Y(n_1511)
);

INVx6_ASAP7_75t_L g1512 ( 
.A(n_1427),
.Y(n_1512)
);

AOI22xp33_ASAP7_75t_L g1513 ( 
.A1(n_1374),
.A2(n_1419),
.B1(n_1440),
.B2(n_1475),
.Y(n_1513)
);

CKINVDCx14_ASAP7_75t_R g1514 ( 
.A(n_1384),
.Y(n_1514)
);

CKINVDCx11_ASAP7_75t_R g1515 ( 
.A(n_1455),
.Y(n_1515)
);

INVx1_ASAP7_75t_SL g1516 ( 
.A(n_1485),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1340),
.Y(n_1517)
);

OAI21xp5_ASAP7_75t_SL g1518 ( 
.A1(n_1335),
.A2(n_1374),
.B(n_1386),
.Y(n_1518)
);

AOI22xp33_ASAP7_75t_L g1519 ( 
.A1(n_1357),
.A2(n_1356),
.B1(n_1344),
.B2(n_1322),
.Y(n_1519)
);

BUFx8_ASAP7_75t_L g1520 ( 
.A(n_1465),
.Y(n_1520)
);

BUFx12f_ASAP7_75t_L g1521 ( 
.A(n_1427),
.Y(n_1521)
);

AOI22xp33_ASAP7_75t_SL g1522 ( 
.A1(n_1357),
.A2(n_1342),
.B1(n_1353),
.B2(n_1376),
.Y(n_1522)
);

BUFx12f_ASAP7_75t_L g1523 ( 
.A(n_1376),
.Y(n_1523)
);

CKINVDCx11_ASAP7_75t_R g1524 ( 
.A(n_1336),
.Y(n_1524)
);

OAI22xp5_ASAP7_75t_L g1525 ( 
.A1(n_1346),
.A2(n_1403),
.B1(n_1347),
.B2(n_1337),
.Y(n_1525)
);

INVx6_ASAP7_75t_L g1526 ( 
.A(n_1350),
.Y(n_1526)
);

BUFx2_ASAP7_75t_SL g1527 ( 
.A(n_1443),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1321),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1480),
.Y(n_1529)
);

INVx3_ASAP7_75t_L g1530 ( 
.A(n_1369),
.Y(n_1530)
);

BUFx10_ASAP7_75t_L g1531 ( 
.A(n_1394),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1370),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1380),
.Y(n_1533)
);

AOI22xp33_ASAP7_75t_L g1534 ( 
.A1(n_1377),
.A2(n_1467),
.B1(n_1392),
.B2(n_1434),
.Y(n_1534)
);

BUFx3_ASAP7_75t_L g1535 ( 
.A(n_1404),
.Y(n_1535)
);

OAI22xp5_ASAP7_75t_L g1536 ( 
.A1(n_1472),
.A2(n_1355),
.B1(n_1383),
.B2(n_1342),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1370),
.Y(n_1537)
);

INVxp67_ASAP7_75t_L g1538 ( 
.A(n_1353),
.Y(n_1538)
);

CKINVDCx5p33_ASAP7_75t_R g1539 ( 
.A(n_1441),
.Y(n_1539)
);

CKINVDCx11_ASAP7_75t_R g1540 ( 
.A(n_1441),
.Y(n_1540)
);

CKINVDCx20_ASAP7_75t_R g1541 ( 
.A(n_1348),
.Y(n_1541)
);

BUFx10_ASAP7_75t_L g1542 ( 
.A(n_1394),
.Y(n_1542)
);

AOI22xp33_ASAP7_75t_L g1543 ( 
.A1(n_1324),
.A2(n_1385),
.B1(n_1460),
.B2(n_1362),
.Y(n_1543)
);

BUFx12f_ASAP7_75t_SL g1544 ( 
.A(n_1407),
.Y(n_1544)
);

AOI22xp33_ASAP7_75t_L g1545 ( 
.A1(n_1324),
.A2(n_1396),
.B1(n_1330),
.B2(n_1390),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1393),
.Y(n_1546)
);

OR2x6_ASAP7_75t_L g1547 ( 
.A(n_1400),
.B(n_1395),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1382),
.Y(n_1548)
);

OAI22xp33_ASAP7_75t_L g1549 ( 
.A1(n_1388),
.A2(n_1368),
.B1(n_1442),
.B2(n_1397),
.Y(n_1549)
);

INVx2_ASAP7_75t_SL g1550 ( 
.A(n_1379),
.Y(n_1550)
);

AOI22xp33_ASAP7_75t_L g1551 ( 
.A1(n_1388),
.A2(n_1442),
.B1(n_1368),
.B2(n_1332),
.Y(n_1551)
);

NAND2x1p5_ASAP7_75t_L g1552 ( 
.A(n_1369),
.B(n_1373),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1445),
.Y(n_1553)
);

AOI22xp33_ASAP7_75t_L g1554 ( 
.A1(n_1366),
.A2(n_1371),
.B1(n_1438),
.B2(n_1478),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1401),
.Y(n_1555)
);

INVx1_ASAP7_75t_SL g1556 ( 
.A(n_1373),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1398),
.B(n_1371),
.Y(n_1557)
);

AOI22xp33_ASAP7_75t_L g1558 ( 
.A1(n_1366),
.A2(n_1438),
.B1(n_1338),
.B2(n_1391),
.Y(n_1558)
);

AOI22xp33_ASAP7_75t_L g1559 ( 
.A1(n_1415),
.A2(n_1484),
.B1(n_1435),
.B2(n_1474),
.Y(n_1559)
);

AOI22xp33_ASAP7_75t_L g1560 ( 
.A1(n_1428),
.A2(n_1454),
.B1(n_1471),
.B2(n_1463),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1367),
.Y(n_1561)
);

CKINVDCx6p67_ASAP7_75t_R g1562 ( 
.A(n_1449),
.Y(n_1562)
);

INVxp67_ASAP7_75t_SL g1563 ( 
.A(n_1422),
.Y(n_1563)
);

AOI22xp33_ASAP7_75t_L g1564 ( 
.A1(n_1360),
.A2(n_1328),
.B1(n_1354),
.B2(n_1389),
.Y(n_1564)
);

INVx3_ASAP7_75t_L g1565 ( 
.A(n_1449),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1378),
.Y(n_1566)
);

AOI22xp33_ASAP7_75t_L g1567 ( 
.A1(n_1354),
.A2(n_1339),
.B1(n_1449),
.B2(n_1451),
.Y(n_1567)
);

INVx8_ASAP7_75t_L g1568 ( 
.A(n_1451),
.Y(n_1568)
);

INVx5_ASAP7_75t_L g1569 ( 
.A(n_1349),
.Y(n_1569)
);

HB1xp67_ASAP7_75t_L g1570 ( 
.A(n_1405),
.Y(n_1570)
);

AOI22xp33_ASAP7_75t_L g1571 ( 
.A1(n_1482),
.A2(n_1345),
.B1(n_1363),
.B2(n_1372),
.Y(n_1571)
);

AOI22xp33_ASAP7_75t_L g1572 ( 
.A1(n_1410),
.A2(n_1456),
.B1(n_1426),
.B2(n_1459),
.Y(n_1572)
);

AOI22xp33_ASAP7_75t_L g1573 ( 
.A1(n_1323),
.A2(n_1327),
.B1(n_1351),
.B2(n_1359),
.Y(n_1573)
);

INVx1_ASAP7_75t_SL g1574 ( 
.A(n_1325),
.Y(n_1574)
);

OAI22xp5_ASAP7_75t_L g1575 ( 
.A1(n_1481),
.A2(n_1364),
.B1(n_1456),
.B2(n_1410),
.Y(n_1575)
);

CKINVDCx11_ASAP7_75t_R g1576 ( 
.A(n_1424),
.Y(n_1576)
);

OAI22xp33_ASAP7_75t_L g1577 ( 
.A1(n_1424),
.A2(n_1459),
.B1(n_1477),
.B2(n_1426),
.Y(n_1577)
);

BUFx10_ASAP7_75t_L g1578 ( 
.A(n_1358),
.Y(n_1578)
);

CKINVDCx11_ASAP7_75t_R g1579 ( 
.A(n_1424),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1426),
.B(n_1459),
.Y(n_1580)
);

AOI22xp33_ASAP7_75t_L g1581 ( 
.A1(n_1425),
.A2(n_1430),
.B1(n_1436),
.B2(n_1479),
.Y(n_1581)
);

CKINVDCx20_ASAP7_75t_R g1582 ( 
.A(n_1456),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1477),
.Y(n_1583)
);

AOI22xp33_ASAP7_75t_L g1584 ( 
.A1(n_1458),
.A2(n_1461),
.B1(n_1464),
.B2(n_1469),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1477),
.B(n_1470),
.Y(n_1585)
);

AOI22xp33_ASAP7_75t_L g1586 ( 
.A1(n_1476),
.A2(n_1225),
.B1(n_1331),
.B2(n_1203),
.Y(n_1586)
);

INVx1_ASAP7_75t_SL g1587 ( 
.A(n_1485),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1387),
.Y(n_1588)
);

AOI22xp33_ASAP7_75t_SL g1589 ( 
.A1(n_1341),
.A2(n_1225),
.B1(n_1203),
.B2(n_602),
.Y(n_1589)
);

AOI22xp33_ASAP7_75t_L g1590 ( 
.A1(n_1476),
.A2(n_1225),
.B1(n_1331),
.B2(n_1203),
.Y(n_1590)
);

OAI22xp5_ASAP7_75t_L g1591 ( 
.A1(n_1418),
.A2(n_1421),
.B1(n_1431),
.B2(n_1412),
.Y(n_1591)
);

OAI22x1_ASAP7_75t_L g1592 ( 
.A1(n_1412),
.A2(n_1437),
.B1(n_1225),
.B2(n_1347),
.Y(n_1592)
);

CKINVDCx11_ASAP7_75t_R g1593 ( 
.A(n_1343),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1387),
.Y(n_1594)
);

AOI22xp5_ASAP7_75t_L g1595 ( 
.A1(n_1476),
.A2(n_1225),
.B1(n_1331),
.B2(n_1418),
.Y(n_1595)
);

INVx1_ASAP7_75t_SL g1596 ( 
.A(n_1485),
.Y(n_1596)
);

INVx6_ASAP7_75t_L g1597 ( 
.A(n_1417),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1387),
.Y(n_1598)
);

AOI22xp33_ASAP7_75t_SL g1599 ( 
.A1(n_1341),
.A2(n_1225),
.B1(n_1203),
.B2(n_602),
.Y(n_1599)
);

INVx8_ASAP7_75t_L g1600 ( 
.A(n_1333),
.Y(n_1600)
);

INVx6_ASAP7_75t_L g1601 ( 
.A(n_1417),
.Y(n_1601)
);

CKINVDCx20_ASAP7_75t_R g1602 ( 
.A(n_1453),
.Y(n_1602)
);

AOI22xp5_ASAP7_75t_L g1603 ( 
.A1(n_1476),
.A2(n_1225),
.B1(n_1331),
.B2(n_1418),
.Y(n_1603)
);

NAND2x1p5_ASAP7_75t_L g1604 ( 
.A(n_1369),
.B(n_1373),
.Y(n_1604)
);

AOI22xp33_ASAP7_75t_L g1605 ( 
.A1(n_1476),
.A2(n_1225),
.B1(n_1331),
.B2(n_1203),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1387),
.Y(n_1606)
);

AOI22x1_ASAP7_75t_SL g1607 ( 
.A1(n_1381),
.A2(n_1448),
.B1(n_1343),
.B2(n_934),
.Y(n_1607)
);

INVx4_ASAP7_75t_L g1608 ( 
.A(n_1417),
.Y(n_1608)
);

AOI22xp33_ASAP7_75t_L g1609 ( 
.A1(n_1476),
.A2(n_1225),
.B1(n_1331),
.B2(n_1203),
.Y(n_1609)
);

CKINVDCx11_ASAP7_75t_R g1610 ( 
.A(n_1343),
.Y(n_1610)
);

BUFx4f_ASAP7_75t_SL g1611 ( 
.A(n_1343),
.Y(n_1611)
);

OAI21xp5_ASAP7_75t_L g1612 ( 
.A1(n_1418),
.A2(n_1431),
.B(n_1421),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_1387),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1387),
.Y(n_1614)
);

AOI22xp33_ASAP7_75t_L g1615 ( 
.A1(n_1476),
.A2(n_1225),
.B1(n_1331),
.B2(n_1203),
.Y(n_1615)
);

CKINVDCx11_ASAP7_75t_R g1616 ( 
.A(n_1343),
.Y(n_1616)
);

BUFx3_ASAP7_75t_L g1617 ( 
.A(n_1406),
.Y(n_1617)
);

BUFx2_ASAP7_75t_L g1618 ( 
.A(n_1402),
.Y(n_1618)
);

OAI22x1_ASAP7_75t_L g1619 ( 
.A1(n_1412),
.A2(n_1437),
.B1(n_1225),
.B2(n_1347),
.Y(n_1619)
);

AOI22xp33_ASAP7_75t_L g1620 ( 
.A1(n_1476),
.A2(n_1225),
.B1(n_1331),
.B2(n_1203),
.Y(n_1620)
);

AOI22xp33_ASAP7_75t_SL g1621 ( 
.A1(n_1341),
.A2(n_1225),
.B1(n_1203),
.B2(n_602),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1416),
.B(n_1420),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1387),
.Y(n_1623)
);

CKINVDCx5p33_ASAP7_75t_R g1624 ( 
.A(n_1361),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1387),
.Y(n_1625)
);

AOI22xp33_ASAP7_75t_SL g1626 ( 
.A1(n_1341),
.A2(n_1225),
.B1(n_1203),
.B2(n_602),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1387),
.Y(n_1627)
);

AOI22xp33_ASAP7_75t_L g1628 ( 
.A1(n_1476),
.A2(n_1225),
.B1(n_1331),
.B2(n_1203),
.Y(n_1628)
);

AOI22xp33_ASAP7_75t_L g1629 ( 
.A1(n_1476),
.A2(n_1225),
.B1(n_1331),
.B2(n_1203),
.Y(n_1629)
);

INVx8_ASAP7_75t_L g1630 ( 
.A(n_1333),
.Y(n_1630)
);

BUFx3_ASAP7_75t_L g1631 ( 
.A(n_1547),
.Y(n_1631)
);

NOR2xp33_ASAP7_75t_L g1632 ( 
.A(n_1524),
.B(n_1540),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1507),
.Y(n_1633)
);

AO21x1_ASAP7_75t_SL g1634 ( 
.A1(n_1612),
.A2(n_1551),
.B(n_1497),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1507),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1580),
.B(n_1490),
.Y(n_1636)
);

OAI21x1_ASAP7_75t_L g1637 ( 
.A1(n_1508),
.A2(n_1584),
.B(n_1581),
.Y(n_1637)
);

OR2x2_ASAP7_75t_L g1638 ( 
.A(n_1538),
.B(n_1536),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1570),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1490),
.B(n_1496),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1570),
.Y(n_1641)
);

OR2x2_ASAP7_75t_L g1642 ( 
.A(n_1538),
.B(n_1497),
.Y(n_1642)
);

INVx3_ASAP7_75t_L g1643 ( 
.A(n_1574),
.Y(n_1643)
);

BUFx2_ASAP7_75t_SL g1644 ( 
.A(n_1569),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1583),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1509),
.B(n_1517),
.Y(n_1646)
);

CKINVDCx5p33_ASAP7_75t_R g1647 ( 
.A(n_1491),
.Y(n_1647)
);

BUFx12f_ASAP7_75t_L g1648 ( 
.A(n_1491),
.Y(n_1648)
);

NOR4xp25_ASAP7_75t_SL g1649 ( 
.A(n_1518),
.B(n_1553),
.C(n_1561),
.D(n_1546),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1532),
.Y(n_1650)
);

OA21x2_ASAP7_75t_L g1651 ( 
.A1(n_1508),
.A2(n_1560),
.B(n_1559),
.Y(n_1651)
);

INVx3_ASAP7_75t_L g1652 ( 
.A(n_1548),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1622),
.B(n_1505),
.Y(n_1653)
);

BUFx3_ASAP7_75t_L g1654 ( 
.A(n_1547),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1537),
.Y(n_1655)
);

AOI221xp5_ASAP7_75t_L g1656 ( 
.A1(n_1589),
.A2(n_1621),
.B1(n_1599),
.B2(n_1626),
.C(n_1615),
.Y(n_1656)
);

BUFx3_ASAP7_75t_L g1657 ( 
.A(n_1547),
.Y(n_1657)
);

BUFx4f_ASAP7_75t_L g1658 ( 
.A(n_1492),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1529),
.Y(n_1659)
);

INVxp67_ASAP7_75t_L g1660 ( 
.A(n_1535),
.Y(n_1660)
);

OAI22xp5_ASAP7_75t_L g1661 ( 
.A1(n_1589),
.A2(n_1599),
.B1(n_1626),
.B2(n_1621),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1528),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1582),
.Y(n_1663)
);

INVx3_ASAP7_75t_L g1664 ( 
.A(n_1578),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1585),
.Y(n_1665)
);

HB1xp67_ASAP7_75t_L g1666 ( 
.A(n_1493),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1578),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1533),
.Y(n_1668)
);

OR2x2_ASAP7_75t_L g1669 ( 
.A(n_1572),
.B(n_1500),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1577),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1576),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1579),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1575),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1563),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1563),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1500),
.B(n_1499),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1588),
.Y(n_1677)
);

OAI21xp5_ASAP7_75t_L g1678 ( 
.A1(n_1615),
.A2(n_1620),
.B(n_1595),
.Y(n_1678)
);

OAI21x1_ASAP7_75t_L g1679 ( 
.A1(n_1573),
.A2(n_1560),
.B(n_1559),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1594),
.Y(n_1680)
);

AOI21xp5_ASAP7_75t_L g1681 ( 
.A1(n_1591),
.A2(n_1486),
.B(n_1551),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1606),
.Y(n_1682)
);

BUFx2_ASAP7_75t_L g1683 ( 
.A(n_1566),
.Y(n_1683)
);

A2O1A1Ixp33_ASAP7_75t_L g1684 ( 
.A1(n_1603),
.A2(n_1620),
.B(n_1586),
.C(n_1628),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1499),
.B(n_1572),
.Y(n_1685)
);

BUFx6f_ASAP7_75t_L g1686 ( 
.A(n_1502),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1614),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1505),
.B(n_1510),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1623),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1545),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1545),
.Y(n_1691)
);

INVx1_ASAP7_75t_SL g1692 ( 
.A(n_1487),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1598),
.Y(n_1693)
);

AOI22xp33_ASAP7_75t_SL g1694 ( 
.A1(n_1525),
.A2(n_1498),
.B1(n_1511),
.B2(n_1629),
.Y(n_1694)
);

OAI21x1_ASAP7_75t_SL g1695 ( 
.A1(n_1489),
.A2(n_1519),
.B(n_1590),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1613),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1522),
.B(n_1510),
.Y(n_1697)
);

HB1xp67_ASAP7_75t_L g1698 ( 
.A(n_1625),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1627),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1567),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1567),
.Y(n_1701)
);

INVx4_ASAP7_75t_L g1702 ( 
.A(n_1569),
.Y(n_1702)
);

AO21x2_ASAP7_75t_L g1703 ( 
.A1(n_1503),
.A2(n_1549),
.B(n_1555),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1549),
.Y(n_1704)
);

INVx3_ASAP7_75t_L g1705 ( 
.A(n_1569),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1522),
.B(n_1605),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1564),
.B(n_1543),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1557),
.Y(n_1708)
);

AO21x1_ASAP7_75t_SL g1709 ( 
.A1(n_1564),
.A2(n_1571),
.B(n_1543),
.Y(n_1709)
);

OAI21x1_ASAP7_75t_L g1710 ( 
.A1(n_1571),
.A2(n_1554),
.B(n_1558),
.Y(n_1710)
);

NOR2xp33_ASAP7_75t_L g1711 ( 
.A(n_1539),
.B(n_1611),
.Y(n_1711)
);

HB1xp67_ASAP7_75t_L g1712 ( 
.A(n_1592),
.Y(n_1712)
);

HB1xp67_ASAP7_75t_L g1713 ( 
.A(n_1619),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1534),
.Y(n_1714)
);

BUFx3_ASAP7_75t_L g1715 ( 
.A(n_1530),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1565),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1565),
.Y(n_1717)
);

INVx1_ASAP7_75t_SL g1718 ( 
.A(n_1617),
.Y(n_1718)
);

AO21x2_ASAP7_75t_L g1719 ( 
.A1(n_1609),
.A2(n_1513),
.B(n_1556),
.Y(n_1719)
);

OR2x2_ASAP7_75t_L g1720 ( 
.A(n_1513),
.B(n_1488),
.Y(n_1720)
);

OAI21x1_ASAP7_75t_L g1721 ( 
.A1(n_1552),
.A2(n_1604),
.B(n_1562),
.Y(n_1721)
);

AOI21x1_ASAP7_75t_L g1722 ( 
.A1(n_1618),
.A2(n_1550),
.B(n_1544),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1526),
.Y(n_1723)
);

HB1xp67_ASAP7_75t_L g1724 ( 
.A(n_1520),
.Y(n_1724)
);

AO221x2_ASAP7_75t_L g1725 ( 
.A1(n_1607),
.A2(n_1616),
.B1(n_1610),
.B2(n_1593),
.C(n_1512),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1568),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1492),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1568),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1568),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1492),
.Y(n_1730)
);

INVxp67_ASAP7_75t_SL g1731 ( 
.A(n_1608),
.Y(n_1731)
);

AND2x4_ASAP7_75t_L g1732 ( 
.A(n_1495),
.B(n_1541),
.Y(n_1732)
);

OAI21x1_ASAP7_75t_L g1733 ( 
.A1(n_1597),
.A2(n_1601),
.B(n_1527),
.Y(n_1733)
);

OAI21x1_ASAP7_75t_L g1734 ( 
.A1(n_1597),
.A2(n_1601),
.B(n_1506),
.Y(n_1734)
);

INVx2_ASAP7_75t_L g1735 ( 
.A(n_1531),
.Y(n_1735)
);

AOI21xp33_ASAP7_75t_L g1736 ( 
.A1(n_1523),
.A2(n_1495),
.B(n_1630),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1531),
.Y(n_1737)
);

HB1xp67_ASAP7_75t_L g1738 ( 
.A(n_1506),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1542),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1542),
.Y(n_1740)
);

BUFx12f_ASAP7_75t_L g1741 ( 
.A(n_1647),
.Y(n_1741)
);

O2A1O1Ixp33_ASAP7_75t_SL g1742 ( 
.A1(n_1661),
.A2(n_1587),
.B(n_1596),
.C(n_1516),
.Y(n_1742)
);

INVx3_ASAP7_75t_L g1743 ( 
.A(n_1722),
.Y(n_1743)
);

HB1xp67_ASAP7_75t_L g1744 ( 
.A(n_1633),
.Y(n_1744)
);

AOI22xp5_ASAP7_75t_L g1745 ( 
.A1(n_1656),
.A2(n_1512),
.B1(n_1521),
.B2(n_1501),
.Y(n_1745)
);

OAI22xp5_ASAP7_75t_L g1746 ( 
.A1(n_1694),
.A2(n_1512),
.B1(n_1611),
.B2(n_1514),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1666),
.B(n_1504),
.Y(n_1747)
);

AO21x1_ASAP7_75t_L g1748 ( 
.A1(n_1681),
.A2(n_1515),
.B(n_1600),
.Y(n_1748)
);

OAI22xp5_ASAP7_75t_L g1749 ( 
.A1(n_1684),
.A2(n_1624),
.B1(n_1600),
.B2(n_1630),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1638),
.B(n_1633),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1646),
.B(n_1494),
.Y(n_1751)
);

AND2x4_ASAP7_75t_L g1752 ( 
.A(n_1715),
.B(n_1602),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1646),
.B(n_1660),
.Y(n_1753)
);

OAI22xp5_ASAP7_75t_L g1754 ( 
.A1(n_1678),
.A2(n_1706),
.B1(n_1704),
.B2(n_1688),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1636),
.B(n_1671),
.Y(n_1755)
);

OA21x2_ASAP7_75t_L g1756 ( 
.A1(n_1637),
.A2(n_1679),
.B(n_1704),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1659),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1635),
.B(n_1653),
.Y(n_1758)
);

AO21x1_ASAP7_75t_L g1759 ( 
.A1(n_1697),
.A2(n_1713),
.B(n_1712),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1642),
.B(n_1650),
.Y(n_1760)
);

A2O1A1Ixp33_ASAP7_75t_L g1761 ( 
.A1(n_1676),
.A2(n_1720),
.B(n_1640),
.C(n_1707),
.Y(n_1761)
);

BUFx3_ASAP7_75t_L g1762 ( 
.A(n_1648),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1671),
.B(n_1672),
.Y(n_1763)
);

A2O1A1Ixp33_ASAP7_75t_L g1764 ( 
.A1(n_1676),
.A2(n_1720),
.B(n_1640),
.C(n_1707),
.Y(n_1764)
);

AOI221xp5_ASAP7_75t_L g1765 ( 
.A1(n_1695),
.A2(n_1691),
.B1(n_1690),
.B2(n_1685),
.C(n_1670),
.Y(n_1765)
);

AOI22xp33_ASAP7_75t_SL g1766 ( 
.A1(n_1695),
.A2(n_1685),
.B1(n_1703),
.B2(n_1719),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1659),
.Y(n_1767)
);

OA21x2_ASAP7_75t_L g1768 ( 
.A1(n_1637),
.A2(n_1710),
.B(n_1701),
.Y(n_1768)
);

A2O1A1Ixp33_ASAP7_75t_L g1769 ( 
.A1(n_1631),
.A2(n_1657),
.B(n_1654),
.C(n_1710),
.Y(n_1769)
);

OAI22xp5_ASAP7_75t_L g1770 ( 
.A1(n_1634),
.A2(n_1669),
.B1(n_1649),
.B2(n_1651),
.Y(n_1770)
);

OR2x6_ASAP7_75t_L g1771 ( 
.A(n_1733),
.B(n_1734),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1650),
.B(n_1655),
.Y(n_1772)
);

OAI22xp5_ASAP7_75t_L g1773 ( 
.A1(n_1634),
.A2(n_1669),
.B1(n_1649),
.B2(n_1651),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1663),
.B(n_1677),
.Y(n_1774)
);

O2A1O1Ixp33_ASAP7_75t_SL g1775 ( 
.A1(n_1724),
.A2(n_1731),
.B(n_1736),
.C(n_1632),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1663),
.B(n_1677),
.Y(n_1776)
);

OA21x2_ASAP7_75t_L g1777 ( 
.A1(n_1700),
.A2(n_1673),
.B(n_1674),
.Y(n_1777)
);

INVxp33_ASAP7_75t_L g1778 ( 
.A(n_1711),
.Y(n_1778)
);

NOR2x1_ASAP7_75t_SL g1779 ( 
.A(n_1644),
.B(n_1709),
.Y(n_1779)
);

O2A1O1Ixp33_ASAP7_75t_SL g1780 ( 
.A1(n_1739),
.A2(n_1740),
.B(n_1738),
.C(n_1725),
.Y(n_1780)
);

O2A1O1Ixp33_ASAP7_75t_L g1781 ( 
.A1(n_1703),
.A2(n_1673),
.B(n_1719),
.C(n_1643),
.Y(n_1781)
);

AND2x4_ASAP7_75t_L g1782 ( 
.A(n_1643),
.B(n_1683),
.Y(n_1782)
);

OR2x2_ASAP7_75t_L g1783 ( 
.A(n_1680),
.B(n_1682),
.Y(n_1783)
);

OA21x2_ASAP7_75t_L g1784 ( 
.A1(n_1675),
.A2(n_1639),
.B(n_1641),
.Y(n_1784)
);

O2A1O1Ixp33_ASAP7_75t_SL g1785 ( 
.A1(n_1725),
.A2(n_1740),
.B(n_1739),
.C(n_1648),
.Y(n_1785)
);

O2A1O1Ixp33_ASAP7_75t_SL g1786 ( 
.A1(n_1725),
.A2(n_1729),
.B(n_1726),
.C(n_1728),
.Y(n_1786)
);

BUFx12f_ASAP7_75t_L g1787 ( 
.A(n_1647),
.Y(n_1787)
);

O2A1O1Ixp33_ASAP7_75t_L g1788 ( 
.A1(n_1703),
.A2(n_1719),
.B(n_1651),
.C(n_1737),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1680),
.B(n_1682),
.Y(n_1789)
);

AOI22xp33_ASAP7_75t_L g1790 ( 
.A1(n_1714),
.A2(n_1725),
.B1(n_1689),
.B2(n_1693),
.Y(n_1790)
);

OAI21x1_ASAP7_75t_L g1791 ( 
.A1(n_1705),
.A2(n_1664),
.B(n_1667),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1692),
.B(n_1718),
.Y(n_1792)
);

INVx3_ASAP7_75t_L g1793 ( 
.A(n_1705),
.Y(n_1793)
);

HB1xp67_ASAP7_75t_L g1794 ( 
.A(n_1665),
.Y(n_1794)
);

NAND3xp33_ASAP7_75t_L g1795 ( 
.A(n_1639),
.B(n_1641),
.C(n_1716),
.Y(n_1795)
);

NAND3xp33_ASAP7_75t_L g1796 ( 
.A(n_1716),
.B(n_1717),
.C(n_1708),
.Y(n_1796)
);

OAI21x1_ASAP7_75t_SL g1797 ( 
.A1(n_1737),
.A2(n_1735),
.B(n_1702),
.Y(n_1797)
);

OAI21xp5_ASAP7_75t_L g1798 ( 
.A1(n_1665),
.A2(n_1721),
.B(n_1717),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1784),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1744),
.Y(n_1800)
);

INVx3_ASAP7_75t_L g1801 ( 
.A(n_1791),
.Y(n_1801)
);

OR2x2_ASAP7_75t_L g1802 ( 
.A(n_1750),
.B(n_1687),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1782),
.B(n_1753),
.Y(n_1803)
);

AOI22xp33_ASAP7_75t_L g1804 ( 
.A1(n_1766),
.A2(n_1693),
.B1(n_1696),
.B2(n_1699),
.Y(n_1804)
);

NOR2xp33_ASAP7_75t_L g1805 ( 
.A(n_1778),
.B(n_1732),
.Y(n_1805)
);

INVx3_ASAP7_75t_L g1806 ( 
.A(n_1793),
.Y(n_1806)
);

INVx3_ASAP7_75t_L g1807 ( 
.A(n_1793),
.Y(n_1807)
);

NOR2x1p5_ASAP7_75t_L g1808 ( 
.A(n_1762),
.B(n_1705),
.Y(n_1808)
);

BUFx2_ASAP7_75t_L g1809 ( 
.A(n_1743),
.Y(n_1809)
);

OR2x2_ASAP7_75t_L g1810 ( 
.A(n_1758),
.B(n_1698),
.Y(n_1810)
);

AND2x2_ASAP7_75t_L g1811 ( 
.A(n_1774),
.B(n_1652),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1794),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1776),
.B(n_1664),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1794),
.B(n_1645),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_SL g1815 ( 
.A(n_1748),
.B(n_1686),
.Y(n_1815)
);

BUFx3_ASAP7_75t_L g1816 ( 
.A(n_1797),
.Y(n_1816)
);

NOR2xp33_ASAP7_75t_L g1817 ( 
.A(n_1752),
.B(n_1741),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1757),
.Y(n_1818)
);

HB1xp67_ASAP7_75t_L g1819 ( 
.A(n_1760),
.Y(n_1819)
);

INVxp67_ASAP7_75t_SL g1820 ( 
.A(n_1788),
.Y(n_1820)
);

HB1xp67_ASAP7_75t_L g1821 ( 
.A(n_1789),
.Y(n_1821)
);

OAI22xp5_ASAP7_75t_L g1822 ( 
.A1(n_1754),
.A2(n_1658),
.B1(n_1732),
.B2(n_1702),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1767),
.Y(n_1823)
);

AOI22xp33_ASAP7_75t_L g1824 ( 
.A1(n_1754),
.A2(n_1727),
.B1(n_1730),
.B2(n_1723),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1772),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1772),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1783),
.Y(n_1827)
);

INVx2_ASAP7_75t_L g1828 ( 
.A(n_1777),
.Y(n_1828)
);

AND2x4_ASAP7_75t_L g1829 ( 
.A(n_1771),
.B(n_1705),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1795),
.Y(n_1830)
);

HB1xp67_ASAP7_75t_L g1831 ( 
.A(n_1796),
.Y(n_1831)
);

AOI22xp33_ASAP7_75t_L g1832 ( 
.A1(n_1765),
.A2(n_1723),
.B1(n_1668),
.B2(n_1662),
.Y(n_1832)
);

INVx2_ASAP7_75t_L g1833 ( 
.A(n_1768),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1800),
.Y(n_1834)
);

OR2x2_ASAP7_75t_L g1835 ( 
.A(n_1830),
.B(n_1756),
.Y(n_1835)
);

INVx3_ASAP7_75t_L g1836 ( 
.A(n_1816),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1800),
.Y(n_1837)
);

OAI21xp5_ASAP7_75t_SL g1838 ( 
.A1(n_1822),
.A2(n_1746),
.B(n_1749),
.Y(n_1838)
);

HB1xp67_ASAP7_75t_L g1839 ( 
.A(n_1830),
.Y(n_1839)
);

HB1xp67_ASAP7_75t_L g1840 ( 
.A(n_1831),
.Y(n_1840)
);

INVx2_ASAP7_75t_L g1841 ( 
.A(n_1799),
.Y(n_1841)
);

NAND4xp25_ASAP7_75t_L g1842 ( 
.A(n_1809),
.B(n_1746),
.C(n_1765),
.D(n_1749),
.Y(n_1842)
);

BUFx2_ASAP7_75t_L g1843 ( 
.A(n_1816),
.Y(n_1843)
);

AOI22xp33_ASAP7_75t_L g1844 ( 
.A1(n_1820),
.A2(n_1770),
.B1(n_1773),
.B2(n_1759),
.Y(n_1844)
);

OR2x6_ASAP7_75t_L g1845 ( 
.A(n_1829),
.B(n_1781),
.Y(n_1845)
);

INVxp67_ASAP7_75t_L g1846 ( 
.A(n_1812),
.Y(n_1846)
);

INVx3_ASAP7_75t_SL g1847 ( 
.A(n_1815),
.Y(n_1847)
);

INVx2_ASAP7_75t_SL g1848 ( 
.A(n_1816),
.Y(n_1848)
);

INVx2_ASAP7_75t_L g1849 ( 
.A(n_1799),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1819),
.B(n_1788),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1811),
.B(n_1768),
.Y(n_1851)
);

AND2x2_ASAP7_75t_L g1852 ( 
.A(n_1813),
.B(n_1755),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1821),
.B(n_1779),
.Y(n_1853)
);

NAND3xp33_ASAP7_75t_SL g1854 ( 
.A(n_1822),
.B(n_1790),
.C(n_1773),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1803),
.B(n_1798),
.Y(n_1855)
);

INVxp67_ASAP7_75t_L g1856 ( 
.A(n_1812),
.Y(n_1856)
);

INVx5_ASAP7_75t_L g1857 ( 
.A(n_1801),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1814),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1825),
.B(n_1826),
.Y(n_1859)
);

AND2x4_ASAP7_75t_L g1860 ( 
.A(n_1829),
.B(n_1798),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1818),
.Y(n_1861)
);

AOI22xp33_ASAP7_75t_SL g1862 ( 
.A1(n_1828),
.A2(n_1770),
.B1(n_1764),
.B2(n_1761),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1825),
.B(n_1769),
.Y(n_1863)
);

NOR3xp33_ASAP7_75t_L g1864 ( 
.A(n_1801),
.B(n_1742),
.C(n_1781),
.Y(n_1864)
);

INVx1_ASAP7_75t_SL g1865 ( 
.A(n_1810),
.Y(n_1865)
);

AOI211xp5_ASAP7_75t_L g1866 ( 
.A1(n_1805),
.A2(n_1742),
.B(n_1780),
.C(n_1786),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_SL g1867 ( 
.A(n_1847),
.B(n_1866),
.Y(n_1867)
);

INVxp67_ASAP7_75t_SL g1868 ( 
.A(n_1840),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1839),
.B(n_1818),
.Y(n_1869)
);

INVx2_ASAP7_75t_L g1870 ( 
.A(n_1841),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1861),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1839),
.B(n_1823),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1861),
.Y(n_1873)
);

AND2x2_ASAP7_75t_L g1874 ( 
.A(n_1851),
.B(n_1801),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1840),
.B(n_1823),
.Y(n_1875)
);

INVx2_ASAP7_75t_L g1876 ( 
.A(n_1841),
.Y(n_1876)
);

INVx2_ASAP7_75t_L g1877 ( 
.A(n_1841),
.Y(n_1877)
);

INVx2_ASAP7_75t_L g1878 ( 
.A(n_1849),
.Y(n_1878)
);

AND2x2_ASAP7_75t_L g1879 ( 
.A(n_1855),
.B(n_1827),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1834),
.Y(n_1880)
);

AND2x2_ASAP7_75t_L g1881 ( 
.A(n_1855),
.B(n_1827),
.Y(n_1881)
);

INVx2_ASAP7_75t_L g1882 ( 
.A(n_1849),
.Y(n_1882)
);

OR2x2_ASAP7_75t_L g1883 ( 
.A(n_1835),
.B(n_1802),
.Y(n_1883)
);

AND2x2_ASAP7_75t_L g1884 ( 
.A(n_1855),
.B(n_1806),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1834),
.Y(n_1885)
);

INVx2_ASAP7_75t_L g1886 ( 
.A(n_1849),
.Y(n_1886)
);

AND2x4_ASAP7_75t_L g1887 ( 
.A(n_1857),
.B(n_1829),
.Y(n_1887)
);

INVxp33_ASAP7_75t_L g1888 ( 
.A(n_1864),
.Y(n_1888)
);

AOI22xp33_ASAP7_75t_L g1889 ( 
.A1(n_1862),
.A2(n_1790),
.B1(n_1832),
.B2(n_1763),
.Y(n_1889)
);

AND2x2_ASAP7_75t_L g1890 ( 
.A(n_1852),
.B(n_1807),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1837),
.Y(n_1891)
);

AND2x4_ASAP7_75t_L g1892 ( 
.A(n_1857),
.B(n_1808),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1837),
.Y(n_1893)
);

OR2x2_ASAP7_75t_L g1894 ( 
.A(n_1835),
.B(n_1810),
.Y(n_1894)
);

AND2x2_ASAP7_75t_L g1895 ( 
.A(n_1852),
.B(n_1807),
.Y(n_1895)
);

AOI22xp33_ASAP7_75t_L g1896 ( 
.A1(n_1862),
.A2(n_1824),
.B1(n_1833),
.B2(n_1804),
.Y(n_1896)
);

INVx1_ASAP7_75t_SL g1897 ( 
.A(n_1847),
.Y(n_1897)
);

AND2x2_ASAP7_75t_L g1898 ( 
.A(n_1897),
.B(n_1847),
.Y(n_1898)
);

AND2x4_ASAP7_75t_L g1899 ( 
.A(n_1892),
.B(n_1864),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1871),
.Y(n_1900)
);

AND2x2_ASAP7_75t_L g1901 ( 
.A(n_1897),
.B(n_1843),
.Y(n_1901)
);

HB1xp67_ASAP7_75t_L g1902 ( 
.A(n_1875),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1871),
.Y(n_1903)
);

OR2x2_ASAP7_75t_L g1904 ( 
.A(n_1894),
.B(n_1865),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1888),
.B(n_1865),
.Y(n_1905)
);

AND2x2_ASAP7_75t_L g1906 ( 
.A(n_1879),
.B(n_1843),
.Y(n_1906)
);

AND2x2_ASAP7_75t_L g1907 ( 
.A(n_1879),
.B(n_1836),
.Y(n_1907)
);

OAI21xp33_ASAP7_75t_SL g1908 ( 
.A1(n_1867),
.A2(n_1842),
.B(n_1848),
.Y(n_1908)
);

OR2x2_ASAP7_75t_L g1909 ( 
.A(n_1894),
.B(n_1858),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1871),
.Y(n_1910)
);

INVx2_ASAP7_75t_L g1911 ( 
.A(n_1870),
.Y(n_1911)
);

OAI21xp33_ASAP7_75t_L g1912 ( 
.A1(n_1888),
.A2(n_1842),
.B(n_1838),
.Y(n_1912)
);

AND2x2_ASAP7_75t_L g1913 ( 
.A(n_1879),
.B(n_1836),
.Y(n_1913)
);

AND2x4_ASAP7_75t_L g1914 ( 
.A(n_1892),
.B(n_1857),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1868),
.B(n_1846),
.Y(n_1915)
);

INVx2_ASAP7_75t_L g1916 ( 
.A(n_1870),
.Y(n_1916)
);

INVx2_ASAP7_75t_L g1917 ( 
.A(n_1870),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1873),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1868),
.B(n_1846),
.Y(n_1919)
);

BUFx2_ASAP7_75t_L g1920 ( 
.A(n_1892),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1873),
.Y(n_1921)
);

INVx2_ASAP7_75t_SL g1922 ( 
.A(n_1894),
.Y(n_1922)
);

AND2x4_ASAP7_75t_L g1923 ( 
.A(n_1892),
.B(n_1857),
.Y(n_1923)
);

AND2x2_ASAP7_75t_L g1924 ( 
.A(n_1879),
.B(n_1836),
.Y(n_1924)
);

HB1xp67_ASAP7_75t_L g1925 ( 
.A(n_1875),
.Y(n_1925)
);

INVx2_ASAP7_75t_L g1926 ( 
.A(n_1870),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1873),
.Y(n_1927)
);

AND2x2_ASAP7_75t_L g1928 ( 
.A(n_1881),
.B(n_1836),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1881),
.B(n_1869),
.Y(n_1929)
);

AND2x2_ASAP7_75t_L g1930 ( 
.A(n_1881),
.B(n_1848),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_L g1931 ( 
.A(n_1881),
.B(n_1859),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1880),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1880),
.Y(n_1933)
);

NOR2xp33_ASAP7_75t_L g1934 ( 
.A(n_1867),
.B(n_1787),
.Y(n_1934)
);

INVx3_ASAP7_75t_L g1935 ( 
.A(n_1892),
.Y(n_1935)
);

AND2x2_ASAP7_75t_L g1936 ( 
.A(n_1884),
.B(n_1848),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1880),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1884),
.B(n_1853),
.Y(n_1938)
);

AND2x4_ASAP7_75t_L g1939 ( 
.A(n_1892),
.B(n_1857),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_L g1940 ( 
.A(n_1869),
.B(n_1856),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1885),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1885),
.Y(n_1942)
);

AND2x2_ASAP7_75t_L g1943 ( 
.A(n_1884),
.B(n_1853),
.Y(n_1943)
);

OAI21xp33_ASAP7_75t_L g1944 ( 
.A1(n_1896),
.A2(n_1838),
.B(n_1844),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1885),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1891),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_L g1947 ( 
.A(n_1872),
.B(n_1856),
.Y(n_1947)
);

AND2x2_ASAP7_75t_L g1948 ( 
.A(n_1884),
.B(n_1853),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1906),
.B(n_1890),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1900),
.Y(n_1950)
);

AND2x2_ASAP7_75t_L g1951 ( 
.A(n_1906),
.B(n_1890),
.Y(n_1951)
);

INVx2_ASAP7_75t_L g1952 ( 
.A(n_1911),
.Y(n_1952)
);

AND2x4_ASAP7_75t_L g1953 ( 
.A(n_1898),
.B(n_1887),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1900),
.Y(n_1954)
);

OAI21xp5_ASAP7_75t_L g1955 ( 
.A1(n_1908),
.A2(n_1889),
.B(n_1896),
.Y(n_1955)
);

AND2x2_ASAP7_75t_L g1956 ( 
.A(n_1898),
.B(n_1890),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1903),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_L g1958 ( 
.A(n_1912),
.B(n_1872),
.Y(n_1958)
);

INVx2_ASAP7_75t_SL g1959 ( 
.A(n_1901),
.Y(n_1959)
);

NOR2xp33_ASAP7_75t_L g1960 ( 
.A(n_1912),
.B(n_1817),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_L g1961 ( 
.A(n_1944),
.B(n_1891),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1944),
.B(n_1891),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1903),
.Y(n_1963)
);

HB1xp67_ASAP7_75t_L g1964 ( 
.A(n_1901),
.Y(n_1964)
);

AND2x2_ASAP7_75t_L g1965 ( 
.A(n_1930),
.B(n_1890),
.Y(n_1965)
);

OR2x2_ASAP7_75t_L g1966 ( 
.A(n_1922),
.B(n_1883),
.Y(n_1966)
);

INVx2_ASAP7_75t_L g1967 ( 
.A(n_1911),
.Y(n_1967)
);

BUFx3_ASAP7_75t_L g1968 ( 
.A(n_1934),
.Y(n_1968)
);

AND2x2_ASAP7_75t_L g1969 ( 
.A(n_1930),
.B(n_1895),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1922),
.B(n_1902),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_L g1971 ( 
.A(n_1925),
.B(n_1893),
.Y(n_1971)
);

AND2x2_ASAP7_75t_L g1972 ( 
.A(n_1899),
.B(n_1895),
.Y(n_1972)
);

OAI21xp33_ASAP7_75t_L g1973 ( 
.A1(n_1908),
.A2(n_1905),
.B(n_1915),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_L g1974 ( 
.A(n_1905),
.B(n_1859),
.Y(n_1974)
);

INVx2_ASAP7_75t_L g1975 ( 
.A(n_1911),
.Y(n_1975)
);

INVx2_ASAP7_75t_L g1976 ( 
.A(n_1916),
.Y(n_1976)
);

INVx2_ASAP7_75t_L g1977 ( 
.A(n_1916),
.Y(n_1977)
);

NOR3xp33_ASAP7_75t_L g1978 ( 
.A(n_1915),
.B(n_1854),
.C(n_1866),
.Y(n_1978)
);

INVx2_ASAP7_75t_SL g1979 ( 
.A(n_1904),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1910),
.Y(n_1980)
);

OR2x2_ASAP7_75t_L g1981 ( 
.A(n_1904),
.B(n_1883),
.Y(n_1981)
);

XNOR2xp5_ASAP7_75t_L g1982 ( 
.A(n_1899),
.B(n_1745),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1910),
.Y(n_1983)
);

NOR2x1_ASAP7_75t_L g1984 ( 
.A(n_1899),
.B(n_1747),
.Y(n_1984)
);

CKINVDCx16_ASAP7_75t_R g1985 ( 
.A(n_1899),
.Y(n_1985)
);

INVx2_ASAP7_75t_L g1986 ( 
.A(n_1916),
.Y(n_1986)
);

INVx2_ASAP7_75t_SL g1987 ( 
.A(n_1920),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1918),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_L g1989 ( 
.A(n_1929),
.B(n_1859),
.Y(n_1989)
);

AOI221xp5_ASAP7_75t_L g1990 ( 
.A1(n_1955),
.A2(n_1889),
.B1(n_1850),
.B2(n_1947),
.C(n_1940),
.Y(n_1990)
);

INVx2_ASAP7_75t_L g1991 ( 
.A(n_1972),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1950),
.Y(n_1992)
);

INVx1_ASAP7_75t_SL g1993 ( 
.A(n_1968),
.Y(n_1993)
);

OAI21xp33_ASAP7_75t_SL g1994 ( 
.A1(n_1955),
.A2(n_1919),
.B(n_1913),
.Y(n_1994)
);

NOR3xp33_ASAP7_75t_L g1995 ( 
.A(n_1973),
.B(n_1920),
.C(n_1935),
.Y(n_1995)
);

AO22x1_ASAP7_75t_L g1996 ( 
.A1(n_1978),
.A2(n_1923),
.B1(n_1939),
.B2(n_1914),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1950),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1954),
.Y(n_1998)
);

AOI22xp5_ASAP7_75t_L g1999 ( 
.A1(n_1973),
.A2(n_1854),
.B1(n_1845),
.B2(n_1850),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1964),
.B(n_1929),
.Y(n_2000)
);

XOR2x2_ASAP7_75t_SL g2001 ( 
.A(n_1961),
.B(n_1919),
.Y(n_2001)
);

AOI21xp5_ASAP7_75t_L g2002 ( 
.A1(n_1961),
.A2(n_1947),
.B(n_1940),
.Y(n_2002)
);

A2O1A1Ixp33_ASAP7_75t_SL g2003 ( 
.A1(n_1958),
.A2(n_1935),
.B(n_1946),
.C(n_1945),
.Y(n_2003)
);

AOI22xp5_ASAP7_75t_L g2004 ( 
.A1(n_1962),
.A2(n_1845),
.B1(n_1863),
.B2(n_1860),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1954),
.Y(n_2005)
);

INVx3_ASAP7_75t_L g2006 ( 
.A(n_1953),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_L g2007 ( 
.A(n_1979),
.B(n_1931),
.Y(n_2007)
);

OA21x2_ASAP7_75t_SL g2008 ( 
.A1(n_1962),
.A2(n_1923),
.B(n_1914),
.Y(n_2008)
);

A2O1A1Ixp33_ASAP7_75t_L g2009 ( 
.A1(n_1958),
.A2(n_1883),
.B(n_1863),
.C(n_1874),
.Y(n_2009)
);

INVx1_ASAP7_75t_SL g2010 ( 
.A(n_1968),
.Y(n_2010)
);

NOR2xp67_ASAP7_75t_SL g2011 ( 
.A(n_1985),
.B(n_1935),
.Y(n_2011)
);

NAND2xp33_ASAP7_75t_SL g2012 ( 
.A(n_1959),
.B(n_1907),
.Y(n_2012)
);

AOI21xp33_ASAP7_75t_SL g2013 ( 
.A1(n_1985),
.A2(n_1923),
.B(n_1914),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1957),
.Y(n_2014)
);

OAI22xp5_ASAP7_75t_L g2015 ( 
.A1(n_1984),
.A2(n_1935),
.B1(n_1948),
.B2(n_1938),
.Y(n_2015)
);

AOI221xp5_ASAP7_75t_L g2016 ( 
.A1(n_1979),
.A2(n_1917),
.B1(n_1926),
.B2(n_1874),
.C(n_1945),
.Y(n_2016)
);

AOI21xp33_ASAP7_75t_L g2017 ( 
.A1(n_1982),
.A2(n_1921),
.B(n_1918),
.Y(n_2017)
);

OAI22xp33_ASAP7_75t_L g2018 ( 
.A1(n_1999),
.A2(n_1845),
.B1(n_1984),
.B2(n_1981),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1992),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_L g2020 ( 
.A(n_1993),
.B(n_1959),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1997),
.Y(n_2021)
);

BUFx2_ASAP7_75t_L g2022 ( 
.A(n_2006),
.Y(n_2022)
);

INVxp33_ASAP7_75t_L g2023 ( 
.A(n_2011),
.Y(n_2023)
);

INVxp67_ASAP7_75t_L g2024 ( 
.A(n_1993),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1998),
.Y(n_2025)
);

OR2x2_ASAP7_75t_L g2026 ( 
.A(n_2010),
.B(n_1970),
.Y(n_2026)
);

OAI21xp5_ASAP7_75t_L g2027 ( 
.A1(n_1994),
.A2(n_1960),
.B(n_1982),
.Y(n_2027)
);

AND2x2_ASAP7_75t_L g2028 ( 
.A(n_2010),
.B(n_1953),
.Y(n_2028)
);

AND2x2_ASAP7_75t_L g2029 ( 
.A(n_2006),
.B(n_1953),
.Y(n_2029)
);

OR2x2_ASAP7_75t_L g2030 ( 
.A(n_2000),
.B(n_1981),
.Y(n_2030)
);

OAI31xp33_ASAP7_75t_L g2031 ( 
.A1(n_2003),
.A2(n_1966),
.A3(n_1970),
.B(n_1967),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_L g2032 ( 
.A(n_1990),
.B(n_2002),
.Y(n_2032)
);

NOR2xp33_ASAP7_75t_L g2033 ( 
.A(n_2017),
.B(n_1968),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_2005),
.Y(n_2034)
);

OR2x2_ASAP7_75t_L g2035 ( 
.A(n_2007),
.B(n_1966),
.Y(n_2035)
);

INVx2_ASAP7_75t_L g2036 ( 
.A(n_2001),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_2014),
.Y(n_2037)
);

OAI21xp5_ASAP7_75t_L g2038 ( 
.A1(n_1995),
.A2(n_1987),
.B(n_1956),
.Y(n_2038)
);

NAND2x1p5_ASAP7_75t_L g2039 ( 
.A(n_1991),
.B(n_1987),
.Y(n_2039)
);

OAI21xp33_ASAP7_75t_SL g2040 ( 
.A1(n_2016),
.A2(n_1972),
.B(n_1956),
.Y(n_2040)
);

NAND2xp5_ASAP7_75t_L g2041 ( 
.A(n_2028),
.B(n_1996),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_2026),
.Y(n_2042)
);

OA22x2_ASAP7_75t_L g2043 ( 
.A1(n_2036),
.A2(n_2004),
.B1(n_2015),
.B2(n_1953),
.Y(n_2043)
);

AO22x2_ASAP7_75t_L g2044 ( 
.A1(n_2036),
.A2(n_2008),
.B1(n_1957),
.B2(n_1980),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_2024),
.Y(n_2045)
);

OAI21xp5_ASAP7_75t_L g2046 ( 
.A1(n_2031),
.A2(n_2009),
.B(n_2013),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_2022),
.Y(n_2047)
);

NOR2x1_ASAP7_75t_L g2048 ( 
.A(n_2033),
.B(n_1963),
.Y(n_2048)
);

INVx2_ASAP7_75t_SL g2049 ( 
.A(n_2028),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_2030),
.Y(n_2050)
);

NAND2xp5_ASAP7_75t_L g2051 ( 
.A(n_2033),
.B(n_1949),
.Y(n_2051)
);

NOR2xp33_ASAP7_75t_SL g2052 ( 
.A(n_2023),
.B(n_2029),
.Y(n_2052)
);

O2A1O1Ixp33_ASAP7_75t_L g2053 ( 
.A1(n_2032),
.A2(n_1971),
.B(n_1967),
.C(n_1952),
.Y(n_2053)
);

OAI21xp5_ASAP7_75t_L g2054 ( 
.A1(n_2027),
.A2(n_2023),
.B(n_2038),
.Y(n_2054)
);

AOI22xp5_ASAP7_75t_L g2055 ( 
.A1(n_2018),
.A2(n_2012),
.B1(n_1967),
.B2(n_1975),
.Y(n_2055)
);

NAND2xp5_ASAP7_75t_L g2056 ( 
.A(n_2049),
.B(n_2030),
.Y(n_2056)
);

NAND2xp33_ASAP7_75t_L g2057 ( 
.A(n_2051),
.B(n_2020),
.Y(n_2057)
);

AND2x2_ASAP7_75t_L g2058 ( 
.A(n_2052),
.B(n_2029),
.Y(n_2058)
);

AND3x2_ASAP7_75t_L g2059 ( 
.A(n_2042),
.B(n_2021),
.C(n_2019),
.Y(n_2059)
);

NOR3xp33_ASAP7_75t_L g2060 ( 
.A(n_2054),
.B(n_2035),
.C(n_2034),
.Y(n_2060)
);

AND2x4_ASAP7_75t_SL g2061 ( 
.A(n_2045),
.B(n_1751),
.Y(n_2061)
);

NOR2xp33_ASAP7_75t_L g2062 ( 
.A(n_2050),
.B(n_2035),
.Y(n_2062)
);

NAND2xp5_ASAP7_75t_SL g2063 ( 
.A(n_2046),
.B(n_2039),
.Y(n_2063)
);

AOI21xp5_ASAP7_75t_L g2064 ( 
.A1(n_2044),
.A2(n_2053),
.B(n_2048),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_2047),
.Y(n_2065)
);

NAND4xp25_ASAP7_75t_L g2066 ( 
.A(n_2041),
.B(n_2037),
.C(n_2025),
.D(n_1971),
.Y(n_2066)
);

NAND4xp25_ASAP7_75t_L g2067 ( 
.A(n_2055),
.B(n_2044),
.C(n_2043),
.D(n_2039),
.Y(n_2067)
);

AOI22xp33_ASAP7_75t_L g2068 ( 
.A1(n_2067),
.A2(n_2064),
.B1(n_2060),
.B2(n_2063),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_2056),
.Y(n_2069)
);

AOI211x1_ASAP7_75t_L g2070 ( 
.A1(n_2058),
.A2(n_1980),
.B(n_1983),
.C(n_1963),
.Y(n_2070)
);

NOR4xp25_ASAP7_75t_L g2071 ( 
.A(n_2065),
.B(n_2040),
.C(n_1975),
.D(n_1976),
.Y(n_2071)
);

AOI221xp5_ASAP7_75t_L g2072 ( 
.A1(n_2062),
.A2(n_1976),
.B1(n_1975),
.B2(n_1986),
.C(n_1952),
.Y(n_2072)
);

NOR3xp33_ASAP7_75t_L g2073 ( 
.A(n_2066),
.B(n_1976),
.C(n_1952),
.Y(n_2073)
);

AOI221xp5_ASAP7_75t_L g2074 ( 
.A1(n_2057),
.A2(n_1986),
.B1(n_1977),
.B2(n_1983),
.C(n_1988),
.Y(n_2074)
);

AOI211xp5_ASAP7_75t_L g2075 ( 
.A1(n_2059),
.A2(n_1785),
.B(n_1988),
.C(n_1923),
.Y(n_2075)
);

NOR3xp33_ASAP7_75t_L g2076 ( 
.A(n_2061),
.B(n_1986),
.C(n_1977),
.Y(n_2076)
);

OAI211xp5_ASAP7_75t_L g2077 ( 
.A1(n_2068),
.A2(n_1974),
.B(n_1951),
.C(n_1949),
.Y(n_2077)
);

OAI211xp5_ASAP7_75t_SL g2078 ( 
.A1(n_2069),
.A2(n_2075),
.B(n_2073),
.C(n_2074),
.Y(n_2078)
);

AOI221xp5_ASAP7_75t_L g2079 ( 
.A1(n_2071),
.A2(n_1977),
.B1(n_1926),
.B2(n_1917),
.C(n_1921),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_2070),
.Y(n_2080)
);

OAI22xp5_ASAP7_75t_L g2081 ( 
.A1(n_2072),
.A2(n_1909),
.B1(n_1989),
.B2(n_1914),
.Y(n_2081)
);

OAI221xp5_ASAP7_75t_L g2082 ( 
.A1(n_2076),
.A2(n_1926),
.B1(n_1917),
.B2(n_1909),
.C(n_1932),
.Y(n_2082)
);

AOI221x1_ASAP7_75t_L g2083 ( 
.A1(n_2069),
.A2(n_1942),
.B1(n_1937),
.B2(n_1941),
.C(n_1927),
.Y(n_2083)
);

A2O1A1Ixp33_ASAP7_75t_SL g2084 ( 
.A1(n_2068),
.A2(n_1937),
.B(n_1927),
.C(n_1941),
.Y(n_2084)
);

AOI222xp33_ASAP7_75t_L g2085 ( 
.A1(n_2068),
.A2(n_1882),
.B1(n_1876),
.B2(n_1878),
.C1(n_1886),
.C2(n_1877),
.Y(n_2085)
);

NOR2xp33_ASAP7_75t_L g2086 ( 
.A(n_2077),
.B(n_1792),
.Y(n_2086)
);

INVx2_ASAP7_75t_L g2087 ( 
.A(n_2080),
.Y(n_2087)
);

NAND2xp5_ASAP7_75t_L g2088 ( 
.A(n_2084),
.B(n_1951),
.Y(n_2088)
);

BUFx2_ASAP7_75t_L g2089 ( 
.A(n_2079),
.Y(n_2089)
);

AOI22xp5_ASAP7_75t_L g2090 ( 
.A1(n_2085),
.A2(n_2078),
.B1(n_2081),
.B2(n_2082),
.Y(n_2090)
);

AND2x4_ASAP7_75t_L g2091 ( 
.A(n_2083),
.B(n_1936),
.Y(n_2091)
);

AND2x4_ASAP7_75t_L g2092 ( 
.A(n_2080),
.B(n_1936),
.Y(n_2092)
);

OR2x2_ASAP7_75t_L g2093 ( 
.A(n_2088),
.B(n_1965),
.Y(n_2093)
);

NAND4xp75_ASAP7_75t_L g2094 ( 
.A(n_2087),
.B(n_1969),
.C(n_1965),
.D(n_1907),
.Y(n_2094)
);

OAI321xp33_ASAP7_75t_L g2095 ( 
.A1(n_2090),
.A2(n_1845),
.A3(n_1946),
.B1(n_1942),
.B2(n_1932),
.C(n_1933),
.Y(n_2095)
);

NOR4xp75_ASAP7_75t_L g2096 ( 
.A(n_2089),
.B(n_1969),
.C(n_1913),
.D(n_1924),
.Y(n_2096)
);

NAND4xp75_ASAP7_75t_L g2097 ( 
.A(n_2086),
.B(n_1928),
.C(n_1924),
.D(n_1948),
.Y(n_2097)
);

BUFx3_ASAP7_75t_L g2098 ( 
.A(n_2093),
.Y(n_2098)
);

INVx2_ASAP7_75t_L g2099 ( 
.A(n_2094),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_2098),
.Y(n_2100)
);

OAI22xp5_ASAP7_75t_L g2101 ( 
.A1(n_2100),
.A2(n_2098),
.B1(n_2092),
.B2(n_2091),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_2100),
.Y(n_2102)
);

AOI22xp5_ASAP7_75t_L g2103 ( 
.A1(n_2101),
.A2(n_2099),
.B1(n_2097),
.B2(n_2095),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_2102),
.Y(n_2104)
);

NAND3xp33_ASAP7_75t_L g2105 ( 
.A(n_2104),
.B(n_2096),
.C(n_1877),
.Y(n_2105)
);

XNOR2xp5_ASAP7_75t_L g2106 ( 
.A(n_2105),
.B(n_2103),
.Y(n_2106)
);

NAND3xp33_ASAP7_75t_L g2107 ( 
.A(n_2106),
.B(n_1933),
.C(n_1877),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_2107),
.Y(n_2108)
);

OAI221xp5_ASAP7_75t_R g2109 ( 
.A1(n_2108),
.A2(n_1939),
.B1(n_1928),
.B2(n_1938),
.C(n_1943),
.Y(n_2109)
);

AOI211xp5_ASAP7_75t_L g2110 ( 
.A1(n_2109),
.A2(n_1775),
.B(n_1780),
.C(n_1786),
.Y(n_2110)
);


endmodule