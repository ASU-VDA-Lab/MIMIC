module real_jpeg_13249_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_216;
wire n_213;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx4_ASAP7_75t_L g84 ( 
.A(n_0),
.Y(n_84)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx4f_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_4),
.A2(n_22),
.B1(n_23),
.B2(n_25),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_4),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_4),
.A2(n_25),
.B1(n_32),
.B2(n_33),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_4),
.A2(n_25),
.B1(n_48),
.B2(n_49),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_4),
.A2(n_25),
.B1(n_43),
.B2(n_45),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_4),
.B(n_30),
.C(n_33),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_4),
.B(n_31),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_4),
.B(n_48),
.C(n_57),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_4),
.B(n_40),
.C(n_45),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_4),
.B(n_204),
.Y(n_203)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_6),
.A2(n_32),
.B1(n_33),
.B2(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_6),
.A2(n_48),
.B1(n_49),
.B2(n_54),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_6),
.A2(n_43),
.B1(n_45),
.B2(n_54),
.Y(n_109)
);

BUFx12_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

BUFx8_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_9),
.A2(n_48),
.B1(n_49),
.B2(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_9),
.A2(n_32),
.B1(n_33),
.B2(n_51),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_9),
.A2(n_43),
.B1(n_45),
.B2(n_51),
.Y(n_86)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

XOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_94),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_SL g12 ( 
.A(n_13),
.B(n_93),
.Y(n_12)
);

INVxp67_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_66),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_15),
.B(n_66),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_63),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_20),
.B1(n_35),
.B2(n_36),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_19),
.A2(n_20),
.B1(n_68),
.B2(n_69),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_19),
.A2(n_79),
.B(n_92),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_19),
.A2(n_20),
.B1(n_81),
.B2(n_92),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_19),
.B(n_112),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_19),
.A2(n_20),
.B1(n_73),
.B2(n_112),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_19),
.A2(n_20),
.B1(n_158),
.B2(n_159),
.Y(n_157)
);

AOI211xp5_ASAP7_75t_SL g168 ( 
.A1(n_19),
.A2(n_110),
.B(n_114),
.C(n_169),
.Y(n_168)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_20),
.B(n_37),
.C(n_64),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_20),
.B(n_73),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_26),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_L g28 ( 
.A1(n_22),
.A2(n_23),
.B1(n_29),
.B2(n_30),
.Y(n_28)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_23),
.B(n_151),
.Y(n_150)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_25),
.B(n_91),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_25),
.B(n_84),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_31),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_31),
.Y(n_27)
);

AO22x1_ASAP7_75t_L g31 ( 
.A1(n_29),
.A2(n_30),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_32),
.A2(n_33),
.B1(n_57),
.B2(n_58),
.Y(n_56)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_33),
.B(n_185),
.Y(n_184)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_37),
.A2(n_52),
.B1(n_61),
.B2(n_62),
.Y(n_36)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_37),
.A2(n_61),
.B1(n_64),
.B2(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_38),
.B(n_50),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_46),
.Y(n_38)
);

NOR2x1_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_47),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_39),
.A2(n_46),
.B1(n_75),
.B2(n_77),
.Y(n_74)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_39),
.Y(n_91)
);

OA21x2_ASAP7_75t_L g110 ( 
.A1(n_39),
.A2(n_46),
.B(n_90),
.Y(n_110)
);

AO22x1_ASAP7_75t_SL g39 ( 
.A1(n_40),
.A2(n_41),
.B1(n_43),
.B2(n_45),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_40),
.A2(n_41),
.B1(n_48),
.B2(n_49),
.Y(n_47)
);

CKINVDCx14_ASAP7_75t_SL g40 ( 
.A(n_41),
.Y(n_40)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx5_ASAP7_75t_SL g45 ( 
.A(n_43),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_43),
.B(n_212),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_45),
.B(n_84),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_48),
.Y(n_49)
);

OA22x2_ASAP7_75t_SL g59 ( 
.A1(n_48),
.A2(n_49),
.B1(n_57),
.B2(n_58),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_48),
.B(n_199),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_55),
.B1(n_59),
.B2(n_60),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_53),
.A2(n_55),
.B1(n_59),
.B2(n_65),
.Y(n_64)
);

AO21x1_ASAP7_75t_L g73 ( 
.A1(n_55),
.A2(n_59),
.B(n_65),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_59),
.Y(n_55)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_57),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_59),
.Y(n_204)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_71),
.C(n_78),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_67),
.A2(n_71),
.B1(n_72),
.B2(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_67),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_72),
.A2(n_73),
.B(n_74),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_73),
.B(n_74),
.Y(n_72)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_73),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_73),
.A2(n_110),
.B1(n_112),
.B2(n_144),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_73),
.B(n_144),
.Y(n_169)
);

A2O1A1Ixp33_ASAP7_75t_L g180 ( 
.A1(n_73),
.A2(n_144),
.B(n_181),
.C(n_186),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_73),
.A2(n_112),
.B1(n_189),
.B2(n_190),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_76),
.A2(n_88),
.B1(n_89),
.B2(n_91),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_97),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_79),
.A2(n_80),
.B1(n_101),
.B2(n_102),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_87),
.Y(n_80)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_81),
.A2(n_87),
.B1(n_92),
.B2(n_124),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_82),
.B(n_86),
.Y(n_81)
);

INVxp33_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_83),
.B(n_129),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_85),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_84),
.A2(n_85),
.B1(n_86),
.B2(n_109),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_84),
.A2(n_85),
.B1(n_109),
.B2(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_87),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_115),
.B(n_236),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_96),
.B(n_99),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_96),
.B(n_99),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_103),
.C(n_105),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_100),
.A2(n_103),
.B1(n_104),
.B2(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_100),
.Y(n_133)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_101),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_105),
.A2(n_106),
.B1(n_131),
.B2(n_132),
.Y(n_130)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_107),
.A2(n_111),
.B(n_113),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_107),
.A2(n_120),
.B1(n_121),
.B2(n_122),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_107),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_110),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_108),
.A2(n_110),
.B1(n_144),
.B2(n_145),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_108),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_110),
.B(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_SL g144 ( 
.A(n_110),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_110),
.A2(n_127),
.B1(n_144),
.B2(n_172),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_110),
.A2(n_144),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_110),
.A2(n_144),
.B1(n_202),
.B2(n_203),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_110),
.A2(n_144),
.B1(n_198),
.B2(n_215),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_110),
.B(n_152),
.C(n_202),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_110),
.B(n_188),
.C(n_192),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_111),
.A2(n_113),
.B(n_126),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_111),
.A2(n_113),
.B(n_148),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_112),
.B(n_152),
.C(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

AO21x1_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_134),
.B(n_235),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_130),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_118),
.B(n_130),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_123),
.C(n_125),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_123),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_120),
.A2(n_121),
.B1(n_126),
.B2(n_141),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_120),
.A2(n_121),
.B1(n_148),
.B2(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_125),
.B(n_137),
.Y(n_136)
);

CKINVDCx14_ASAP7_75t_R g141 ( 
.A(n_126),
.Y(n_141)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_127),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_154),
.B(n_234),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_136),
.B(n_138),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_136),
.B(n_138),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_142),
.C(n_146),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_139),
.A2(n_140),
.B1(n_142),
.B2(n_143),
.Y(n_232)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_144),
.B(n_198),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_146),
.A2(n_147),
.B1(n_231),
.B2(n_232),
.Y(n_230)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_148),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_152),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_149),
.A2(n_150),
.B1(n_152),
.B2(n_153),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_152),
.A2(n_153),
.B1(n_183),
.B2(n_184),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_152),
.A2(n_153),
.B1(n_163),
.B2(n_164),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_152),
.B(n_183),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_152),
.A2(n_153),
.B1(n_201),
.B2(n_205),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_152),
.B(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_152),
.B(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g152 ( 
.A(n_153),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_153),
.B(n_214),
.Y(n_213)
);

O2A1O1Ixp33_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_175),
.B(n_228),
.C(n_233),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_165),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_156),
.B(n_165),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_160),
.C(n_162),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_157),
.B(n_224),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_158),
.A2(n_159),
.B1(n_181),
.B2(n_182),
.Y(n_218)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_160),
.A2(n_161),
.B1(n_162),
.B2(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_162),
.Y(n_225)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_173),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_170),
.B2(n_171),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_167),
.B(n_171),
.C(n_173),
.Y(n_229)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_169),
.Y(n_186)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_222),
.B(n_227),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_194),
.B(n_221),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_187),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_180),
.B(n_187),
.Y(n_221)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_191),
.Y(n_187)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_189),
.Y(n_190)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_195),
.A2(n_217),
.B(n_220),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_196),
.A2(n_206),
.B(n_216),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_200),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_197),
.B(n_200),
.Y(n_216)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_198),
.Y(n_215)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_201),
.Y(n_205)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_213),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_210),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_218),
.B(n_219),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_223),
.B(n_226),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_223),
.B(n_226),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_229),
.B(n_230),
.Y(n_233)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);


endmodule