module fake_jpeg_5977_n_178 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_178);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_178;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_122;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx14_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

INVx6_ASAP7_75t_SL g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_15),
.B(n_1),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_30),
.B(n_31),
.Y(n_46)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_22),
.B(n_1),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_36),
.Y(n_50)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_23),
.Y(n_52)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_36),
.A2(n_27),
.B1(n_25),
.B2(n_18),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_39),
.B(n_42),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_35),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_40),
.B(n_18),
.Y(n_60)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_34),
.A2(n_26),
.B(n_14),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_44),
.A2(n_49),
.B(n_22),
.Y(n_71)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_48),
.Y(n_70)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_38),
.A2(n_26),
.B(n_20),
.Y(n_49)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_52),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_20),
.Y(n_53)
);

NAND3xp33_ASAP7_75t_L g82 ( 
.A(n_53),
.B(n_65),
.C(n_55),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_50),
.B(n_30),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_55),
.A2(n_71),
.B(n_16),
.Y(n_77)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_56),
.B(n_57),
.Y(n_84)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_20),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_58),
.B(n_21),
.C(n_17),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_38),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_59),
.B(n_66),
.Y(n_79)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_46),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_61),
.B(n_63),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_19),
.Y(n_64)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_49),
.B(n_15),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_19),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_22),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_67),
.B(n_69),
.Y(n_90)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_72),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_45),
.B(n_33),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_73),
.Y(n_95)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_74),
.A2(n_48),
.B1(n_47),
.B2(n_41),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_16),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_76),
.B(n_81),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_77),
.B(n_92),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_78),
.B(n_87),
.Y(n_109)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_82),
.A2(n_67),
.B1(n_56),
.B2(n_72),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_71),
.A2(n_36),
.B1(n_24),
.B2(n_27),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_83),
.A2(n_53),
.B1(n_54),
.B2(n_60),
.Y(n_111)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_85),
.Y(n_96)
);

AO22x1_ASAP7_75t_L g86 ( 
.A1(n_65),
.A2(n_33),
.B1(n_37),
.B2(n_31),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_86),
.A2(n_94),
.B1(n_66),
.B2(n_64),
.Y(n_110)
);

NOR3xp33_ASAP7_75t_SL g87 ( 
.A(n_65),
.B(n_37),
.C(n_25),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_69),
.B(n_33),
.C(n_21),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_93),
.B(n_58),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_68),
.A2(n_24),
.B1(n_17),
.B2(n_23),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_97),
.B(n_98),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_91),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_79),
.B(n_59),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_99),
.B(n_100),
.Y(n_121)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_94),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_101),
.B(n_102),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_76),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_93),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_103),
.B(n_111),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_90),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_104),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_86),
.A2(n_54),
.B(n_57),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_105),
.A2(n_108),
.B(n_95),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_77),
.B(n_53),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_110),
.A2(n_92),
.B1(n_88),
.B2(n_89),
.Y(n_116)
);

BUFx24_ASAP7_75t_SL g112 ( 
.A(n_89),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_112),
.B(n_113),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_86),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_114),
.B(n_29),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_116),
.A2(n_129),
.B1(n_111),
.B2(n_104),
.Y(n_135)
);

A2O1A1O1Ixp25_ASAP7_75t_L g119 ( 
.A1(n_105),
.A2(n_87),
.B(n_70),
.C(n_95),
.D(n_29),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_119),
.B(n_110),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_103),
.B(n_74),
.C(n_80),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_120),
.B(n_128),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_107),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_122),
.B(n_123),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_97),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_124),
.A2(n_126),
.B(n_106),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_106),
.B(n_85),
.C(n_81),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_113),
.A2(n_75),
.B1(n_24),
.B2(n_23),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_96),
.B(n_75),
.Y(n_130)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_130),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_117),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_131),
.B(n_120),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_132),
.B(n_143),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_115),
.A2(n_101),
.B1(n_108),
.B2(n_98),
.Y(n_133)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_133),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_121),
.B(n_100),
.Y(n_134)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_134),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_135),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_138),
.A2(n_142),
.B(n_124),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_129),
.B(n_118),
.Y(n_139)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_139),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_128),
.B(n_109),
.Y(n_140)
);

NOR2xp67_ASAP7_75t_SL g152 ( 
.A(n_140),
.B(n_12),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_126),
.A2(n_102),
.B(n_63),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_125),
.Y(n_143)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_146),
.Y(n_154)
);

OAI321xp33_ASAP7_75t_L g149 ( 
.A1(n_142),
.A2(n_124),
.A3(n_119),
.B1(n_116),
.B2(n_127),
.C(n_29),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_149),
.A2(n_151),
.B(n_141),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_152),
.B(n_136),
.C(n_8),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_133),
.B(n_2),
.Y(n_153)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_153),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_148),
.A2(n_138),
.B1(n_137),
.B2(n_132),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_155),
.A2(n_157),
.B1(n_3),
.B2(n_4),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_156),
.B(n_158),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_144),
.A2(n_136),
.B1(n_140),
.B2(n_4),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_150),
.B(n_12),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_160),
.B(n_3),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_151),
.B(n_9),
.C(n_10),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_153),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_162),
.B(n_165),
.Y(n_169)
);

AOI322xp5_ASAP7_75t_L g164 ( 
.A1(n_154),
.A2(n_145),
.A3(n_144),
.B1(n_147),
.B2(n_5),
.C1(n_2),
.C2(n_4),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_164),
.A2(n_167),
.B(n_5),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_166),
.B(n_3),
.Y(n_170)
);

OR2x2_ASAP7_75t_L g167 ( 
.A(n_159),
.B(n_7),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_167),
.A2(n_161),
.B1(n_157),
.B2(n_158),
.Y(n_168)
);

AO21x1_ASAP7_75t_SL g172 ( 
.A1(n_168),
.A2(n_164),
.B(n_163),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_170),
.B(n_171),
.Y(n_173)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_172),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_169),
.B(n_5),
.Y(n_174)
);

BUFx24_ASAP7_75t_SL g175 ( 
.A(n_174),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_176),
.A2(n_173),
.B(n_7),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_175),
.Y(n_178)
);


endmodule