module fake_jpeg_15462_n_319 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_319);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_319;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx8_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx3_ASAP7_75t_SL g65 ( 
.A(n_34),
.Y(n_65)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_23),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_23),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_39),
.B(n_29),
.Y(n_44)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_43),
.A2(n_16),
.B1(n_20),
.B2(n_19),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_47),
.A2(n_51),
.B1(n_28),
.B2(n_23),
.Y(n_68)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_48),
.B(n_52),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_43),
.A2(n_16),
.B1(n_19),
.B2(n_20),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_50),
.A2(n_24),
.B1(n_25),
.B2(n_29),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_42),
.A2(n_16),
.B1(n_20),
.B2(n_19),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_34),
.Y(n_54)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_36),
.B(n_29),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_56),
.B(n_58),
.Y(n_81)
);

AND2x4_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_33),
.Y(n_57)
);

NAND2xp67_ASAP7_75t_L g80 ( 
.A(n_57),
.B(n_33),
.Y(n_80)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVxp33_ASAP7_75t_L g92 ( 
.A(n_60),
.Y(n_92)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_66),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_55),
.A2(n_19),
.B1(n_20),
.B2(n_28),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_67),
.A2(n_86),
.B1(n_88),
.B2(n_65),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_68),
.A2(n_83),
.B1(n_18),
.B2(n_27),
.Y(n_112)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_71),
.Y(n_103)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_73),
.Y(n_109)
);

INVx2_ASAP7_75t_SL g76 ( 
.A(n_57),
.Y(n_76)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_76),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_49),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_77),
.B(n_24),
.Y(n_108)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_80),
.B(n_0),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_58),
.B(n_66),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_60),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_57),
.A2(n_35),
.B1(n_41),
.B2(n_37),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_87),
.B(n_33),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_62),
.A2(n_35),
.B1(n_41),
.B2(n_37),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_55),
.A2(n_25),
.B1(n_24),
.B2(n_27),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_90),
.Y(n_102)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_91),
.Y(n_104)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_93),
.B(n_97),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_76),
.A2(n_62),
.B1(n_63),
.B2(n_51),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_94),
.A2(n_100),
.B1(n_106),
.B2(n_112),
.Y(n_132)
);

OA22x2_ASAP7_75t_L g95 ( 
.A1(n_76),
.A2(n_65),
.B1(n_45),
.B2(n_40),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_95),
.A2(n_116),
.B1(n_74),
.B2(n_91),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_96),
.B(n_99),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_25),
.Y(n_99)
);

AO22x1_ASAP7_75t_SL g100 ( 
.A1(n_87),
.A2(n_65),
.B1(n_40),
.B2(n_64),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_85),
.A2(n_45),
.B1(n_41),
.B2(n_48),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_107),
.A2(n_117),
.B(n_22),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_108),
.B(n_110),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_69),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_84),
.Y(n_113)
);

INVx1_ASAP7_75t_SL g145 ( 
.A(n_113),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_81),
.B(n_40),
.C(n_46),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_115),
.B(n_118),
.C(n_88),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_86),
.A2(n_53),
.B1(n_64),
.B2(n_46),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_70),
.B(n_64),
.C(n_46),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_84),
.Y(n_119)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_119),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_120),
.B(n_121),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_109),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_102),
.Y(n_123)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_123),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_124),
.B(n_130),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_114),
.A2(n_70),
.B(n_22),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_126),
.A2(n_148),
.B(n_18),
.Y(n_155)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_102),
.Y(n_128)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_128),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_129),
.A2(n_31),
.B1(n_32),
.B2(n_21),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_115),
.B(n_73),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_131),
.B(n_135),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_93),
.B(n_68),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_133),
.B(n_146),
.C(n_33),
.Y(n_170)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_98),
.Y(n_134)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_134),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_105),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_117),
.B(n_82),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_136),
.B(n_138),
.Y(n_172)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_103),
.Y(n_137)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_137),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_117),
.B(n_111),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_114),
.A2(n_74),
.B1(n_79),
.B2(n_71),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_140),
.Y(n_156)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_101),
.Y(n_141)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_141),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_106),
.B(n_75),
.Y(n_142)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_142),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_118),
.B(n_103),
.Y(n_143)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_143),
.Y(n_179)
);

AOI22x1_ASAP7_75t_L g144 ( 
.A1(n_95),
.A2(n_92),
.B1(n_72),
.B2(n_84),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_144),
.A2(n_100),
.B1(n_105),
.B2(n_113),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_94),
.B(n_26),
.C(n_30),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_104),
.B(n_90),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_147),
.B(n_101),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_95),
.A2(n_18),
.B(n_27),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_129),
.A2(n_97),
.B1(n_116),
.B2(n_95),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_153),
.A2(n_154),
.B1(n_176),
.B2(n_142),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_127),
.A2(n_100),
.B1(n_72),
.B2(n_78),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_155),
.A2(n_33),
.B(n_17),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_122),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_157),
.B(n_158),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_140),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_144),
.A2(n_135),
.B1(n_145),
.B2(n_137),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_161),
.A2(n_166),
.B1(n_158),
.B2(n_156),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_122),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_162),
.B(n_141),
.Y(n_190)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_134),
.Y(n_165)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_165),
.Y(n_185)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_123),
.Y(n_168)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_168),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_169),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_170),
.B(n_174),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_145),
.B(n_119),
.Y(n_171)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_171),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_133),
.B(n_30),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_173),
.B(n_174),
.C(n_175),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_131),
.B(n_30),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_130),
.B(n_30),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_144),
.A2(n_32),
.B1(n_21),
.B2(n_31),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_177),
.A2(n_120),
.B1(n_128),
.B2(n_121),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_136),
.B(n_33),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_178),
.B(n_124),
.C(n_26),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_157),
.Y(n_180)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_180),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_166),
.B(n_138),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_182),
.A2(n_179),
.B(n_155),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_184),
.A2(n_187),
.B1(n_153),
.B2(n_172),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_163),
.B(n_139),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_186),
.B(n_188),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_149),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_189),
.B(n_191),
.C(n_197),
.Y(n_223)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_190),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_151),
.B(n_125),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_168),
.B(n_125),
.Y(n_192)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_192),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_164),
.B(n_132),
.Y(n_194)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_194),
.Y(n_230)
);

BUFx12f_ASAP7_75t_L g196 ( 
.A(n_162),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_196),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_151),
.B(n_126),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_150),
.A2(n_132),
.B1(n_146),
.B2(n_148),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_198),
.A2(n_203),
.B1(n_200),
.B2(n_187),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_199),
.B(n_204),
.C(n_17),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_200),
.A2(n_152),
.B(n_159),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_202),
.A2(n_176),
.B1(n_154),
.B2(n_178),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_156),
.A2(n_32),
.B1(n_31),
.B2(n_26),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_173),
.B(n_26),
.Y(n_204)
);

BUFx2_ASAP7_75t_L g205 ( 
.A(n_165),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_205),
.Y(n_214)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_160),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_206),
.Y(n_225)
);

OR2x2_ASAP7_75t_L g207 ( 
.A(n_183),
.B(n_167),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_207),
.B(n_196),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_189),
.B(n_170),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_208),
.B(n_211),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_L g241 ( 
.A1(n_210),
.A2(n_212),
.B1(n_193),
.B2(n_185),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_197),
.B(n_175),
.Y(n_211)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_215),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_216),
.A2(n_221),
.B1(n_227),
.B2(n_199),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_181),
.B(n_191),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_217),
.B(n_219),
.C(n_226),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_195),
.B(n_32),
.Y(n_218)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_218),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_181),
.B(n_17),
.Y(n_219)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_220),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_182),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_204),
.B(n_17),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_182),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_201),
.B(n_3),
.Y(n_229)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_229),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_231),
.B(n_196),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_224),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_232),
.B(n_239),
.Y(n_260)
);

OAI22x1_ASAP7_75t_L g235 ( 
.A1(n_207),
.A2(n_184),
.B1(n_198),
.B2(n_203),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_235),
.A2(n_247),
.B1(n_252),
.B2(n_215),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_213),
.B(n_180),
.Y(n_238)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_238),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_222),
.Y(n_239)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_240),
.Y(n_264)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_241),
.Y(n_266)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_222),
.Y(n_242)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_242),
.Y(n_268)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_218),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_244),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_228),
.B(n_205),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_245),
.B(n_250),
.Y(n_255)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_229),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_246),
.B(n_251),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_249),
.B(n_208),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_225),
.B(n_10),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_214),
.B(n_17),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_230),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_248),
.A2(n_235),
.B1(n_234),
.B2(n_242),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_254),
.A2(n_220),
.B1(n_240),
.B2(n_252),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_SL g274 ( 
.A(n_257),
.B(n_259),
.Y(n_274)
);

FAx1_ASAP7_75t_L g258 ( 
.A(n_234),
.B(n_216),
.CI(n_227),
.CON(n_258),
.SN(n_258)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_258),
.B(n_3),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_249),
.B(n_223),
.Y(n_259)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_261),
.Y(n_277)
);

FAx1_ASAP7_75t_SL g263 ( 
.A(n_233),
.B(n_211),
.CI(n_223),
.CON(n_263),
.SN(n_263)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_263),
.B(n_243),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_233),
.B(n_217),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_267),
.C(n_17),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_243),
.B(n_219),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_255),
.B(n_246),
.Y(n_269)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_269),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_270),
.B(n_278),
.C(n_282),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_260),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_271),
.B(n_273),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_264),
.A2(n_237),
.B1(n_244),
.B2(n_236),
.Y(n_272)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_272),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_253),
.B(n_237),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_256),
.A2(n_236),
.B(n_212),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_275),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_276),
.B(n_279),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_266),
.A2(n_209),
.B1(n_231),
.B2(n_221),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_262),
.B(n_226),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_280),
.B(n_281),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_263),
.B(n_10),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_275),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_286),
.B(n_292),
.Y(n_303)
);

OAI21xp33_ASAP7_75t_L g287 ( 
.A1(n_277),
.A2(n_258),
.B(n_268),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_287),
.A2(n_289),
.B(n_274),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_SL g288 ( 
.A(n_274),
.B(n_257),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_288),
.B(n_12),
.C(n_7),
.Y(n_301)
);

A2O1A1Ixp33_ASAP7_75t_L g289 ( 
.A1(n_281),
.A2(n_258),
.B(n_259),
.C(n_267),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_271),
.A2(n_265),
.B(n_7),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_294),
.B(n_282),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_295),
.B(n_296),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_283),
.A2(n_289),
.B(n_287),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_297),
.A2(n_301),
.B(n_302),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_291),
.B(n_11),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_298),
.A2(n_9),
.B(n_13),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_285),
.B(n_11),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_299),
.B(n_300),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_293),
.B(n_12),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_290),
.A2(n_284),
.B(n_286),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_303),
.B(n_8),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_305),
.B(n_306),
.Y(n_313)
);

OAI21x1_ASAP7_75t_SL g306 ( 
.A1(n_303),
.A2(n_288),
.B(n_8),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_308),
.B(n_310),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_299),
.B(n_9),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_309),
.B(n_9),
.C(n_13),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_311),
.B(n_304),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_313),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_315),
.B(n_307),
.C(n_312),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_14),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_15),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_318),
.A2(n_6),
.B1(n_15),
.B2(n_237),
.Y(n_319)
);


endmodule