module fake_aes_5666_n_49 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_14, n_7, n_10, n_8, n_0, n_49);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_14;
input n_7;
input n_10;
input n_8;
input n_0;
output n_49;
wire n_45;
wire n_20;
wire n_38;
wire n_44;
wire n_36;
wire n_47;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_46;
wire n_48;
wire n_30;
wire n_16;
wire n_26;
wire n_25;
wire n_33;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_17;
wire n_15;
wire n_42;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_43;
wire n_40;
wire n_27;
wire n_39;
INVx2_ASAP7_75t_L g15 ( .A(n_5), .Y(n_15) );
CKINVDCx20_ASAP7_75t_R g16 ( .A(n_6), .Y(n_16) );
INVx2_ASAP7_75t_SL g17 ( .A(n_4), .Y(n_17) );
INVx2_ASAP7_75t_L g18 ( .A(n_9), .Y(n_18) );
CKINVDCx5p33_ASAP7_75t_R g19 ( .A(n_3), .Y(n_19) );
BUFx6f_ASAP7_75t_L g20 ( .A(n_3), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_14), .Y(n_21) );
OAI22xp5_ASAP7_75t_SL g22 ( .A1(n_1), .A2(n_13), .B1(n_12), .B2(n_7), .Y(n_22) );
BUFx6f_ASAP7_75t_L g23 ( .A(n_11), .Y(n_23) );
AND2x4_ASAP7_75t_L g24 ( .A(n_17), .B(n_0), .Y(n_24) );
CKINVDCx20_ASAP7_75t_R g25 ( .A(n_16), .Y(n_25) );
HB1xp67_ASAP7_75t_L g26 ( .A(n_19), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_15), .Y(n_27) );
AOI22xp5_ASAP7_75t_L g28 ( .A1(n_16), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_28) );
AOI222xp33_ASAP7_75t_L g29 ( .A1(n_27), .A2(n_22), .B1(n_20), .B2(n_21), .C1(n_18), .C2(n_23), .Y(n_29) );
OAI22xp5_ASAP7_75t_L g30 ( .A1(n_26), .A2(n_20), .B1(n_23), .B2(n_5), .Y(n_30) );
OAI21x1_ASAP7_75t_L g31 ( .A1(n_26), .A2(n_23), .B(n_8), .Y(n_31) );
INVx1_ASAP7_75t_L g32 ( .A(n_30), .Y(n_32) );
INVx2_ASAP7_75t_L g33 ( .A(n_31), .Y(n_33) );
AND2x2_ASAP7_75t_L g34 ( .A(n_32), .B(n_25), .Y(n_34) );
NAND2xp5_ASAP7_75t_L g35 ( .A(n_33), .B(n_29), .Y(n_35) );
INVx1_ASAP7_75t_SL g36 ( .A(n_34), .Y(n_36) );
A2O1A1Ixp33_ASAP7_75t_L g37 ( .A1(n_35), .A2(n_31), .B(n_24), .C(n_33), .Y(n_37) );
OR2x2_ASAP7_75t_L g38 ( .A(n_34), .B(n_28), .Y(n_38) );
NOR2xp33_ASAP7_75t_L g39 ( .A(n_38), .B(n_24), .Y(n_39) );
NOR2x1p5_ASAP7_75t_L g40 ( .A(n_36), .B(n_20), .Y(n_40) );
AOI21xp5_ASAP7_75t_L g41 ( .A1(n_37), .A2(n_23), .B(n_20), .Y(n_41) );
INVx1_ASAP7_75t_L g42 ( .A(n_40), .Y(n_42) );
AND2x4_ASAP7_75t_L g43 ( .A(n_41), .B(n_2), .Y(n_43) );
NAND2x1p5_ASAP7_75t_L g44 ( .A(n_39), .B(n_4), .Y(n_44) );
INVx1_ASAP7_75t_L g45 ( .A(n_42), .Y(n_45) );
INVx2_ASAP7_75t_L g46 ( .A(n_43), .Y(n_46) );
BUFx2_ASAP7_75t_L g47 ( .A(n_42), .Y(n_47) );
OAI22xp33_ASAP7_75t_L g48 ( .A1(n_46), .A2(n_44), .B1(n_43), .B2(n_10), .Y(n_48) );
AOI22xp5_ASAP7_75t_SL g49 ( .A1(n_48), .A2(n_46), .B1(n_47), .B2(n_45), .Y(n_49) );
endmodule