module fake_jpeg_8486_n_79 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_79);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_79;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

BUFx12f_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_4),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx4f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_0),
.B(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_16),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_22),
.A2(n_25),
.B1(n_14),
.B2(n_11),
.Y(n_35)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_24),
.Y(n_29)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_11),
.A2(n_0),
.B1(n_4),
.B2(n_5),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_26),
.B(n_15),
.Y(n_30)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_10),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_37),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_12),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_36),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_35),
.A2(n_18),
.B1(n_21),
.B2(n_19),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_23),
.B(n_20),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_22),
.B(n_26),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_35),
.A2(n_24),
.B1(n_27),
.B2(n_14),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_38),
.A2(n_40),
.B1(n_42),
.B2(n_46),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_37),
.A2(n_25),
.B1(n_24),
.B2(n_27),
.Y(n_40)
);

NAND2xp33_ASAP7_75t_SL g41 ( 
.A(n_32),
.B(n_24),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_43),
.Y(n_51)
);

MAJx2_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_28),
.C(n_10),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_28),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_15),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_31),
.A2(n_28),
.B1(n_13),
.B2(n_19),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_31),
.A2(n_15),
.B1(n_10),
.B2(n_4),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_48),
.Y(n_55)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_33),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_50),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_53),
.Y(n_61)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_54),
.A2(n_48),
.B1(n_43),
.B2(n_50),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_47),
.Y(n_56)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_56),
.Y(n_59)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_58),
.A2(n_39),
.B1(n_46),
.B2(n_42),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_60),
.A2(n_54),
.B1(n_53),
.B2(n_55),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_62),
.A2(n_63),
.B(n_52),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_39),
.C(n_49),
.Y(n_63)
);

BUFx12_ASAP7_75t_L g65 ( 
.A(n_64),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_65),
.A2(n_67),
.B1(n_68),
.B2(n_61),
.Y(n_70)
);

A2O1A1O1Ixp25_ASAP7_75t_L g71 ( 
.A1(n_66),
.A2(n_63),
.B(n_59),
.C(n_64),
.D(n_9),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_61),
.A2(n_51),
.B(n_44),
.Y(n_68)
);

AO22x1_ASAP7_75t_SL g69 ( 
.A1(n_67),
.A2(n_59),
.B1(n_60),
.B2(n_62),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_69),
.A2(n_59),
.B(n_65),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_70),
.B(n_71),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_69),
.B(n_63),
.C(n_65),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_73),
.B(n_6),
.C(n_7),
.Y(n_76)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_74),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_72),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_77),
.A2(n_75),
.B(n_8),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_78),
.B(n_6),
.Y(n_79)
);


endmodule