module fake_ibex_1969_n_214 (n_7, n_20, n_40, n_17, n_25, n_36, n_41, n_43, n_18, n_3, n_22, n_28, n_32, n_39, n_4, n_33, n_5, n_11, n_30, n_6, n_29, n_13, n_2, n_8, n_26, n_35, n_14, n_0, n_9, n_34, n_12, n_38, n_42, n_15, n_37, n_24, n_31, n_44, n_10, n_23, n_21, n_27, n_45, n_19, n_16, n_1, n_214);

input n_7;
input n_20;
input n_40;
input n_17;
input n_25;
input n_36;
input n_41;
input n_43;
input n_18;
input n_3;
input n_22;
input n_28;
input n_32;
input n_39;
input n_4;
input n_33;
input n_5;
input n_11;
input n_30;
input n_6;
input n_29;
input n_13;
input n_2;
input n_8;
input n_26;
input n_35;
input n_14;
input n_0;
input n_9;
input n_34;
input n_12;
input n_38;
input n_42;
input n_15;
input n_37;
input n_24;
input n_31;
input n_44;
input n_10;
input n_23;
input n_21;
input n_27;
input n_45;
input n_19;
input n_16;
input n_1;

output n_214;

wire n_151;
wire n_147;
wire n_85;
wire n_167;
wire n_128;
wire n_208;
wire n_84;
wire n_64;
wire n_73;
wire n_152;
wire n_171;
wire n_145;
wire n_65;
wire n_103;
wire n_95;
wire n_205;
wire n_204;
wire n_139;
wire n_55;
wire n_130;
wire n_63;
wire n_98;
wire n_129;
wire n_161;
wire n_143;
wire n_106;
wire n_177;
wire n_203;
wire n_148;
wire n_76;
wire n_118;
wire n_183;
wire n_67;
wire n_209;
wire n_164;
wire n_198;
wire n_124;
wire n_110;
wire n_193;
wire n_47;
wire n_169;
wire n_108;
wire n_82;
wire n_165;
wire n_78;
wire n_60;
wire n_86;
wire n_70;
wire n_87;
wire n_69;
wire n_75;
wire n_109;
wire n_121;
wire n_127;
wire n_175;
wire n_137;
wire n_48;
wire n_57;
wire n_59;
wire n_125;
wire n_191;
wire n_178;
wire n_62;
wire n_71;
wire n_153;
wire n_173;
wire n_120;
wire n_93;
wire n_168;
wire n_155;
wire n_162;
wire n_180;
wire n_194;
wire n_122;
wire n_116;
wire n_61;
wire n_201;
wire n_94;
wire n_134;
wire n_77;
wire n_112;
wire n_150;
wire n_88;
wire n_133;
wire n_142;
wire n_51;
wire n_46;
wire n_80;
wire n_172;
wire n_49;
wire n_66;
wire n_90;
wire n_74;
wire n_176;
wire n_58;
wire n_192;
wire n_140;
wire n_136;
wire n_119;
wire n_100;
wire n_179;
wire n_72;
wire n_206;
wire n_166;
wire n_195;
wire n_163;
wire n_212;
wire n_188;
wire n_200;
wire n_114;
wire n_199;
wire n_97;
wire n_102;
wire n_197;
wire n_181;
wire n_131;
wire n_123;
wire n_52;
wire n_189;
wire n_99;
wire n_156;
wire n_105;
wire n_135;
wire n_126;
wire n_187;
wire n_154;
wire n_182;
wire n_111;
wire n_196;
wire n_104;
wire n_141;
wire n_89;
wire n_83;
wire n_53;
wire n_107;
wire n_115;
wire n_149;
wire n_54;
wire n_186;
wire n_50;
wire n_92;
wire n_144;
wire n_170;
wire n_213;
wire n_101;
wire n_190;
wire n_113;
wire n_138;
wire n_96;
wire n_185;
wire n_68;
wire n_117;
wire n_79;
wire n_81;
wire n_159;
wire n_202;
wire n_158;
wire n_211;
wire n_132;
wire n_174;
wire n_210;
wire n_157;
wire n_160;
wire n_184;
wire n_56;
wire n_146;
wire n_91;
wire n_207;

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_21),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_17),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

CKINVDCx5p33_ASAP7_75t_R g50 ( 
.A(n_38),
.Y(n_50)
);

CKINVDCx5p33_ASAP7_75t_R g51 ( 
.A(n_9),
.Y(n_51)
);

CKINVDCx5p33_ASAP7_75t_R g52 ( 
.A(n_3),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_1),
.Y(n_53)
);

NOR2xp67_ASAP7_75t_L g54 ( 
.A(n_35),
.B(n_36),
.Y(n_54)
);

CKINVDCx5p33_ASAP7_75t_R g55 ( 
.A(n_7),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_8),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_14),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_34),
.Y(n_60)
);

CKINVDCx5p33_ASAP7_75t_R g61 ( 
.A(n_7),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_12),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_16),
.Y(n_63)
);

INVxp67_ASAP7_75t_SL g64 ( 
.A(n_5),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_6),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

INVxp67_ASAP7_75t_SL g67 ( 
.A(n_5),
.Y(n_67)
);

CKINVDCx5p33_ASAP7_75t_R g68 ( 
.A(n_11),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_33),
.Y(n_70)
);

NOR2xp67_ASAP7_75t_L g71 ( 
.A(n_9),
.B(n_27),
.Y(n_71)
);

CKINVDCx5p33_ASAP7_75t_R g72 ( 
.A(n_32),
.Y(n_72)
);

INVxp33_ASAP7_75t_SL g73 ( 
.A(n_30),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_42),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_19),
.Y(n_76)
);

CKINVDCx5p33_ASAP7_75t_R g77 ( 
.A(n_26),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_6),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_15),
.Y(n_80)
);

CKINVDCx5p33_ASAP7_75t_R g81 ( 
.A(n_10),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_23),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_37),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_1),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_29),
.Y(n_85)
);

INVxp33_ASAP7_75t_SL g86 ( 
.A(n_13),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

CKINVDCx5p33_ASAP7_75t_R g88 ( 
.A(n_0),
.Y(n_88)
);

CKINVDCx5p33_ASAP7_75t_R g89 ( 
.A(n_22),
.Y(n_89)
);

CKINVDCx5p33_ASAP7_75t_R g90 ( 
.A(n_3),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_49),
.B(n_79),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_57),
.B(n_0),
.Y(n_93)
);

AND2x2_ASAP7_75t_SL g94 ( 
.A(n_46),
.B(n_2),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_2),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_60),
.B(n_4),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_58),
.B(n_4),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_59),
.B(n_20),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_66),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_L g101 ( 
.A1(n_65),
.A2(n_40),
.B1(n_41),
.B2(n_67),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_75),
.B(n_78),
.Y(n_103)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_80),
.B(n_82),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_85),
.B(n_87),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_64),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_53),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_70),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_52),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_86),
.A2(n_73),
.B1(n_88),
.B2(n_90),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_50),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_55),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_61),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_68),
.B(n_72),
.Y(n_116)
);

AND2x6_ASAP7_75t_L g117 ( 
.A(n_54),
.B(n_89),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_65),
.B(n_81),
.Y(n_118)
);

OR2x6_ASAP7_75t_L g119 ( 
.A(n_71),
.B(n_48),
.Y(n_119)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_77),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_48),
.Y(n_121)
);

OR2x6_ASAP7_75t_L g122 ( 
.A(n_62),
.B(n_63),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_62),
.B(n_63),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_83),
.A2(n_57),
.B1(n_65),
.B2(n_76),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_74),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_74),
.Y(n_126)
);

AND2x6_ASAP7_75t_L g127 ( 
.A(n_76),
.B(n_83),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_57),
.B(n_56),
.Y(n_128)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_46),
.Y(n_129)
);

AND2x6_ASAP7_75t_L g130 ( 
.A(n_47),
.B(n_58),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_57),
.A2(n_65),
.B1(n_48),
.B2(n_74),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_47),
.Y(n_132)
);

OAI21x1_ASAP7_75t_L g133 ( 
.A1(n_99),
.A2(n_107),
.B(n_98),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_107),
.A2(n_111),
.B(n_114),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_103),
.A2(n_106),
.B(n_91),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_115),
.A2(n_109),
.B(n_92),
.Y(n_136)
);

OAI321xp33_ASAP7_75t_L g137 ( 
.A1(n_96),
.A2(n_98),
.A3(n_108),
.B1(n_92),
.B2(n_101),
.C(n_110),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_129),
.B(n_116),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_109),
.A2(n_100),
.B(n_102),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_109),
.A2(n_95),
.B(n_132),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_129),
.B(n_128),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_130),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_112),
.A2(n_105),
.B1(n_119),
.B2(n_125),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_130),
.A2(n_117),
.B(n_96),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_129),
.B(n_120),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_129),
.A2(n_104),
.B(n_97),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_97),
.A2(n_112),
.B(n_113),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_105),
.A2(n_119),
.B1(n_121),
.B2(n_124),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_118),
.B(n_122),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_120),
.B(n_117),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_113),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_113),
.A2(n_101),
.B(n_93),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_117),
.B(n_130),
.Y(n_153)
);

O2A1O1Ixp5_ASAP7_75t_L g154 ( 
.A1(n_130),
.A2(n_117),
.B(n_126),
.C(n_123),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_94),
.B(n_119),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_124),
.A2(n_131),
.B1(n_122),
.B2(n_127),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_131),
.B(n_122),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_127),
.B(n_110),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_127),
.B(n_110),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_127),
.B(n_128),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_104),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_128),
.B(n_104),
.Y(n_162)
);

AND3x2_ASAP7_75t_L g163 ( 
.A(n_118),
.B(n_128),
.C(n_126),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_109),
.B(n_107),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_91),
.B(n_110),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_109),
.B(n_107),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_162),
.B(n_161),
.Y(n_167)
);

NOR3xp33_ASAP7_75t_L g168 ( 
.A(n_156),
.B(n_148),
.C(n_157),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_143),
.B(n_157),
.Y(n_169)
);

AND2x4_ASAP7_75t_L g170 ( 
.A(n_147),
.B(n_166),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_142),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_165),
.B(n_141),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_134),
.B(n_135),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_144),
.A2(n_153),
.B(n_136),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_149),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_164),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_165),
.B(n_166),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_164),
.A2(n_146),
.B(n_150),
.Y(n_178)
);

INVx3_ASAP7_75t_SL g179 ( 
.A(n_160),
.Y(n_179)
);

NAND2x1p5_ASAP7_75t_L g180 ( 
.A(n_133),
.B(n_142),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_140),
.B(n_152),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_155),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_158),
.A2(n_159),
.B1(n_139),
.B2(n_133),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_138),
.A2(n_137),
.B1(n_145),
.B2(n_151),
.Y(n_184)
);

OR2x2_ASAP7_75t_SL g185 ( 
.A(n_163),
.B(n_154),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_173),
.Y(n_186)
);

OAI21x1_ASAP7_75t_L g187 ( 
.A1(n_180),
.A2(n_142),
.B(n_174),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_172),
.B(n_142),
.Y(n_188)
);

NAND3xp33_ASAP7_75t_L g189 ( 
.A(n_168),
.B(n_169),
.C(n_184),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_170),
.Y(n_190)
);

AND2x6_ASAP7_75t_L g191 ( 
.A(n_170),
.B(n_171),
.Y(n_191)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_170),
.Y(n_192)
);

AO21x2_ASAP7_75t_L g193 ( 
.A1(n_178),
.A2(n_181),
.B(n_177),
.Y(n_193)
);

AO21x2_ASAP7_75t_L g194 ( 
.A1(n_176),
.A2(n_172),
.B(n_185),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_171),
.Y(n_195)
);

OAI221xp5_ASAP7_75t_L g196 ( 
.A1(n_190),
.A2(n_175),
.B1(n_167),
.B2(n_182),
.C(n_179),
.Y(n_196)
);

AND2x2_ASAP7_75t_SL g197 ( 
.A(n_188),
.B(n_167),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_189),
.A2(n_175),
.B1(n_182),
.B2(n_179),
.Y(n_198)
);

OAI221xp5_ASAP7_75t_L g199 ( 
.A1(n_190),
.A2(n_180),
.B1(n_183),
.B2(n_185),
.C(n_192),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_188),
.B(n_189),
.Y(n_200)
);

NAND3xp33_ASAP7_75t_L g201 ( 
.A(n_186),
.B(n_180),
.C(n_188),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_192),
.B(n_186),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_192),
.B(n_194),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_192),
.B(n_194),
.Y(n_204)
);

NOR2x1p5_ASAP7_75t_SL g205 ( 
.A(n_199),
.B(n_195),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_205),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_206),
.B(n_204),
.Y(n_207)
);

NOR2x1_ASAP7_75t_L g208 ( 
.A(n_207),
.B(n_201),
.Y(n_208)
);

NOR2x1_ASAP7_75t_L g209 ( 
.A(n_208),
.B(n_203),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_209),
.B(n_198),
.Y(n_210)
);

AOI221xp5_ASAP7_75t_L g211 ( 
.A1(n_210),
.A2(n_196),
.B1(n_203),
.B2(n_200),
.C(n_192),
.Y(n_211)
);

OAI21x1_ASAP7_75t_L g212 ( 
.A1(n_211),
.A2(n_187),
.B(n_202),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_212),
.Y(n_213)
);

OAI221xp5_ASAP7_75t_R g214 ( 
.A1(n_213),
.A2(n_197),
.B1(n_194),
.B2(n_191),
.C(n_193),
.Y(n_214)
);


endmodule