module real_jpeg_30430_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_705, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_705;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_661;
wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_663;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_648;
wire n_541;
wire n_441;
wire n_696;
wire n_657;
wire n_643;
wire n_656;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_669;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_679;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_640;
wire n_666;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_685;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_680;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_678;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_578;
wire n_456;
wire n_620;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_668;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_605;
wire n_483;
wire n_367;
wire n_639;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_682;
wire n_317;
wire n_658;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_674;
wire n_252;
wire n_601;
wire n_655;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_611;
wire n_104;
wire n_153;
wire n_634;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_684;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_646;
wire n_214;
wire n_671;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_631;
wire n_673;
wire n_175;
wire n_338;
wire n_653;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_650;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_219;
wire n_372;
wire n_122;
wire n_262;
wire n_652;
wire n_334;
wire n_647;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_703;
wire n_110;
wire n_195;
wire n_533;
wire n_592;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_651;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_689;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_615;
wire n_212;
wire n_697;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_672;
wire n_59;
wire n_452;
wire n_213;
wire n_670;
wire n_511;
wire n_524;
wire n_589;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_644;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_693;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_692;
wire n_49;
wire n_514;
wire n_68;
wire n_638;
wire n_497;
wire n_633;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_596;
wire n_312;
wire n_617;
wire n_325;
wire n_307;
wire n_316;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_604;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_688;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_572;
wire n_586;
wire n_548;
wire n_319;
wire n_664;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_637;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_698;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_635;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_642;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_654;
wire n_377;
wire n_616;
wire n_109;
wire n_503;
wire n_686;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_699;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_667;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_683;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_537;
wire n_318;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_691;
wire n_458;
wire n_677;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_701;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_675;
wire n_695;
wire n_138;
wire n_662;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_649;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_702;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_681;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_636;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_597;
wire n_618;
wire n_609;
wire n_700;
wire n_94;
wire n_645;
wire n_687;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_694;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_641;
wire n_225;
wire n_43;
wire n_438;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_690;
wire n_24;
wire n_92;
wire n_676;
wire n_187;
wire n_436;
wire n_629;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_659;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_660;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_625;
wire n_96;
wire n_665;
wire n_308;
wire n_433;
wire n_364;

BUFx12f_ASAP7_75t_L g208 ( 
.A(n_0),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_0),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_0),
.Y(n_279)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_0),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_0),
.Y(n_585)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_1),
.A2(n_243),
.B1(n_244),
.B2(n_246),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_1),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_1),
.A2(n_243),
.B1(n_419),
.B2(n_421),
.Y(n_418)
);

AOI22xp33_ASAP7_75t_SL g532 ( 
.A1(n_1),
.A2(n_243),
.B1(n_533),
.B2(n_537),
.Y(n_532)
);

AOI22xp33_ASAP7_75t_SL g570 ( 
.A1(n_1),
.A2(n_243),
.B1(n_571),
.B2(n_573),
.Y(n_570)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_2),
.A2(n_57),
.B1(n_63),
.B2(n_64),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_2),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_2),
.A2(n_63),
.B1(n_232),
.B2(n_239),
.Y(n_238)
);

OAI22xp33_ASAP7_75t_SL g317 ( 
.A1(n_2),
.A2(n_63),
.B1(n_142),
.B2(n_318),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_L g393 ( 
.A1(n_2),
.A2(n_63),
.B1(n_394),
.B2(n_397),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_4),
.A2(n_44),
.B1(n_49),
.B2(n_50),
.Y(n_43)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_4),
.A2(n_49),
.B1(n_211),
.B2(n_215),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_4),
.A2(n_49),
.B1(n_287),
.B2(n_290),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_4),
.A2(n_49),
.B1(n_335),
.B2(n_336),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g703 ( 
.A(n_5),
.Y(n_703)
);

OAI22x1_ASAP7_75t_SL g263 ( 
.A1(n_6),
.A2(n_264),
.B1(n_267),
.B2(n_268),
.Y(n_263)
);

INVx2_ASAP7_75t_SL g267 ( 
.A(n_6),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_6),
.A2(n_51),
.B1(n_267),
.B2(n_312),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_6),
.A2(n_267),
.B1(n_438),
.B2(n_440),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_6),
.A2(n_267),
.B1(n_495),
.B2(n_497),
.Y(n_494)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_7),
.Y(n_73)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_8),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_8),
.Y(n_136)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_9),
.Y(n_90)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_9),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_9),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_9),
.Y(n_283)
);

AO22x1_ASAP7_75t_L g162 ( 
.A1(n_10),
.A2(n_163),
.B1(n_167),
.B2(n_168),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_10),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_10),
.A2(n_167),
.B1(n_175),
.B2(n_178),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_10),
.A2(n_167),
.B1(n_221),
.B2(n_223),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_10),
.A2(n_167),
.B1(n_293),
.B2(n_295),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_11),
.A2(n_226),
.B1(n_231),
.B2(n_232),
.Y(n_225)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_11),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_11),
.A2(n_231),
.B1(n_257),
.B2(n_260),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_11),
.A2(n_187),
.B1(n_231),
.B2(n_347),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_11),
.A2(n_231),
.B1(n_463),
.B2(n_466),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_12),
.B(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_12),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_12),
.B(n_29),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_12),
.B(n_501),
.Y(n_500)
);

AOI22xp33_ASAP7_75t_SL g523 ( 
.A1(n_12),
.A2(n_432),
.B1(n_524),
.B2(n_527),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_12),
.B(n_125),
.Y(n_549)
);

OAI21xp33_ASAP7_75t_L g579 ( 
.A1(n_12),
.A2(n_202),
.B(n_559),
.Y(n_579)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_13),
.Y(n_94)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_13),
.Y(n_98)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_14),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_14),
.B(n_703),
.Y(n_702)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_15),
.A2(n_114),
.B1(n_120),
.B2(n_121),
.Y(n_113)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_15),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_15),
.A2(n_120),
.B1(n_141),
.B2(n_146),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_15),
.A2(n_120),
.B1(n_186),
.B2(n_190),
.Y(n_185)
);

AO22x1_ASAP7_75t_SL g280 ( 
.A1(n_15),
.A2(n_120),
.B1(n_281),
.B2(n_284),
.Y(n_280)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_16),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_16),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_16),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_16),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_17),
.A2(n_178),
.B1(n_249),
.B2(n_250),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_17),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_17),
.A2(n_249),
.B1(n_363),
.B2(n_365),
.Y(n_362)
);

AOI22xp33_ASAP7_75t_SL g483 ( 
.A1(n_17),
.A2(n_249),
.B1(n_484),
.B2(n_488),
.Y(n_483)
);

AOI22xp33_ASAP7_75t_SL g551 ( 
.A1(n_17),
.A2(n_249),
.B1(n_552),
.B2(n_557),
.Y(n_551)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_18),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_18),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_700),
.B(n_702),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_193),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_192),
.Y(n_21)
);

OR2x2_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_184),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_23),
.B(n_184),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_172),
.C(n_182),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g688 ( 
.A(n_24),
.B(n_689),
.Y(n_688)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_82),
.C(n_124),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

XNOR2x1_ASAP7_75t_L g678 ( 
.A(n_26),
.B(n_679),
.Y(n_678)
);

OA22x2_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_43),
.B1(n_55),
.B2(n_66),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_28),
.A2(n_67),
.B1(n_173),
.B2(n_174),
.Y(n_172)
);

AOI22x1_ASAP7_75t_L g184 ( 
.A1(n_28),
.A2(n_67),
.B1(n_174),
.B2(n_185),
.Y(n_184)
);

AO22x2_ASAP7_75t_L g662 ( 
.A1(n_28),
.A2(n_56),
.B1(n_68),
.B2(n_346),
.Y(n_662)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

AO22x1_ASAP7_75t_SL g241 ( 
.A1(n_29),
.A2(n_68),
.B1(n_242),
.B2(n_248),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_29),
.B(n_311),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_29),
.B(n_346),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_29),
.B(n_242),
.Y(n_360)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_30),
.B(n_69),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_34),
.B1(n_38),
.B2(n_41),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_33),
.Y(n_76)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_33),
.Y(n_81)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_33),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_33),
.Y(n_387)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_36),
.Y(n_320)
);

INVx2_ASAP7_75t_SL g424 ( 
.A(n_36),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_37),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_37),
.Y(n_271)
);

BUFx5_ASAP7_75t_L g384 ( 
.A(n_37),
.Y(n_384)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_40),
.Y(n_526)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_43),
.Y(n_173)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_45),
.Y(n_380)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_47),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_48),
.Y(n_181)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_54),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_54),
.Y(n_247)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_54),
.Y(n_350)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_68),
.B(n_248),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_68),
.B(n_311),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_68),
.B(n_427),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_74),
.B1(n_77),
.B2(n_79),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_73),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_73),
.Y(n_191)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_78),
.Y(n_314)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

XOR2x2_ASAP7_75t_L g658 ( 
.A(n_83),
.B(n_659),
.Y(n_658)
);

MAJIxp5_ASAP7_75t_L g675 ( 
.A(n_83),
.B(n_659),
.C(n_661),
.Y(n_675)
);

XNOR2xp5_ASAP7_75t_L g679 ( 
.A(n_83),
.B(n_124),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_113),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_103),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_85),
.A2(n_103),
.B1(n_225),
.B2(n_238),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_85),
.A2(n_103),
.B1(n_286),
.B2(n_292),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_85),
.A2(n_103),
.B1(n_238),
.B2(n_286),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_85),
.Y(n_330)
);

OAI22xp33_ASAP7_75t_L g531 ( 
.A1(n_85),
.A2(n_103),
.B1(n_483),
.B2(n_532),
.Y(n_531)
);

OAI21xp5_ASAP7_75t_L g546 ( 
.A1(n_85),
.A2(n_532),
.B(n_547),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_SL g568 ( 
.A(n_85),
.B(n_432),
.Y(n_568)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_86),
.A2(n_331),
.B1(n_436),
.B2(n_437),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_86),
.B(n_437),
.Y(n_489)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_104),
.Y(n_103)
);

OAI22x1_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_91),
.B1(n_95),
.B2(n_99),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_88),
.Y(n_223)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx4_ASAP7_75t_L g396 ( 
.A(n_89),
.Y(n_396)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_90),
.Y(n_214)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_90),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_90),
.Y(n_601)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_96),
.Y(n_108)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx6_ASAP7_75t_L g606 ( 
.A(n_97),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g498 ( 
.A(n_100),
.Y(n_498)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_103),
.Y(n_331)
);

OAI21xp33_ASAP7_75t_SL g482 ( 
.A1(n_103),
.A2(n_483),
.B(n_489),
.Y(n_482)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_108),
.B1(n_109),
.B2(n_111),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_106),
.Y(n_240)
);

BUFx5_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_107),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_107),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_111),
.Y(n_296)
);

INVx2_ASAP7_75t_SL g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_112),
.Y(n_487)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_112),
.Y(n_627)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_113),
.A2(n_330),
.B1(n_331),
.B2(n_332),
.Y(n_329)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_118),
.Y(n_291)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_118),
.Y(n_443)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_119),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_119),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g509 ( 
.A(n_123),
.Y(n_509)
);

AO22x1_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_140),
.B1(n_150),
.B2(n_162),
.Y(n_124)
);

OAI21xp33_ASAP7_75t_SL g183 ( 
.A1(n_125),
.A2(n_140),
.B(n_150),
.Y(n_183)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_125),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_125),
.A2(n_150),
.B1(n_256),
.B2(n_317),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_SL g333 ( 
.A1(n_125),
.A2(n_150),
.B1(n_317),
.B2(n_334),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_125),
.B(n_263),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_125),
.A2(n_150),
.B1(n_417),
.B2(n_418),
.Y(n_416)
);

AO22x1_ASAP7_75t_L g659 ( 
.A1(n_125),
.A2(n_150),
.B1(n_162),
.B2(n_334),
.Y(n_659)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

AND2x4_ASAP7_75t_L g150 ( 
.A(n_126),
.B(n_151),
.Y(n_150)
);

AOI22x1_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_130),
.B1(n_133),
.B2(n_137),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_129),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_136),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_136),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g515 ( 
.A(n_136),
.Y(n_515)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_144),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_145),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_145),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_145),
.Y(n_372)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVxp67_ASAP7_75t_SL g147 ( 
.A(n_148),
.Y(n_147)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_148),
.Y(n_261)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_149),
.Y(n_159)
);

INVx2_ASAP7_75t_SL g272 ( 
.A(n_150),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_150),
.B(n_263),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_155),
.B1(n_158),
.B2(n_160),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx3_ASAP7_75t_SL g163 ( 
.A(n_164),
.Y(n_163)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx5_ASAP7_75t_L g266 ( 
.A(n_165),
.Y(n_266)
);

INVx8_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_166),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_166),
.Y(n_364)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_171),
.Y(n_511)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_171),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_SL g689 ( 
.A1(n_172),
.A2(n_182),
.B1(n_183),
.B2(n_690),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_172),
.Y(n_690)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_181),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_181),
.Y(n_251)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx4_ASAP7_75t_SL g188 ( 
.A(n_189),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g375 ( 
.A(n_189),
.Y(n_375)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_693),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_649),
.B(n_691),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_470),
.B(n_640),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_406),
.Y(n_196)
);

AOI21x1_ASAP7_75t_L g640 ( 
.A1(n_197),
.A2(n_641),
.B(n_645),
.Y(n_640)
);

OA21x2_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_321),
.B(n_352),
.Y(n_197)
);

NOR2x1_ASAP7_75t_SL g646 ( 
.A(n_198),
.B(n_321),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_198),
.B(n_321),
.Y(n_648)
);

MAJx2_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_273),
.C(n_298),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_199),
.B(n_354),
.Y(n_353)
);

MAJx2_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_241),
.C(n_252),
.Y(n_199)
);

XNOR2x1_ASAP7_75t_L g403 ( 
.A(n_200),
.B(n_404),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_224),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_201),
.B(n_224),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_209),
.B1(n_217),
.B2(n_220),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_202),
.A2(n_220),
.B(n_302),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_202),
.A2(n_278),
.B1(n_393),
.B2(n_462),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_L g550 ( 
.A1(n_202),
.A2(n_551),
.B(n_559),
.Y(n_550)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_203),
.Y(n_202)
);

OA21x2_ASAP7_75t_L g276 ( 
.A1(n_203),
.A2(n_277),
.B(n_280),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_203),
.A2(n_210),
.B1(n_389),
.B2(n_392),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_203),
.B(n_494),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g590 ( 
.A1(n_203),
.A2(n_591),
.B1(n_592),
.B2(n_593),
.Y(n_590)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_207),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_204),
.Y(n_222)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

BUFx2_ASAP7_75t_L g216 ( 
.A(n_205),
.Y(n_216)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_205),
.Y(n_284)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_205),
.Y(n_398)
);

INVx6_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_206),
.Y(n_467)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_206),
.Y(n_616)
);

INVx8_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx8_ASAP7_75t_L g561 ( 
.A(n_208),
.Y(n_561)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_211),
.Y(n_558)
);

BUFx3_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

BUFx12f_ASAP7_75t_L g496 ( 
.A(n_214),
.Y(n_496)
);

BUFx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

BUFx4f_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_225),
.Y(n_436)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_227),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_229),
.Y(n_294)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_230),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_230),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g621 ( 
.A(n_230),
.Y(n_621)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

BUFx2_ASAP7_75t_L g488 ( 
.A(n_234),
.Y(n_488)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_236),
.Y(n_611)
);

INVx5_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_241),
.B(n_253),
.Y(n_404)
);

INVx2_ASAP7_75t_SL g244 ( 
.A(n_245),
.Y(n_244)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_255),
.B1(n_262),
.B2(n_272),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g458 ( 
.A1(n_254),
.A2(n_459),
.B(n_460),
.Y(n_458)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

BUFx2_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_269),
.Y(n_366)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

OA21x2_ASAP7_75t_L g361 ( 
.A1(n_272),
.A2(n_362),
.B(n_367),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_SL g522 ( 
.A1(n_272),
.A2(n_367),
.B(n_523),
.Y(n_522)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_274),
.B(n_299),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_276),
.B1(n_285),
.B2(n_297),
.Y(n_274)
);

OA21x2_ASAP7_75t_SL g653 ( 
.A1(n_275),
.A2(n_351),
.B(n_654),
.Y(n_653)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_276),
.B(n_343),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_276),
.B(n_285),
.Y(n_351)
);

INVx4_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx5_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g592 ( 
.A(n_279),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_280),
.B(n_303),
.Y(n_302)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_283),
.Y(n_556)
);

BUFx2_ASAP7_75t_L g572 ( 
.A(n_283),
.Y(n_572)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_285),
.Y(n_297)
);

BUFx2_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx4_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_291),
.Y(n_439)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_291),
.Y(n_503)
);

INVxp67_ASAP7_75t_SL g332 ( 
.A(n_292),
.Y(n_332)
);

BUFx6f_ASAP7_75t_SL g293 ( 
.A(n_294),
.Y(n_293)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVxp33_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_308),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_300),
.B(n_323),
.C(n_325),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_307),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_301),
.B(n_401),
.Y(n_400)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_303),
.Y(n_492)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_306),
.Y(n_391)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_306),
.Y(n_577)
);

HB1xp67_ASAP7_75t_L g401 ( 
.A(n_307),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_316),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_309),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_315),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_310),
.B(n_426),
.Y(n_425)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVxp33_ASAP7_75t_L g326 ( 
.A(n_316),
.Y(n_326)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

XNOR2x1_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_327),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g668 ( 
.A1(n_322),
.A2(n_669),
.B(n_671),
.Y(n_668)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_341),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g669 ( 
.A(n_328),
.B(n_670),
.Y(n_669)
);

NAND2xp33_ASAP7_75t_R g671 ( 
.A(n_328),
.B(n_670),
.Y(n_671)
);

OA21x2_ASAP7_75t_SL g328 ( 
.A1(n_329),
.A2(n_333),
.B(n_340),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_329),
.B(n_333),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_331),
.B(n_437),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_331),
.B(n_624),
.Y(n_623)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_339),
.Y(n_420)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_339),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_R g660 ( 
.A(n_340),
.B(n_661),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_340),
.B(n_662),
.Y(n_663)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_340),
.Y(n_666)
);

INVxp33_ASAP7_75t_L g670 ( 
.A(n_341),
.Y(n_670)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_351),
.Y(n_341)
);

HB1xp67_ASAP7_75t_L g654 ( 
.A(n_343),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_345),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_344),
.B(n_360),
.Y(n_359)
);

INVx3_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx4_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_355),
.Y(n_352)
);

OR2x2_ASAP7_75t_L g647 ( 
.A(n_353),
.B(n_355),
.Y(n_647)
);

OAI21x1_ASAP7_75t_L g355 ( 
.A1(n_356),
.A2(n_402),
.B(n_405),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_399),
.Y(n_356)
);

OR2x2_ASAP7_75t_L g405 ( 
.A(n_357),
.B(n_399),
.Y(n_405)
);

XOR2x1_ASAP7_75t_L g445 ( 
.A(n_357),
.B(n_446),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_361),
.C(n_368),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_358),
.A2(n_359),
.B1(n_361),
.B2(n_412),
.Y(n_411)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_361),
.Y(n_412)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_362),
.Y(n_417)
);

INVx8_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_368),
.B(n_411),
.Y(n_410)
);

OR2x2_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_388),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_369),
.B(n_388),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_370),
.A2(n_373),
.B1(n_379),
.B2(n_381),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_376),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

BUFx2_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_379),
.Y(n_433)
);

NAND2xp33_ASAP7_75t_SL g381 ( 
.A(n_382),
.B(n_385),
.Y(n_381)
);

HB1xp67_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx2_ASAP7_75t_SL g386 ( 
.A(n_387),
.Y(n_386)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx2_ASAP7_75t_SL g390 ( 
.A(n_391),
.Y(n_390)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx2_ASAP7_75t_SL g394 ( 
.A(n_395),
.Y(n_394)
);

INVx3_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_400),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

XNOR2x1_ASAP7_75t_L g446 ( 
.A(n_403),
.B(n_447),
.Y(n_446)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_SL g407 ( 
.A1(n_408),
.A2(n_445),
.B(n_448),
.Y(n_407)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_408),
.Y(n_643)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_413),
.C(n_444),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_409),
.A2(n_410),
.B1(n_450),
.B2(n_451),
.Y(n_449)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

HB1xp67_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_414),
.B(n_444),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_415),
.B(n_425),
.C(n_434),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_416),
.B(n_435),
.Y(n_454)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_418),
.Y(n_459)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx2_ASAP7_75t_SL g422 ( 
.A(n_423),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_SL g453 ( 
.A(n_425),
.B(n_454),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_SL g427 ( 
.A1(n_428),
.A2(n_432),
.B(n_433),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx2_ASAP7_75t_SL g429 ( 
.A(n_430),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

OR2x2_ASAP7_75t_L g507 ( 
.A(n_432),
.B(n_508),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_432),
.B(n_582),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_432),
.B(n_609),
.Y(n_608)
);

OAI21xp33_ASAP7_75t_SL g624 ( 
.A1(n_432),
.A2(n_608),
.B(n_625),
.Y(n_624)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_445),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_452),
.Y(n_448)
);

OR2x2_ASAP7_75t_L g642 ( 
.A(n_449),
.B(n_452),
.Y(n_642)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_450),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_455),
.C(n_456),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_453),
.B(n_473),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_455),
.A2(n_456),
.B1(n_457),
.B2(n_474),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_455),
.Y(n_474)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_458),
.B(n_461),
.C(n_468),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_SL g478 ( 
.A(n_458),
.B(n_479),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_461),
.A2(n_468),
.B1(n_469),
.B2(n_480),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_461),
.Y(n_480)
);

OA21x2_ASAP7_75t_L g491 ( 
.A1(n_462),
.A2(n_492),
.B(n_493),
.Y(n_491)
);

BUFx2_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_465),
.Y(n_587)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

AOI21x1_ASAP7_75t_L g470 ( 
.A1(n_471),
.A2(n_516),
.B(n_638),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_475),
.Y(n_471)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_472),
.Y(n_639)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_476),
.B(n_639),
.Y(n_638)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_477),
.B(n_481),
.C(n_490),
.Y(n_476)
);

INVxp67_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g518 ( 
.A(n_478),
.B(n_519),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_L g519 ( 
.A1(n_481),
.A2(n_482),
.B1(n_490),
.B2(n_520),
.Y(n_519)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

INVx3_ASAP7_75t_SL g484 ( 
.A(n_485),
.Y(n_484)
);

INVx4_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

INVx4_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_489),
.B(n_623),
.Y(n_622)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_490),
.Y(n_520)
);

OR2x2_ASAP7_75t_L g490 ( 
.A(n_491),
.B(n_499),
.Y(n_490)
);

XNOR2x1_ASAP7_75t_L g541 ( 
.A(n_491),
.B(n_499),
.Y(n_541)
);

OAI21xp5_ASAP7_75t_SL g569 ( 
.A1(n_493),
.A2(n_570),
.B(n_574),
.Y(n_569)
);

NAND2xp33_ASAP7_75t_SL g559 ( 
.A(n_494),
.B(n_560),
.Y(n_559)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

INVx3_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_500),
.A2(n_504),
.B1(n_507),
.B2(n_510),
.Y(n_499)
);

BUFx3_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

BUFx2_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

INVx1_ASAP7_75t_SL g508 ( 
.A(n_509),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_511),
.B(n_512),
.Y(n_510)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

AO21x2_ASAP7_75t_L g516 ( 
.A1(n_517),
.A2(n_542),
.B(n_637),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_518),
.B(n_521),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_518),
.B(n_521),
.Y(n_637)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_522),
.B(n_530),
.C(n_540),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g564 ( 
.A(n_522),
.B(n_531),
.Y(n_564)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_525),
.Y(n_524)
);

INVx3_ASAP7_75t_SL g525 ( 
.A(n_526),
.Y(n_525)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_528),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_529),
.Y(n_528)
);

HB1xp67_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);

INVx4_ASAP7_75t_L g533 ( 
.A(n_534),
.Y(n_533)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_535),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_536),
.Y(n_535)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_538),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_539),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_L g562 ( 
.A1(n_540),
.A2(n_541),
.B1(n_563),
.B2(n_564),
.Y(n_562)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_541),
.Y(n_540)
);

OAI321xp33_ASAP7_75t_L g542 ( 
.A1(n_543),
.A2(n_565),
.A3(n_629),
.B1(n_635),
.B2(n_636),
.C(n_705),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_544),
.B(n_562),
.Y(n_543)
);

OR2x2_ASAP7_75t_L g636 ( 
.A(n_544),
.B(n_562),
.Y(n_636)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_545),
.B(n_548),
.C(n_550),
.Y(n_544)
);

HB1xp67_ASAP7_75t_L g545 ( 
.A(n_546),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_L g633 ( 
.A1(n_546),
.A2(n_548),
.B1(n_549),
.B2(n_634),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_546),
.Y(n_634)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_549),
.Y(n_548)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_550),
.Y(n_632)
);

INVxp33_ASAP7_75t_SL g591 ( 
.A(n_551),
.Y(n_591)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_553),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_554),
.Y(n_553)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_554),
.Y(n_573)
);

INVx4_ASAP7_75t_L g554 ( 
.A(n_555),
.Y(n_554)
);

INVx4_ASAP7_75t_L g555 ( 
.A(n_556),
.Y(n_555)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_558),
.Y(n_557)
);

INVx5_ASAP7_75t_L g560 ( 
.A(n_561),
.Y(n_560)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_564),
.Y(n_563)
);

AOI21xp5_ASAP7_75t_L g565 ( 
.A1(n_566),
.A2(n_589),
.B(n_628),
.Y(n_565)
);

OAI21xp5_ASAP7_75t_SL g566 ( 
.A1(n_567),
.A2(n_578),
.B(n_588),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_568),
.B(n_569),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_568),
.B(n_569),
.Y(n_588)
);

INVxp67_ASAP7_75t_L g593 ( 
.A(n_570),
.Y(n_593)
);

INVx2_ASAP7_75t_SL g571 ( 
.A(n_572),
.Y(n_571)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_575),
.Y(n_574)
);

INVx4_ASAP7_75t_L g575 ( 
.A(n_576),
.Y(n_575)
);

INVx2_ASAP7_75t_SL g576 ( 
.A(n_577),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_579),
.B(n_580),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_SL g580 ( 
.A(n_581),
.B(n_586),
.Y(n_580)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_583),
.Y(n_582)
);

BUFx2_ASAP7_75t_L g583 ( 
.A(n_584),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_585),
.Y(n_584)
);

INVx5_ASAP7_75t_L g586 ( 
.A(n_587),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_590),
.B(n_594),
.Y(n_589)
);

NOR2xp67_ASAP7_75t_L g628 ( 
.A(n_590),
.B(n_594),
.Y(n_628)
);

XNOR2xp5_ASAP7_75t_L g594 ( 
.A(n_595),
.B(n_622),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_595),
.B(n_622),
.Y(n_630)
);

AOI22xp5_ASAP7_75t_L g595 ( 
.A1(n_596),
.A2(n_607),
.B1(n_612),
.B2(n_617),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_597),
.B(n_602),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_598),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_599),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_600),
.Y(n_599)
);

HB1xp67_ASAP7_75t_L g600 ( 
.A(n_601),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_602),
.B(n_618),
.Y(n_617)
);

BUFx2_ASAP7_75t_L g602 ( 
.A(n_603),
.Y(n_602)
);

HB1xp67_ASAP7_75t_L g603 ( 
.A(n_604),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_605),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_606),
.Y(n_605)
);

INVxp67_ASAP7_75t_L g607 ( 
.A(n_608),
.Y(n_607)
);

INVx3_ASAP7_75t_L g609 ( 
.A(n_610),
.Y(n_609)
);

BUFx6f_ASAP7_75t_L g610 ( 
.A(n_611),
.Y(n_610)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_613),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_614),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_615),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_616),
.Y(n_615)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_619),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_620),
.Y(n_619)
);

INVx4_ASAP7_75t_L g620 ( 
.A(n_621),
.Y(n_620)
);

BUFx4f_ASAP7_75t_SL g625 ( 
.A(n_626),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_627),
.Y(n_626)
);

NOR2xp67_ASAP7_75t_L g629 ( 
.A(n_630),
.B(n_631),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_630),
.B(n_631),
.Y(n_635)
);

XNOR2xp5_ASAP7_75t_L g631 ( 
.A(n_632),
.B(n_633),
.Y(n_631)
);

MAJIxp5_ASAP7_75t_L g641 ( 
.A(n_642),
.B(n_643),
.C(n_644),
.Y(n_641)
);

OAI21xp5_ASAP7_75t_L g645 ( 
.A1(n_646),
.A2(n_647),
.B(n_648),
.Y(n_645)
);

NOR3xp33_ASAP7_75t_L g649 ( 
.A(n_650),
.B(n_672),
.C(n_684),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_651),
.Y(n_650)
);

NAND2xp33_ASAP7_75t_L g651 ( 
.A(n_652),
.B(n_668),
.Y(n_651)
);

NOR2xp67_ASAP7_75t_L g697 ( 
.A(n_652),
.B(n_668),
.Y(n_697)
);

XOR2xp5_ASAP7_75t_L g652 ( 
.A(n_653),
.B(n_655),
.Y(n_652)
);

MAJIxp5_ASAP7_75t_L g680 ( 
.A(n_653),
.B(n_681),
.C(n_682),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_656),
.B(n_664),
.Y(n_655)
);

AOI22xp33_ASAP7_75t_L g656 ( 
.A1(n_657),
.A2(n_658),
.B1(n_660),
.B2(n_663),
.Y(n_656)
);

AOI22xp5_ASAP7_75t_L g664 ( 
.A1(n_657),
.A2(n_658),
.B1(n_665),
.B2(n_667),
.Y(n_664)
);

OAI22xp33_ASAP7_75t_L g681 ( 
.A1(n_657),
.A2(n_658),
.B1(n_661),
.B2(n_662),
.Y(n_681)
);

INVx1_ASAP7_75t_SL g657 ( 
.A(n_658),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_661),
.B(n_666),
.Y(n_665)
);

AOI22xp5_ASAP7_75t_SL g676 ( 
.A1(n_661),
.A2(n_662),
.B1(n_677),
.B2(n_678),
.Y(n_676)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_662),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_662),
.B(n_666),
.Y(n_667)
);

MAJIxp5_ASAP7_75t_L g686 ( 
.A(n_662),
.B(n_678),
.C(n_687),
.Y(n_686)
);

BUFx2_ASAP7_75t_L g683 ( 
.A(n_666),
.Y(n_683)
);

OAI21xp5_ASAP7_75t_L g695 ( 
.A1(n_672),
.A2(n_696),
.B(n_698),
.Y(n_695)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_673),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_674),
.B(n_680),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_674),
.B(n_680),
.Y(n_699)
);

XNOR2xp5_ASAP7_75t_L g674 ( 
.A(n_675),
.B(n_676),
.Y(n_674)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_675),
.Y(n_687)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_678),
.Y(n_677)
);

CKINVDCx14_ASAP7_75t_R g682 ( 
.A(n_683),
.Y(n_682)
);

INVxp67_ASAP7_75t_SL g694 ( 
.A(n_684),
.Y(n_694)
);

INVxp67_ASAP7_75t_SL g684 ( 
.A(n_685),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_686),
.B(n_688),
.Y(n_685)
);

OR2x2_ASAP7_75t_L g692 ( 
.A(n_686),
.B(n_688),
.Y(n_692)
);

INVxp67_ASAP7_75t_L g691 ( 
.A(n_692),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_694),
.B(n_695),
.Y(n_693)
);

INVx1_ASAP7_75t_SL g696 ( 
.A(n_697),
.Y(n_696)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_699),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_701),
.Y(n_700)
);


endmodule