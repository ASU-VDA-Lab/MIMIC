module real_jpeg_32286_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_548;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_546;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_537;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx2_ASAP7_75t_L g82 ( 
.A(n_0),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_0),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_0),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_0),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_1),
.A2(n_61),
.B1(n_65),
.B2(n_66),
.Y(n_60)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_1),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_1),
.A2(n_65),
.B1(n_214),
.B2(n_217),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_1),
.A2(n_65),
.B1(n_149),
.B2(n_272),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_2),
.A2(n_230),
.B1(n_235),
.B2(n_236),
.Y(n_229)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_2),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g344 ( 
.A1(n_2),
.A2(n_235),
.B1(n_345),
.B2(n_350),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_2),
.A2(n_235),
.B1(n_423),
.B2(n_424),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_2),
.A2(n_235),
.B1(n_478),
.B2(n_479),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_3),
.A2(n_262),
.B1(n_263),
.B2(n_265),
.Y(n_261)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_3),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_4),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_4),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_4),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_5),
.A2(n_111),
.B1(n_117),
.B2(n_118),
.Y(n_110)
);

INVx2_ASAP7_75t_R g117 ( 
.A(n_5),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_5),
.A2(n_117),
.B1(n_241),
.B2(n_244),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_5),
.A2(n_117),
.B1(n_371),
.B2(n_374),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_5),
.A2(n_117),
.B1(n_442),
.B2(n_446),
.Y(n_441)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_6),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_6),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_7),
.Y(n_157)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_7),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_8),
.A2(n_133),
.B1(n_136),
.B2(n_138),
.Y(n_132)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_8),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g328 ( 
.A1(n_8),
.A2(n_138),
.B1(n_329),
.B2(n_330),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_L g458 ( 
.A1(n_8),
.A2(n_138),
.B1(n_423),
.B2(n_459),
.Y(n_458)
);

AOI22xp33_ASAP7_75t_SL g466 ( 
.A1(n_8),
.A2(n_138),
.B1(n_467),
.B2(n_468),
.Y(n_466)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_9),
.A2(n_85),
.B1(n_88),
.B2(n_89),
.Y(n_84)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_9),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g290 ( 
.A1(n_9),
.A2(n_89),
.B1(n_291),
.B2(n_293),
.Y(n_290)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_10),
.Y(n_64)
);

AOI21x1_ASAP7_75t_L g27 ( 
.A1(n_11),
.A2(n_28),
.B(n_34),
.Y(n_27)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_11),
.A2(n_35),
.B1(n_171),
.B2(n_175),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_11),
.A2(n_35),
.B1(n_358),
.B2(n_359),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_12),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_13),
.B(n_209),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_13),
.A2(n_208),
.B(n_313),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_13),
.B(n_363),
.Y(n_362)
);

OAI32xp33_ASAP7_75t_L g379 ( 
.A1(n_13),
.A2(n_152),
.A3(n_380),
.B1(n_383),
.B2(n_389),
.Y(n_379)
);

INVx1_ASAP7_75t_SL g390 ( 
.A(n_13),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_13),
.B(n_179),
.Y(n_455)
);

OAI22xp33_ASAP7_75t_SL g484 ( 
.A1(n_13),
.A2(n_256),
.B1(n_477),
.B2(n_485),
.Y(n_484)
);

AOI22xp33_ASAP7_75t_L g502 ( 
.A1(n_13),
.A2(n_390),
.B1(n_503),
.B2(n_508),
.Y(n_502)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_15),
.A2(n_141),
.B1(n_148),
.B2(n_149),
.Y(n_140)
);

INVx2_ASAP7_75t_R g148 ( 
.A(n_15),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_15),
.A2(n_148),
.B1(n_281),
.B2(n_283),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_SL g319 ( 
.A1(n_15),
.A2(n_148),
.B1(n_320),
.B2(n_323),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_15),
.A2(n_148),
.B1(n_397),
.B2(n_401),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_16),
.Y(n_102)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_16),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_16),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_16),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_17),
.A2(n_72),
.B1(n_74),
.B2(n_75),
.Y(n_71)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_17),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_17),
.A2(n_74),
.B1(n_251),
.B2(n_252),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_304),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_302),
.Y(n_19)
);

HB1xp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_266),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_22),
.B(n_266),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_182),
.C(n_248),
.Y(n_22)
);

HB1xp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g545 ( 
.A(n_24),
.B(n_546),
.Y(n_545)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_94),
.Y(n_24)
);

MAJx2_ASAP7_75t_L g300 ( 
.A(n_25),
.B(n_181),
.C(n_301),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_70),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g531 ( 
.A(n_26),
.B(n_70),
.Y(n_531)
);

OAI22x1_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_39),
.B1(n_60),
.B2(n_68),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_27),
.A2(n_39),
.B1(n_68),
.B2(n_319),
.Y(n_318)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_32),
.A2(n_166),
.B1(n_167),
.B2(n_169),
.Y(n_165)
);

INVx4_ASAP7_75t_L g394 ( 
.A(n_32),
.Y(n_394)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_33),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_36),
.Y(n_34)
);

BUFx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g254 ( 
.A(n_37),
.Y(n_254)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_37),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_38),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_38),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_39),
.A2(n_60),
.B1(n_68),
.B2(n_250),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_39),
.A2(n_68),
.B1(n_250),
.B2(n_290),
.Y(n_289)
);

OAI22xp33_ASAP7_75t_SL g368 ( 
.A1(n_39),
.A2(n_68),
.B1(n_319),
.B2(n_369),
.Y(n_368)
);

OAI22x1_ASAP7_75t_L g456 ( 
.A1(n_39),
.A2(n_68),
.B1(n_457),
.B2(n_458),
.Y(n_456)
);

AO21x2_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_47),
.B(n_52),
.Y(n_39)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_40),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_44),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_46),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_46),
.Y(n_376)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_46),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g419 ( 
.A(n_47),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_50),
.Y(n_47)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

INVxp67_ASAP7_75t_SL g420 ( 
.A(n_52),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_53),
.A2(n_55),
.B1(n_58),
.B2(n_59),
.Y(n_52)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_54),
.Y(n_58)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_54),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_54),
.Y(n_445)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_54),
.Y(n_449)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_57),
.Y(n_437)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

BUFx4f_ASAP7_75t_SL g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_64),
.Y(n_373)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g292 ( 
.A(n_67),
.Y(n_292)
);

INVx4_ASAP7_75t_L g425 ( 
.A(n_67),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_SL g482 ( 
.A(n_68),
.B(n_390),
.Y(n_482)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_68),
.Y(n_513)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_71),
.A2(n_78),
.B1(n_84),
.B2(n_90),
.Y(n_70)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_71),
.Y(n_222)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_73),
.Y(n_264)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_78),
.Y(n_212)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_78),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_78),
.A2(n_466),
.B1(n_477),
.B2(n_480),
.Y(n_476)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_83),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_82),
.Y(n_260)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_83),
.Y(n_216)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_83),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_84),
.A2(n_256),
.B1(n_257),
.B2(n_261),
.Y(n_255)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_86),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g360 ( 
.A(n_86),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx6_ASAP7_75t_L g430 ( 
.A(n_87),
.Y(n_430)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_87),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_87),
.Y(n_492)
);

INVx2_ASAP7_75t_SL g262 ( 
.A(n_88),
.Y(n_262)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_91),
.A2(n_356),
.B1(n_465),
.B2(n_472),
.Y(n_464)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx8_ASAP7_75t_L g298 ( 
.A(n_93),
.Y(n_298)
);

INVx4_ASAP7_75t_SL g485 ( 
.A(n_93),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_96),
.B1(n_139),
.B2(n_181),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVxp67_ASAP7_75t_SL g301 ( 
.A(n_96),
.Y(n_301)
);

OAI22x1_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_110),
.B1(n_120),
.B2(n_132),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_L g311 ( 
.A1(n_97),
.A2(n_120),
.B1(n_229),
.B2(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_97),
.Y(n_363)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_98),
.Y(n_227)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_98),
.Y(n_278)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_99),
.B(n_122),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_103),
.B1(n_106),
.B2(n_108),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_101),
.Y(n_177)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_102),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_102),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_102),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_102),
.Y(n_507)
);

INVx2_ASAP7_75t_SL g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_105),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_105),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_105),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_105),
.Y(n_194)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_105),
.Y(n_203)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_107),
.Y(n_150)
);

INVx2_ASAP7_75t_SL g243 ( 
.A(n_107),
.Y(n_243)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_110),
.A2(n_120),
.B1(n_277),
.B2(n_279),
.Y(n_276)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_115),
.Y(n_119)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_115),
.Y(n_137)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_115),
.Y(n_189)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_116),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_116),
.Y(n_135)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_116),
.Y(n_316)
);

HB1xp67_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_119),
.Y(n_209)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_121),
.A2(n_225),
.B1(n_226),
.B2(n_228),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_125),
.B1(n_128),
.B2(n_130),
.Y(n_122)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_129),
.Y(n_282)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_132),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

HB1xp67_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_139),
.Y(n_181)
);

OAI22x1_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_151),
.B1(n_170),
.B2(n_178),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_140),
.A2(n_151),
.B1(n_178),
.B2(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_146),
.Y(n_198)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_146),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_147),
.Y(n_247)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_SL g275 ( 
.A(n_151),
.Y(n_275)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_151),
.Y(n_343)
);

AO21x2_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_158),
.B(n_165),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_155),
.Y(n_152)
);

INVx1_ASAP7_75t_SL g329 ( 
.A(n_153),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_154),
.Y(n_206)
);

INVx8_ASAP7_75t_L g273 ( 
.A(n_154),
.Y(n_273)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_157),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_162),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

BUFx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx8_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_164),
.Y(n_331)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_165),
.Y(n_180)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_166),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_167),
.Y(n_251)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_170),
.Y(n_274)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_178),
.A2(n_240),
.B1(n_327),
.B2(n_328),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_178),
.A2(n_328),
.B1(n_342),
.B2(n_344),
.Y(n_341)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_179),
.A2(n_271),
.B1(n_274),
.B2(n_275),
.Y(n_270)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_180),
.A2(n_327),
.B1(n_344),
.B2(n_502),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_223),
.C(n_237),
.Y(n_182)
);

MAJx2_ASAP7_75t_L g544 ( 
.A(n_183),
.B(n_223),
.C(n_237),
.Y(n_544)
);

INVxp33_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g535 ( 
.A(n_184),
.B(n_536),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_210),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_185),
.A2(n_210),
.B1(n_211),
.B2(n_334),
.Y(n_333)
);

OAI32xp33_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_190),
.A3(n_195),
.B1(n_199),
.B2(n_207),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

OAI32xp33_ASAP7_75t_L g335 ( 
.A1(n_190),
.A2(n_195),
.A3(n_199),
.B1(n_207),
.B2(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_192),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_200),
.B(n_204),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_213),
.B1(n_220),
.B2(n_222),
.Y(n_211)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_212),
.Y(n_256)
);

OA21x2_ASAP7_75t_L g296 ( 
.A1(n_212),
.A2(n_297),
.B(n_299),
.Y(n_296)
);

AO22x1_ASAP7_75t_L g395 ( 
.A1(n_212),
.A2(n_220),
.B1(n_357),
.B2(n_396),
.Y(n_395)
);

AO22x1_ASAP7_75t_SL g351 ( 
.A1(n_213),
.A2(n_352),
.B1(n_356),
.B2(n_357),
.Y(n_351)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_224),
.A2(n_238),
.B1(n_239),
.B2(n_537),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_224),
.Y(n_537)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_232),
.Y(n_284)
);

INVx6_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_233),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx2_ASAP7_75t_SL g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx2_ASAP7_75t_SL g246 ( 
.A(n_247),
.Y(n_246)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_247),
.Y(n_382)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_248),
.Y(n_546)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_255),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_249),
.B(n_255),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_253),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx4_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx2_ASAP7_75t_SL g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_261),
.Y(n_299)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_287),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

OAI22xp33_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_276),
.B1(n_285),
.B2(n_286),
.Y(n_269)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_270),
.Y(n_286)
);

INVx5_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx5_ASAP7_75t_L g350 ( 
.A(n_273),
.Y(n_350)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_275),
.Y(n_327)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_276),
.Y(n_285)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_300),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_SL g288 ( 
.A(n_289),
.B(n_296),
.Y(n_288)
);

INVx2_ASAP7_75t_SL g291 ( 
.A(n_292),
.Y(n_291)
);

BUFx6f_ASAP7_75t_SL g293 ( 
.A(n_294),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx4_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

AOI21x1_ASAP7_75t_L g304 ( 
.A1(n_305),
.A2(n_524),
.B(n_547),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

AOI21x1_ASAP7_75t_L g306 ( 
.A1(n_307),
.A2(n_405),
.B(n_523),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_308),
.B(n_364),
.Y(n_307)
);

NOR2xp67_ASAP7_75t_SL g523 ( 
.A(n_308),
.B(n_364),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_SL g308 ( 
.A(n_309),
.B(n_332),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_309),
.B(n_333),
.C(n_340),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_SL g309 ( 
.A(n_310),
.B(n_317),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_311),
.B(n_318),
.C(n_326),
.Y(n_530)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_314),
.Y(n_313)
);

BUFx2_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_315),
.Y(n_339)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_326),
.Y(n_317)
);

INVx2_ASAP7_75t_SL g320 ( 
.A(n_321),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_340),
.Y(n_332)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx2_ASAP7_75t_SL g336 ( 
.A(n_337),
.Y(n_336)
);

BUFx3_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_351),
.C(n_361),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_341),
.B(n_366),
.Y(n_365)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

BUFx3_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx3_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx4_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_351),
.B(n_362),
.Y(n_366)
);

INVx3_ASAP7_75t_SL g352 ( 
.A(n_353),
.Y(n_352)
);

INVx8_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_355),
.Y(n_452)
);

HB1xp67_ASAP7_75t_L g481 ( 
.A(n_355),
.Y(n_481)
);

BUFx3_ASAP7_75t_L g489 ( 
.A(n_355),
.Y(n_489)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_356),
.Y(n_440)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_367),
.C(n_377),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_SL g518 ( 
.A(n_365),
.B(n_519),
.Y(n_518)
);

AOI21xp5_ASAP7_75t_L g519 ( 
.A1(n_367),
.A2(n_378),
.B(n_520),
.Y(n_519)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_SL g520 ( 
.A(n_368),
.B(n_378),
.Y(n_520)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_370),
.A2(n_417),
.B1(n_512),
.B2(n_513),
.Y(n_511)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx4_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx5_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_376),
.Y(n_414)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_395),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_SL g499 ( 
.A(n_379),
.B(n_395),
.Y(n_499)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

BUFx3_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVxp67_ASAP7_75t_SL g416 ( 
.A(n_386),
.Y(n_416)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

BUFx3_ASAP7_75t_L g423 ( 
.A(n_387),
.Y(n_423)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_391),
.Y(n_389)
);

OAI21xp33_ASAP7_75t_SL g412 ( 
.A1(n_390),
.A2(n_413),
.B(n_415),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_390),
.B(n_416),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_390),
.B(n_488),
.Y(n_487)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx3_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_396),
.Y(n_453)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx5_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx4_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVx4_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_404),
.Y(n_434)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_404),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_L g405 ( 
.A1(n_406),
.A2(n_517),
.B(n_522),
.Y(n_405)
);

AOI21x1_ASAP7_75t_L g406 ( 
.A1(n_407),
.A2(n_496),
.B(n_516),
.Y(n_406)
);

OAI21x1_ASAP7_75t_L g407 ( 
.A1(n_408),
.A2(n_462),
.B(n_495),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_438),
.Y(n_408)
);

OR2x2_ASAP7_75t_L g495 ( 
.A(n_409),
.B(n_438),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_410),
.B(n_426),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_410),
.A2(n_411),
.B1(n_426),
.B2(n_427),
.Y(n_473)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_412),
.A2(n_417),
.B1(n_421),
.B2(n_422),
.Y(n_411)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g431 ( 
.A1(n_415),
.A2(n_432),
.B(n_435),
.Y(n_431)
);

OA21x2_ASAP7_75t_SL g417 ( 
.A1(n_418),
.A2(n_419),
.B(n_420),
.Y(n_417)
);

AOI21xp33_ASAP7_75t_L g427 ( 
.A1(n_419),
.A2(n_428),
.B(n_431),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_420),
.Y(n_421)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_422),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

BUFx2_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

BUFx2_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVx1_ASAP7_75t_SL g432 ( 
.A(n_433),
.Y(n_432)
);

BUFx2_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

BUFx2_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_439),
.B(n_454),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_439),
.B(n_456),
.C(n_460),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_L g439 ( 
.A1(n_440),
.A2(n_441),
.B1(n_450),
.B2(n_453),
.Y(n_439)
);

INVxp67_ASAP7_75t_L g472 ( 
.A(n_441),
.Y(n_472)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

BUFx3_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_444),
.Y(n_467)
);

INVx6_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

BUFx3_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

INVx4_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

BUFx2_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_L g454 ( 
.A1(n_455),
.A2(n_456),
.B1(n_460),
.B2(n_461),
.Y(n_454)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_455),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_456),
.Y(n_461)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_458),
.Y(n_512)
);

AOI21xp5_ASAP7_75t_L g462 ( 
.A1(n_463),
.A2(n_474),
.B(n_494),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_473),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_464),
.B(n_473),
.Y(n_494)
);

INVxp67_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_467),
.Y(n_479)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

OAI21xp5_ASAP7_75t_SL g474 ( 
.A1(n_475),
.A2(n_483),
.B(n_493),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_482),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_476),
.B(n_482),
.Y(n_493)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_484),
.B(n_486),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_R g486 ( 
.A(n_487),
.B(n_490),
.Y(n_486)
);

INVx3_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

HB1xp67_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_497),
.B(n_498),
.Y(n_496)
);

NOR2x1_ASAP7_75t_SL g516 ( 
.A(n_497),
.B(n_498),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_499),
.B(n_500),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_499),
.B(n_511),
.C(n_515),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_501),
.A2(n_511),
.B1(n_514),
.B2(n_515),
.Y(n_500)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_501),
.Y(n_515)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

BUFx3_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_511),
.Y(n_514)
);

NOR2x1_ASAP7_75t_SL g517 ( 
.A(n_518),
.B(n_521),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_518),
.B(n_521),
.Y(n_522)
);

NOR2xp67_ASAP7_75t_L g524 ( 
.A(n_525),
.B(n_538),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_526),
.Y(n_525)
);

OR2x2_ASAP7_75t_L g526 ( 
.A(n_527),
.B(n_528),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_527),
.B(n_528),
.Y(n_549)
);

XNOR2xp5_ASAP7_75t_L g528 ( 
.A(n_529),
.B(n_534),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_L g529 ( 
.A1(n_530),
.A2(n_531),
.B1(n_532),
.B2(n_533),
.Y(n_529)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_530),
.Y(n_532)
);

INVxp33_ASAP7_75t_L g542 ( 
.A(n_530),
.Y(n_542)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_531),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_533),
.B(n_535),
.C(n_542),
.Y(n_541)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_535),
.Y(n_534)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_539),
.Y(n_538)
);

HB1xp67_ASAP7_75t_L g539 ( 
.A(n_540),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_541),
.B(n_543),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_541),
.B(n_543),
.C(n_549),
.Y(n_548)
);

XNOR2xp5_ASAP7_75t_L g543 ( 
.A(n_544),
.B(n_545),
.Y(n_543)
);

HB1xp67_ASAP7_75t_L g547 ( 
.A(n_548),
.Y(n_547)
);


endmodule