module fake_netlist_6_152_n_5895 (n_52, n_591, n_435, n_1, n_91, n_326, n_256, n_440, n_587, n_695, n_507, n_580, n_209, n_367, n_465, n_680, n_590, n_625, n_63, n_661, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_607, n_671, n_316, n_419, n_28, n_304, n_212, n_700, n_50, n_694, n_7, n_578, n_703, n_144, n_365, n_125, n_168, n_384, n_297, n_595, n_627, n_524, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_575, n_677, n_396, n_495, n_350, n_78, n_84, n_585, n_568, n_392, n_442, n_480, n_142, n_143, n_382, n_673, n_180, n_62, n_628, n_557, n_349, n_643, n_233, n_617, n_698, n_255, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_38, n_471, n_289, n_421, n_424, n_615, n_59, n_181, n_182, n_238, n_573, n_202, n_320, n_108, n_639, n_676, n_327, n_369, n_597, n_685, n_280, n_287, n_353, n_610, n_555, n_389, n_415, n_65, n_230, n_605, n_461, n_141, n_383, n_669, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_667, n_71, n_74, n_229, n_542, n_644, n_682, n_621, n_305, n_72, n_532, n_173, n_535, n_691, n_250, n_372, n_468, n_544, n_111, n_504, n_314, n_378, n_413, n_377, n_35, n_183, n_510, n_79, n_375, n_601, n_338, n_522, n_466, n_704, n_506, n_56, n_360, n_603, n_119, n_235, n_536, n_622, n_147, n_191, n_340, n_710, n_387, n_452, n_616, n_658, n_39, n_344, n_73, n_581, n_428, n_609, n_432, n_641, n_693, n_101, n_167, n_631, n_174, n_127, n_516, n_153, n_525, n_611, n_156, n_491, n_145, n_42, n_133, n_656, n_96, n_8, n_666, n_371, n_567, n_189, n_405, n_213, n_538, n_294, n_302, n_499, n_380, n_129, n_705, n_647, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_539, n_493, n_397, n_155, n_109, n_614, n_529, n_445, n_425, n_684, n_122, n_45, n_454, n_34, n_218, n_638, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_653, n_112, n_172, n_713, n_648, n_657, n_576, n_472, n_270, n_239, n_126, n_414, n_97, n_563, n_58, n_490, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_708, n_196, n_402, n_352, n_668, n_478, n_626, n_574, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_662, n_89, n_374, n_659, n_709, n_366, n_407, n_450, n_103, n_272, n_526, n_185, n_712, n_348, n_711, n_579, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_559, n_53, n_370, n_44, n_458, n_232, n_650, n_16, n_163, n_46, n_330, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_551, n_154, n_699, n_456, n_564, n_98, n_260, n_265, n_313, n_451, n_624, n_279, n_686, n_252, n_228, n_565, n_594, n_356, n_577, n_166, n_184, n_552, n_619, n_216, n_455, n_83, n_521, n_363, n_572, n_395, n_592, n_654, n_323, n_606, n_393, n_411, n_503, n_716, n_152, n_623, n_92, n_599, n_513, n_321, n_645, n_331, n_105, n_227, n_132, n_570, n_406, n_483, n_102, n_204, n_482, n_474, n_527, n_261, n_608, n_620, n_420, n_683, n_630, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_476, n_714, n_2, n_291, n_219, n_543, n_357, n_150, n_264, n_263, n_589, n_481, n_325, n_329, n_464, n_600, n_561, n_33, n_477, n_549, n_533, n_408, n_61, n_237, n_584, n_244, n_399, n_76, n_243, n_124, n_548, n_94, n_282, n_436, n_116, n_211, n_523, n_117, n_175, n_322, n_707, n_345, n_409, n_231, n_354, n_689, n_40, n_505, n_240, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_558, n_635, n_95, n_311, n_10, n_403, n_253, n_634, n_583, n_596, n_123, n_136, n_546, n_562, n_249, n_201, n_386, n_556, n_159, n_157, n_162, n_692, n_115, n_487, n_550, n_128, n_241, n_30, n_275, n_553, n_43, n_652, n_560, n_642, n_276, n_569, n_441, n_221, n_444, n_586, n_423, n_146, n_318, n_303, n_511, n_715, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_418, n_113, n_618, n_582, n_4, n_199, n_138, n_266, n_296, n_674, n_571, n_268, n_271, n_404, n_651, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_679, n_5, n_453, n_612, n_633, n_665, n_333, n_588, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_632, n_702, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_672, n_534, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_675, n_85, n_99, n_257, n_655, n_13, n_706, n_670, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_690, n_29, n_75, n_401, n_324, n_335, n_430, n_463, n_545, n_489, n_205, n_604, n_120, n_251, n_301, n_274, n_636, n_681, n_110, n_151, n_412, n_640, n_81, n_660, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_598, n_422, n_696, n_688, n_135, n_165, n_351, n_437, n_259, n_177, n_540, n_593, n_514, n_646, n_528, n_391, n_457, n_687, n_697, n_364, n_637, n_295, n_385, n_701, n_629, n_388, n_190, n_262, n_484, n_613, n_187, n_501, n_531, n_60, n_361, n_508, n_663, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_566, n_554, n_602, n_194, n_664, n_171, n_678, n_192, n_57, n_169, n_51, n_649, n_283, n_5895);

input n_52;
input n_591;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_587;
input n_695;
input n_507;
input n_580;
input n_209;
input n_367;
input n_465;
input n_680;
input n_590;
input n_625;
input n_63;
input n_661;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_607;
input n_671;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_700;
input n_50;
input n_694;
input n_7;
input n_578;
input n_703;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_595;
input n_627;
input n_524;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_575;
input n_677;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_585;
input n_568;
input n_392;
input n_442;
input n_480;
input n_142;
input n_143;
input n_382;
input n_673;
input n_180;
input n_62;
input n_628;
input n_557;
input n_349;
input n_643;
input n_233;
input n_617;
input n_698;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_471;
input n_289;
input n_421;
input n_424;
input n_615;
input n_59;
input n_181;
input n_182;
input n_238;
input n_573;
input n_202;
input n_320;
input n_108;
input n_639;
input n_676;
input n_327;
input n_369;
input n_597;
input n_685;
input n_280;
input n_287;
input n_353;
input n_610;
input n_555;
input n_389;
input n_415;
input n_65;
input n_230;
input n_605;
input n_461;
input n_141;
input n_383;
input n_669;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_667;
input n_71;
input n_74;
input n_229;
input n_542;
input n_644;
input n_682;
input n_621;
input n_305;
input n_72;
input n_532;
input n_173;
input n_535;
input n_691;
input n_250;
input n_372;
input n_468;
input n_544;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_510;
input n_79;
input n_375;
input n_601;
input n_338;
input n_522;
input n_466;
input n_704;
input n_506;
input n_56;
input n_360;
input n_603;
input n_119;
input n_235;
input n_536;
input n_622;
input n_147;
input n_191;
input n_340;
input n_710;
input n_387;
input n_452;
input n_616;
input n_658;
input n_39;
input n_344;
input n_73;
input n_581;
input n_428;
input n_609;
input n_432;
input n_641;
input n_693;
input n_101;
input n_167;
input n_631;
input n_174;
input n_127;
input n_516;
input n_153;
input n_525;
input n_611;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_656;
input n_96;
input n_8;
input n_666;
input n_371;
input n_567;
input n_189;
input n_405;
input n_213;
input n_538;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_705;
input n_647;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_109;
input n_614;
input n_529;
input n_445;
input n_425;
input n_684;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_638;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_653;
input n_112;
input n_172;
input n_713;
input n_648;
input n_657;
input n_576;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_563;
input n_58;
input n_490;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_708;
input n_196;
input n_402;
input n_352;
input n_668;
input n_478;
input n_626;
input n_574;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_662;
input n_89;
input n_374;
input n_659;
input n_709;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_526;
input n_185;
input n_712;
input n_348;
input n_711;
input n_579;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_559;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_650;
input n_16;
input n_163;
input n_46;
input n_330;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_551;
input n_154;
input n_699;
input n_456;
input n_564;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_624;
input n_279;
input n_686;
input n_252;
input n_228;
input n_565;
input n_594;
input n_356;
input n_577;
input n_166;
input n_184;
input n_552;
input n_619;
input n_216;
input n_455;
input n_83;
input n_521;
input n_363;
input n_572;
input n_395;
input n_592;
input n_654;
input n_323;
input n_606;
input n_393;
input n_411;
input n_503;
input n_716;
input n_152;
input n_623;
input n_92;
input n_599;
input n_513;
input n_321;
input n_645;
input n_331;
input n_105;
input n_227;
input n_132;
input n_570;
input n_406;
input n_483;
input n_102;
input n_204;
input n_482;
input n_474;
input n_527;
input n_261;
input n_608;
input n_620;
input n_420;
input n_683;
input n_630;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_476;
input n_714;
input n_2;
input n_291;
input n_219;
input n_543;
input n_357;
input n_150;
input n_264;
input n_263;
input n_589;
input n_481;
input n_325;
input n_329;
input n_464;
input n_600;
input n_561;
input n_33;
input n_477;
input n_549;
input n_533;
input n_408;
input n_61;
input n_237;
input n_584;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_548;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_707;
input n_345;
input n_409;
input n_231;
input n_354;
input n_689;
input n_40;
input n_505;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_558;
input n_635;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_634;
input n_583;
input n_596;
input n_123;
input n_136;
input n_546;
input n_562;
input n_249;
input n_201;
input n_386;
input n_556;
input n_159;
input n_157;
input n_162;
input n_692;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_30;
input n_275;
input n_553;
input n_43;
input n_652;
input n_560;
input n_642;
input n_276;
input n_569;
input n_441;
input n_221;
input n_444;
input n_586;
input n_423;
input n_146;
input n_318;
input n_303;
input n_511;
input n_715;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_418;
input n_113;
input n_618;
input n_582;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_674;
input n_571;
input n_268;
input n_271;
input n_404;
input n_651;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_679;
input n_5;
input n_453;
input n_612;
input n_633;
input n_665;
input n_333;
input n_588;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_632;
input n_702;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_672;
input n_534;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_675;
input n_85;
input n_99;
input n_257;
input n_655;
input n_13;
input n_706;
input n_670;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_690;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_463;
input n_545;
input n_489;
input n_205;
input n_604;
input n_120;
input n_251;
input n_301;
input n_274;
input n_636;
input n_681;
input n_110;
input n_151;
input n_412;
input n_640;
input n_81;
input n_660;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_598;
input n_422;
input n_696;
input n_688;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_540;
input n_593;
input n_514;
input n_646;
input n_528;
input n_391;
input n_457;
input n_687;
input n_697;
input n_364;
input n_637;
input n_295;
input n_385;
input n_701;
input n_629;
input n_388;
input n_190;
input n_262;
input n_484;
input n_613;
input n_187;
input n_501;
input n_531;
input n_60;
input n_361;
input n_508;
input n_663;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_566;
input n_554;
input n_602;
input n_194;
input n_664;
input n_171;
input n_678;
input n_192;
input n_57;
input n_169;
input n_51;
input n_649;
input n_283;

output n_5895;

wire n_5643;
wire n_2542;
wire n_1671;
wire n_2817;
wire n_801;
wire n_4452;
wire n_2576;
wire n_5172;
wire n_4649;
wire n_1674;
wire n_5315;
wire n_741;
wire n_1351;
wire n_5254;
wire n_1212;
wire n_5362;
wire n_4251;
wire n_2157;
wire n_5019;
wire n_2332;
wire n_3849;
wire n_5138;
wire n_4388;
wire n_4395;
wire n_1061;
wire n_3089;
wire n_783;
wire n_5653;
wire n_4978;
wire n_5409;
wire n_5301;
wire n_1854;
wire n_3088;
wire n_3257;
wire n_1342;
wire n_4829;
wire n_5393;
wire n_1387;
wire n_3222;
wire n_4699;
wire n_1151;
wire n_4686;
wire n_2317;
wire n_5524;
wire n_5345;
wire n_1975;
wire n_1930;
wire n_3706;
wire n_5818;
wire n_2179;
wire n_5055;
wire n_1547;
wire n_3376;
wire n_4868;
wire n_893;
wire n_3801;
wire n_5267;
wire n_4249;
wire n_1192;
wire n_3564;
wire n_1844;
wire n_1555;
wire n_5548;
wire n_5057;
wire n_3030;
wire n_830;
wire n_5838;
wire n_5725;
wire n_2838;
wire n_5229;
wire n_5325;
wire n_3427;
wire n_852;
wire n_5101;
wire n_2628;
wire n_3071;
wire n_2926;
wire n_1078;
wire n_4273;
wire n_5545;
wire n_2321;
wire n_2019;
wire n_5102;
wire n_3345;
wire n_2074;
wire n_2919;
wire n_4501;
wire n_2129;
wire n_4724;
wire n_945;
wire n_5598;
wire n_4997;
wire n_2399;
wire n_4843;
wire n_1232;
wire n_4696;
wire n_4347;
wire n_5259;
wire n_5819;
wire n_2480;
wire n_3877;
wire n_3929;
wire n_3048;
wire n_1455;
wire n_5279;
wire n_2786;
wire n_5894;
wire n_5239;
wire n_1971;
wire n_1781;
wire n_5354;
wire n_5332;
wire n_2004;
wire n_1106;
wire n_4814;
wire n_953;
wire n_3979;
wire n_3077;
wire n_2873;
wire n_3452;
wire n_3107;
wire n_4956;
wire n_1421;
wire n_3664;
wire n_1936;
wire n_5337;
wire n_5129;
wire n_5420;
wire n_1660;
wire n_5070;
wire n_3047;
wire n_4414;
wire n_1400;
wire n_2625;
wire n_4646;
wire n_2843;
wire n_3760;
wire n_1560;
wire n_4262;
wire n_734;
wire n_1088;
wire n_1894;
wire n_3347;
wire n_5136;
wire n_907;
wire n_5638;
wire n_4110;
wire n_1658;
wire n_4950;
wire n_4729;
wire n_4268;
wire n_1967;
wire n_3999;
wire n_3928;
wire n_2613;
wire n_3535;
wire n_4751;
wire n_2708;
wire n_1648;
wire n_5151;
wire n_1911;
wire n_2011;
wire n_5684;
wire n_5729;
wire n_5680;
wire n_4102;
wire n_1641;
wire n_3871;
wire n_2735;
wire n_4662;
wire n_4671;
wire n_3959;
wire n_2268;
wire n_1367;
wire n_5504;
wire n_1336;
wire n_5522;
wire n_5828;
wire n_4314;
wire n_2080;
wire n_5099;
wire n_1381;
wire n_1699;
wire n_2093;
wire n_4296;
wire n_2770;
wire n_2101;
wire n_4507;
wire n_3484;
wire n_4677;
wire n_792;
wire n_5063;
wire n_1328;
wire n_2917;
wire n_2616;
wire n_5275;
wire n_5306;
wire n_3923;
wire n_3900;
wire n_3488;
wire n_939;
wire n_2811;
wire n_3732;
wire n_2832;
wire n_4226;
wire n_5493;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_3980;
wire n_2998;
wire n_5346;
wire n_4366;
wire n_3446;
wire n_5252;
wire n_5309;
wire n_1895;
wire n_4294;
wire n_4698;
wire n_4445;
wire n_4810;
wire n_3859;
wire n_2692;
wire n_3914;
wire n_4456;
wire n_3397;
wire n_3575;
wire n_2469;
wire n_3927;
wire n_5452;
wire n_3888;
wire n_764;
wire n_5476;
wire n_2764;
wire n_2895;
wire n_733;
wire n_2922;
wire n_3882;
wire n_4856;
wire n_3492;
wire n_4369;
wire n_2068;
wire n_4331;
wire n_4972;
wire n_1290;
wire n_4993;
wire n_5536;
wire n_2072;
wire n_1354;
wire n_4375;
wire n_1701;
wire n_2678;
wire n_3935;
wire n_5130;
wire n_4291;
wire n_5532;
wire n_1726;
wire n_4613;
wire n_2434;
wire n_2878;
wire n_3012;
wire n_3875;
wire n_5609;
wire n_1167;
wire n_2428;
wire n_4717;
wire n_4877;
wire n_3247;
wire n_871;
wire n_2641;
wire n_5658;
wire n_4731;
wire n_3052;
wire n_5046;
wire n_2749;
wire n_3298;
wire n_2254;
wire n_5058;
wire n_1926;
wire n_3273;
wire n_4467;
wire n_1747;
wire n_5667;
wire n_780;
wire n_2624;
wire n_5865;
wire n_2350;
wire n_5042;
wire n_5305;
wire n_4681;
wire n_4072;
wire n_4752;
wire n_4220;
wire n_835;
wire n_928;
wire n_5281;
wire n_2092;
wire n_1654;
wire n_1750;
wire n_1462;
wire n_2514;
wire n_5314;
wire n_1588;
wire n_3942;
wire n_3997;
wire n_2468;
wire n_4381;
wire n_5144;
wire n_2096;
wire n_3968;
wire n_4466;
wire n_4418;
wire n_3434;
wire n_4510;
wire n_5795;
wire n_4473;
wire n_5552;
wire n_5226;
wire n_890;
wire n_5457;
wire n_2812;
wire n_4518;
wire n_1709;
wire n_2393;
wire n_2657;
wire n_5291;
wire n_2921;
wire n_2136;
wire n_2409;
wire n_2252;
wire n_3237;
wire n_949;
wire n_3500;
wire n_3834;
wire n_4589;
wire n_2075;
wire n_2972;
wire n_3542;
wire n_2763;
wire n_2762;
wire n_3192;
wire n_760;
wire n_1546;
wire n_4394;
wire n_2279;
wire n_1296;
wire n_3352;
wire n_3073;
wire n_5343;
wire n_2150;
wire n_1294;
wire n_3696;
wire n_1420;
wire n_4082;
wire n_1779;
wire n_4921;
wire n_1858;
wire n_4329;
wire n_5135;
wire n_3021;
wire n_2558;
wire n_1164;
wire n_4697;
wire n_4288;
wire n_4289;
wire n_3763;
wire n_2712;
wire n_5529;
wire n_3733;
wire n_1487;
wire n_3614;
wire n_874;
wire n_5183;
wire n_2145;
wire n_898;
wire n_4964;
wire n_4228;
wire n_3423;
wire n_1932;
wire n_925;
wire n_1101;
wire n_4636;
wire n_4322;
wire n_3644;
wire n_1249;
wire n_4946;
wire n_2706;
wire n_4767;
wire n_4287;
wire n_2693;
wire n_4137;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_963;
wire n_2767;
wire n_4576;
wire n_4615;
wire n_5787;
wire n_1139;
wire n_3179;
wire n_1018;
wire n_3400;
wire n_1521;
wire n_1366;
wire n_4000;
wire n_5445;
wire n_2897;
wire n_4389;
wire n_3970;
wire n_5342;
wire n_5501;
wire n_4345;
wire n_996;
wire n_1376;
wire n_4664;
wire n_2170;
wire n_4156;
wire n_948;
wire n_977;
wire n_3158;
wire n_1788;
wire n_4873;
wire n_2643;
wire n_5748;
wire n_3782;
wire n_1835;
wire n_3470;
wire n_5076;
wire n_5870;
wire n_4713;
wire n_4098;
wire n_5026;
wire n_4476;
wire n_3700;
wire n_4995;
wire n_3166;
wire n_3104;
wire n_3435;
wire n_842;
wire n_5636;
wire n_2239;
wire n_4310;
wire n_1432;
wire n_5212;
wire n_989;
wire n_2689;
wire n_1473;
wire n_5286;
wire n_2191;
wire n_1246;
wire n_4528;
wire n_5811;
wire n_899;
wire n_1035;
wire n_4914;
wire n_4939;
wire n_1426;
wire n_3418;
wire n_1004;
wire n_1529;
wire n_5530;
wire n_2473;
wire n_5397;
wire n_4634;
wire n_2069;
wire n_2362;
wire n_4096;
wire n_2539;
wire n_2698;
wire n_4123;
wire n_5595;
wire n_3119;
wire n_5427;
wire n_3735;
wire n_2297;
wire n_4379;
wire n_5388;
wire n_4718;
wire n_1448;
wire n_3631;
wire n_5599;
wire n_2445;
wire n_5324;
wire n_2057;
wire n_2103;
wire n_3770;
wire n_2772;
wire n_4440;
wire n_4402;
wire n_927;
wire n_5052;
wire n_4541;
wire n_5009;
wire n_4872;
wire n_929;
wire n_4551;
wire n_2857;
wire n_5326;
wire n_1183;
wire n_4627;
wire n_4079;
wire n_2494;
wire n_5300;
wire n_3342;
wire n_998;
wire n_5035;
wire n_717;
wire n_1383;
wire n_3390;
wire n_3656;
wire n_1424;
wire n_1000;
wire n_3025;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_2482;
wire n_3810;
wire n_4798;
wire n_2532;
wire n_1388;
wire n_3006;
wire n_912;
wire n_5010;
wire n_2296;
wire n_3633;
wire n_5352;
wire n_5089;
wire n_2849;
wire n_1398;
wire n_1201;
wire n_884;
wire n_5394;
wire n_4592;
wire n_1395;
wire n_2199;
wire n_2661;
wire n_731;
wire n_5359;
wire n_1955;
wire n_931;
wire n_1791;
wire n_958;
wire n_5137;
wire n_3331;
wire n_5104;
wire n_1897;
wire n_2064;
wire n_5741;
wire n_2773;
wire n_5405;
wire n_5288;
wire n_3606;
wire n_1310;
wire n_819;
wire n_1334;
wire n_3591;
wire n_2788;
wire n_964;
wire n_4756;
wire n_2797;
wire n_4746;
wire n_3892;
wire n_4970;
wire n_4069;
wire n_2748;
wire n_5194;
wire n_1834;
wire n_2331;
wire n_2292;
wire n_3441;
wire n_3534;
wire n_3964;
wire n_2416;
wire n_1877;
wire n_3944;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_2209;
wire n_3605;
wire n_1602;
wire n_4633;
wire n_3306;
wire n_3026;
wire n_4584;
wire n_3090;
wire n_5232;
wire n_3724;
wire n_4276;
wire n_5116;
wire n_2990;
wire n_3847;
wire n_1773;
wire n_5001;
wire n_2552;
wire n_1053;
wire n_5176;
wire n_4428;
wire n_1533;
wire n_3323;
wire n_2274;
wire n_5761;
wire n_4618;
wire n_4679;
wire n_1745;
wire n_914;
wire n_3479;
wire n_4496;
wire n_4805;
wire n_1679;
wire n_3454;
wire n_2160;
wire n_5760;
wire n_2146;
wire n_2131;
wire n_5472;
wire n_3547;
wire n_5679;
wire n_2575;
wire n_5100;
wire n_4410;
wire n_1933;
wire n_1179;
wire n_3816;
wire n_4807;
wire n_4411;
wire n_3214;
wire n_1243;
wire n_2928;
wire n_5166;
wire n_1917;
wire n_1580;
wire n_2822;
wire n_4180;
wire n_1281;
wire n_3109;
wire n_3354;
wire n_2572;
wire n_1520;
wire n_3126;
wire n_3663;
wire n_2863;
wire n_1419;
wire n_3299;
wire n_5688;
wire n_5740;
wire n_1731;
wire n_5820;
wire n_5648;
wire n_2135;
wire n_5745;
wire n_4707;
wire n_1645;
wire n_1832;
wire n_4676;
wire n_5180;
wire n_858;
wire n_2049;
wire n_5182;
wire n_956;
wire n_5534;
wire n_4880;
wire n_3566;
wire n_2781;
wire n_4126;
wire n_2829;
wire n_1696;
wire n_3845;
wire n_1594;
wire n_1869;
wire n_3804;
wire n_4207;
wire n_5196;
wire n_2016;
wire n_5171;
wire n_4470;
wire n_4813;
wire n_5542;
wire n_1030;
wire n_3901;
wire n_1937;
wire n_1790;
wire n_5261;
wire n_4014;
wire n_4704;
wire n_1744;
wire n_828;
wire n_2142;
wire n_4252;
wire n_4028;
wire n_2448;
wire n_4048;
wire n_4596;
wire n_4444;
wire n_5255;
wire n_3756;
wire n_3406;
wire n_820;
wire n_951;
wire n_952;
wire n_3919;
wire n_2263;
wire n_5185;
wire n_974;
wire n_4952;
wire n_2656;
wire n_5023;
wire n_2375;
wire n_1934;
wire n_5660;
wire n_1434;
wire n_1573;
wire n_3981;
wire n_3973;
wire n_2756;
wire n_5334;
wire n_807;
wire n_4761;
wire n_1275;
wire n_2884;
wire n_1510;
wire n_5783;
wire n_3120;
wire n_5821;
wire n_3797;
wire n_2024;
wire n_1595;
wire n_4770;
wire n_1749;
wire n_3474;
wire n_2549;
wire n_4690;
wire n_1669;
wire n_1024;
wire n_3864;
wire n_5556;
wire n_4932;
wire n_5456;
wire n_2302;
wire n_1667;
wire n_1037;
wire n_5143;
wire n_3592;
wire n_5500;
wire n_4230;
wire n_2637;
wire n_1639;
wire n_3967;
wire n_3195;
wire n_2526;
wire n_4274;
wire n_5215;
wire n_3277;
wire n_2548;
wire n_5386;
wire n_991;
wire n_4189;
wire n_3817;
wire n_1108;
wire n_3659;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_5003;
wire n_4827;
wire n_1601;
wire n_1960;
wire n_2694;
wire n_3648;
wire n_1686;
wire n_3042;
wire n_5094;
wire n_4610;
wire n_4472;
wire n_5433;
wire n_3228;
wire n_3657;
wire n_3081;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_5618;
wire n_1586;
wire n_2264;
wire n_3464;
wire n_3723;
wire n_1190;
wire n_4380;
wire n_4990;
wire n_4996;
wire n_5247;
wire n_4398;
wire n_2498;
wire n_4515;
wire n_5031;
wire n_1891;
wire n_1213;
wire n_2235;
wire n_4193;
wire n_3570;
wire n_5082;
wire n_1673;
wire n_5338;
wire n_3828;
wire n_2392;
wire n_3424;
wire n_4131;
wire n_2298;
wire n_2326;
wire n_1539;
wire n_3594;
wire n_5689;
wire n_1043;
wire n_4090;
wire n_4165;
wire n_2305;
wire n_2120;
wire n_4626;
wire n_4144;
wire n_2964;
wire n_2169;
wire n_3485;
wire n_4077;
wire n_2371;
wire n_1361;
wire n_3262;
wire n_4008;
wire n_3356;
wire n_5221;
wire n_5641;
wire n_1642;
wire n_3210;
wire n_937;
wire n_4689;
wire n_1682;
wire n_4547;
wire n_5731;
wire n_3329;
wire n_3826;
wire n_4905;
wire n_1406;
wire n_4601;
wire n_962;
wire n_3647;
wire n_3681;
wire n_1883;
wire n_4300;
wire n_1288;
wire n_1186;
wire n_4623;
wire n_5007;
wire n_3320;
wire n_2518;
wire n_5883;
wire n_5754;
wire n_3988;
wire n_1720;
wire n_3476;
wire n_4842;
wire n_5629;
wire n_3439;
wire n_4135;
wire n_2688;
wire n_1845;
wire n_1489;
wire n_942;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_1964;
wire n_1920;
wire n_2753;
wire n_1496;
wire n_3292;
wire n_2007;
wire n_2039;
wire n_5434;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_1846;
wire n_3437;
wire n_4111;
wire n_3712;
wire n_4608;
wire n_879;
wire n_2310;
wire n_2506;
wire n_4859;
wire n_2626;
wire n_5880;
wire n_1567;
wire n_4037;
wire n_3562;
wire n_5852;
wire n_2973;
wire n_5218;
wire n_3665;
wire n_3007;
wire n_3528;
wire n_4571;
wire n_3698;
wire n_5358;
wire n_3355;
wire n_2454;
wire n_2114;
wire n_3174;
wire n_5321;
wire n_1066;
wire n_1948;
wire n_4215;
wire n_2154;
wire n_1484;
wire n_5290;
wire n_4185;
wire n_3752;
wire n_2283;
wire n_5145;
wire n_4219;
wire n_1229;
wire n_1373;
wire n_3958;
wire n_3985;
wire n_2427;
wire n_4196;
wire n_1447;
wire n_4774;
wire n_2056;
wire n_5210;
wire n_4242;
wire n_5109;
wire n_3389;
wire n_4232;
wire n_4190;
wire n_4902;
wire n_3000;
wire n_5149;
wire n_5571;
wire n_2680;
wire n_1047;
wire n_3375;
wire n_3899;
wire n_1385;
wire n_3713;
wire n_1931;
wire n_2668;
wire n_1257;
wire n_3197;
wire n_4987;
wire n_2128;
wire n_5512;
wire n_4736;
wire n_2398;
wire n_1725;
wire n_3743;
wire n_834;
wire n_5033;
wire n_2695;
wire n_4035;
wire n_3818;
wire n_3124;
wire n_1741;
wire n_1002;
wire n_1949;
wire n_3759;
wire n_2671;
wire n_4516;
wire n_2715;
wire n_1804;
wire n_2508;
wire n_3511;
wire n_2054;
wire n_1337;
wire n_1477;
wire n_2614;
wire n_4492;
wire n_2833;
wire n_2758;
wire n_5607;
wire n_3694;
wire n_2937;
wire n_4789;
wire n_4376;
wire n_1001;
wire n_2241;
wire n_4708;
wire n_4657;
wire n_1690;
wire n_5341;
wire n_1191;
wire n_1076;
wire n_4512;
wire n_1378;
wire n_855;
wire n_1377;
wire n_4081;
wire n_1542;
wire n_4542;
wire n_4462;
wire n_1716;
wire n_4931;
wire n_4536;
wire n_5562;
wire n_3303;
wire n_978;
wire n_4324;
wire n_1976;
wire n_4382;
wire n_2905;
wire n_1291;
wire n_749;
wire n_1824;
wire n_3954;
wire n_2122;
wire n_5622;
wire n_2140;
wire n_3503;
wire n_3160;
wire n_1065;
wire n_5577;
wire n_1255;
wire n_5124;
wire n_3951;
wire n_823;
wire n_1074;
wire n_3569;
wire n_739;
wire n_3874;
wire n_2528;
wire n_5123;
wire n_4639;
wire n_5413;
wire n_1338;
wire n_1097;
wire n_3027;
wire n_781;
wire n_4083;
wire n_1810;
wire n_1583;
wire n_4480;
wire n_1730;
wire n_2295;
wire n_2746;
wire n_814;
wire n_5779;
wire n_2020;
wire n_1643;
wire n_4171;
wire n_3652;
wire n_4023;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_3617;
wire n_2076;
wire n_3567;
wire n_1598;
wire n_4344;
wire n_2935;
wire n_4705;
wire n_4046;
wire n_3807;
wire n_918;
wire n_1114;
wire n_4027;
wire n_763;
wire n_3154;
wire n_1227;
wire n_2485;
wire n_3898;
wire n_3520;
wire n_4391;
wire n_946;
wire n_1303;
wire n_4095;
wire n_2881;
wire n_1116;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_3551;
wire n_4947;
wire n_3064;
wire n_1780;
wire n_3897;
wire n_1689;
wire n_5591;
wire n_3372;
wire n_1944;
wire n_1347;
wire n_795;
wire n_1221;
wire n_1245;
wire n_3215;
wire n_3853;
wire n_4740;
wire n_4631;
wire n_1561;
wire n_1112;
wire n_5518;
wire n_2081;
wire n_2168;
wire n_5068;
wire n_5847;
wire n_1460;
wire n_911;
wire n_5159;
wire n_2862;
wire n_2615;
wire n_4068;
wire n_4625;
wire n_2474;
wire n_3703;
wire n_2437;
wire n_2444;
wire n_3962;
wire n_2743;
wire n_4766;
wire n_4863;
wire n_2267;
wire n_3035;
wire n_4166;
wire n_1821;
wire n_1058;
wire n_3378;
wire n_3745;
wire n_3362;
wire n_4744;
wire n_4188;
wire n_5357;
wire n_2934;
wire n_3667;
wire n_3523;
wire n_2222;
wire n_3176;
wire n_5541;
wire n_5568;
wire n_2505;
wire n_4817;
wire n_4115;
wire n_2999;
wire n_2014;
wire n_1239;
wire n_3697;
wire n_1584;
wire n_3680;
wire n_5381;
wire n_2408;
wire n_5723;
wire n_3468;
wire n_5045;
wire n_1972;
wire n_4383;
wire n_4491;
wire n_5696;
wire n_4486;
wire n_1816;
wire n_5848;
wire n_3024;
wire n_4612;
wire n_5673;
wire n_5443;
wire n_2531;
wire n_5163;
wire n_4529;
wire n_3361;
wire n_3478;
wire n_3936;
wire n_1349;
wire n_2723;
wire n_5485;
wire n_5823;
wire n_2800;
wire n_3496;
wire n_5473;
wire n_4390;
wire n_3096;
wire n_2651;
wire n_2095;
wire n_3239;
wire n_3161;
wire n_2799;
wire n_5537;
wire n_3902;
wire n_4062;
wire n_3295;
wire n_4396;
wire n_1998;
wire n_3101;
wire n_1574;
wire n_756;
wire n_1981;
wire n_4233;
wire n_1606;
wire n_3374;
wire n_2640;
wire n_1552;
wire n_3288;
wire n_2918;
wire n_4307;
wire n_3992;
wire n_3876;
wire n_3125;
wire n_4293;
wire n_941;
wire n_3552;
wire n_1031;
wire n_849;
wire n_4684;
wire n_3116;
wire n_4091;
wire n_1753;
wire n_5027;
wire n_3095;
wire n_2471;
wire n_4412;
wire n_2807;
wire n_1921;
wire n_3618;
wire n_4580;
wire n_1055;
wire n_2217;
wire n_2197;
wire n_4758;
wire n_5630;
wire n_4781;
wire n_4148;
wire n_2461;
wire n_4057;
wire n_1170;
wire n_5379;
wire n_5335;
wire n_3444;
wire n_1040;
wire n_3059;
wire n_2634;
wire n_1761;
wire n_5424;
wire n_1890;
wire n_3017;
wire n_1805;
wire n_2477;
wire n_5505;
wire n_5868;
wire n_2308;
wire n_2333;
wire n_3001;
wire n_1089;
wire n_3795;
wire n_3852;
wire n_1365;
wire n_4138;
wire n_5289;
wire n_5018;
wire n_3896;
wire n_3815;
wire n_5274;
wire n_3274;
wire n_5401;
wire n_4457;
wire n_4093;
wire n_1616;
wire n_1862;
wire n_4928;
wire n_5769;
wire n_4794;
wire n_722;
wire n_5613;
wire n_5612;
wire n_2223;
wire n_4197;
wire n_4482;
wire n_1621;
wire n_2547;
wire n_2415;
wire n_5073;
wire n_827;
wire n_4834;
wire n_4762;
wire n_5581;
wire n_3113;
wire n_992;
wire n_3813;
wire n_3660;
wire n_3766;
wire n_1613;
wire n_1458;
wire n_5303;
wire n_1027;
wire n_3266;
wire n_3574;
wire n_1189;
wire n_4154;
wire n_4907;
wire n_5077;
wire n_5034;
wire n_726;
wire n_4504;
wire n_3844;
wire n_1237;
wire n_2534;
wire n_4975;
wire n_3741;
wire n_5375;
wire n_2451;
wire n_5370;
wire n_2243;
wire n_4815;
wire n_4898;
wire n_5601;
wire n_5784;
wire n_3443;
wire n_4819;
wire n_1209;
wire n_5248;
wire n_1708;
wire n_805;
wire n_2051;
wire n_4370;
wire n_2359;
wire n_5112;
wire n_1402;
wire n_1691;
wire n_3332;
wire n_4134;
wire n_1238;
wire n_2570;
wire n_4092;
wire n_4645;
wire n_3668;
wire n_2491;
wire n_1264;
wire n_4755;
wire n_4359;
wire n_4960;
wire n_4087;
wire n_1700;
wire n_5635;
wire n_4933;
wire n_5091;
wire n_3487;
wire n_4591;
wire n_5528;
wire n_4302;
wire n_5111;
wire n_3340;
wire n_5227;
wire n_873;
wire n_3946;
wire n_2989;
wire n_5778;
wire n_3395;
wire n_4474;
wire n_5665;
wire n_2509;
wire n_2513;
wire n_3757;
wire n_5363;
wire n_4178;
wire n_5165;
wire n_1704;
wire n_2247;
wire n_1711;
wire n_4884;
wire n_1579;
wire n_3275;
wire n_836;
wire n_3678;
wire n_3440;
wire n_2094;
wire n_1511;
wire n_2356;
wire n_1422;
wire n_1772;
wire n_4692;
wire n_3165;
wire n_1119;
wire n_5788;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2739;
wire n_1735;
wire n_3890;
wire n_1541;
wire n_1300;
wire n_3750;
wire n_1313;
wire n_3607;
wire n_3316;
wire n_2418;
wire n_2864;
wire n_4311;
wire n_1180;
wire n_2703;
wire n_3371;
wire n_4722;
wire n_4606;
wire n_3261;
wire n_4187;
wire n_940;
wire n_2058;
wire n_2660;
wire n_5317;
wire n_1094;
wire n_5430;
wire n_4962;
wire n_4563;
wire n_5056;
wire n_4820;
wire n_2394;
wire n_5540;
wire n_3532;
wire n_5716;
wire n_3948;
wire n_2124;
wire n_4619;
wire n_5762;
wire n_4327;
wire n_1961;
wire n_5211;
wire n_5336;
wire n_3765;
wire n_5447;
wire n_4125;
wire n_5036;
wire n_4221;
wire n_3297;
wire n_976;
wire n_3067;
wire n_2155;
wire n_2686;
wire n_5327;
wire n_2364;
wire n_4392;
wire n_2996;
wire n_3803;
wire n_2085;
wire n_917;
wire n_5014;
wire n_5747;
wire n_3639;
wire n_5192;
wire n_4334;
wire n_3351;
wire n_808;
wire n_5519;
wire n_4047;
wire n_5753;
wire n_3413;
wire n_1193;
wire n_5233;
wire n_3412;
wire n_3791;
wire n_3164;
wire n_4575;
wire n_4320;
wire n_3884;
wire n_5808;
wire n_5436;
wire n_5139;
wire n_757;
wire n_5231;
wire n_2190;
wire n_3438;
wire n_4141;
wire n_5193;
wire n_2850;
wire n_1481;
wire n_1441;
wire n_3373;
wire n_5789;
wire n_2104;
wire n_3883;
wire n_5866;
wire n_3728;
wire n_2925;
wire n_4499;
wire n_5822;
wire n_5195;
wire n_3949;
wire n_5726;
wire n_2792;
wire n_5364;
wire n_3315;
wire n_5533;
wire n_3798;
wire n_788;
wire n_1543;
wire n_1599;
wire n_4257;
wire n_4458;
wire n_2674;
wire n_5103;
wire n_4641;
wire n_4720;
wire n_4893;
wire n_3857;
wire n_1876;
wire n_4107;
wire n_1873;
wire n_3630;
wire n_3518;
wire n_1866;
wire n_2130;
wire n_1413;
wire n_1330;
wire n_3714;
wire n_2228;
wire n_5039;
wire n_2455;
wire n_2876;
wire n_4772;
wire n_3099;
wire n_5198;
wire n_4468;
wire n_5718;
wire n_4161;
wire n_1663;
wire n_4172;
wire n_3403;
wire n_2714;
wire n_2245;
wire n_4961;
wire n_4454;
wire n_1107;
wire n_2457;
wire n_3294;
wire n_4119;
wire n_3686;
wire n_4502;
wire n_2971;
wire n_1713;
wire n_4277;
wire n_4526;
wire n_1265;
wire n_3490;
wire n_4849;
wire n_4319;
wire n_3369;
wire n_5792;
wire n_3581;
wire n_3069;
wire n_2028;
wire n_3715;
wire n_1069;
wire n_3725;
wire n_3933;
wire n_5554;
wire n_1175;
wire n_2311;
wire n_1012;
wire n_3691;
wire n_5553;
wire n_4485;
wire n_4066;
wire n_903;
wire n_4146;
wire n_5711;
wire n_1802;
wire n_1504;
wire n_4340;
wire n_5790;
wire n_3961;
wire n_4855;
wire n_1801;
wire n_2347;
wire n_3917;
wire n_816;
wire n_1188;
wire n_2206;
wire n_4004;
wire n_2967;
wire n_5404;
wire n_2916;
wire n_5739;
wire n_4292;
wire n_2467;
wire n_5549;
wire n_3145;
wire n_1124;
wire n_1624;
wire n_3983;
wire n_4940;
wire n_5444;
wire n_3538;
wire n_3280;
wire n_5757;
wire n_1515;
wire n_961;
wire n_4356;
wire n_3510;
wire n_2824;
wire n_2377;
wire n_950;
wire n_3009;
wire n_5824;
wire n_3719;
wire n_2525;
wire n_4361;
wire n_5488;
wire n_3827;
wire n_891;
wire n_5154;
wire n_2067;
wire n_3889;
wire n_2687;
wire n_1630;
wire n_2887;
wire n_4245;
wire n_4136;
wire n_3526;
wire n_2194;
wire n_2619;
wire n_5329;
wire n_4367;
wire n_5637;
wire n_1987;
wire n_968;
wire n_2271;
wire n_1008;
wire n_2583;
wire n_4560;
wire n_2606;
wire n_4899;
wire n_5728;
wire n_5471;
wire n_1052;
wire n_1033;
wire n_2794;
wire n_5164;
wire n_2391;
wire n_2431;
wire n_5843;
wire n_2078;
wire n_2932;
wire n_1767;
wire n_3431;
wire n_3450;
wire n_4663;
wire n_2893;
wire n_1208;
wire n_5484;
wire n_2954;
wire n_2728;
wire n_1072;
wire n_815;
wire n_3421;
wire n_3183;
wire n_2493;
wire n_4802;
wire n_2705;
wire n_5523;
wire n_1067;
wire n_3405;
wire n_5423;
wire n_1952;
wire n_5074;
wire n_4044;
wire n_3436;
wire n_1026;
wire n_1880;
wire n_3442;
wire n_3366;
wire n_2631;
wire n_3937;
wire n_1293;
wire n_3159;
wire n_4701;
wire n_794;
wire n_727;
wire n_894;
wire n_3240;
wire n_3576;
wire n_1863;
wire n_3385;
wire n_4851;
wire n_3293;
wire n_872;
wire n_3922;
wire n_5204;
wire n_5333;
wire n_847;
wire n_851;
wire n_4991;
wire n_5594;
wire n_2554;
wire n_5422;
wire n_1513;
wire n_1913;
wire n_4934;
wire n_837;
wire n_5087;
wire n_5526;
wire n_5292;
wire n_2517;
wire n_2713;
wire n_5000;
wire n_2765;
wire n_5403;
wire n_2590;
wire n_5551;
wire n_3150;
wire n_2060;
wire n_4479;
wire n_2608;
wire n_4011;
wire n_5131;
wire n_1959;
wire n_3133;
wire n_5257;
wire n_765;
wire n_1492;
wire n_1340;
wire n_4753;
wire n_4688;
wire n_4058;
wire n_2262;
wire n_3611;
wire n_3082;
wire n_4848;
wire n_5059;
wire n_5887;
wire n_843;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_3799;
wire n_2574;
wire n_4475;
wire n_5242;
wire n_5219;
wire n_2675;
wire n_5631;
wire n_3537;
wire n_4443;
wire n_3887;
wire n_1022;
wire n_5854;
wire n_2667;
wire n_5460;
wire n_4587;
wire n_1615;
wire n_4114;
wire n_1474;
wire n_1571;
wire n_2948;
wire n_1577;
wire n_2119;
wire n_947;
wire n_1117;
wire n_1992;
wire n_5686;
wire n_3223;
wire n_3140;
wire n_3185;
wire n_4749;
wire n_2605;
wire n_5155;
wire n_926;
wire n_3654;
wire n_1849;
wire n_2848;
wire n_919;
wire n_1698;
wire n_4100;
wire n_4264;
wire n_3788;
wire n_4891;
wire n_777;
wire n_1299;
wire n_5339;
wire n_3837;
wire n_2718;
wire n_1436;
wire n_1384;
wire n_3325;
wire n_2238;
wire n_4085;
wire n_4464;
wire n_4624;
wire n_4818;
wire n_4659;
wire n_3600;
wire n_5217;
wire n_5465;
wire n_5015;
wire n_4339;
wire n_1178;
wire n_2338;
wire n_3324;
wire n_796;
wire n_1195;
wire n_1811;
wire n_3987;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_1284;
wire n_1604;
wire n_4487;
wire n_4889;
wire n_4866;
wire n_1142;
wire n_1048;
wire n_5721;
wire n_3638;
wire n_4816;
wire n_2110;
wire n_5719;
wire n_1502;
wire n_5773;
wire n_1659;
wire n_5482;
wire n_3393;
wire n_3451;
wire n_1418;
wire n_1250;
wire n_4937;
wire n_5277;
wire n_3615;
wire n_3072;
wire n_3087;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_4222;
wire n_4874;
wire n_4401;
wire n_889;
wire n_2710;
wire n_3142;
wire n_4015;
wire n_1966;
wire n_5793;
wire n_1110;
wire n_4709;
wire n_2213;
wire n_4976;
wire n_2389;
wire n_2132;
wire n_2892;
wire n_4120;
wire n_1564;
wire n_5578;
wire n_4658;
wire n_2860;
wire n_2330;
wire n_5296;
wire n_1457;
wire n_3718;
wire n_5893;
wire n_1787;
wire n_1993;
wire n_2281;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_5742;
wire n_5207;
wire n_3705;
wire n_3211;
wire n_3909;
wire n_5676;
wire n_1220;
wire n_1893;
wire n_2301;
wire n_4665;
wire n_3582;
wire n_4223;
wire n_2387;
wire n_5674;
wire n_3270;
wire n_5539;
wire n_2846;
wire n_5282;
wire n_970;
wire n_2488;
wire n_1980;
wire n_5464;
wire n_2237;
wire n_1060;
wire n_1951;
wire n_4362;
wire n_1252;
wire n_3311;
wire n_3913;
wire n_1223;
wire n_5121;
wire n_1286;
wire n_2115;
wire n_4430;
wire n_3302;
wire n_4348;
wire n_5013;
wire n_1597;
wire n_4489;
wire n_4839;
wire n_2596;
wire n_3163;
wire n_775;
wire n_4404;
wire n_1153;
wire n_5589;
wire n_1531;
wire n_2828;
wire n_2384;
wire n_4261;
wire n_4204;
wire n_759;
wire n_2724;
wire n_2585;
wire n_5628;
wire n_4825;
wire n_2352;
wire n_1625;
wire n_3986;
wire n_5006;
wire n_4513;
wire n_4006;
wire n_2226;
wire n_2801;
wire n_1901;
wire n_3869;
wire n_2556;
wire n_4747;
wire n_1647;
wire n_5251;
wire n_3753;
wire n_2306;
wire n_1614;
wire n_1892;
wire n_3742;
wire n_3683;
wire n_4801;
wire n_3260;
wire n_2550;
wire n_3175;
wire n_3736;
wire n_5475;
wire n_5807;
wire n_4448;
wire n_1096;
wire n_2227;
wire n_5216;
wire n_3284;
wire n_4869;
wire n_2159;
wire n_4386;
wire n_2315;
wire n_1077;
wire n_4132;
wire n_2995;
wire n_5273;
wire n_1437;
wire n_4438;
wire n_4844;
wire n_4836;
wire n_5439;
wire n_4955;
wire n_4149;
wire n_4355;
wire n_3234;
wire n_2276;
wire n_856;
wire n_2803;
wire n_1668;
wire n_2777;
wire n_3202;
wire n_2830;
wire n_3220;
wire n_1129;
wire n_2181;
wire n_2911;
wire n_4655;
wire n_1429;
wire n_5706;
wire n_2826;
wire n_3429;
wire n_2379;
wire n_3554;
wire n_1593;
wire n_1202;
wire n_1635;
wire n_5431;
wire n_4067;
wire n_4357;
wire n_3462;
wire n_2851;
wire n_4374;
wire n_5132;
wire n_2420;
wire n_5627;
wire n_5774;
wire n_3722;
wire n_4400;
wire n_4846;
wire n_5798;
wire n_2984;
wire n_5187;
wire n_5875;
wire n_4024;
wire n_1508;
wire n_5621;
wire n_5608;
wire n_732;
wire n_2983;
wire n_2240;
wire n_2538;
wire n_724;
wire n_3250;
wire n_1042;
wire n_4582;
wire n_1728;
wire n_1871;
wire n_4860;
wire n_845;
wire n_5844;
wire n_3414;
wire n_1549;
wire n_4870;
wire n_768;
wire n_3651;
wire n_2102;
wire n_2563;
wire n_4989;
wire n_3449;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_1187;
wire n_4304;
wire n_4558;
wire n_1403;
wire n_4488;
wire n_3767;
wire n_2544;
wire n_3550;
wire n_4211;
wire n_1206;
wire n_4016;
wire n_5867;
wire n_750;
wire n_5508;
wire n_4656;
wire n_3839;
wire n_2823;
wire n_5597;
wire n_4915;
wire n_4328;
wire n_1057;
wire n_2785;
wire n_5515;
wire n_1997;
wire n_5662;
wire n_2636;
wire n_3131;
wire n_1818;
wire n_3730;
wire n_1298;
wire n_5862;
wire n_4397;
wire n_3399;
wire n_2088;
wire n_1611;
wire n_5050;
wire n_2740;
wire n_746;
wire n_4808;
wire n_5697;
wire n_3416;
wire n_3498;
wire n_5767;
wire n_2401;
wire n_1589;
wire n_4712;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_1740;
wire n_2737;
wire n_3994;
wire n_5462;
wire n_1497;
wire n_3672;
wire n_5318;
wire n_3533;
wire n_1622;
wire n_4725;
wire n_4406;
wire n_1694;
wire n_1535;
wire n_3382;
wire n_3132;
wire n_5498;
wire n_2571;
wire n_3138;
wire n_5053;
wire n_2171;
wire n_2988;
wire n_4908;
wire n_3136;
wire n_1350;
wire n_4192;
wire n_4109;
wire n_4824;
wire n_2037;
wire n_2808;
wire n_4567;
wire n_5150;
wire n_782;
wire n_809;
wire n_3819;
wire n_4778;
wire n_5477;
wire n_1797;
wire n_5175;
wire n_986;
wire n_2050;
wire n_4595;
wire n_2164;
wire n_4174;
wire n_1870;
wire n_1171;
wire n_5179;
wire n_1827;
wire n_4904;
wire n_2187;
wire n_1152;
wire n_3544;
wire n_4150;
wire n_2904;
wire n_5585;
wire n_3105;
wire n_2872;
wire n_3692;
wire n_4616;
wire n_4982;
wire n_1695;
wire n_2046;
wire n_2272;
wire n_2760;
wire n_1979;
wire n_4643;
wire n_2738;
wire n_972;
wire n_5348;
wire n_1332;
wire n_5480;
wire n_4323;
wire n_2346;
wire n_4831;
wire n_936;
wire n_3045;
wire n_3821;
wire n_885;
wire n_2342;
wire n_2167;
wire n_2970;
wire n_3676;
wire n_4896;
wire n_2882;
wire n_3675;
wire n_3666;
wire n_4017;
wire n_4260;
wire n_4916;
wire n_2541;
wire n_2940;
wire n_4739;
wire n_1974;
wire n_4122;
wire n_934;
wire n_4209;
wire n_2768;
wire n_3858;
wire n_1341;
wire n_5284;
wire n_4298;
wire n_2314;
wire n_3502;
wire n_5461;
wire n_3003;
wire n_4128;
wire n_5147;
wire n_4271;
wire n_4644;
wire n_1355;
wire n_2258;
wire n_5503;
wire n_5845;
wire n_804;
wire n_2390;
wire n_959;
wire n_2562;
wire n_4716;
wire n_4312;
wire n_1343;
wire n_1522;
wire n_2734;
wire n_1782;
wire n_5600;
wire n_5755;
wire n_1900;
wire n_5048;
wire n_3246;
wire n_1548;
wire n_3381;
wire n_1155;
wire n_2195;
wire n_3208;
wire n_4944;
wire n_5245;
wire n_4343;
wire n_4715;
wire n_4935;
wire n_4694;
wire n_4672;
wire n_5054;
wire n_2962;
wire n_5448;
wire n_2939;
wire n_5749;
wire n_1672;
wire n_1925;
wire n_4407;
wire n_737;
wire n_3517;
wire n_4045;
wire n_2945;
wire n_4598;
wire n_3061;
wire n_3893;
wire n_3932;
wire n_3469;
wire n_2960;
wire n_3258;
wire n_4524;
wire n_3143;
wire n_4084;
wire n_3149;
wire n_3365;
wire n_3379;
wire n_4850;
wire n_4424;
wire n_3008;
wire n_1751;
wire n_2840;
wire n_3939;
wire n_4776;
wire n_1375;
wire n_3972;
wire n_4153;
wire n_1650;
wire n_3506;
wire n_1962;
wire n_3855;
wire n_1928;
wire n_3091;
wire n_4317;
wire n_4723;
wire n_4269;
wire n_5418;
wire n_4088;
wire n_3398;
wire n_5685;
wire n_2761;
wire n_2793;
wire n_3776;
wire n_3711;
wire n_4235;
wire n_5459;
wire n_1019;
wire n_4143;
wire n_4170;
wire n_729;
wire n_876;
wire n_774;
wire n_3642;
wire n_2845;
wire n_4650;
wire n_4719;
wire n_5173;
wire n_1860;
wire n_5016;
wire n_1904;
wire n_2874;
wire n_1200;
wire n_2588;
wire n_1353;
wire n_1777;
wire n_4967;
wire n_3308;
wire n_1600;
wire n_1113;
wire n_2253;
wire n_2366;
wire n_4912;
wire n_4799;
wire n_2261;
wire n_4423;
wire n_5086;
wire n_5283;
wire n_2210;
wire n_4735;
wire n_3602;
wire n_3300;
wire n_2978;
wire n_2516;
wire n_1050;
wire n_1411;
wire n_5170;
wire n_2827;
wire n_1177;
wire n_3515;
wire n_1150;
wire n_1023;
wire n_2951;
wire n_1118;
wire n_2949;
wire n_1807;
wire n_5028;
wire n_5839;
wire n_1814;
wire n_1631;
wire n_1879;
wire n_3806;
wire n_5514;
wire n_2931;
wire n_2569;
wire n_3866;
wire n_5351;
wire n_4543;
wire n_740;
wire n_4157;
wire n_4229;
wire n_5293;
wire n_3865;
wire n_4073;
wire n_1324;
wire n_3629;
wire n_1435;
wire n_5400;
wire n_3920;
wire n_969;
wire n_4892;
wire n_3255;
wire n_1401;
wire n_1516;
wire n_3846;
wire n_3512;
wire n_5201;
wire n_2029;
wire n_5890;
wire n_4439;
wire n_1394;
wire n_1326;
wire n_4783;
wire n_1379;
wire n_935;
wire n_4910;
wire n_1130;
wire n_3083;
wire n_832;
wire n_3049;
wire n_5389;
wire n_5142;
wire n_3830;
wire n_3679;
wire n_5891;
wire n_3541;
wire n_3117;
wire n_4930;
wire n_5623;
wire n_1283;
wire n_2385;
wire n_4112;
wire n_2149;
wire n_2396;
wire n_4557;
wire n_4917;
wire n_895;
wire n_2450;
wire n_3739;
wire n_4432;
wire n_2284;
wire n_4352;
wire n_4416;
wire n_4593;
wire n_2769;
wire n_4465;
wire n_3622;
wire n_5114;
wire n_4980;
wire n_1392;
wire n_5693;
wire n_4495;
wire n_5117;
wire n_1924;
wire n_5663;
wire n_2463;
wire n_3363;
wire n_1677;
wire n_3721;
wire n_3062;
wire n_2679;
wire n_5024;
wire n_4559;
wire n_838;
wire n_3969;
wire n_3336;
wire n_4160;
wire n_4231;
wire n_2952;
wire n_5647;
wire n_1017;
wire n_4256;
wire n_2779;
wire n_4938;
wire n_5396;
wire n_5203;
wire n_930;
wire n_2620;
wire n_5162;
wire n_1945;
wire n_5426;
wire n_1656;
wire n_5803;
wire n_2112;
wire n_1464;
wire n_2430;
wire n_1414;
wire n_5285;
wire n_2721;
wire n_944;
wire n_4335;
wire n_2034;
wire n_2683;
wire n_5365;
wire n_2744;
wire n_1011;
wire n_4521;
wire n_1566;
wire n_990;
wire n_3204;
wire n_1104;
wire n_5715;
wire n_4920;
wire n_870;
wire n_5395;
wire n_1253;
wire n_5709;
wire n_1693;
wire n_3256;
wire n_3802;
wire n_2118;
wire n_2111;
wire n_2915;
wire n_1148;
wire n_2188;
wire n_1989;
wire n_2802;
wire n_3643;
wire n_2425;
wire n_4265;
wire n_2950;
wire n_5634;
wire n_5672;
wire n_719;
wire n_3060;
wire n_3098;
wire n_4105;
wire n_1851;
wire n_1090;
wire n_4861;
wire n_5799;
wire n_4064;
wire n_4926;
wire n_1518;
wire n_1362;
wire n_3123;
wire n_3380;
wire n_5617;
wire n_1829;
wire n_5266;
wire n_5580;
wire n_1450;
wire n_4828;
wire n_1638;
wire n_3038;
wire n_1789;
wire n_2523;
wire n_5450;
wire n_2413;
wire n_3769;
wire n_1482;
wire n_5310;
wire n_3863;
wire n_3669;
wire n_3130;
wire n_4316;
wire n_5722;
wire n_4640;
wire n_5122;
wire n_5390;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_2805;
wire n_5593;
wire n_4769;
wire n_5764;
wire n_2282;
wire n_4628;
wire n_2047;
wire n_5385;
wire n_1609;
wire n_3344;
wire n_5237;
wire n_2334;
wire n_5133;
wire n_1763;
wire n_5322;
wire n_3989;
wire n_2490;
wire n_4460;
wire n_4108;
wire n_3786;
wire n_3841;
wire n_4254;
wire n_1996;
wire n_2867;
wire n_1442;
wire n_2726;
wire n_4303;
wire n_5853;
wire n_1158;
wire n_2248;
wire n_5011;
wire n_2662;
wire n_3147;
wire n_4909;
wire n_753;
wire n_3925;
wire n_3180;
wire n_2795;
wire n_3472;
wire n_5376;
wire n_5106;
wire n_1479;
wire n_4768;
wire n_1675;
wire n_3717;
wire n_5561;
wire n_5410;
wire n_2215;
wire n_1884;
wire n_2055;
wire n_5156;
wire n_2553;
wire n_2038;
wire n_4447;
wire n_4826;
wire n_3445;
wire n_1833;
wire n_3903;
wire n_1494;
wire n_2325;
wire n_1850;
wire n_5304;
wire n_3854;
wire n_3235;
wire n_5378;
wire n_1417;
wire n_3673;
wire n_4281;
wire n_4648;
wire n_3094;
wire n_965;
wire n_1428;
wire n_1576;
wire n_1856;
wire n_2077;
wire n_5691;
wire n_1059;
wire n_4951;
wire n_4957;
wire n_3079;
wire n_4360;
wire n_4039;
wire n_3070;
wire n_3800;
wire n_4566;
wire n_3263;
wire n_4853;
wire n_1748;
wire n_3504;
wire n_4272;
wire n_2930;
wire n_5615;
wire n_1025;
wire n_3111;
wire n_1885;
wire n_5269;
wire n_3054;
wire n_1538;
wire n_1240;
wire n_5468;
wire n_4730;
wire n_5399;
wire n_1234;
wire n_5262;
wire n_3254;
wire n_3684;
wire n_4670;
wire n_4882;
wire n_4620;
wire n_3152;
wire n_4738;
wire n_3579;
wire n_5421;
wire n_3335;
wire n_4177;
wire n_3783;
wire n_1307;
wire n_3178;
wire n_4127;
wire n_5206;
wire n_1003;
wire n_5713;
wire n_5256;
wire n_2353;
wire n_4099;
wire n_4517;
wire n_4168;
wire n_5188;
wire n_1738;
wire n_4490;
wire n_1575;
wire n_1923;
wire n_2260;
wire n_3952;
wire n_5550;
wire n_3911;
wire n_1688;
wire n_4285;
wire n_3465;
wire n_1743;
wire n_2997;
wire n_1991;
wire n_2386;
wire n_5161;
wire n_5373;
wire n_1724;
wire n_3708;
wire n_4078;
wire n_3046;
wire n_2956;
wire n_5573;
wire n_1553;
wire n_5509;
wire n_5382;
wire n_5659;
wire n_3619;
wire n_1415;
wire n_5881;
wire n_1370;
wire n_1786;
wire n_4198;
wire n_2382;
wire n_3754;
wire n_2291;
wire n_1371;
wire n_2886;
wire n_2974;
wire n_4213;
wire n_2184;
wire n_2982;
wire n_1803;
wire n_4065;
wire n_5863;
wire n_2645;
wire n_3904;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_2630;
wire n_1444;
wire n_1603;
wire n_2470;
wire n_4446;
wire n_1263;
wire n_4417;
wire n_5466;
wire n_4733;
wire n_4764;
wire n_1261;
wire n_3879;
wire n_2286;
wire n_4743;
wire n_2018;
wire n_3080;
wire n_1903;
wire n_1143;
wire n_1874;
wire n_2865;
wire n_2825;
wire n_2013;
wire n_2044;
wire n_3023;
wire n_3232;
wire n_1056;
wire n_758;
wire n_5851;
wire n_2256;
wire n_943;
wire n_4060;
wire n_5110;
wire n_4879;
wire n_5796;
wire n_772;
wire n_2806;
wire n_770;
wire n_3028;
wire n_3662;
wire n_2981;
wire n_3076;
wire n_886;
wire n_3624;
wire n_1345;
wire n_1820;
wire n_4556;
wire n_4117;
wire n_4687;
wire n_2836;
wire n_1404;
wire n_5492;
wire n_2378;
wire n_887;
wire n_2655;
wire n_4600;
wire n_1467;
wire n_4250;
wire n_5829;
wire n_3906;
wire n_4954;
wire n_5191;
wire n_1231;
wire n_2599;
wire n_3963;
wire n_3368;
wire n_2370;
wire n_2612;
wire n_2591;
wire n_4881;
wire n_1815;
wire n_2214;
wire n_4253;
wire n_913;
wire n_5734;
wire n_2593;
wire n_4255;
wire n_867;
wire n_4071;
wire n_3568;
wire n_1230;
wire n_3850;
wire n_5770;
wire n_1333;
wire n_2496;
wire n_5705;
wire n_3313;
wire n_4605;
wire n_3189;
wire n_5525;
wire n_1644;
wire n_2725;
wire n_2277;
wire n_4691;
wire n_1558;
wire n_1732;
wire n_2300;
wire n_3943;
wire n_4305;
wire n_824;
wire n_4297;
wire n_2907;
wire n_5374;
wire n_5575;
wire n_1843;
wire n_5675;
wire n_4227;
wire n_2778;
wire n_1909;
wire n_5020;
wire n_5297;
wire n_1309;
wire n_1123;
wire n_2961;
wire n_916;
wire n_3934;
wire n_4033;
wire n_4415;
wire n_1970;
wire n_2059;
wire n_2669;
wire n_4094;
wire n_4765;
wire n_2546;
wire n_3193;
wire n_2522;
wire n_4364;
wire n_1957;
wire n_4354;
wire n_4732;
wire n_3912;
wire n_3118;
wire n_3720;
wire n_1907;
wire n_2529;
wire n_860;
wire n_1530;
wire n_4745;
wire n_938;
wire n_1302;
wire n_5642;
wire n_4581;
wire n_4377;
wire n_2143;
wire n_905;
wire n_4792;
wire n_1680;
wire n_3842;
wire n_993;
wire n_2031;
wire n_4878;
wire n_1605;
wire n_3514;
wire n_4979;
wire n_1988;
wire n_2654;
wire n_3036;
wire n_5302;
wire n_966;
wire n_4511;
wire n_2908;
wire n_3357;
wire n_5639;
wire n_5781;
wire n_1233;
wire n_3895;
wire n_4520;
wire n_5299;
wire n_3455;
wire n_4118;
wire n_4503;
wire n_2176;
wire n_2459;
wire n_1111;
wire n_3599;
wire n_5543;
wire n_1251;
wire n_5361;
wire n_2711;
wire n_4199;
wire n_5885;
wire n_1912;
wire n_5356;
wire n_4441;
wire n_1982;
wire n_3872;
wire n_3772;
wire n_5458;
wire n_1312;
wire n_5668;
wire n_5038;
wire n_1760;
wire n_5330;
wire n_4585;
wire n_2664;
wire n_1722;
wire n_1664;
wire n_5463;
wire n_3022;
wire n_5489;
wire n_1165;
wire n_5892;
wire n_4773;
wire n_5654;
wire n_2008;
wire n_2192;
wire n_3281;
wire n_2345;
wire n_1386;
wire n_4427;
wire n_5113;
wire n_5479;
wire n_3549;
wire n_5714;
wire n_2804;
wire n_2453;
wire n_2676;
wire n_5510;
wire n_3940;
wire n_4822;
wire n_1214;
wire n_850;
wire n_5692;
wire n_4800;
wire n_1157;
wire n_3453;
wire n_5555;
wire n_3410;
wire n_1752;
wire n_1813;
wire n_3768;
wire n_4958;
wire n_2810;
wire n_4043;
wire n_2319;
wire n_5441;
wire n_825;
wire n_3785;
wire n_2963;
wire n_5366;
wire n_2602;
wire n_3873;
wire n_2980;
wire n_4886;
wire n_1082;
wire n_1317;
wire n_3227;
wire n_2733;
wire n_3289;
wire n_4055;
wire n_2178;
wire n_2644;
wire n_2036;
wire n_3326;
wire n_4200;
wire n_3460;
wire n_2411;
wire n_1796;
wire n_2082;
wire n_3519;
wire n_5078;
wire n_3707;
wire n_3578;
wire n_909;
wire n_4737;
wire n_4925;
wire n_4116;
wire n_5415;
wire n_5419;
wire n_1990;
wire n_3805;
wire n_2943;
wire n_5205;
wire n_1634;
wire n_3252;
wire n_3253;
wire n_1465;
wire n_2622;
wire n_2658;
wire n_2665;
wire n_2133;
wire n_1712;
wire n_4603;
wire n_1523;
wire n_1627;
wire n_5080;
wire n_3128;
wire n_1527;
wire n_5732;
wire n_5372;
wire n_2691;
wire n_840;
wire n_2913;
wire n_4471;
wire n_2230;
wire n_1969;
wire n_2690;
wire n_5208;
wire n_1565;
wire n_1493;
wire n_5690;
wire n_2573;
wire n_2646;
wire n_2535;
wire n_1364;
wire n_3078;
wire n_2436;
wire n_3838;
wire n_5371;
wire n_4651;
wire n_3941;
wire n_3793;
wire n_4854;
wire n_5071;
wire n_3789;
wire n_1514;
wire n_5801;
wire n_3037;
wire n_1646;
wire n_3729;
wire n_4994;
wire n_2537;
wire n_4483;
wire n_5347;
wire n_5168;
wire n_4661;
wire n_1308;
wire n_4988;
wire n_3171;
wire n_3608;
wire n_4540;
wire n_2097;
wire n_3459;
wire n_2853;
wire n_1808;
wire n_3053;
wire n_3358;
wire n_3499;
wire n_4284;
wire n_1005;
wire n_1947;
wire n_3426;
wire n_4971;
wire n_5656;
wire n_1469;
wire n_5125;
wire n_5857;
wire n_2650;
wire n_5652;
wire n_987;
wire n_5499;
wire n_720;
wire n_3229;
wire n_3348;
wire n_1707;
wire n_5228;
wire n_797;
wire n_2933;
wire n_2717;
wire n_1723;
wire n_1878;
wire n_738;
wire n_2012;
wire n_3497;
wire n_5066;
wire n_2842;
wire n_3580;
wire n_2335;
wire n_2307;
wire n_3704;
wire n_5507;
wire n_1809;
wire n_5569;
wire n_4280;
wire n_1181;
wire n_5190;
wire n_3173;
wire n_3677;
wire n_3996;
wire n_1049;
wire n_4097;
wire n_1666;
wire n_803;
wire n_4218;
wire n_5392;
wire n_1717;
wire n_1817;
wire n_2449;
wire n_3880;
wire n_3685;
wire n_2868;
wire n_2231;
wire n_3609;
wire n_1228;
wire n_5455;
wire n_5442;
wire n_4459;
wire n_4545;
wire n_2896;
wire n_3019;
wire n_2639;
wire n_3471;
wire n_5511;
wire n_2898;
wire n_5295;
wire n_2368;
wire n_4175;
wire n_5490;
wire n_3200;
wire n_4771;
wire n_3259;
wire n_2524;
wire n_3167;
wire n_2460;
wire n_5836;
wire n_3867;
wire n_3593;
wire n_4455;
wire n_1073;
wire n_4514;
wire n_5834;
wire n_3191;
wire n_5584;
wire n_4140;
wire n_2481;
wire n_3561;
wire n_4806;
wire n_2682;
wire n_3032;
wire n_5160;
wire n_2877;
wire n_5098;
wire n_1021;
wire n_811;
wire n_1207;
wire n_5707;
wire n_5140;
wire n_4992;
wire n_5197;
wire n_5497;
wire n_880;
wire n_3505;
wire n_3540;
wire n_3577;
wire n_2432;
wire n_1478;
wire n_4796;
wire n_3598;
wire n_4442;
wire n_2581;
wire n_1363;
wire n_3641;
wire n_3777;
wire n_4203;
wire n_767;
wire n_1837;
wire n_2218;
wire n_4533;
wire n_831;
wire n_5481;
wire n_3590;
wire n_2435;
wire n_5344;
wire n_954;
wire n_4419;
wire n_5308;
wire n_1410;
wire n_5184;
wire n_5794;
wire n_1382;
wire n_5408;
wire n_1736;
wire n_4053;
wire n_1483;
wire n_3848;
wire n_1372;
wire n_3327;
wire n_1719;
wire n_2701;
wire n_2511;
wire n_4167;
wire n_1427;
wire n_2745;
wire n_1080;
wire n_5271;
wire n_2323;
wire n_2784;
wire n_5494;
wire n_5234;
wire n_4431;
wire n_2421;
wire n_1136;
wire n_4387;
wire n_2618;
wire n_3265;
wire n_2464;
wire n_1125;
wire n_3755;
wire n_4042;
wire n_5128;
wire n_2224;
wire n_2329;
wire n_1092;
wire n_5467;
wire n_4299;
wire n_4890;
wire n_1784;
wire n_3571;
wire n_1775;
wire n_2410;
wire n_1093;
wire n_1783;
wire n_2929;
wire n_4176;
wire n_5827;
wire n_5199;
wire n_3407;
wire n_5313;
wire n_1185;
wire n_3856;
wire n_4236;
wire n_3425;
wire n_3894;
wire n_3127;
wire n_1831;
wire n_2621;
wire n_3623;
wire n_5312;
wire n_5079;
wire n_1453;
wire n_2502;
wire n_3646;
wire n_5513;
wire n_5614;
wire n_4830;
wire n_4706;
wire n_1315;
wire n_5225;
wire n_4570;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_3188;
wire n_1459;
wire n_2462;
wire n_3243;
wire n_1135;
wire n_2889;
wire n_4034;
wire n_4056;
wire n_4622;
wire n_3960;
wire n_1470;
wire n_4887;
wire n_2732;
wire n_4693;
wire n_4206;
wire n_2249;
wire n_1091;
wire n_2000;
wire n_3862;
wire n_4267;
wire n_5835;
wire n_2270;
wire n_1425;
wire n_5049;
wire n_983;
wire n_5846;
wire n_906;
wire n_1390;
wire n_2289;
wire n_1733;
wire n_2955;
wire n_5592;
wire n_2158;
wire n_4609;
wire n_1855;
wire n_3051;
wire n_3367;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_2859;
wire n_2202;
wire n_1331;
wire n_736;
wire n_5278;
wire n_3314;
wire n_3525;
wire n_2100;
wire n_5157;
wire n_3016;
wire n_4754;
wire n_2993;
wire n_4647;
wire n_1134;
wire n_3688;
wire n_4003;
wire n_5708;
wire n_1995;
wire n_3751;
wire n_5223;
wire n_4894;
wire n_5474;
wire n_4113;
wire n_1889;
wire n_4760;
wire n_5649;
wire n_1905;
wire n_3466;
wire n_762;
wire n_5704;
wire n_4983;
wire n_1778;
wire n_5287;
wire n_1079;
wire n_2139;
wire n_5083;
wire n_4509;
wire n_2875;
wire n_1103;
wire n_3907;
wire n_3338;
wire n_4217;
wire n_4906;
wire n_2219;
wire n_1203;
wire n_3636;
wire n_2327;
wire n_999;
wire n_5516;
wire n_1254;
wire n_2841;
wire n_4897;
wire n_3539;
wire n_3291;
wire n_4399;
wire n_2304;
wire n_2487;
wire n_5698;
wire n_3276;
wire n_2597;
wire n_3194;
wire n_5084;
wire n_5771;
wire n_3572;
wire n_3886;
wire n_4710;
wire n_4420;
wire n_892;
wire n_3637;
wire n_4574;
wire n_1468;
wire n_2855;
wire n_1859;
wire n_2156;
wire n_1718;
wire n_5174;
wire n_4234;
wire n_5538;
wire n_4101;
wire n_3548;
wire n_5017;
wire n_1768;
wire n_3974;
wire n_1847;
wire n_3634;
wire n_1397;
wire n_3236;
wire n_901;
wire n_5096;
wire n_2755;
wire n_3141;
wire n_923;
wire n_1841;
wire n_4660;
wire n_5241;
wire n_1623;
wire n_1015;
wire n_3112;
wire n_4797;
wire n_3108;
wire n_4270;
wire n_5428;
wire n_4151;
wire n_4945;
wire n_3417;
wire n_5677;
wire n_4124;
wire n_5570;
wire n_785;
wire n_5153;
wire n_4611;
wire n_5435;
wire n_2337;
wire n_1356;
wire n_3213;
wire n_4333;
wire n_3820;
wire n_5200;
wire n_2607;
wire n_2890;
wire n_1168;
wire n_5115;
wire n_1943;
wire n_5566;
wire n_3249;
wire n_1320;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_2499;
wire n_4152;
wire n_5487;
wire n_5486;
wire n_1596;
wire n_5092;
wire n_5244;
wire n_1734;
wire n_3172;
wire n_4832;
wire n_2902;
wire n_5889;
wire n_3217;
wire n_1983;
wire n_5391;
wire n_1938;
wire n_2472;
wire n_3394;
wire n_1715;
wire n_3536;
wire n_1443;
wire n_1272;
wire n_2894;
wire n_3957;
wire n_3710;
wire n_4195;
wire n_5849;
wire n_4554;
wire n_3040;
wire n_3279;
wire n_5240;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_1692;
wire n_1084;
wire n_1864;
wire n_2006;
wire n_3402;
wire n_3501;
wire n_3475;
wire n_1705;
wire n_3905;
wire n_4680;
wire n_3013;
wire n_921;
wire n_2789;
wire n_5152;
wire n_5265;
wire n_2257;
wire n_4927;
wire n_5574;
wire n_4258;
wire n_1828;
wire n_2699;
wire n_2200;
wire n_1940;
wire n_4548;
wire n_4862;
wire n_1405;
wire n_2376;
wire n_5469;
wire n_3878;
wire n_2670;
wire n_2700;
wire n_1041;
wire n_5804;
wire n_3134;
wire n_1569;
wire n_3115;
wire n_1062;
wire n_896;
wire n_4553;
wire n_3278;
wire n_2084;
wire n_4875;
wire n_5682;
wire n_5387;
wire n_5557;
wire n_2458;
wire n_1222;
wire n_3050;
wire n_2673;
wire n_2456;
wire n_2527;
wire n_2635;
wire n_3307;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_2871;
wire n_4321;
wire n_4183;
wire n_5681;
wire n_1271;
wire n_4901;
wire n_1545;
wire n_4145;
wire n_3121;
wire n_4821;
wire n_1640;
wire n_4040;
wire n_2406;
wire n_806;
wire n_2141;
wire n_5316;
wire n_5703;
wire n_833;
wire n_3930;
wire n_4943;
wire n_799;
wire n_3044;
wire n_4757;
wire n_2196;
wire n_2629;
wire n_2809;
wire n_787;
wire n_2172;
wire n_4682;
wire n_5564;
wire n_5620;
wire n_4530;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_4942;
wire n_1086;
wire n_5406;
wire n_2125;
wire n_2561;
wire n_4604;
wire n_1906;
wire n_3305;
wire n_2992;
wire n_5724;
wire n_1241;
wire n_3157;
wire n_4841;
wire n_1758;
wire n_3221;
wire n_3267;
wire n_2422;
wire n_1914;
wire n_1318;
wire n_5806;
wire n_4338;
wire n_3457;
wire n_3762;
wire n_5738;
wire n_3005;
wire n_3151;
wire n_3411;
wire n_4840;
wire n_1029;
wire n_4519;
wire n_3779;
wire n_2388;
wire n_5355;
wire n_3984;
wire n_5320;
wire n_5353;
wire n_1706;
wire n_5186;
wire n_5710;
wire n_1498;
wire n_2417;
wire n_1210;
wire n_5093;
wire n_1556;
wire n_4052;
wire n_3558;
wire n_1984;
wire n_2236;
wire n_5438;
wire n_4326;
wire n_1269;
wire n_2083;
wire n_2834;
wire n_5517;
wire n_3207;
wire n_5605;
wire n_2441;
wire n_3401;
wire n_3242;
wire n_3613;
wire n_4726;
wire n_1045;
wire n_786;
wire n_1559;
wire n_1872;
wire n_5040;
wire n_1325;
wire n_3761;
wire n_4315;
wire n_2923;
wire n_2888;
wire n_1727;
wire n_4301;
wire n_3744;
wire n_4788;
wire n_2041;
wire n_1360;
wire n_3814;
wire n_3781;
wire n_1908;
wire n_2484;
wire n_2126;
wire n_3843;
wire n_1098;
wire n_5746;
wire n_2045;
wire n_817;
wire n_5451;
wire n_3687;
wire n_2216;
wire n_5402;
wire n_3543;
wire n_3621;
wire n_2903;
wire n_3216;
wire n_3808;
wire n_4365;
wire n_1882;
wire n_3726;
wire n_1007;
wire n_1929;
wire n_2369;
wire n_1592;
wire n_2719;
wire n_3758;
wire n_5417;
wire n_2587;
wire n_3199;
wire n_3339;
wire n_4923;
wire n_2400;
wire n_5864;
wire n_1953;
wire n_4741;
wire n_3343;
wire n_2752;
wire n_4885;
wire n_751;
wire n_5432;
wire n_1399;
wire n_4550;
wire n_4652;
wire n_2358;
wire n_5453;
wire n_3658;
wire n_4900;
wire n_2163;
wire n_2186;
wire n_2815;
wire n_3034;
wire n_4408;
wire n_4577;
wire n_4748;
wire n_5842;
wire n_5814;
wire n_2814;
wire n_5253;
wire n_5209;
wire n_789;
wire n_3231;
wire n_4212;
wire n_2979;
wire n_5699;
wire n_5531;
wire n_5765;
wire n_2953;
wire n_4295;
wire n_2946;
wire n_2500;
wire n_3430;
wire n_2269;
wire n_1729;
wire n_5777;
wire n_4225;
wire n_747;
wire n_2565;
wire n_5495;
wire n_1389;
wire n_3583;
wire n_3860;
wire n_3851;
wire n_5655;
wire n_5064;
wire n_5610;
wire n_3015;
wire n_2175;
wire n_2182;
wire n_4009;
wire n_1848;
wire n_5002;
wire n_5759;
wire n_1506;
wire n_3473;
wire n_1652;
wire n_1994;
wire n_957;
wire n_2566;
wire n_744;
wire n_971;
wire n_2702;
wire n_3241;
wire n_2906;
wire n_4342;
wire n_4568;
wire n_1205;
wire n_5559;
wire n_1258;
wire n_2438;
wire n_2914;
wire n_5786;
wire n_3100;
wire n_2180;
wire n_2858;
wire n_5377;
wire n_3573;
wire n_1016;
wire n_4106;
wire n_5737;
wire n_1501;
wire n_3604;
wire n_4373;
wire n_4711;
wire n_3068;
wire n_2685;
wire n_1083;
wire n_5768;
wire n_3553;
wire n_2275;
wire n_2465;
wire n_2568;
wire n_2022;
wire n_3811;
wire n_910;
wire n_1721;
wire n_3494;
wire n_1737;
wire n_3486;
wire n_4086;
wire n_752;
wire n_908;
wire n_1028;
wire n_2106;
wire n_2265;
wire n_5350;
wire n_5470;
wire n_2032;
wire n_4812;
wire n_4409;
wire n_5872;
wire n_5858;
wire n_4629;
wire n_4638;
wire n_1973;
wire n_3181;
wire n_5700;
wire n_1500;
wire n_3699;
wire n_854;
wire n_4913;
wire n_2312;
wire n_5874;
wire n_904;
wire n_1266;
wire n_2242;
wire n_3328;
wire n_3868;
wire n_1276;
wire n_4266;
wire n_2466;
wire n_2530;
wire n_5873;
wire n_1085;
wire n_2042;
wire n_771;
wire n_924;
wire n_1582;
wire n_5588;
wire n_2318;
wire n_3286;
wire n_4012;
wire n_1149;
wire n_3170;
wire n_3645;
wire n_5075;
wire n_3682;
wire n_3304;
wire n_2592;
wire n_4968;
wire n_3771;
wire n_2666;
wire n_1585;
wire n_1799;
wire n_2564;
wire n_5085;
wire n_5736;
wire n_4259;
wire n_2433;
wire n_829;
wire n_2035;
wire n_3422;
wire n_4572;
wire n_859;
wire n_3086;
wire n_2033;
wire n_4104;
wire n_4845;
wire n_1770;
wire n_878;
wire n_5120;
wire n_3285;
wire n_4208;
wire n_981;
wire n_4089;
wire n_5478;
wire n_1144;
wire n_2071;
wire n_3219;
wire n_3702;
wire n_2233;
wire n_4779;
wire n_3233;
wire n_4599;
wire n_997;
wire n_4437;
wire n_5222;
wire n_3310;
wire n_1306;
wire n_3264;
wire n_2010;
wire n_1198;
wire n_4061;
wire n_2174;
wire n_3881;
wire n_4508;
wire n_4727;
wire n_4594;
wire n_2426;
wire n_2478;
wire n_1133;
wire n_4429;
wire n_4642;
wire n_4051;
wire n_1051;
wire n_4865;
wire n_1039;
wire n_2043;
wire n_1480;
wire n_5832;
wire n_3206;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_4562;
wire n_3383;
wire n_4903;
wire n_3709;
wire n_3738;
wire n_4186;
wire n_5812;
wire n_2540;
wire n_973;
wire n_5743;
wire n_3610;
wire n_4998;
wire n_3330;
wire n_2065;
wire n_2879;
wire n_967;
wire n_4522;
wire n_2001;
wire n_4341;
wire n_1629;
wire n_5368;
wire n_4263;
wire n_1260;
wire n_1819;
wire n_3555;
wire n_915;
wire n_812;
wire n_1131;
wire n_3155;
wire n_1006;
wire n_3110;
wire n_1632;
wire n_1888;
wire n_1311;
wire n_4780;
wire n_2697;
wire n_3908;
wire n_4973;
wire n_3467;
wire n_1887;
wire n_1587;
wire n_3916;
wire n_3527;
wire n_4803;
wire n_2512;
wire n_3950;
wire n_1242;
wire n_2086;
wire n_2927;
wire n_4750;
wire n_3039;
wire n_1226;
wire n_3740;
wire n_2166;
wire n_2899;
wire n_3186;
wire n_1322;
wire n_1958;
wire n_1197;
wire n_3065;
wire n_2632;
wire n_4984;
wire n_2579;
wire n_2105;
wire n_1423;
wire n_3387;
wire n_5782;
wire n_3420;
wire n_5041;
wire n_1915;
wire n_4275;
wire n_4283;
wire n_4959;
wire n_900;
wire n_4426;
wire n_2912;
wire n_2659;
wire n_4425;
wire n_3409;
wire n_4449;
wire n_2116;
wire n_2320;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_3002;
wire n_1612;
wire n_4809;
wire n_1199;
wire n_3392;
wire n_3773;
wire n_2003;
wire n_1038;
wire n_1581;
wire n_3301;
wire n_1357;
wire n_4241;
wire n_1853;
wire n_798;
wire n_2324;
wire n_5563;
wire n_1348;
wire n_2977;
wire n_1739;
wire n_5840;
wire n_1380;
wire n_2847;
wire n_2557;
wire n_1009;
wire n_2405;
wire n_4050;
wire n_1160;
wire n_883;
wire n_2647;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_5717;
wire n_2521;
wire n_1099;
wire n_4578;
wire n_2211;
wire n_4777;
wire n_5720;
wire n_2672;
wire n_4702;
wire n_2299;
wire n_4179;
wire n_4895;
wire n_5871;
wire n_1285;
wire n_1985;
wire n_1172;
wire n_4026;
wire n_4531;
wire n_3282;
wire n_1590;
wire n_3626;
wire n_1532;
wire n_2313;
wire n_5072;
wire n_3106;
wire n_1140;
wire n_1670;
wire n_2344;
wire n_2365;
wire n_4666;
wire n_3031;
wire n_4029;
wire n_2447;
wire n_4617;
wire n_2340;
wire n_4010;
wire n_1649;
wire n_4555;
wire n_5882;
wire n_5650;
wire n_4969;
wire n_5105;
wire n_1572;
wire n_4308;
wire n_5021;
wire n_3463;
wire n_5263;
wire n_2510;
wire n_1954;
wire n_822;
wire n_2791;
wire n_4325;
wire n_3251;
wire n_4602;
wire n_5044;
wire n_5134;
wire n_2212;
wire n_3063;
wire n_2729;
wire n_1163;
wire n_2582;
wire n_1798;
wire n_1550;
wire n_3998;
wire n_1591;
wire n_3632;
wire n_3122;
wire n_5567;
wire n_1344;
wire n_2730;
wire n_2495;
wire n_5249;
wire n_2090;
wire n_2603;
wire n_3829;
wire n_4164;
wire n_2173;
wire n_5625;
wire n_1471;
wire n_4919;
wire n_3737;
wire n_3655;
wire n_3825;
wire n_3225;
wire n_2880;
wire n_2108;
wire n_5158;
wire n_1211;
wire n_5022;
wire n_5670;
wire n_1280;
wire n_3296;
wire n_5276;
wire n_1445;
wire n_2551;
wire n_1526;
wire n_5047;
wire n_2985;
wire n_1978;
wire n_3792;
wire n_4202;
wire n_1446;
wire n_3938;
wire n_4791;
wire n_3507;
wire n_5879;
wire n_4403;
wire n_5238;
wire n_5855;
wire n_3269;
wire n_3531;
wire n_1054;
wire n_1956;
wire n_4139;
wire n_4549;
wire n_1986;
wire n_2397;
wire n_3931;
wire n_4349;
wire n_5141;
wire n_2113;
wire n_1918;
wire n_3603;
wire n_5429;
wire n_813;
wire n_3822;
wire n_4163;
wire n_818;
wire n_5535;
wire n_3812;
wire n_3910;
wire n_2633;
wire n_2207;
wire n_4948;
wire n_5268;
wire n_2696;
wire n_3482;
wire n_4080;
wire n_2198;
wire n_3319;
wire n_2073;
wire n_2273;
wire n_3748;
wire n_3272;
wire n_4941;
wire n_5506;
wire n_5298;
wire n_3396;
wire n_4393;
wire n_1162;
wire n_4372;
wire n_821;
wire n_1068;
wire n_982;
wire n_5640;
wire n_932;
wire n_2831;
wire n_4318;
wire n_4158;
wire n_3317;
wire n_3978;
wire n_5560;
wire n_2123;
wire n_1697;
wire n_979;
wire n_4074;
wire n_3716;
wire n_4795;
wire n_5544;
wire n_4918;
wire n_3824;
wire n_5067;
wire n_5744;
wire n_4013;
wire n_5384;
wire n_4544;
wire n_3248;
wire n_5841;
wire n_2941;
wire n_1278;
wire n_5108;
wire n_4032;
wire n_1064;
wire n_1396;
wire n_2355;
wire n_4147;
wire n_4477;
wire n_3168;
wire n_2751;
wire n_4337;
wire n_4130;
wire n_2009;
wire n_1793;
wire n_3601;
wire n_5611;
wire n_3092;
wire n_1289;
wire n_3055;
wire n_3966;
wire n_2866;
wire n_4742;
wire n_3734;
wire n_1014;
wire n_1703;
wire n_2580;
wire n_882;
wire n_3649;
wire n_2821;
wire n_1875;
wire n_1865;
wire n_5701;
wire n_3746;
wire n_3384;
wire n_1950;
wire n_1563;
wire n_3419;
wire n_1297;
wire n_1662;
wire n_4478;
wire n_1359;
wire n_2818;
wire n_5367;
wire n_3794;
wire n_3921;
wire n_922;
wire n_1335;
wire n_1927;
wire n_4838;
wire n_5202;
wire n_4965;
wire n_3346;
wire n_1896;
wire n_2965;
wire n_3058;
wire n_3861;
wire n_1540;
wire n_1977;
wire n_3891;
wire n_2193;
wire n_4523;
wire n_1655;
wire n_1886;
wire n_4371;
wire n_2994;
wire n_5502;
wire n_3428;
wire n_3153;
wire n_4552;
wire n_3689;
wire n_877;
wire n_5850;
wire n_4673;
wire n_2519;
wire n_728;
wire n_3415;
wire n_1063;
wire n_4607;
wire n_4041;
wire n_2947;
wire n_3918;
wire n_5876;
wire n_5521;
wire n_1965;
wire n_4837;
wire n_2476;
wire n_4169;
wire n_3271;
wire n_5088;
wire n_4248;
wire n_2976;
wire n_2152;
wire n_2652;
wire n_1825;
wire n_1757;
wire n_1792;
wire n_5856;
wire n_1412;
wire n_2497;
wire n_3809;
wire n_3139;
wire n_4070;
wire n_3545;
wire n_3885;
wire n_1369;
wire n_881;
wire n_3993;
wire n_4685;
wire n_4031;
wire n_5837;
wire n_4675;
wire n_2663;
wire n_5825;
wire n_4018;
wire n_5491;
wire n_2987;
wire n_2938;
wire n_3780;
wire n_5496;
wire n_5802;
wire n_3337;
wire n_4002;
wire n_3209;
wire n_5178;
wire n_1044;
wire n_2165;
wire n_5547;
wire n_1391;
wire n_2750;
wire n_2775;
wire n_1295;
wire n_3477;
wire n_2349;
wire n_5596;
wire n_2684;
wire n_3146;
wire n_1495;
wire n_1438;
wire n_3953;
wire n_4588;
wire n_1100;
wire n_4653;
wire n_4435;
wire n_5604;
wire n_1756;
wire n_1128;
wire n_5411;
wire n_4019;
wire n_1071;
wire n_1968;
wire n_4728;
wire n_4999;
wire n_4385;
wire n_4922;
wire n_865;
wire n_3616;
wire n_5815;
wire n_4191;
wire n_5695;
wire n_2870;
wire n_2151;
wire n_1839;
wire n_2341;
wire n_1765;
wire n_3727;
wire n_5235;
wire n_2707;
wire n_826;
wire n_4350;
wire n_3747;
wire n_1714;
wire n_718;
wire n_5331;
wire n_4330;
wire n_5311;
wire n_2089;
wire n_3522;
wire n_2747;
wire n_3924;
wire n_791;
wire n_4621;
wire n_4216;
wire n_5797;
wire n_4240;
wire n_3491;
wire n_5572;
wire n_1488;
wire n_2148;
wire n_4162;
wire n_5565;
wire n_2339;
wire n_2861;
wire n_1999;
wire n_2731;
wire n_5520;
wire n_3353;
wire n_3018;
wire n_3975;
wire n_5800;
wire n_1838;
wire n_2638;
wire n_4785;
wire n_4683;
wire n_1776;
wire n_1766;
wire n_2002;
wire n_2138;
wire n_4021;
wire n_2414;
wire n_3014;
wire n_1771;
wire n_2316;
wire n_4103;
wire n_5060;
wire n_3148;
wire n_4022;
wire n_4986;
wire n_5888;
wire n_5669;
wire n_5772;
wire n_2208;
wire n_4775;
wire n_5884;
wire n_4864;
wire n_5758;
wire n_4674;
wire n_4481;
wire n_1304;
wire n_3775;
wire n_4669;
wire n_2134;
wire n_1176;
wire n_5603;
wire n_1431;
wire n_3312;
wire n_3835;
wire n_4286;
wire n_5763;
wire n_2958;
wire n_3731;
wire n_1822;
wire n_2936;
wire n_3224;
wire n_2489;
wire n_1087;
wire n_5751;
wire n_2771;
wire n_3020;
wire n_5264;
wire n_4525;
wire n_1505;
wire n_5712;
wire n_3557;
wire n_2610;
wire n_3129;
wire n_3620;
wire n_3832;
wire n_2520;
wire n_4484;
wire n_3693;
wire n_4497;
wire n_1568;
wire n_2372;
wire n_1490;
wire n_2251;
wire n_3674;
wire n_2959;
wire n_2501;
wire n_3203;
wire n_5694;
wire n_4871;
wire n_1070;
wire n_2403;
wire n_2837;
wire n_4700;
wire n_4883;
wire n_1665;
wire n_4306;
wire n_4224;
wire n_2127;
wire n_3341;
wire n_4453;
wire n_3559;
wire n_5449;
wire n_4005;
wire n_3546;
wire n_1358;
wire n_3661;
wire n_4564;
wire n_5146;
wire n_3056;
wire n_745;
wire n_2424;
wire n_3201;
wire n_3447;
wire n_3971;
wire n_1475;
wire n_1774;
wire n_2354;
wire n_3103;
wire n_4573;
wire n_5398;
wire n_5860;
wire n_2589;
wire n_4535;
wire n_755;
wire n_2442;
wire n_3627;
wire n_3480;
wire n_1368;
wire n_1137;
wire n_3612;
wire n_4695;
wire n_2545;
wire n_3509;
wire n_4368;
wire n_2966;
wire n_2294;
wire n_1942;
wire n_1314;
wire n_3196;
wire n_864;
wire n_5319;
wire n_2504;
wire n_2623;
wire n_1440;
wire n_5270;
wire n_2063;
wire n_1534;
wire n_5005;
wire n_1339;
wire n_2475;
wire n_5181;
wire n_723;
wire n_3144;
wire n_3244;
wire n_1141;
wire n_1268;
wire n_3287;
wire n_3322;
wire n_1755;
wire n_5043;
wire n_2025;
wire n_2357;
wire n_5583;
wire n_4654;
wire n_3640;
wire n_1159;
wire n_995;
wire n_3481;
wire n_2250;
wire n_3033;
wire n_5775;
wire n_2374;
wire n_1681;
wire n_4597;
wire n_3364;
wire n_3226;
wire n_2780;
wire n_4020;
wire n_5220;
wire n_1618;
wire n_4867;
wire n_5061;
wire n_1653;
wire n_4063;
wire n_4237;
wire n_2601;
wire n_5029;
wire n_5127;
wire n_2920;
wire n_773;
wire n_920;
wire n_1374;
wire n_2648;
wire n_3212;
wire n_1169;
wire n_1617;
wire n_3370;
wire n_3386;
wire n_4721;
wire n_3093;
wire n_848;
wire n_4247;
wire n_3169;
wire n_3205;
wire n_1881;
wire n_1267;
wire n_1806;
wire n_2023;
wire n_2204;
wire n_2720;
wire n_4614;
wire n_3360;
wire n_2087;
wire n_1636;
wire n_3956;
wire n_4001;
wire n_1323;
wire n_2627;
wire n_4422;
wire n_960;
wire n_778;
wire n_3004;
wire n_3870;
wire n_5177;
wire n_5483;
wire n_3625;
wire n_1764;
wire n_4632;
wire n_1610;
wire n_3084;
wire n_5785;
wire n_2343;
wire n_793;
wire n_4546;
wire n_4583;
wire n_4963;
wire n_3749;
wire n_2942;
wire n_4966;
wire n_5780;
wire n_4714;
wire n_5037;
wire n_2515;
wire n_1551;
wire n_4847;
wire n_4054;
wire n_2555;
wire n_3586;
wire n_3653;
wire n_2201;
wire n_725;
wire n_3349;
wire n_4668;
wire n_5213;
wire n_4635;
wire n_994;
wire n_5735;
wire n_2278;
wire n_1020;
wire n_1273;
wire n_4214;
wire n_3448;
wire n_2924;
wire n_1036;
wire n_3595;
wire n_1138;
wire n_5752;
wire n_1661;
wire n_5360;
wire n_3991;
wire n_3516;
wire n_3926;
wire n_1095;
wire n_1270;
wire n_4405;
wire n_4413;
wire n_1852;
wire n_4036;
wire n_4759;
wire n_2153;
wire n_3670;
wire n_2381;
wire n_2052;
wire n_4667;
wire n_5081;
wire n_4182;
wire n_3230;
wire n_1279;
wire n_1115;
wire n_1499;
wire n_1409;
wire n_5877;
wire n_5189;
wire n_1503;
wire n_2819;
wire n_3041;
wire n_4637;
wire n_2423;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_5869;
wire n_2439;
wire n_2404;
wire n_1182;
wire n_3635;
wire n_5118;
wire n_4155;
wire n_4238;
wire n_3011;
wire n_2061;
wire n_2757;
wire n_4977;
wire n_5632;
wire n_5582;
wire n_5425;
wire n_5886;
wire n_1216;
wire n_2716;
wire n_2452;
wire n_3650;
wire n_5446;
wire n_3010;
wire n_3043;
wire n_5224;
wire n_4590;
wire n_2543;
wire n_5090;
wire n_3137;
wire n_2486;
wire n_3560;
wire n_3177;
wire n_4929;
wire n_5678;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_3238;
wire n_3529;
wire n_4835;
wire n_2232;
wire n_4038;
wire n_2790;
wire n_4565;
wire n_5414;
wire n_4159;
wire n_3784;
wire n_5437;
wire n_4586;
wire n_1608;
wire n_2373;
wire n_1472;
wire n_3628;
wire n_5454;
wire n_800;
wire n_4734;
wire n_1491;
wire n_1840;
wire n_4434;
wire n_5307;
wire n_2244;
wire n_4290;
wire n_2586;
wire n_1684;
wire n_2446;
wire n_1346;
wire n_1352;
wire n_5407;
wire n_2017;
wire n_3029;
wire n_3597;
wire n_1046;
wire n_2560;
wire n_2704;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_3790;
wire n_2766;
wire n_3318;
wire n_4833;
wire n_5062;
wire n_5230;
wire n_4888;
wire n_776;
wire n_1823;
wire n_2479;
wire n_3350;
wire n_2782;
wire n_3977;
wire n_3588;
wire n_4279;
wire n_5008;
wire n_1456;
wire n_5004;
wire n_5294;
wire n_2229;
wire n_4133;
wire n_4527;
wire n_2288;
wire n_2099;
wire n_5323;
wire n_3388;
wire n_4790;
wire n_1946;
wire n_4181;
wire n_3184;
wire n_5810;
wire n_4561;
wire n_4461;
wire n_3245;
wire n_3075;
wire n_4007;
wire n_4949;
wire n_2642;
wire n_4239;
wire n_2383;
wire n_4184;
wire n_1676;
wire n_1830;
wire n_2351;
wire n_1319;
wire n_5069;
wire n_2986;
wire n_5702;
wire n_2536;
wire n_3915;
wire n_1633;
wire n_3489;
wire n_2835;
wire n_5243;
wire n_1416;
wire n_2820;
wire n_2293;
wire n_5250;
wire n_3074;
wire n_3102;
wire n_5590;
wire n_2026;
wire n_1282;
wire n_5260;
wire n_3321;
wire n_2567;
wire n_5809;
wire n_2322;
wire n_2727;
wire n_3377;
wire n_4782;
wire n_1321;
wire n_2533;
wire n_3530;
wire n_2869;
wire n_4378;
wire n_5349;
wire n_1235;
wire n_2759;
wire n_2361;
wire n_1292;
wire n_2266;
wire n_4876;
wire n_5813;
wire n_790;
wire n_5833;
wire n_2611;
wire n_2901;
wire n_4358;
wire n_5616;
wire n_5805;
wire n_2653;
wire n_1248;
wire n_902;
wire n_2189;
wire n_2246;
wire n_4469;
wire n_5169;
wire n_5816;
wire n_3156;
wire n_1941;
wire n_3483;
wire n_5416;
wire n_1794;
wire n_1236;
wire n_4493;
wire n_4924;
wire n_743;
wire n_766;
wire n_1746;
wire n_3524;
wire n_2885;
wire n_3097;
wire n_2062;
wire n_4539;
wire n_2975;
wire n_4421;
wire n_2839;
wire n_2856;
wire n_4793;
wire n_4498;
wire n_2070;
wire n_1607;
wire n_1454;
wire n_4953;
wire n_2348;
wire n_2944;
wire n_3831;
wire n_869;
wire n_1154;
wire n_1329;
wire n_5167;
wire n_5661;
wire n_5830;
wire n_3589;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_3391;
wire n_1800;
wire n_1463;
wire n_3458;
wire n_4505;
wire n_3190;
wire n_1562;
wire n_5558;
wire n_1826;
wire n_5687;
wire n_5383;
wire n_5126;
wire n_1759;
wire n_5051;
wire n_5587;
wire n_5236;
wire n_853;
wire n_875;
wire n_5012;
wire n_1678;
wire n_3787;
wire n_1256;
wire n_3585;
wire n_3565;
wire n_4450;
wire n_5025;
wire n_933;
wire n_4173;
wire n_3135;
wire n_5651;
wire n_4630;
wire n_1217;
wire n_5645;
wire n_3990;
wire n_1628;
wire n_5766;
wire n_2109;
wire n_988;
wire n_2796;
wire n_2507;
wire n_5878;
wire n_5671;
wire n_4534;
wire n_1536;
wire n_1204;
wire n_1132;
wire n_1327;
wire n_955;
wire n_2787;
wire n_2969;
wire n_2395;
wire n_1554;
wire n_4494;
wire n_5412;
wire n_769;
wire n_2380;
wire n_4786;
wire n_1120;
wire n_4579;
wire n_2290;
wire n_4811;
wire n_2048;
wire n_2005;
wire n_4857;
wire n_3432;
wire n_2736;
wire n_2883;
wire n_1408;
wire n_4282;
wire n_1196;
wire n_3493;
wire n_863;
wire n_3774;
wire n_5733;
wire n_2910;
wire n_748;
wire n_3268;
wire n_1785;
wire n_1147;
wire n_1754;
wire n_3057;
wire n_3701;
wire n_5148;
wire n_2584;
wire n_1812;
wire n_866;
wire n_2287;
wire n_5791;
wire n_5727;
wire n_761;
wire n_2492;
wire n_3778;
wire n_5328;
wire n_5657;
wire n_1173;
wire n_4974;
wire n_4911;
wire n_4436;
wire n_5119;
wire n_4569;
wire n_1174;
wire n_3334;
wire n_5602;
wire n_5097;
wire n_844;
wire n_4985;
wire n_2117;
wire n_2234;
wire n_3823;
wire n_4384;
wire n_2741;
wire n_3114;
wire n_888;
wire n_2203;
wire n_2255;
wire n_3584;
wire n_5246;
wire n_4858;
wire n_4678;
wire n_2649;
wire n_3556;
wire n_3836;
wire n_5579;
wire n_1922;
wire n_5750;
wire n_4823;
wire n_5831;
wire n_4309;
wire n_4363;
wire n_1215;
wire n_839;
wire n_5107;
wire n_3456;
wire n_5095;
wire n_779;
wire n_1537;
wire n_2205;
wire n_4243;
wire n_4025;
wire n_3404;
wire n_1122;
wire n_5666;
wire n_4059;
wire n_1509;
wire n_4121;
wire n_3290;
wire n_1109;
wire n_4313;
wire n_3309;
wire n_3671;
wire n_4142;
wire n_2015;
wire n_3982;
wire n_2609;
wire n_1161;
wire n_5546;
wire n_3796;
wire n_3840;
wire n_3461;
wire n_3408;
wire n_4246;
wire n_3513;
wire n_3690;
wire n_1184;
wire n_2483;
wire n_4532;
wire n_1525;
wire n_3995;
wire n_4076;
wire n_2594;
wire n_4244;
wire n_2147;
wire n_2503;
wire n_4049;
wire n_1156;
wire n_2600;
wire n_984;
wire n_5626;
wire n_3508;
wire n_868;
wire n_4353;
wire n_735;
wire n_4787;
wire n_5633;
wire n_1218;
wire n_5664;
wire n_3596;
wire n_4537;
wire n_4346;
wire n_4351;
wire n_2429;
wire n_985;
wire n_2440;
wire n_3521;
wire n_802;
wire n_980;
wire n_2681;
wire n_1651;
wire n_2360;
wire n_3764;
wire n_4784;
wire n_4075;
wire n_5340;
wire n_3947;
wire n_1244;
wire n_1685;
wire n_3066;
wire n_2844;
wire n_2303;
wire n_1619;
wire n_2285;
wire n_5280;
wire n_4451;
wire n_4332;
wire n_810;
wire n_1194;
wire n_4538;
wire n_4506;
wire n_2742;
wire n_3695;
wire n_3976;
wire n_3563;
wire n_2367;
wire n_3198;
wire n_3495;
wire n_1034;
wire n_2909;
wire n_754;
wire n_5369;
wire n_975;
wire n_5730;
wire n_5576;
wire n_3359;
wire n_5272;
wire n_3187;
wire n_3218;
wire n_861;
wire n_857;
wire n_2107;
wire n_2040;
wire n_2968;
wire n_4201;
wire n_4336;
wire n_2221;
wire n_5646;
wire n_5624;
wire n_4852;
wire n_1010;
wire n_4210;
wire n_4981;
wire n_1166;
wire n_5440;
wire n_2891;
wire n_2709;
wire n_1578;
wire n_1861;
wire n_3955;
wire n_1557;
wire n_2280;
wire n_3945;
wire n_730;
wire n_5817;
wire n_5214;
wire n_1898;
wire n_2443;
wire n_4936;
wire n_4205;
wire n_2162;
wire n_1868;
wire n_2079;
wire n_4763;
wire n_3587;
wire n_4278;
wire n_5586;
wire n_3433;
wire n_4463;
wire n_2185;
wire n_5861;
wire n_3833;
wire n_1836;
wire n_2774;
wire n_3162;
wire n_1274;
wire n_1486;
wire n_3333;
wire n_4129;
wire n_5258;
wire n_5032;
wire n_1899;
wire n_784;
wire n_4804;
wire n_5619;
wire n_3965;
wire n_5859;
wire n_5380;
wire n_4500;
wire n_5065;
wire n_862;
wire n_5776;
wire n_2098;
wire n_3085;
wire n_4433;
wire n_5606;
wire n_5644;
wire n_2813;
wire n_1935;
wire n_5826;
wire n_2027;
wire n_2091;
wire n_2991;
wire n_5030;
wire n_4194;
wire n_1449;
wire n_4703;
wire n_2419;
wire n_5683;
wire n_2677;
wire n_3182;
wire n_5756;
wire n_3283;
wire n_5527;
wire n_1742;
wire n_4030;

INVx1_ASAP7_75t_L g717 ( 
.A(n_408),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_550),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_709),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_577),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_453),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_568),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_213),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_118),
.Y(n_724)
);

CKINVDCx20_ASAP7_75t_R g725 ( 
.A(n_0),
.Y(n_725)
);

CKINVDCx20_ASAP7_75t_R g726 ( 
.A(n_630),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_201),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_92),
.Y(n_728)
);

CKINVDCx20_ASAP7_75t_R g729 ( 
.A(n_263),
.Y(n_729)
);

BUFx10_ASAP7_75t_L g730 ( 
.A(n_502),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_310),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_441),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_636),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_1),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_108),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_657),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_193),
.Y(n_737)
);

BUFx6f_ASAP7_75t_L g738 ( 
.A(n_92),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_705),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_63),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_692),
.Y(n_741)
);

INVxp67_ASAP7_75t_L g742 ( 
.A(n_79),
.Y(n_742)
);

BUFx2_ASAP7_75t_L g743 ( 
.A(n_303),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_701),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_710),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_697),
.Y(n_746)
);

INVx2_ASAP7_75t_SL g747 ( 
.A(n_609),
.Y(n_747)
);

BUFx2_ASAP7_75t_L g748 ( 
.A(n_631),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_504),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_114),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_351),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_432),
.Y(n_752)
);

BUFx10_ASAP7_75t_L g753 ( 
.A(n_229),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_333),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_164),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_231),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_585),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_459),
.Y(n_758)
);

BUFx2_ASAP7_75t_L g759 ( 
.A(n_687),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_704),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_459),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_8),
.Y(n_762)
);

CKINVDCx16_ASAP7_75t_R g763 ( 
.A(n_689),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_517),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_550),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_134),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_558),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_488),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_190),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_590),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_591),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_7),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_532),
.Y(n_773)
);

CKINVDCx20_ASAP7_75t_R g774 ( 
.A(n_60),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_4),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_114),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_119),
.Y(n_777)
);

INVx2_ASAP7_75t_SL g778 ( 
.A(n_52),
.Y(n_778)
);

BUFx6f_ASAP7_75t_L g779 ( 
.A(n_454),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_154),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_207),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_310),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_504),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_406),
.Y(n_784)
);

CKINVDCx20_ASAP7_75t_R g785 ( 
.A(n_15),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_377),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_445),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_166),
.Y(n_788)
);

BUFx6f_ASAP7_75t_L g789 ( 
.A(n_676),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_213),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_242),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_495),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_17),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_603),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_393),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_268),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_461),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_534),
.Y(n_798)
);

CKINVDCx20_ASAP7_75t_R g799 ( 
.A(n_589),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_486),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_621),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_488),
.Y(n_802)
);

CKINVDCx20_ASAP7_75t_R g803 ( 
.A(n_318),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_259),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_165),
.Y(n_805)
);

BUFx10_ASAP7_75t_L g806 ( 
.A(n_679),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_396),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_236),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_77),
.Y(n_809)
);

BUFx10_ASAP7_75t_L g810 ( 
.A(n_632),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_305),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_526),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_163),
.Y(n_813)
);

BUFx10_ASAP7_75t_L g814 ( 
.A(n_399),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_389),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_224),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_162),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_422),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_321),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_699),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_144),
.Y(n_821)
);

BUFx10_ASAP7_75t_L g822 ( 
.A(n_526),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_151),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_580),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_534),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_325),
.Y(n_826)
);

INVxp67_ASAP7_75t_L g827 ( 
.A(n_443),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_522),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_324),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_623),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_143),
.Y(n_831)
);

CKINVDCx20_ASAP7_75t_R g832 ( 
.A(n_537),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_228),
.Y(n_833)
);

INVx1_ASAP7_75t_SL g834 ( 
.A(n_66),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_183),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_431),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_44),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_202),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_378),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_448),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_707),
.Y(n_841)
);

CKINVDCx20_ASAP7_75t_R g842 ( 
.A(n_360),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_357),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_277),
.Y(n_844)
);

CKINVDCx20_ASAP7_75t_R g845 ( 
.A(n_437),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_90),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_118),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_160),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_81),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_117),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_13),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_108),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_413),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_473),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_484),
.Y(n_855)
);

BUFx2_ASAP7_75t_L g856 ( 
.A(n_506),
.Y(n_856)
);

CKINVDCx16_ASAP7_75t_R g857 ( 
.A(n_604),
.Y(n_857)
);

BUFx6f_ASAP7_75t_L g858 ( 
.A(n_485),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_17),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_512),
.Y(n_860)
);

BUFx10_ASAP7_75t_L g861 ( 
.A(n_252),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_397),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_423),
.Y(n_863)
);

BUFx6f_ASAP7_75t_L g864 ( 
.A(n_346),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_431),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_456),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_127),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_242),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_629),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_599),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_712),
.Y(n_871)
);

CKINVDCx20_ASAP7_75t_R g872 ( 
.A(n_585),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_122),
.Y(n_873)
);

BUFx2_ASAP7_75t_L g874 ( 
.A(n_570),
.Y(n_874)
);

BUFx3_ASAP7_75t_L g875 ( 
.A(n_591),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_437),
.Y(n_876)
);

BUFx3_ASAP7_75t_L g877 ( 
.A(n_649),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_680),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_208),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_352),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_168),
.Y(n_881)
);

CKINVDCx20_ASAP7_75t_R g882 ( 
.A(n_237),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_421),
.Y(n_883)
);

BUFx6f_ASAP7_75t_L g884 ( 
.A(n_614),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_11),
.Y(n_885)
);

CKINVDCx20_ASAP7_75t_R g886 ( 
.A(n_300),
.Y(n_886)
);

INVx1_ASAP7_75t_SL g887 ( 
.A(n_597),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_408),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_194),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_271),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_349),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_395),
.Y(n_892)
);

INVx1_ASAP7_75t_SL g893 ( 
.A(n_539),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_652),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_514),
.Y(n_895)
);

CKINVDCx20_ASAP7_75t_R g896 ( 
.A(n_76),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_227),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_130),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_153),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_634),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_198),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_112),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_14),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_518),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_548),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_425),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_294),
.Y(n_907)
);

INVx1_ASAP7_75t_SL g908 ( 
.A(n_141),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_566),
.Y(n_909)
);

CKINVDCx20_ASAP7_75t_R g910 ( 
.A(n_224),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_377),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_535),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_319),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_714),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_61),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_693),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_460),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_566),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_428),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_248),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_644),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_482),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_611),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_170),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_106),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_110),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_662),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_180),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_12),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_616),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_354),
.Y(n_931)
);

CKINVDCx20_ASAP7_75t_R g932 ( 
.A(n_563),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_579),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_93),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_338),
.Y(n_935)
);

BUFx3_ASAP7_75t_L g936 ( 
.A(n_31),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_327),
.Y(n_937)
);

BUFx10_ASAP7_75t_L g938 ( 
.A(n_677),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_70),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_326),
.Y(n_940)
);

INVxp67_ASAP7_75t_SL g941 ( 
.A(n_72),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_539),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_170),
.Y(n_943)
);

CKINVDCx20_ASAP7_75t_R g944 ( 
.A(n_61),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_486),
.Y(n_945)
);

BUFx6f_ASAP7_75t_L g946 ( 
.A(n_601),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_670),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_33),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_463),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_96),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_572),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_453),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_240),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_212),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_387),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_35),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_233),
.Y(n_957)
);

BUFx3_ASAP7_75t_L g958 ( 
.A(n_119),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_85),
.Y(n_959)
);

CKINVDCx20_ASAP7_75t_R g960 ( 
.A(n_350),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_237),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_329),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_304),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_267),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_590),
.Y(n_965)
);

BUFx3_ASAP7_75t_L g966 ( 
.A(n_438),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_162),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_264),
.Y(n_968)
);

BUFx3_ASAP7_75t_L g969 ( 
.A(n_97),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_522),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_21),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_93),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_335),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_65),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_87),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_382),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_357),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_147),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_596),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_641),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_344),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_683),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_140),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_563),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_222),
.Y(n_985)
);

INVx1_ASAP7_75t_SL g986 ( 
.A(n_24),
.Y(n_986)
);

INVxp67_ASAP7_75t_SL g987 ( 
.A(n_577),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_510),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_33),
.Y(n_989)
);

CKINVDCx20_ASAP7_75t_R g990 ( 
.A(n_667),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_14),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_243),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_306),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_548),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_691),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_643),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_178),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_530),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_695),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_369),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_449),
.Y(n_1001)
);

CKINVDCx20_ASAP7_75t_R g1002 ( 
.A(n_94),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_523),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_440),
.Y(n_1004)
);

CKINVDCx20_ASAP7_75t_R g1005 ( 
.A(n_419),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_251),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_307),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_675),
.Y(n_1008)
);

INVx1_ASAP7_75t_SL g1009 ( 
.A(n_678),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_716),
.Y(n_1010)
);

INVx1_ASAP7_75t_SL g1011 ( 
.A(n_538),
.Y(n_1011)
);

BUFx6f_ASAP7_75t_L g1012 ( 
.A(n_354),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_50),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_379),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_216),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_416),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_85),
.Y(n_1017)
);

INVx2_ASAP7_75t_SL g1018 ( 
.A(n_286),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_514),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_264),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_382),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_250),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_196),
.Y(n_1023)
);

INVx2_ASAP7_75t_SL g1024 ( 
.A(n_650),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_622),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_446),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_485),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_686),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_702),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_694),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_246),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_635),
.Y(n_1032)
);

BUFx10_ASAP7_75t_L g1033 ( 
.A(n_161),
.Y(n_1033)
);

CKINVDCx20_ASAP7_75t_R g1034 ( 
.A(n_659),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_639),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_576),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_373),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_703),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_410),
.Y(n_1039)
);

INVx2_ASAP7_75t_SL g1040 ( 
.A(n_706),
.Y(n_1040)
);

INVx1_ASAP7_75t_SL g1041 ( 
.A(n_188),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_435),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_385),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_445),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_120),
.Y(n_1045)
);

CKINVDCx20_ASAP7_75t_R g1046 ( 
.A(n_201),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_479),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_560),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_262),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_255),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_222),
.Y(n_1051)
);

CKINVDCx20_ASAP7_75t_R g1052 ( 
.A(n_146),
.Y(n_1052)
);

BUFx2_ASAP7_75t_SL g1053 ( 
.A(n_524),
.Y(n_1053)
);

BUFx3_ASAP7_75t_L g1054 ( 
.A(n_461),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_421),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_420),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_265),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_537),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_665),
.Y(n_1059)
);

BUFx10_ASAP7_75t_L g1060 ( 
.A(n_545),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_94),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_575),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_292),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_598),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_536),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_183),
.Y(n_1066)
);

CKINVDCx20_ASAP7_75t_R g1067 ( 
.A(n_529),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_105),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_128),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_672),
.Y(n_1070)
);

CKINVDCx20_ASAP7_75t_R g1071 ( 
.A(n_101),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_150),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_669),
.Y(n_1073)
);

INVxp67_ASAP7_75t_L g1074 ( 
.A(n_711),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_317),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_380),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_172),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_412),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_394),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_579),
.Y(n_1080)
);

INVxp67_ASAP7_75t_L g1081 ( 
.A(n_148),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_681),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_465),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_384),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_444),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_90),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_18),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_59),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_335),
.Y(n_1089)
);

CKINVDCx16_ASAP7_75t_R g1090 ( 
.A(n_356),
.Y(n_1090)
);

BUFx10_ASAP7_75t_L g1091 ( 
.A(n_389),
.Y(n_1091)
);

BUFx3_ASAP7_75t_L g1092 ( 
.A(n_82),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_168),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_473),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_220),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_243),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_660),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_551),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_36),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_5),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_196),
.Y(n_1101)
);

CKINVDCx20_ASAP7_75t_R g1102 ( 
.A(n_387),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_178),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_544),
.Y(n_1104)
);

BUFx10_ASAP7_75t_L g1105 ( 
.A(n_215),
.Y(n_1105)
);

INVx2_ASAP7_75t_SL g1106 ( 
.A(n_460),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_399),
.Y(n_1107)
);

BUFx6f_ASAP7_75t_L g1108 ( 
.A(n_575),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_334),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_122),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_133),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_220),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_696),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_20),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_296),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_217),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_52),
.Y(n_1117)
);

CKINVDCx20_ASAP7_75t_R g1118 ( 
.A(n_238),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_713),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_181),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_166),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_637),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_81),
.Y(n_1123)
);

BUFx3_ASAP7_75t_L g1124 ( 
.A(n_176),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_661),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_531),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_261),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_470),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_332),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_440),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_521),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_651),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_76),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_228),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_319),
.Y(n_1135)
);

CKINVDCx20_ASAP7_75t_R g1136 ( 
.A(n_372),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_156),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_150),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_255),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_518),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_433),
.Y(n_1141)
);

INVxp67_ASAP7_75t_SL g1142 ( 
.A(n_429),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_100),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_715),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_564),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_463),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_89),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_59),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_216),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_136),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_658),
.Y(n_1151)
);

CKINVDCx14_ASAP7_75t_R g1152 ( 
.A(n_214),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_684),
.Y(n_1153)
);

INVx1_ASAP7_75t_SL g1154 ( 
.A(n_475),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_449),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_471),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_227),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_223),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_290),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_65),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_682),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_369),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_342),
.Y(n_1163)
);

BUFx6f_ASAP7_75t_L g1164 ( 
.A(n_543),
.Y(n_1164)
);

INVx1_ASAP7_75t_SL g1165 ( 
.A(n_111),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_673),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_458),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_688),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_208),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_509),
.Y(n_1170)
);

INVx2_ASAP7_75t_SL g1171 ( 
.A(n_230),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_308),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_322),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_690),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_441),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_581),
.Y(n_1176)
);

INVx1_ASAP7_75t_SL g1177 ( 
.A(n_312),
.Y(n_1177)
);

BUFx5_ASAP7_75t_L g1178 ( 
.A(n_29),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_278),
.Y(n_1179)
);

BUFx10_ASAP7_75t_L g1180 ( 
.A(n_232),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_533),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_619),
.Y(n_1182)
);

CKINVDCx16_ASAP7_75t_R g1183 ( 
.A(n_348),
.Y(n_1183)
);

CKINVDCx14_ASAP7_75t_R g1184 ( 
.A(n_350),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_171),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_256),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_321),
.Y(n_1187)
);

BUFx2_ASAP7_75t_L g1188 ( 
.A(n_542),
.Y(n_1188)
);

INVx1_ASAP7_75t_SL g1189 ( 
.A(n_24),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_351),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_700),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_646),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_402),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_80),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_326),
.Y(n_1195)
);

BUFx3_ASAP7_75t_L g1196 ( 
.A(n_469),
.Y(n_1196)
);

INVxp67_ASAP7_75t_L g1197 ( 
.A(n_270),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_44),
.Y(n_1198)
);

BUFx6f_ASAP7_75t_L g1199 ( 
.A(n_358),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_656),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_322),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_248),
.Y(n_1202)
);

BUFx3_ASAP7_75t_L g1203 ( 
.A(n_229),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_41),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_234),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_645),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_501),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_685),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_355),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_204),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_360),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_708),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_188),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_664),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_474),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_368),
.Y(n_1216)
);

INVx2_ASAP7_75t_SL g1217 ( 
.A(n_258),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_373),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_238),
.Y(n_1219)
);

INVx4_ASAP7_75t_R g1220 ( 
.A(n_490),
.Y(n_1220)
);

INVxp67_ASAP7_75t_L g1221 ( 
.A(n_63),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_120),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_497),
.Y(n_1223)
);

BUFx8_ASAP7_75t_SL g1224 ( 
.A(n_562),
.Y(n_1224)
);

INVx2_ASAP7_75t_L g1225 ( 
.A(n_138),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_558),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_328),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_523),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_149),
.Y(n_1229)
);

CKINVDCx20_ASAP7_75t_R g1230 ( 
.A(n_551),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_648),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_274),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_330),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_278),
.Y(n_1234)
);

BUFx3_ASAP7_75t_L g1235 ( 
.A(n_138),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_448),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_25),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_300),
.Y(n_1238)
);

CKINVDCx20_ASAP7_75t_R g1239 ( 
.A(n_71),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_95),
.Y(n_1240)
);

CKINVDCx20_ASAP7_75t_R g1241 ( 
.A(n_531),
.Y(n_1241)
);

CKINVDCx5p33_ASAP7_75t_R g1242 ( 
.A(n_323),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_26),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_583),
.Y(n_1244)
);

BUFx10_ASAP7_75t_L g1245 ( 
.A(n_606),
.Y(n_1245)
);

BUFx10_ASAP7_75t_L g1246 ( 
.A(n_594),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_698),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_38),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_74),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_415),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_315),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_542),
.Y(n_1252)
);

CKINVDCx20_ASAP7_75t_R g1253 ( 
.A(n_125),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_223),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1178),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_1224),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1178),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1178),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_1152),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1178),
.Y(n_1260)
);

BUFx3_ASAP7_75t_L g1261 ( 
.A(n_877),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1178),
.Y(n_1262)
);

INVx2_ASAP7_75t_L g1263 ( 
.A(n_1178),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1178),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1178),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1178),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_738),
.Y(n_1267)
);

BUFx3_ASAP7_75t_L g1268 ( 
.A(n_877),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_733),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_733),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_741),
.Y(n_1271)
);

INVxp33_ASAP7_75t_L g1272 ( 
.A(n_743),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_738),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_741),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_745),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_745),
.Y(n_1276)
);

CKINVDCx20_ASAP7_75t_R g1277 ( 
.A(n_725),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_738),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_760),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_760),
.Y(n_1280)
);

BUFx3_ASAP7_75t_L g1281 ( 
.A(n_806),
.Y(n_1281)
);

INVxp33_ASAP7_75t_L g1282 ( 
.A(n_743),
.Y(n_1282)
);

INVxp33_ASAP7_75t_L g1283 ( 
.A(n_856),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_794),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_794),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_738),
.Y(n_1286)
);

CKINVDCx20_ASAP7_75t_R g1287 ( 
.A(n_729),
.Y(n_1287)
);

BUFx3_ASAP7_75t_L g1288 ( 
.A(n_806),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_801),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_801),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_830),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_830),
.Y(n_1292)
);

INVx2_ASAP7_75t_SL g1293 ( 
.A(n_730),
.Y(n_1293)
);

BUFx6f_ASAP7_75t_L g1294 ( 
.A(n_789),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_841),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_841),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_870),
.Y(n_1297)
);

INVx1_ASAP7_75t_SL g1298 ( 
.A(n_856),
.Y(n_1298)
);

CKINVDCx20_ASAP7_75t_R g1299 ( 
.A(n_774),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_870),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_1184),
.Y(n_1301)
);

INVxp33_ASAP7_75t_L g1302 ( 
.A(n_874),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_871),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_871),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_900),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_719),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_900),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_916),
.Y(n_1308)
);

INVx1_ASAP7_75t_SL g1309 ( 
.A(n_874),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_738),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_916),
.Y(n_1311)
);

INVx1_ASAP7_75t_SL g1312 ( 
.A(n_1188),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_923),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_923),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_930),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_930),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_996),
.Y(n_1317)
);

INVx2_ASAP7_75t_SL g1318 ( 
.A(n_730),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_996),
.Y(n_1319)
);

CKINVDCx20_ASAP7_75t_R g1320 ( 
.A(n_785),
.Y(n_1320)
);

CKINVDCx5p33_ASAP7_75t_R g1321 ( 
.A(n_1090),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1025),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1025),
.Y(n_1323)
);

INVx2_ASAP7_75t_L g1324 ( 
.A(n_779),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1028),
.Y(n_1325)
);

INVxp33_ASAP7_75t_L g1326 ( 
.A(n_1188),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_1183),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_718),
.Y(n_1328)
);

INVxp33_ASAP7_75t_L g1329 ( 
.A(n_717),
.Y(n_1329)
);

CKINVDCx20_ASAP7_75t_R g1330 ( 
.A(n_799),
.Y(n_1330)
);

CKINVDCx5p33_ASAP7_75t_R g1331 ( 
.A(n_720),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1028),
.Y(n_1332)
);

INVxp67_ASAP7_75t_SL g1333 ( 
.A(n_748),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1035),
.Y(n_1334)
);

INVxp67_ASAP7_75t_SL g1335 ( 
.A(n_748),
.Y(n_1335)
);

CKINVDCx14_ASAP7_75t_R g1336 ( 
.A(n_759),
.Y(n_1336)
);

INVxp67_ASAP7_75t_SL g1337 ( 
.A(n_759),
.Y(n_1337)
);

CKINVDCx16_ASAP7_75t_R g1338 ( 
.A(n_763),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1035),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1070),
.Y(n_1340)
);

INVxp33_ASAP7_75t_L g1341 ( 
.A(n_717),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1070),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1073),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_721),
.Y(n_1344)
);

INVxp67_ASAP7_75t_L g1345 ( 
.A(n_1053),
.Y(n_1345)
);

CKINVDCx5p33_ASAP7_75t_R g1346 ( 
.A(n_722),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_723),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1073),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_779),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_779),
.Y(n_1350)
);

INVxp67_ASAP7_75t_L g1351 ( 
.A(n_1053),
.Y(n_1351)
);

INVxp33_ASAP7_75t_SL g1352 ( 
.A(n_727),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1097),
.Y(n_1353)
);

BUFx6f_ASAP7_75t_L g1354 ( 
.A(n_789),
.Y(n_1354)
);

INVxp67_ASAP7_75t_SL g1355 ( 
.A(n_1074),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1097),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1122),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_779),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1122),
.Y(n_1359)
);

CKINVDCx20_ASAP7_75t_R g1360 ( 
.A(n_803),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1125),
.Y(n_1361)
);

BUFx2_ASAP7_75t_L g1362 ( 
.A(n_875),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1125),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1153),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1153),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1174),
.Y(n_1366)
);

CKINVDCx20_ASAP7_75t_R g1367 ( 
.A(n_832),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1174),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_779),
.Y(n_1369)
);

CKINVDCx16_ASAP7_75t_R g1370 ( 
.A(n_857),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1208),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1208),
.Y(n_1372)
);

CKINVDCx20_ASAP7_75t_R g1373 ( 
.A(n_842),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_875),
.Y(n_1374)
);

INVxp33_ASAP7_75t_L g1375 ( 
.A(n_724),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_936),
.Y(n_1376)
);

BUFx3_ASAP7_75t_L g1377 ( 
.A(n_806),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_936),
.Y(n_1378)
);

BUFx5_ASAP7_75t_L g1379 ( 
.A(n_806),
.Y(n_1379)
);

CKINVDCx20_ASAP7_75t_R g1380 ( 
.A(n_845),
.Y(n_1380)
);

CKINVDCx20_ASAP7_75t_R g1381 ( 
.A(n_872),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_958),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_958),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_966),
.Y(n_1384)
);

BUFx10_ASAP7_75t_L g1385 ( 
.A(n_858),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_966),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_969),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_969),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1054),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1054),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1092),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1092),
.Y(n_1392)
);

NOR2xp33_ASAP7_75t_L g1393 ( 
.A(n_747),
.B(n_1),
.Y(n_1393)
);

CKINVDCx16_ASAP7_75t_R g1394 ( 
.A(n_730),
.Y(n_1394)
);

INVxp33_ASAP7_75t_L g1395 ( 
.A(n_724),
.Y(n_1395)
);

BUFx3_ASAP7_75t_L g1396 ( 
.A(n_810),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1124),
.Y(n_1397)
);

INVx2_ASAP7_75t_L g1398 ( 
.A(n_858),
.Y(n_1398)
);

INVxp67_ASAP7_75t_SL g1399 ( 
.A(n_858),
.Y(n_1399)
);

INVxp33_ASAP7_75t_SL g1400 ( 
.A(n_734),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1124),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1196),
.Y(n_1402)
);

INVxp33_ASAP7_75t_L g1403 ( 
.A(n_731),
.Y(n_1403)
);

INVxp33_ASAP7_75t_L g1404 ( 
.A(n_731),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1196),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1203),
.Y(n_1406)
);

INVx1_ASAP7_75t_SL g1407 ( 
.A(n_882),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1203),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1235),
.Y(n_1409)
);

HB1xp67_ASAP7_75t_L g1410 ( 
.A(n_735),
.Y(n_1410)
);

INVxp33_ASAP7_75t_L g1411 ( 
.A(n_740),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1235),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_858),
.Y(n_1413)
);

CKINVDCx5p33_ASAP7_75t_R g1414 ( 
.A(n_737),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_858),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_864),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_864),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_864),
.Y(n_1418)
);

CKINVDCx14_ASAP7_75t_R g1419 ( 
.A(n_810),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_864),
.Y(n_1420)
);

HB1xp67_ASAP7_75t_L g1421 ( 
.A(n_749),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_864),
.Y(n_1422)
);

NOR2xp67_ASAP7_75t_L g1423 ( 
.A(n_742),
.B(n_0),
.Y(n_1423)
);

BUFx6f_ASAP7_75t_L g1424 ( 
.A(n_789),
.Y(n_1424)
);

INVx4_ASAP7_75t_R g1425 ( 
.A(n_747),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1012),
.Y(n_1426)
);

INVxp67_ASAP7_75t_SL g1427 ( 
.A(n_1012),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1012),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1012),
.Y(n_1429)
);

CKINVDCx5p33_ASAP7_75t_R g1430 ( 
.A(n_736),
.Y(n_1430)
);

CKINVDCx5p33_ASAP7_75t_R g1431 ( 
.A(n_739),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1012),
.Y(n_1432)
);

CKINVDCx20_ASAP7_75t_R g1433 ( 
.A(n_886),
.Y(n_1433)
);

BUFx3_ASAP7_75t_L g1434 ( 
.A(n_810),
.Y(n_1434)
);

INVxp67_ASAP7_75t_SL g1435 ( 
.A(n_1108),
.Y(n_1435)
);

CKINVDCx5p33_ASAP7_75t_R g1436 ( 
.A(n_746),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1108),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1108),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1108),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1108),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1164),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1164),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1164),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1164),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1164),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_1199),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1199),
.Y(n_1447)
);

CKINVDCx20_ASAP7_75t_R g1448 ( 
.A(n_896),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1199),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1199),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1199),
.Y(n_1451)
);

INVx1_ASAP7_75t_SL g1452 ( 
.A(n_910),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_728),
.Y(n_1453)
);

INVxp33_ASAP7_75t_SL g1454 ( 
.A(n_752),
.Y(n_1454)
);

INVxp33_ASAP7_75t_SL g1455 ( 
.A(n_754),
.Y(n_1455)
);

OR2x2_ASAP7_75t_L g1456 ( 
.A(n_778),
.B(n_1018),
.Y(n_1456)
);

INVxp33_ASAP7_75t_SL g1457 ( 
.A(n_755),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_732),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_732),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_873),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_876),
.Y(n_1461)
);

CKINVDCx20_ASAP7_75t_R g1462 ( 
.A(n_932),
.Y(n_1462)
);

INVx1_ASAP7_75t_SL g1463 ( 
.A(n_944),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_883),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_740),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_750),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_750),
.Y(n_1467)
);

INVxp67_ASAP7_75t_SL g1468 ( 
.A(n_744),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_757),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_751),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_757),
.Y(n_1471)
);

INVxp67_ASAP7_75t_SL g1472 ( 
.A(n_744),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_751),
.Y(n_1473)
);

CKINVDCx5p33_ASAP7_75t_R g1474 ( 
.A(n_756),
.Y(n_1474)
);

INVxp67_ASAP7_75t_SL g1475 ( 
.A(n_1030),
.Y(n_1475)
);

CKINVDCx5p33_ASAP7_75t_R g1476 ( 
.A(n_758),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_762),
.Y(n_1477)
);

INVx1_ASAP7_75t_SL g1478 ( 
.A(n_960),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_762),
.Y(n_1479)
);

CKINVDCx5p33_ASAP7_75t_R g1480 ( 
.A(n_761),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_764),
.Y(n_1481)
);

BUFx6f_ASAP7_75t_L g1482 ( 
.A(n_789),
.Y(n_1482)
);

INVxp33_ASAP7_75t_L g1483 ( 
.A(n_764),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_765),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_765),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_767),
.Y(n_1486)
);

BUFx2_ASAP7_75t_L g1487 ( 
.A(n_766),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_767),
.Y(n_1488)
);

CKINVDCx14_ASAP7_75t_R g1489 ( 
.A(n_810),
.Y(n_1489)
);

INVxp33_ASAP7_75t_SL g1490 ( 
.A(n_773),
.Y(n_1490)
);

INVxp33_ASAP7_75t_SL g1491 ( 
.A(n_776),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_768),
.Y(n_1492)
);

INVxp67_ASAP7_75t_SL g1493 ( 
.A(n_1030),
.Y(n_1493)
);

INVxp33_ASAP7_75t_L g1494 ( 
.A(n_768),
.Y(n_1494)
);

INVxp33_ASAP7_75t_L g1495 ( 
.A(n_769),
.Y(n_1495)
);

INVx3_ASAP7_75t_L g1496 ( 
.A(n_1166),
.Y(n_1496)
);

BUFx3_ASAP7_75t_L g1497 ( 
.A(n_938),
.Y(n_1497)
);

INVxp33_ASAP7_75t_SL g1498 ( 
.A(n_780),
.Y(n_1498)
);

BUFx2_ASAP7_75t_SL g1499 ( 
.A(n_726),
.Y(n_1499)
);

BUFx3_ASAP7_75t_L g1500 ( 
.A(n_938),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_769),
.Y(n_1501)
);

INVxp33_ASAP7_75t_L g1502 ( 
.A(n_770),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_771),
.Y(n_1503)
);

INVxp67_ASAP7_75t_L g1504 ( 
.A(n_770),
.Y(n_1504)
);

CKINVDCx5p33_ASAP7_75t_R g1505 ( 
.A(n_782),
.Y(n_1505)
);

INVxp33_ASAP7_75t_L g1506 ( 
.A(n_772),
.Y(n_1506)
);

NAND2xp33_ASAP7_75t_R g1507 ( 
.A(n_820),
.B(n_2),
.Y(n_1507)
);

CKINVDCx5p33_ASAP7_75t_R g1508 ( 
.A(n_783),
.Y(n_1508)
);

CKINVDCx5p33_ASAP7_75t_R g1509 ( 
.A(n_784),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_772),
.Y(n_1510)
);

CKINVDCx20_ASAP7_75t_R g1511 ( 
.A(n_1002),
.Y(n_1511)
);

CKINVDCx5p33_ASAP7_75t_R g1512 ( 
.A(n_787),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_775),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_771),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_781),
.Y(n_1515)
);

NOR2xp67_ASAP7_75t_L g1516 ( 
.A(n_827),
.B(n_2),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_775),
.Y(n_1517)
);

HB1xp67_ASAP7_75t_L g1518 ( 
.A(n_790),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_777),
.Y(n_1519)
);

CKINVDCx20_ASAP7_75t_R g1520 ( 
.A(n_1005),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_777),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_788),
.Y(n_1522)
);

CKINVDCx5p33_ASAP7_75t_R g1523 ( 
.A(n_791),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_788),
.Y(n_1524)
);

INVxp67_ASAP7_75t_L g1525 ( 
.A(n_802),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_802),
.Y(n_1526)
);

INVxp67_ASAP7_75t_SL g1527 ( 
.A(n_1166),
.Y(n_1527)
);

INVxp67_ASAP7_75t_L g1528 ( 
.A(n_805),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_805),
.Y(n_1529)
);

CKINVDCx5p33_ASAP7_75t_R g1530 ( 
.A(n_793),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_811),
.Y(n_1531)
);

CKINVDCx5p33_ASAP7_75t_R g1532 ( 
.A(n_795),
.Y(n_1532)
);

INVxp67_ASAP7_75t_SL g1533 ( 
.A(n_1081),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_811),
.Y(n_1534)
);

CKINVDCx20_ASAP7_75t_R g1535 ( 
.A(n_1046),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_823),
.Y(n_1536)
);

CKINVDCx5p33_ASAP7_75t_R g1537 ( 
.A(n_796),
.Y(n_1537)
);

CKINVDCx5p33_ASAP7_75t_R g1538 ( 
.A(n_869),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_823),
.Y(n_1539)
);

CKINVDCx20_ASAP7_75t_R g1540 ( 
.A(n_1052),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_835),
.Y(n_1541)
);

CKINVDCx5p33_ASAP7_75t_R g1542 ( 
.A(n_797),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_781),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_835),
.Y(n_1544)
);

HB1xp67_ASAP7_75t_L g1545 ( 
.A(n_798),
.Y(n_1545)
);

CKINVDCx5p33_ASAP7_75t_R g1546 ( 
.A(n_804),
.Y(n_1546)
);

CKINVDCx16_ASAP7_75t_R g1547 ( 
.A(n_730),
.Y(n_1547)
);

INVxp67_ASAP7_75t_SL g1548 ( 
.A(n_1197),
.Y(n_1548)
);

INVx2_ASAP7_75t_SL g1549 ( 
.A(n_753),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_836),
.Y(n_1550)
);

NOR2xp67_ASAP7_75t_L g1551 ( 
.A(n_1221),
.B(n_3),
.Y(n_1551)
);

CKINVDCx16_ASAP7_75t_R g1552 ( 
.A(n_753),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_836),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_838),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_838),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_843),
.Y(n_1556)
);

BUFx2_ASAP7_75t_SL g1557 ( 
.A(n_990),
.Y(n_1557)
);

CKINVDCx20_ASAP7_75t_R g1558 ( 
.A(n_1067),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_843),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_847),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_847),
.Y(n_1561)
);

CKINVDCx14_ASAP7_75t_R g1562 ( 
.A(n_938),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_848),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_848),
.Y(n_1564)
);

CKINVDCx16_ASAP7_75t_R g1565 ( 
.A(n_753),
.Y(n_1565)
);

INVxp33_ASAP7_75t_SL g1566 ( 
.A(n_807),
.Y(n_1566)
);

BUFx3_ASAP7_75t_L g1567 ( 
.A(n_938),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_849),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_849),
.Y(n_1569)
);

HB1xp67_ASAP7_75t_L g1570 ( 
.A(n_808),
.Y(n_1570)
);

BUFx3_ASAP7_75t_L g1571 ( 
.A(n_1245),
.Y(n_1571)
);

CKINVDCx5p33_ASAP7_75t_R g1572 ( 
.A(n_809),
.Y(n_1572)
);

INVxp33_ASAP7_75t_SL g1573 ( 
.A(n_812),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_852),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_852),
.Y(n_1575)
);

INVxp33_ASAP7_75t_L g1576 ( 
.A(n_898),
.Y(n_1576)
);

BUFx3_ASAP7_75t_L g1577 ( 
.A(n_1245),
.Y(n_1577)
);

BUFx3_ASAP7_75t_L g1578 ( 
.A(n_1245),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_898),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_901),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_901),
.Y(n_1581)
);

CKINVDCx5p33_ASAP7_75t_R g1582 ( 
.A(n_878),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_902),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_902),
.Y(n_1584)
);

CKINVDCx5p33_ASAP7_75t_R g1585 ( 
.A(n_894),
.Y(n_1585)
);

CKINVDCx16_ASAP7_75t_R g1586 ( 
.A(n_753),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_906),
.Y(n_1587)
);

INVxp67_ASAP7_75t_SL g1588 ( 
.A(n_1024),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_786),
.Y(n_1589)
);

INVxp67_ASAP7_75t_SL g1590 ( 
.A(n_1024),
.Y(n_1590)
);

BUFx6f_ASAP7_75t_L g1591 ( 
.A(n_789),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_786),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_906),
.Y(n_1593)
);

HB1xp67_ASAP7_75t_L g1594 ( 
.A(n_813),
.Y(n_1594)
);

CKINVDCx20_ASAP7_75t_R g1595 ( 
.A(n_1071),
.Y(n_1595)
);

CKINVDCx5p33_ASAP7_75t_R g1596 ( 
.A(n_815),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_912),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_912),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_920),
.Y(n_1599)
);

INVxp67_ASAP7_75t_SL g1600 ( 
.A(n_1040),
.Y(n_1600)
);

HB1xp67_ASAP7_75t_SL g1601 ( 
.A(n_914),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_SL g1602 ( 
.A(n_1245),
.B(n_3),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_792),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_920),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_922),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_922),
.Y(n_1606)
);

BUFx4f_ASAP7_75t_SL g1607 ( 
.A(n_1034),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_792),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_926),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_926),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_934),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_800),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_934),
.Y(n_1613)
);

BUFx3_ASAP7_75t_L g1614 ( 
.A(n_921),
.Y(n_1614)
);

BUFx3_ASAP7_75t_L g1615 ( 
.A(n_927),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_939),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_800),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_939),
.Y(n_1618)
);

CKINVDCx5p33_ASAP7_75t_R g1619 ( 
.A(n_816),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_948),
.Y(n_1620)
);

INVxp33_ASAP7_75t_L g1621 ( 
.A(n_948),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_950),
.Y(n_1622)
);

INVxp67_ASAP7_75t_SL g1623 ( 
.A(n_1040),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_950),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_954),
.Y(n_1625)
);

CKINVDCx5p33_ASAP7_75t_R g1626 ( 
.A(n_817),
.Y(n_1626)
);

INVxp67_ASAP7_75t_SL g1627 ( 
.A(n_884),
.Y(n_1627)
);

CKINVDCx5p33_ASAP7_75t_R g1628 ( 
.A(n_818),
.Y(n_1628)
);

CKINVDCx5p33_ASAP7_75t_R g1629 ( 
.A(n_947),
.Y(n_1629)
);

CKINVDCx5p33_ASAP7_75t_R g1630 ( 
.A(n_821),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_954),
.Y(n_1631)
);

INVxp67_ASAP7_75t_L g1632 ( 
.A(n_956),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_956),
.Y(n_1633)
);

INVx1_ASAP7_75t_SL g1634 ( 
.A(n_1102),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_963),
.Y(n_1635)
);

INVxp67_ASAP7_75t_L g1636 ( 
.A(n_963),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_967),
.Y(n_1637)
);

CKINVDCx20_ASAP7_75t_R g1638 ( 
.A(n_1118),
.Y(n_1638)
);

INVx1_ASAP7_75t_SL g1639 ( 
.A(n_1136),
.Y(n_1639)
);

INVxp67_ASAP7_75t_SL g1640 ( 
.A(n_884),
.Y(n_1640)
);

CKINVDCx20_ASAP7_75t_R g1641 ( 
.A(n_1230),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_967),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_971),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_971),
.Y(n_1644)
);

INVx2_ASAP7_75t_SL g1645 ( 
.A(n_814),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_978),
.Y(n_1646)
);

INVx2_ASAP7_75t_SL g1647 ( 
.A(n_814),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_978),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_984),
.Y(n_1649)
);

BUFx2_ASAP7_75t_SL g1650 ( 
.A(n_1009),
.Y(n_1650)
);

CKINVDCx20_ASAP7_75t_R g1651 ( 
.A(n_1239),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_984),
.Y(n_1652)
);

INVxp33_ASAP7_75t_SL g1653 ( 
.A(n_824),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_989),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_989),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_993),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_993),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_998),
.Y(n_1658)
);

CKINVDCx5p33_ASAP7_75t_R g1659 ( 
.A(n_825),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_998),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1001),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1001),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1006),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1006),
.Y(n_1664)
);

CKINVDCx5p33_ASAP7_75t_R g1665 ( 
.A(n_826),
.Y(n_1665)
);

CKINVDCx5p33_ASAP7_75t_R g1666 ( 
.A(n_828),
.Y(n_1666)
);

INVxp67_ASAP7_75t_SL g1667 ( 
.A(n_884),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1007),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1007),
.Y(n_1669)
);

INVxp67_ASAP7_75t_SL g1670 ( 
.A(n_884),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1016),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1016),
.Y(n_1672)
);

BUFx6f_ASAP7_75t_L g1673 ( 
.A(n_884),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_819),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1021),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1021),
.Y(n_1676)
);

INVxp33_ASAP7_75t_SL g1677 ( 
.A(n_829),
.Y(n_1677)
);

INVxp33_ASAP7_75t_L g1678 ( 
.A(n_1036),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1036),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1043),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1043),
.Y(n_1681)
);

INVxp67_ASAP7_75t_L g1682 ( 
.A(n_1048),
.Y(n_1682)
);

CKINVDCx16_ASAP7_75t_R g1683 ( 
.A(n_814),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1048),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1049),
.Y(n_1685)
);

INVxp67_ASAP7_75t_L g1686 ( 
.A(n_1049),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1051),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1051),
.Y(n_1688)
);

BUFx6f_ASAP7_75t_L g1689 ( 
.A(n_946),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1055),
.Y(n_1690)
);

BUFx3_ASAP7_75t_L g1691 ( 
.A(n_980),
.Y(n_1691)
);

CKINVDCx5p33_ASAP7_75t_R g1692 ( 
.A(n_831),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1055),
.Y(n_1693)
);

INVxp67_ASAP7_75t_SL g1694 ( 
.A(n_946),
.Y(n_1694)
);

CKINVDCx5p33_ASAP7_75t_R g1695 ( 
.A(n_982),
.Y(n_1695)
);

INVxp33_ASAP7_75t_L g1696 ( 
.A(n_1056),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_819),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1056),
.Y(n_1698)
);

CKINVDCx14_ASAP7_75t_R g1699 ( 
.A(n_995),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1062),
.Y(n_1700)
);

NOR2xp33_ASAP7_75t_L g1701 ( 
.A(n_1588),
.B(n_778),
.Y(n_1701)
);

NOR2xp33_ASAP7_75t_SL g1702 ( 
.A(n_1298),
.B(n_814),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1267),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_SL g1704 ( 
.A(n_1379),
.B(n_822),
.Y(n_1704)
);

HB1xp67_ASAP7_75t_L g1705 ( 
.A(n_1362),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1399),
.Y(n_1706)
);

BUFx12f_ASAP7_75t_L g1707 ( 
.A(n_1256),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1336),
.B(n_822),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1267),
.Y(n_1709)
);

BUFx3_ASAP7_75t_L g1710 ( 
.A(n_1385),
.Y(n_1710)
);

BUFx12f_ASAP7_75t_L g1711 ( 
.A(n_1256),
.Y(n_1711)
);

INVx5_ASAP7_75t_L g1712 ( 
.A(n_1294),
.Y(n_1712)
);

INVx3_ASAP7_75t_L g1713 ( 
.A(n_1385),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1427),
.B(n_999),
.Y(n_1714)
);

HB1xp67_ASAP7_75t_L g1715 ( 
.A(n_1309),
.Y(n_1715)
);

BUFx6f_ASAP7_75t_L g1716 ( 
.A(n_1294),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1435),
.B(n_1008),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_SL g1718 ( 
.A(n_1379),
.B(n_822),
.Y(n_1718)
);

INVx4_ASAP7_75t_L g1719 ( 
.A(n_1306),
.Y(n_1719)
);

INVx2_ASAP7_75t_L g1720 ( 
.A(n_1273),
.Y(n_1720)
);

BUFx6f_ASAP7_75t_L g1721 ( 
.A(n_1294),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1336),
.B(n_822),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1415),
.Y(n_1723)
);

BUFx6f_ASAP7_75t_L g1724 ( 
.A(n_1294),
.Y(n_1724)
);

AND2x4_ASAP7_75t_L g1725 ( 
.A(n_1614),
.B(n_1018),
.Y(n_1725)
);

BUFx2_ASAP7_75t_L g1726 ( 
.A(n_1321),
.Y(n_1726)
);

AND2x4_ASAP7_75t_L g1727 ( 
.A(n_1614),
.B(n_1106),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1416),
.Y(n_1728)
);

INVx5_ASAP7_75t_L g1729 ( 
.A(n_1354),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1627),
.B(n_1010),
.Y(n_1730)
);

INVx2_ASAP7_75t_SL g1731 ( 
.A(n_1328),
.Y(n_1731)
);

BUFx8_ASAP7_75t_L g1732 ( 
.A(n_1293),
.Y(n_1732)
);

AND2x4_ASAP7_75t_L g1733 ( 
.A(n_1615),
.B(n_1106),
.Y(n_1733)
);

NOR2xp33_ASAP7_75t_SL g1734 ( 
.A(n_1312),
.B(n_861),
.Y(n_1734)
);

CKINVDCx5p33_ASAP7_75t_R g1735 ( 
.A(n_1430),
.Y(n_1735)
);

BUFx8_ASAP7_75t_SL g1736 ( 
.A(n_1277),
.Y(n_1736)
);

INVx3_ASAP7_75t_L g1737 ( 
.A(n_1385),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1640),
.B(n_1029),
.Y(n_1738)
);

BUFx6f_ASAP7_75t_L g1739 ( 
.A(n_1354),
.Y(n_1739)
);

BUFx6f_ASAP7_75t_L g1740 ( 
.A(n_1354),
.Y(n_1740)
);

BUFx6f_ASAP7_75t_L g1741 ( 
.A(n_1354),
.Y(n_1741)
);

AND2x4_ASAP7_75t_L g1742 ( 
.A(n_1615),
.B(n_1171),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_1273),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1417),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1667),
.B(n_1032),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1650),
.B(n_861),
.Y(n_1746)
);

AND2x4_ASAP7_75t_L g1747 ( 
.A(n_1691),
.B(n_1171),
.Y(n_1747)
);

BUFx6f_ASAP7_75t_L g1748 ( 
.A(n_1424),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1278),
.Y(n_1749)
);

AND2x4_ASAP7_75t_L g1750 ( 
.A(n_1691),
.B(n_1217),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1410),
.B(n_1421),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1518),
.B(n_861),
.Y(n_1752)
);

NOR2xp33_ASAP7_75t_L g1753 ( 
.A(n_1590),
.B(n_1217),
.Y(n_1753)
);

BUFx2_ASAP7_75t_L g1754 ( 
.A(n_1321),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1278),
.Y(n_1755)
);

INVx2_ASAP7_75t_L g1756 ( 
.A(n_1286),
.Y(n_1756)
);

NOR2xp33_ASAP7_75t_SL g1757 ( 
.A(n_1394),
.B(n_861),
.Y(n_1757)
);

BUFx8_ASAP7_75t_SL g1758 ( 
.A(n_1277),
.Y(n_1758)
);

CKINVDCx6p67_ASAP7_75t_R g1759 ( 
.A(n_1547),
.Y(n_1759)
);

BUFx6f_ASAP7_75t_L g1760 ( 
.A(n_1424),
.Y(n_1760)
);

BUFx6f_ASAP7_75t_L g1761 ( 
.A(n_1424),
.Y(n_1761)
);

NOR2xp33_ASAP7_75t_L g1762 ( 
.A(n_1600),
.B(n_833),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1670),
.B(n_1038),
.Y(n_1763)
);

AND2x4_ASAP7_75t_L g1764 ( 
.A(n_1281),
.B(n_863),
.Y(n_1764)
);

INVx4_ASAP7_75t_L g1765 ( 
.A(n_1431),
.Y(n_1765)
);

BUFx6f_ASAP7_75t_L g1766 ( 
.A(n_1482),
.Y(n_1766)
);

BUFx8_ASAP7_75t_SL g1767 ( 
.A(n_1287),
.Y(n_1767)
);

BUFx6f_ASAP7_75t_L g1768 ( 
.A(n_1482),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1545),
.B(n_1033),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1420),
.Y(n_1770)
);

INVxp67_ASAP7_75t_L g1771 ( 
.A(n_1570),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1286),
.Y(n_1772)
);

AND2x4_ASAP7_75t_L g1773 ( 
.A(n_1281),
.B(n_863),
.Y(n_1773)
);

BUFx12f_ASAP7_75t_L g1774 ( 
.A(n_1327),
.Y(n_1774)
);

INVx3_ASAP7_75t_L g1775 ( 
.A(n_1482),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1310),
.Y(n_1776)
);

NOR2xp33_ASAP7_75t_L g1777 ( 
.A(n_1623),
.B(n_1393),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1694),
.B(n_1059),
.Y(n_1778)
);

BUFx6f_ASAP7_75t_L g1779 ( 
.A(n_1482),
.Y(n_1779)
);

BUFx6f_ASAP7_75t_L g1780 ( 
.A(n_1591),
.Y(n_1780)
);

BUFx8_ASAP7_75t_SL g1781 ( 
.A(n_1287),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1310),
.Y(n_1782)
);

NOR2xp33_ASAP7_75t_L g1783 ( 
.A(n_1333),
.B(n_837),
.Y(n_1783)
);

NOR2xp33_ASAP7_75t_L g1784 ( 
.A(n_1335),
.B(n_839),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1422),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_SL g1786 ( 
.A(n_1379),
.B(n_1033),
.Y(n_1786)
);

BUFx6f_ASAP7_75t_L g1787 ( 
.A(n_1591),
.Y(n_1787)
);

AND2x6_ASAP7_75t_L g1788 ( 
.A(n_1263),
.B(n_946),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1468),
.B(n_1064),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1594),
.B(n_1033),
.Y(n_1790)
);

BUFx6f_ASAP7_75t_L g1791 ( 
.A(n_1673),
.Y(n_1791)
);

BUFx12f_ASAP7_75t_L g1792 ( 
.A(n_1327),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_1324),
.Y(n_1793)
);

NOR2xp33_ASAP7_75t_SL g1794 ( 
.A(n_1552),
.B(n_1033),
.Y(n_1794)
);

BUFx12f_ASAP7_75t_L g1795 ( 
.A(n_1259),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1472),
.B(n_1082),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1475),
.B(n_1113),
.Y(n_1797)
);

XNOR2xp5_ASAP7_75t_L g1798 ( 
.A(n_1299),
.B(n_1241),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1493),
.B(n_1119),
.Y(n_1799)
);

BUFx2_ASAP7_75t_L g1800 ( 
.A(n_1328),
.Y(n_1800)
);

INVx2_ASAP7_75t_L g1801 ( 
.A(n_1324),
.Y(n_1801)
);

INVx3_ASAP7_75t_L g1802 ( 
.A(n_1673),
.Y(n_1802)
);

NOR2xp33_ASAP7_75t_L g1803 ( 
.A(n_1337),
.B(n_840),
.Y(n_1803)
);

AND2x4_ASAP7_75t_L g1804 ( 
.A(n_1288),
.B(n_915),
.Y(n_1804)
);

INVx2_ASAP7_75t_L g1805 ( 
.A(n_1349),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1487),
.B(n_1060),
.Y(n_1806)
);

BUFx12f_ASAP7_75t_L g1807 ( 
.A(n_1259),
.Y(n_1807)
);

BUFx2_ASAP7_75t_L g1808 ( 
.A(n_1331),
.Y(n_1808)
);

NOR2xp33_ASAP7_75t_L g1809 ( 
.A(n_1527),
.B(n_844),
.Y(n_1809)
);

BUFx6f_ASAP7_75t_L g1810 ( 
.A(n_1673),
.Y(n_1810)
);

AND2x6_ASAP7_75t_L g1811 ( 
.A(n_1263),
.B(n_946),
.Y(n_1811)
);

BUFx6f_ASAP7_75t_L g1812 ( 
.A(n_1689),
.Y(n_1812)
);

BUFx6f_ASAP7_75t_L g1813 ( 
.A(n_1689),
.Y(n_1813)
);

INVx2_ASAP7_75t_L g1814 ( 
.A(n_1349),
.Y(n_1814)
);

CKINVDCx6p67_ASAP7_75t_R g1815 ( 
.A(n_1565),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1350),
.Y(n_1816)
);

BUFx6f_ASAP7_75t_L g1817 ( 
.A(n_1689),
.Y(n_1817)
);

BUFx6f_ASAP7_75t_L g1818 ( 
.A(n_1689),
.Y(n_1818)
);

INVx5_ASAP7_75t_L g1819 ( 
.A(n_1496),
.Y(n_1819)
);

BUFx6f_ASAP7_75t_L g1820 ( 
.A(n_1350),
.Y(n_1820)
);

BUFx3_ASAP7_75t_L g1821 ( 
.A(n_1261),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1426),
.B(n_1132),
.Y(n_1822)
);

AND2x4_ASAP7_75t_L g1823 ( 
.A(n_1288),
.B(n_915),
.Y(n_1823)
);

BUFx12f_ASAP7_75t_L g1824 ( 
.A(n_1301),
.Y(n_1824)
);

HB1xp67_ASAP7_75t_L g1825 ( 
.A(n_1261),
.Y(n_1825)
);

BUFx6f_ASAP7_75t_L g1826 ( 
.A(n_1358),
.Y(n_1826)
);

AND2x4_ASAP7_75t_L g1827 ( 
.A(n_1377),
.B(n_1396),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1428),
.Y(n_1828)
);

CKINVDCx5p33_ASAP7_75t_R g1829 ( 
.A(n_1436),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_SL g1830 ( 
.A(n_1379),
.B(n_1060),
.Y(n_1830)
);

INVx2_ASAP7_75t_L g1831 ( 
.A(n_1358),
.Y(n_1831)
);

NOR2xp33_ASAP7_75t_L g1832 ( 
.A(n_1355),
.B(n_846),
.Y(n_1832)
);

NOR2xp33_ASAP7_75t_L g1833 ( 
.A(n_1345),
.B(n_850),
.Y(n_1833)
);

BUFx6f_ASAP7_75t_L g1834 ( 
.A(n_1369),
.Y(n_1834)
);

INVx3_ASAP7_75t_L g1835 ( 
.A(n_1369),
.Y(n_1835)
);

INVx5_ASAP7_75t_L g1836 ( 
.A(n_1496),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1429),
.B(n_1144),
.Y(n_1837)
);

BUFx12f_ASAP7_75t_L g1838 ( 
.A(n_1301),
.Y(n_1838)
);

BUFx6f_ASAP7_75t_L g1839 ( 
.A(n_1398),
.Y(n_1839)
);

INVx5_ASAP7_75t_L g1840 ( 
.A(n_1496),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1432),
.B(n_1151),
.Y(n_1841)
);

NOR2xp33_ASAP7_75t_L g1842 ( 
.A(n_1351),
.B(n_1352),
.Y(n_1842)
);

NOR2xp33_ASAP7_75t_L g1843 ( 
.A(n_1352),
.B(n_1400),
.Y(n_1843)
);

INVx2_ASAP7_75t_SL g1844 ( 
.A(n_1331),
.Y(n_1844)
);

INVx6_ASAP7_75t_L g1845 ( 
.A(n_1268),
.Y(n_1845)
);

INVx2_ASAP7_75t_L g1846 ( 
.A(n_1398),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1419),
.B(n_1060),
.Y(n_1847)
);

INVx3_ASAP7_75t_L g1848 ( 
.A(n_1413),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1437),
.B(n_1161),
.Y(n_1849)
);

INVx4_ASAP7_75t_L g1850 ( 
.A(n_1538),
.Y(n_1850)
);

BUFx6f_ASAP7_75t_L g1851 ( 
.A(n_1413),
.Y(n_1851)
);

BUFx6f_ASAP7_75t_L g1852 ( 
.A(n_1418),
.Y(n_1852)
);

INVx2_ASAP7_75t_L g1853 ( 
.A(n_1418),
.Y(n_1853)
);

BUFx6f_ASAP7_75t_L g1854 ( 
.A(n_1438),
.Y(n_1854)
);

CKINVDCx5p33_ASAP7_75t_R g1855 ( 
.A(n_1582),
.Y(n_1855)
);

AND2x2_ASAP7_75t_L g1856 ( 
.A(n_1419),
.B(n_1060),
.Y(n_1856)
);

BUFx6f_ASAP7_75t_L g1857 ( 
.A(n_1438),
.Y(n_1857)
);

HB1xp67_ASAP7_75t_L g1858 ( 
.A(n_1268),
.Y(n_1858)
);

AND2x4_ASAP7_75t_L g1859 ( 
.A(n_1377),
.B(n_931),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1440),
.Y(n_1860)
);

BUFx6f_ASAP7_75t_L g1861 ( 
.A(n_1439),
.Y(n_1861)
);

INVx2_ASAP7_75t_SL g1862 ( 
.A(n_1344),
.Y(n_1862)
);

INVx3_ASAP7_75t_L g1863 ( 
.A(n_1439),
.Y(n_1863)
);

BUFx12f_ASAP7_75t_L g1864 ( 
.A(n_1344),
.Y(n_1864)
);

AND2x4_ASAP7_75t_L g1865 ( 
.A(n_1396),
.B(n_1434),
.Y(n_1865)
);

INVxp67_ASAP7_75t_L g1866 ( 
.A(n_1601),
.Y(n_1866)
);

INVx5_ASAP7_75t_L g1867 ( 
.A(n_1441),
.Y(n_1867)
);

BUFx8_ASAP7_75t_SL g1868 ( 
.A(n_1299),
.Y(n_1868)
);

INVx2_ASAP7_75t_L g1869 ( 
.A(n_1441),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1442),
.Y(n_1870)
);

BUFx6f_ASAP7_75t_L g1871 ( 
.A(n_1446),
.Y(n_1871)
);

BUFx6f_ASAP7_75t_L g1872 ( 
.A(n_1446),
.Y(n_1872)
);

BUFx8_ASAP7_75t_L g1873 ( 
.A(n_1293),
.Y(n_1873)
);

BUFx6f_ASAP7_75t_L g1874 ( 
.A(n_1443),
.Y(n_1874)
);

AND2x4_ASAP7_75t_L g1875 ( 
.A(n_1434),
.B(n_931),
.Y(n_1875)
);

NOR2xp33_ASAP7_75t_L g1876 ( 
.A(n_1400),
.B(n_851),
.Y(n_1876)
);

INVxp67_ASAP7_75t_L g1877 ( 
.A(n_1533),
.Y(n_1877)
);

BUFx6f_ASAP7_75t_L g1878 ( 
.A(n_1444),
.Y(n_1878)
);

INVx6_ASAP7_75t_L g1879 ( 
.A(n_1456),
.Y(n_1879)
);

AND2x2_ASAP7_75t_L g1880 ( 
.A(n_1489),
.B(n_1091),
.Y(n_1880)
);

INVx5_ASAP7_75t_L g1881 ( 
.A(n_1458),
.Y(n_1881)
);

HB1xp67_ASAP7_75t_L g1882 ( 
.A(n_1346),
.Y(n_1882)
);

INVx3_ASAP7_75t_L g1883 ( 
.A(n_1458),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1445),
.Y(n_1884)
);

BUFx6f_ASAP7_75t_L g1885 ( 
.A(n_1447),
.Y(n_1885)
);

BUFx12f_ASAP7_75t_L g1886 ( 
.A(n_1346),
.Y(n_1886)
);

BUFx3_ASAP7_75t_L g1887 ( 
.A(n_1374),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1489),
.B(n_1091),
.Y(n_1888)
);

HB1xp67_ASAP7_75t_L g1889 ( 
.A(n_1347),
.Y(n_1889)
);

BUFx6f_ASAP7_75t_L g1890 ( 
.A(n_1449),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1450),
.Y(n_1891)
);

INVx2_ASAP7_75t_L g1892 ( 
.A(n_1451),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1269),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_L g1894 ( 
.A(n_1255),
.B(n_1168),
.Y(n_1894)
);

BUFx8_ASAP7_75t_SL g1895 ( 
.A(n_1320),
.Y(n_1895)
);

HB1xp67_ASAP7_75t_L g1896 ( 
.A(n_1347),
.Y(n_1896)
);

AND2x4_ASAP7_75t_L g1897 ( 
.A(n_1497),
.B(n_937),
.Y(n_1897)
);

AND2x2_ASAP7_75t_L g1898 ( 
.A(n_1562),
.B(n_1091),
.Y(n_1898)
);

BUFx6f_ASAP7_75t_L g1899 ( 
.A(n_1459),
.Y(n_1899)
);

INVxp67_ASAP7_75t_L g1900 ( 
.A(n_1548),
.Y(n_1900)
);

BUFx12f_ASAP7_75t_L g1901 ( 
.A(n_1414),
.Y(n_1901)
);

AND2x4_ASAP7_75t_L g1902 ( 
.A(n_1497),
.B(n_937),
.Y(n_1902)
);

CKINVDCx14_ASAP7_75t_R g1903 ( 
.A(n_1562),
.Y(n_1903)
);

INVx3_ASAP7_75t_L g1904 ( 
.A(n_1459),
.Y(n_1904)
);

BUFx3_ASAP7_75t_L g1905 ( 
.A(n_1376),
.Y(n_1905)
);

AND2x4_ASAP7_75t_L g1906 ( 
.A(n_1500),
.B(n_964),
.Y(n_1906)
);

BUFx12f_ASAP7_75t_L g1907 ( 
.A(n_1414),
.Y(n_1907)
);

BUFx6f_ASAP7_75t_L g1908 ( 
.A(n_1469),
.Y(n_1908)
);

BUFx3_ASAP7_75t_L g1909 ( 
.A(n_1378),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_SL g1910 ( 
.A(n_1379),
.B(n_1091),
.Y(n_1910)
);

AND2x2_ASAP7_75t_L g1911 ( 
.A(n_1500),
.B(n_1105),
.Y(n_1911)
);

INVx2_ASAP7_75t_L g1912 ( 
.A(n_1257),
.Y(n_1912)
);

INVx2_ASAP7_75t_L g1913 ( 
.A(n_1258),
.Y(n_1913)
);

BUFx12f_ASAP7_75t_L g1914 ( 
.A(n_1474),
.Y(n_1914)
);

CKINVDCx5p33_ASAP7_75t_R g1915 ( 
.A(n_1585),
.Y(n_1915)
);

HB1xp67_ASAP7_75t_L g1916 ( 
.A(n_1474),
.Y(n_1916)
);

CKINVDCx5p33_ASAP7_75t_R g1917 ( 
.A(n_1629),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_L g1918 ( 
.A(n_1260),
.B(n_1262),
.Y(n_1918)
);

NOR2xp33_ASAP7_75t_L g1919 ( 
.A(n_1454),
.B(n_853),
.Y(n_1919)
);

HB1xp67_ASAP7_75t_L g1920 ( 
.A(n_1476),
.Y(n_1920)
);

BUFx6f_ASAP7_75t_L g1921 ( 
.A(n_1469),
.Y(n_1921)
);

AND2x4_ASAP7_75t_L g1922 ( 
.A(n_1567),
.B(n_964),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1270),
.Y(n_1923)
);

BUFx2_ASAP7_75t_L g1924 ( 
.A(n_1476),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_SL g1925 ( 
.A(n_1379),
.B(n_1105),
.Y(n_1925)
);

INVx5_ASAP7_75t_L g1926 ( 
.A(n_1471),
.Y(n_1926)
);

NOR2xp33_ASAP7_75t_L g1927 ( 
.A(n_1454),
.B(n_854),
.Y(n_1927)
);

INVx5_ASAP7_75t_L g1928 ( 
.A(n_1471),
.Y(n_1928)
);

BUFx6f_ASAP7_75t_L g1929 ( 
.A(n_1503),
.Y(n_1929)
);

NOR2xp33_ASAP7_75t_SL g1930 ( 
.A(n_1586),
.B(n_1105),
.Y(n_1930)
);

NOR2xp33_ASAP7_75t_L g1931 ( 
.A(n_1455),
.B(n_855),
.Y(n_1931)
);

INVx2_ASAP7_75t_L g1932 ( 
.A(n_1264),
.Y(n_1932)
);

CKINVDCx6p67_ASAP7_75t_R g1933 ( 
.A(n_1683),
.Y(n_1933)
);

INVx3_ASAP7_75t_L g1934 ( 
.A(n_1503),
.Y(n_1934)
);

AND2x2_ASAP7_75t_L g1935 ( 
.A(n_1567),
.B(n_1571),
.Y(n_1935)
);

BUFx12f_ASAP7_75t_L g1936 ( 
.A(n_1480),
.Y(n_1936)
);

BUFx6f_ASAP7_75t_L g1937 ( 
.A(n_1514),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1271),
.Y(n_1938)
);

CKINVDCx5p33_ASAP7_75t_R g1939 ( 
.A(n_1695),
.Y(n_1939)
);

INVx2_ASAP7_75t_L g1940 ( 
.A(n_1265),
.Y(n_1940)
);

CKINVDCx5p33_ASAP7_75t_R g1941 ( 
.A(n_1499),
.Y(n_1941)
);

BUFx12f_ASAP7_75t_L g1942 ( 
.A(n_1480),
.Y(n_1942)
);

BUFx2_ASAP7_75t_L g1943 ( 
.A(n_1505),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_L g1944 ( 
.A(n_1266),
.B(n_1182),
.Y(n_1944)
);

INVx2_ASAP7_75t_L g1945 ( 
.A(n_1514),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1274),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_L g1947 ( 
.A(n_1379),
.B(n_1191),
.Y(n_1947)
);

INVx2_ASAP7_75t_L g1948 ( 
.A(n_1515),
.Y(n_1948)
);

AND2x4_ASAP7_75t_L g1949 ( 
.A(n_1571),
.B(n_974),
.Y(n_1949)
);

INVx5_ASAP7_75t_L g1950 ( 
.A(n_1515),
.Y(n_1950)
);

BUFx6f_ASAP7_75t_L g1951 ( 
.A(n_1543),
.Y(n_1951)
);

BUFx6f_ASAP7_75t_L g1952 ( 
.A(n_1543),
.Y(n_1952)
);

HB1xp67_ASAP7_75t_L g1953 ( 
.A(n_1505),
.Y(n_1953)
);

BUFx6f_ASAP7_75t_L g1954 ( 
.A(n_1589),
.Y(n_1954)
);

AND2x2_ASAP7_75t_L g1955 ( 
.A(n_1577),
.B(n_1105),
.Y(n_1955)
);

AND2x2_ASAP7_75t_L g1956 ( 
.A(n_1577),
.B(n_1180),
.Y(n_1956)
);

BUFx6f_ASAP7_75t_L g1957 ( 
.A(n_1589),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_L g1958 ( 
.A(n_1275),
.B(n_1192),
.Y(n_1958)
);

BUFx6f_ASAP7_75t_L g1959 ( 
.A(n_1592),
.Y(n_1959)
);

BUFx6f_ASAP7_75t_L g1960 ( 
.A(n_1592),
.Y(n_1960)
);

BUFx6f_ASAP7_75t_L g1961 ( 
.A(n_1603),
.Y(n_1961)
);

INVx5_ASAP7_75t_L g1962 ( 
.A(n_1603),
.Y(n_1962)
);

NOR2xp33_ASAP7_75t_L g1963 ( 
.A(n_1455),
.B(n_859),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1276),
.Y(n_1964)
);

NOR2xp33_ASAP7_75t_L g1965 ( 
.A(n_1457),
.B(n_1490),
.Y(n_1965)
);

AND2x2_ASAP7_75t_L g1966 ( 
.A(n_1578),
.B(n_1180),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1279),
.Y(n_1967)
);

AND2x6_ASAP7_75t_L g1968 ( 
.A(n_1280),
.B(n_946),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1284),
.B(n_1200),
.Y(n_1969)
);

INVx2_ASAP7_75t_L g1970 ( 
.A(n_1608),
.Y(n_1970)
);

BUFx3_ASAP7_75t_L g1971 ( 
.A(n_1382),
.Y(n_1971)
);

NOR2xp33_ASAP7_75t_SL g1972 ( 
.A(n_1338),
.B(n_1180),
.Y(n_1972)
);

NOR2xp33_ASAP7_75t_L g1973 ( 
.A(n_1457),
.B(n_1490),
.Y(n_1973)
);

NOR2xp33_ASAP7_75t_L g1974 ( 
.A(n_1491),
.B(n_860),
.Y(n_1974)
);

INVx5_ASAP7_75t_L g1975 ( 
.A(n_1608),
.Y(n_1975)
);

AND2x4_ASAP7_75t_L g1976 ( 
.A(n_1578),
.B(n_974),
.Y(n_1976)
);

BUFx12f_ASAP7_75t_L g1977 ( 
.A(n_1508),
.Y(n_1977)
);

AND2x4_ASAP7_75t_L g1978 ( 
.A(n_1318),
.B(n_1549),
.Y(n_1978)
);

BUFx8_ASAP7_75t_L g1979 ( 
.A(n_1318),
.Y(n_1979)
);

INVx3_ASAP7_75t_L g1980 ( 
.A(n_1612),
.Y(n_1980)
);

AND2x6_ASAP7_75t_L g1981 ( 
.A(n_1285),
.B(n_976),
.Y(n_1981)
);

INVx5_ASAP7_75t_L g1982 ( 
.A(n_1612),
.Y(n_1982)
);

BUFx6f_ASAP7_75t_L g1983 ( 
.A(n_1617),
.Y(n_1983)
);

INVx5_ASAP7_75t_L g1984 ( 
.A(n_1617),
.Y(n_1984)
);

BUFx8_ASAP7_75t_SL g1985 ( 
.A(n_1320),
.Y(n_1985)
);

INVx5_ASAP7_75t_L g1986 ( 
.A(n_1674),
.Y(n_1986)
);

BUFx6f_ASAP7_75t_L g1987 ( 
.A(n_1674),
.Y(n_1987)
);

BUFx2_ASAP7_75t_L g1988 ( 
.A(n_1508),
.Y(n_1988)
);

AND2x4_ASAP7_75t_L g1989 ( 
.A(n_1549),
.B(n_1645),
.Y(n_1989)
);

AND2x2_ASAP7_75t_L g1990 ( 
.A(n_1509),
.B(n_1180),
.Y(n_1990)
);

BUFx8_ASAP7_75t_L g1991 ( 
.A(n_1645),
.Y(n_1991)
);

BUFx8_ASAP7_75t_SL g1992 ( 
.A(n_1330),
.Y(n_1992)
);

INVx5_ASAP7_75t_L g1993 ( 
.A(n_1697),
.Y(n_1993)
);

NOR2xp33_ASAP7_75t_L g1994 ( 
.A(n_1491),
.B(n_862),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1289),
.B(n_1206),
.Y(n_1995)
);

BUFx8_ASAP7_75t_SL g1996 ( 
.A(n_1330),
.Y(n_1996)
);

AND2x4_ASAP7_75t_L g1997 ( 
.A(n_1647),
.B(n_976),
.Y(n_1997)
);

BUFx2_ASAP7_75t_L g1998 ( 
.A(n_1509),
.Y(n_1998)
);

AND2x6_ASAP7_75t_L g1999 ( 
.A(n_1290),
.B(n_997),
.Y(n_1999)
);

NOR2x1_ASAP7_75t_L g2000 ( 
.A(n_1291),
.B(n_997),
.Y(n_2000)
);

AND2x4_ASAP7_75t_L g2001 ( 
.A(n_1647),
.B(n_1013),
.Y(n_2001)
);

NOR2xp33_ASAP7_75t_SL g2002 ( 
.A(n_1370),
.B(n_1246),
.Y(n_2002)
);

INVx5_ASAP7_75t_L g2003 ( 
.A(n_1697),
.Y(n_2003)
);

AND2x4_ASAP7_75t_L g2004 ( 
.A(n_1383),
.B(n_1013),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1292),
.Y(n_2005)
);

NOR2xp33_ASAP7_75t_L g2006 ( 
.A(n_1498),
.B(n_865),
.Y(n_2006)
);

AND2x4_ASAP7_75t_L g2007 ( 
.A(n_1384),
.B(n_1027),
.Y(n_2007)
);

HB1xp67_ASAP7_75t_L g2008 ( 
.A(n_1512),
.Y(n_2008)
);

INVx2_ASAP7_75t_L g2009 ( 
.A(n_1453),
.Y(n_2009)
);

INVx3_ASAP7_75t_L g2010 ( 
.A(n_1465),
.Y(n_2010)
);

AND2x2_ASAP7_75t_L g2011 ( 
.A(n_1512),
.B(n_1246),
.Y(n_2011)
);

INVx5_ASAP7_75t_L g2012 ( 
.A(n_1425),
.Y(n_2012)
);

BUFx6f_ASAP7_75t_L g2013 ( 
.A(n_1466),
.Y(n_2013)
);

AND2x6_ASAP7_75t_L g2014 ( 
.A(n_1295),
.B(n_1027),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_L g2015 ( 
.A(n_1296),
.B(n_1212),
.Y(n_2015)
);

AND2x2_ASAP7_75t_L g2016 ( 
.A(n_1523),
.B(n_1246),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1297),
.Y(n_2017)
);

BUFx6f_ASAP7_75t_L g2018 ( 
.A(n_1467),
.Y(n_2018)
);

CKINVDCx5p33_ASAP7_75t_R g2019 ( 
.A(n_1557),
.Y(n_2019)
);

BUFx8_ASAP7_75t_L g2020 ( 
.A(n_1386),
.Y(n_2020)
);

BUFx6f_ASAP7_75t_L g2021 ( 
.A(n_1470),
.Y(n_2021)
);

INVx5_ASAP7_75t_L g2022 ( 
.A(n_1699),
.Y(n_2022)
);

BUFx8_ASAP7_75t_SL g2023 ( 
.A(n_1360),
.Y(n_2023)
);

BUFx6f_ASAP7_75t_L g2024 ( 
.A(n_1473),
.Y(n_2024)
);

BUFx6f_ASAP7_75t_L g2025 ( 
.A(n_1477),
.Y(n_2025)
);

INVx5_ASAP7_75t_L g2026 ( 
.A(n_1699),
.Y(n_2026)
);

INVx5_ASAP7_75t_L g2027 ( 
.A(n_1300),
.Y(n_2027)
);

BUFx6f_ASAP7_75t_L g2028 ( 
.A(n_1479),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_L g2029 ( 
.A(n_1303),
.B(n_1304),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1305),
.Y(n_2030)
);

AND2x2_ASAP7_75t_L g2031 ( 
.A(n_1523),
.B(n_1246),
.Y(n_2031)
);

HB1xp67_ASAP7_75t_L g2032 ( 
.A(n_1530),
.Y(n_2032)
);

BUFx3_ASAP7_75t_L g2033 ( 
.A(n_1387),
.Y(n_2033)
);

BUFx8_ASAP7_75t_SL g2034 ( 
.A(n_1360),
.Y(n_2034)
);

BUFx12f_ASAP7_75t_L g2035 ( 
.A(n_1530),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_1307),
.B(n_1214),
.Y(n_2036)
);

INVx2_ASAP7_75t_L g2037 ( 
.A(n_1460),
.Y(n_2037)
);

INVx2_ASAP7_75t_L g2038 ( 
.A(n_1461),
.Y(n_2038)
);

AND2x2_ASAP7_75t_L g2039 ( 
.A(n_1532),
.B(n_941),
.Y(n_2039)
);

NOR2xp33_ASAP7_75t_L g2040 ( 
.A(n_1498),
.B(n_866),
.Y(n_2040)
);

INVx5_ASAP7_75t_L g2041 ( 
.A(n_1308),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_L g2042 ( 
.A(n_1311),
.B(n_1231),
.Y(n_2042)
);

INVx3_ASAP7_75t_L g2043 ( 
.A(n_1481),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_L g2044 ( 
.A(n_1313),
.B(n_1314),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_L g2045 ( 
.A(n_1315),
.B(n_1247),
.Y(n_2045)
);

BUFx6f_ASAP7_75t_L g2046 ( 
.A(n_1484),
.Y(n_2046)
);

INVx5_ASAP7_75t_L g2047 ( 
.A(n_1316),
.Y(n_2047)
);

BUFx6f_ASAP7_75t_L g2048 ( 
.A(n_1485),
.Y(n_2048)
);

INVx2_ASAP7_75t_L g2049 ( 
.A(n_1464),
.Y(n_2049)
);

BUFx6f_ASAP7_75t_L g2050 ( 
.A(n_1486),
.Y(n_2050)
);

BUFx12f_ASAP7_75t_L g2051 ( 
.A(n_1532),
.Y(n_2051)
);

NOR2xp33_ASAP7_75t_L g2052 ( 
.A(n_1566),
.B(n_867),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1317),
.Y(n_2053)
);

BUFx6f_ASAP7_75t_L g2054 ( 
.A(n_1488),
.Y(n_2054)
);

BUFx6f_ASAP7_75t_L g2055 ( 
.A(n_1492),
.Y(n_2055)
);

NAND2xp5_ASAP7_75t_L g2056 ( 
.A(n_1319),
.B(n_1322),
.Y(n_2056)
);

AND2x2_ASAP7_75t_L g2057 ( 
.A(n_1537),
.B(n_987),
.Y(n_2057)
);

AND2x4_ASAP7_75t_L g2058 ( 
.A(n_1388),
.B(n_1112),
.Y(n_2058)
);

OR2x2_ASAP7_75t_L g2059 ( 
.A(n_1389),
.B(n_1390),
.Y(n_2059)
);

NOR2xp33_ASAP7_75t_L g2060 ( 
.A(n_1566),
.B(n_868),
.Y(n_2060)
);

INVx2_ASAP7_75t_L g2061 ( 
.A(n_1501),
.Y(n_2061)
);

BUFx6f_ASAP7_75t_L g2062 ( 
.A(n_1510),
.Y(n_2062)
);

AND2x4_ASAP7_75t_L g2063 ( 
.A(n_1391),
.B(n_1112),
.Y(n_2063)
);

BUFx6f_ASAP7_75t_L g2064 ( 
.A(n_1716),
.Y(n_2064)
);

INVx2_ASAP7_75t_L g2065 ( 
.A(n_1703),
.Y(n_2065)
);

INVxp67_ASAP7_75t_L g2066 ( 
.A(n_1715),
.Y(n_2066)
);

NAND2xp5_ASAP7_75t_L g2067 ( 
.A(n_1730),
.B(n_1323),
.Y(n_2067)
);

INVx2_ASAP7_75t_L g2068 ( 
.A(n_1709),
.Y(n_2068)
);

AND2x4_ASAP7_75t_L g2069 ( 
.A(n_1821),
.B(n_1827),
.Y(n_2069)
);

BUFx6f_ASAP7_75t_L g2070 ( 
.A(n_1716),
.Y(n_2070)
);

BUFx2_ASAP7_75t_L g2071 ( 
.A(n_1715),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_1893),
.Y(n_2072)
);

INVx3_ASAP7_75t_L g2073 ( 
.A(n_1716),
.Y(n_2073)
);

AND2x2_ASAP7_75t_L g2074 ( 
.A(n_1746),
.B(n_1272),
.Y(n_2074)
);

BUFx6f_ASAP7_75t_L g2075 ( 
.A(n_1721),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_1923),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_L g2077 ( 
.A(n_1730),
.B(n_1325),
.Y(n_2077)
);

INVx3_ASAP7_75t_L g2078 ( 
.A(n_1721),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_1938),
.Y(n_2079)
);

BUFx6f_ASAP7_75t_L g2080 ( 
.A(n_1721),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_L g2081 ( 
.A(n_1738),
.B(n_1332),
.Y(n_2081)
);

AND2x4_ASAP7_75t_L g2082 ( 
.A(n_1821),
.B(n_1334),
.Y(n_2082)
);

HB1xp67_ASAP7_75t_L g2083 ( 
.A(n_1705),
.Y(n_2083)
);

BUFx6f_ASAP7_75t_L g2084 ( 
.A(n_1724),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_1946),
.Y(n_2085)
);

AND3x1_ASAP7_75t_L g2086 ( 
.A(n_1702),
.B(n_1063),
.C(n_1062),
.Y(n_2086)
);

AND3x2_ASAP7_75t_L g2087 ( 
.A(n_1757),
.B(n_1930),
.C(n_1794),
.Y(n_2087)
);

HB1xp67_ASAP7_75t_L g2088 ( 
.A(n_1705),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_1964),
.Y(n_2089)
);

AND2x4_ASAP7_75t_L g2090 ( 
.A(n_1764),
.B(n_1339),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_1967),
.Y(n_2091)
);

INVx2_ASAP7_75t_L g2092 ( 
.A(n_1720),
.Y(n_2092)
);

INVx2_ASAP7_75t_L g2093 ( 
.A(n_1743),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_2005),
.Y(n_2094)
);

INVx5_ASAP7_75t_L g2095 ( 
.A(n_1788),
.Y(n_2095)
);

BUFx6f_ASAP7_75t_L g2096 ( 
.A(n_1724),
.Y(n_2096)
);

AND2x6_ASAP7_75t_L g2097 ( 
.A(n_1847),
.B(n_1340),
.Y(n_2097)
);

INVx2_ASAP7_75t_L g2098 ( 
.A(n_1749),
.Y(n_2098)
);

OR2x6_ASAP7_75t_L g2099 ( 
.A(n_1774),
.B(n_1602),
.Y(n_2099)
);

INVx3_ASAP7_75t_L g2100 ( 
.A(n_1724),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_SL g2101 ( 
.A(n_2012),
.B(n_1537),
.Y(n_2101)
);

BUFx6f_ASAP7_75t_L g2102 ( 
.A(n_1739),
.Y(n_2102)
);

INVx6_ASAP7_75t_L g2103 ( 
.A(n_1845),
.Y(n_2103)
);

BUFx6f_ASAP7_75t_L g2104 ( 
.A(n_1739),
.Y(n_2104)
);

AND2x2_ASAP7_75t_L g2105 ( 
.A(n_1978),
.B(n_1272),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_L g2106 ( 
.A(n_1738),
.B(n_1342),
.Y(n_2106)
);

AND2x4_ASAP7_75t_L g2107 ( 
.A(n_1827),
.B(n_1392),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_2017),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_2030),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_2053),
.Y(n_2110)
);

AND2x2_ASAP7_75t_L g2111 ( 
.A(n_1978),
.B(n_1282),
.Y(n_2111)
);

INVx2_ASAP7_75t_L g2112 ( 
.A(n_1755),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_1887),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_1887),
.Y(n_2114)
);

AND2x4_ASAP7_75t_L g2115 ( 
.A(n_1865),
.B(n_1397),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_1905),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_1905),
.Y(n_2117)
);

BUFx8_ASAP7_75t_L g2118 ( 
.A(n_1795),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_1909),
.Y(n_2119)
);

INVx3_ASAP7_75t_L g2120 ( 
.A(n_1739),
.Y(n_2120)
);

BUFx6f_ASAP7_75t_L g2121 ( 
.A(n_1740),
.Y(n_2121)
);

NAND2xp33_ASAP7_75t_L g2122 ( 
.A(n_1981),
.B(n_1542),
.Y(n_2122)
);

INVx1_ASAP7_75t_SL g2123 ( 
.A(n_1736),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_1909),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_1971),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_1971),
.Y(n_2126)
);

NAND2xp5_ASAP7_75t_L g2127 ( 
.A(n_1745),
.B(n_1343),
.Y(n_2127)
);

AND2x2_ASAP7_75t_L g2128 ( 
.A(n_1989),
.B(n_1282),
.Y(n_2128)
);

BUFx6f_ASAP7_75t_L g2129 ( 
.A(n_1740),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_2033),
.Y(n_2130)
);

HB1xp67_ASAP7_75t_L g2131 ( 
.A(n_1825),
.Y(n_2131)
);

NOR2xp33_ASAP7_75t_L g2132 ( 
.A(n_1877),
.B(n_1573),
.Y(n_2132)
);

INVx3_ASAP7_75t_L g2133 ( 
.A(n_1740),
.Y(n_2133)
);

NAND2xp5_ASAP7_75t_L g2134 ( 
.A(n_1745),
.B(n_1348),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_2033),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_L g2136 ( 
.A(n_1763),
.B(n_1353),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_1912),
.Y(n_2137)
);

INVx2_ASAP7_75t_L g2138 ( 
.A(n_1756),
.Y(n_2138)
);

BUFx6f_ASAP7_75t_L g2139 ( 
.A(n_1741),
.Y(n_2139)
);

AND2x4_ASAP7_75t_L g2140 ( 
.A(n_1865),
.B(n_1401),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_1913),
.Y(n_2141)
);

INVx3_ASAP7_75t_L g2142 ( 
.A(n_1741),
.Y(n_2142)
);

NAND2xp5_ASAP7_75t_L g2143 ( 
.A(n_1763),
.B(n_1356),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_1932),
.Y(n_2144)
);

BUFx6f_ASAP7_75t_L g2145 ( 
.A(n_1741),
.Y(n_2145)
);

NAND2xp5_ASAP7_75t_L g2146 ( 
.A(n_1778),
.B(n_1357),
.Y(n_2146)
);

INVx3_ASAP7_75t_L g2147 ( 
.A(n_1748),
.Y(n_2147)
);

INVx2_ASAP7_75t_L g2148 ( 
.A(n_1772),
.Y(n_2148)
);

INVx6_ASAP7_75t_L g2149 ( 
.A(n_1845),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_1940),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_1706),
.Y(n_2151)
);

INVx2_ASAP7_75t_L g2152 ( 
.A(n_1776),
.Y(n_2152)
);

BUFx6f_ASAP7_75t_L g2153 ( 
.A(n_1748),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_2013),
.Y(n_2154)
);

INVx2_ASAP7_75t_L g2155 ( 
.A(n_1782),
.Y(n_2155)
);

INVx6_ASAP7_75t_L g2156 ( 
.A(n_1845),
.Y(n_2156)
);

INVx2_ASAP7_75t_SL g2157 ( 
.A(n_1879),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_2013),
.Y(n_2158)
);

NAND2xp33_ASAP7_75t_L g2159 ( 
.A(n_1981),
.B(n_1542),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_2013),
.Y(n_2160)
);

INVx2_ASAP7_75t_L g2161 ( 
.A(n_1793),
.Y(n_2161)
);

AND2x2_ASAP7_75t_L g2162 ( 
.A(n_1989),
.B(n_1283),
.Y(n_2162)
);

NAND2xp5_ASAP7_75t_L g2163 ( 
.A(n_1778),
.B(n_1359),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_2018),
.Y(n_2164)
);

OA21x2_ASAP7_75t_L g2165 ( 
.A1(n_1918),
.A2(n_1363),
.B(n_1361),
.Y(n_2165)
);

INVx2_ASAP7_75t_L g2166 ( 
.A(n_1801),
.Y(n_2166)
);

CKINVDCx5p33_ASAP7_75t_R g2167 ( 
.A(n_1736),
.Y(n_2167)
);

NAND2xp33_ASAP7_75t_L g2168 ( 
.A(n_1981),
.B(n_1546),
.Y(n_2168)
);

BUFx6f_ASAP7_75t_L g2169 ( 
.A(n_1748),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_2018),
.Y(n_2170)
);

AND2x4_ASAP7_75t_L g2171 ( 
.A(n_1935),
.B(n_1825),
.Y(n_2171)
);

BUFx6f_ASAP7_75t_L g2172 ( 
.A(n_1760),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_2018),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_2021),
.Y(n_2174)
);

AND2x2_ASAP7_75t_L g2175 ( 
.A(n_1708),
.B(n_1283),
.Y(n_2175)
);

AND2x4_ASAP7_75t_L g2176 ( 
.A(n_1858),
.B(n_1402),
.Y(n_2176)
);

INVx2_ASAP7_75t_L g2177 ( 
.A(n_1805),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_2021),
.Y(n_2178)
);

BUFx6f_ASAP7_75t_L g2179 ( 
.A(n_1760),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_2021),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_2024),
.Y(n_2181)
);

AND3x2_ASAP7_75t_L g2182 ( 
.A(n_1757),
.B(n_1068),
.C(n_1063),
.Y(n_2182)
);

BUFx3_ASAP7_75t_L g2183 ( 
.A(n_1710),
.Y(n_2183)
);

INVx2_ASAP7_75t_L g2184 ( 
.A(n_1814),
.Y(n_2184)
);

NAND2xp5_ASAP7_75t_L g2185 ( 
.A(n_1714),
.B(n_1364),
.Y(n_2185)
);

INVx3_ASAP7_75t_L g2186 ( 
.A(n_1760),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_2024),
.Y(n_2187)
);

INVx2_ASAP7_75t_L g2188 ( 
.A(n_1816),
.Y(n_2188)
);

NOR2xp33_ASAP7_75t_L g2189 ( 
.A(n_1877),
.B(n_1573),
.Y(n_2189)
);

BUFx6f_ASAP7_75t_L g2190 ( 
.A(n_1761),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_2024),
.Y(n_2191)
);

INVxp67_ASAP7_75t_L g2192 ( 
.A(n_1809),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_2025),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_2025),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_2025),
.Y(n_2195)
);

BUFx6f_ASAP7_75t_L g2196 ( 
.A(n_1761),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_2028),
.Y(n_2197)
);

NAND2xp33_ASAP7_75t_SL g2198 ( 
.A(n_1722),
.B(n_1302),
.Y(n_2198)
);

INVx3_ASAP7_75t_L g2199 ( 
.A(n_1761),
.Y(n_2199)
);

CKINVDCx16_ASAP7_75t_R g2200 ( 
.A(n_1972),
.Y(n_2200)
);

NAND2xp5_ASAP7_75t_L g2201 ( 
.A(n_1714),
.B(n_1365),
.Y(n_2201)
);

INVx2_ASAP7_75t_L g2202 ( 
.A(n_1831),
.Y(n_2202)
);

AND2x2_ASAP7_75t_L g2203 ( 
.A(n_1903),
.B(n_1302),
.Y(n_2203)
);

INVx2_ASAP7_75t_L g2204 ( 
.A(n_1846),
.Y(n_2204)
);

AND2x4_ASAP7_75t_L g2205 ( 
.A(n_1858),
.B(n_1405),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_2028),
.Y(n_2206)
);

INVx2_ASAP7_75t_L g2207 ( 
.A(n_1853),
.Y(n_2207)
);

AND2x4_ASAP7_75t_L g2208 ( 
.A(n_1764),
.B(n_1406),
.Y(n_2208)
);

NAND2xp5_ASAP7_75t_L g2209 ( 
.A(n_1717),
.B(n_1366),
.Y(n_2209)
);

INVx2_ASAP7_75t_SL g2210 ( 
.A(n_1879),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_2028),
.Y(n_2211)
);

HB1xp67_ASAP7_75t_L g2212 ( 
.A(n_1773),
.Y(n_2212)
);

INVx2_ASAP7_75t_L g2213 ( 
.A(n_1869),
.Y(n_2213)
);

INVxp67_ASAP7_75t_L g2214 ( 
.A(n_1809),
.Y(n_2214)
);

NOR2xp67_ASAP7_75t_L g2215 ( 
.A(n_2012),
.B(n_1692),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_2046),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_2046),
.Y(n_2217)
);

INVx2_ASAP7_75t_L g2218 ( 
.A(n_1921),
.Y(n_2218)
);

NAND2xp5_ASAP7_75t_SL g2219 ( 
.A(n_2012),
.B(n_1546),
.Y(n_2219)
);

HB1xp67_ASAP7_75t_L g2220 ( 
.A(n_1773),
.Y(n_2220)
);

INVx2_ASAP7_75t_L g2221 ( 
.A(n_1921),
.Y(n_2221)
);

INVx2_ASAP7_75t_L g2222 ( 
.A(n_1921),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_2046),
.Y(n_2223)
);

INVx2_ASAP7_75t_L g2224 ( 
.A(n_1921),
.Y(n_2224)
);

NAND2xp5_ASAP7_75t_L g2225 ( 
.A(n_1717),
.B(n_1368),
.Y(n_2225)
);

INVxp33_ASAP7_75t_SL g2226 ( 
.A(n_1794),
.Y(n_2226)
);

INVx2_ASAP7_75t_L g2227 ( 
.A(n_1929),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_2048),
.Y(n_2228)
);

AND2x2_ASAP7_75t_L g2229 ( 
.A(n_1903),
.B(n_1326),
.Y(n_2229)
);

NAND2xp5_ASAP7_75t_SL g2230 ( 
.A(n_2012),
.B(n_1572),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_2048),
.Y(n_2231)
);

AND3x2_ASAP7_75t_L g2232 ( 
.A(n_1930),
.B(n_1069),
.C(n_1068),
.Y(n_2232)
);

AND2x4_ASAP7_75t_L g2233 ( 
.A(n_1804),
.B(n_1408),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_2048),
.Y(n_2234)
);

AND2x4_ASAP7_75t_L g2235 ( 
.A(n_1804),
.B(n_1409),
.Y(n_2235)
);

INVx2_ASAP7_75t_L g2236 ( 
.A(n_1929),
.Y(n_2236)
);

INVx2_ASAP7_75t_L g2237 ( 
.A(n_1929),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_2050),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_2050),
.Y(n_2239)
);

INVx2_ASAP7_75t_L g2240 ( 
.A(n_1929),
.Y(n_2240)
);

HB1xp67_ASAP7_75t_L g2241 ( 
.A(n_1823),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_2050),
.Y(n_2242)
);

NAND2xp5_ASAP7_75t_L g2243 ( 
.A(n_1777),
.B(n_1371),
.Y(n_2243)
);

OA21x2_ASAP7_75t_L g2244 ( 
.A1(n_1918),
.A2(n_1944),
.B(n_1894),
.Y(n_2244)
);

NAND2xp5_ASAP7_75t_L g2245 ( 
.A(n_1777),
.B(n_1713),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_2054),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_2054),
.Y(n_2247)
);

NAND2xp5_ASAP7_75t_L g2248 ( 
.A(n_1713),
.B(n_1372),
.Y(n_2248)
);

AOI22xp5_ASAP7_75t_L g2249 ( 
.A1(n_1842),
.A2(n_1677),
.B1(n_1653),
.B2(n_1572),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_2054),
.Y(n_2250)
);

NOR2xp33_ASAP7_75t_L g2251 ( 
.A(n_1900),
.B(n_1653),
.Y(n_2251)
);

AND2x4_ASAP7_75t_L g2252 ( 
.A(n_1823),
.B(n_1412),
.Y(n_2252)
);

INVx2_ASAP7_75t_L g2253 ( 
.A(n_1899),
.Y(n_2253)
);

BUFx6f_ASAP7_75t_L g2254 ( 
.A(n_1766),
.Y(n_2254)
);

INVx2_ASAP7_75t_L g2255 ( 
.A(n_1899),
.Y(n_2255)
);

HB1xp67_ASAP7_75t_L g2256 ( 
.A(n_1859),
.Y(n_2256)
);

INVx2_ASAP7_75t_L g2257 ( 
.A(n_1899),
.Y(n_2257)
);

AND2x2_ASAP7_75t_L g2258 ( 
.A(n_1856),
.B(n_1326),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_2055),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_2055),
.Y(n_2260)
);

INVx3_ASAP7_75t_L g2261 ( 
.A(n_1766),
.Y(n_2261)
);

INVx3_ASAP7_75t_L g2262 ( 
.A(n_1766),
.Y(n_2262)
);

INVx2_ASAP7_75t_L g2263 ( 
.A(n_1908),
.Y(n_2263)
);

HB1xp67_ASAP7_75t_L g2264 ( 
.A(n_1859),
.Y(n_2264)
);

INVx2_ASAP7_75t_L g2265 ( 
.A(n_1908),
.Y(n_2265)
);

INVxp67_ASAP7_75t_L g2266 ( 
.A(n_1832),
.Y(n_2266)
);

BUFx6f_ASAP7_75t_L g2267 ( 
.A(n_1768),
.Y(n_2267)
);

NAND2xp5_ASAP7_75t_L g2268 ( 
.A(n_1737),
.B(n_1596),
.Y(n_2268)
);

CKINVDCx20_ASAP7_75t_R g2269 ( 
.A(n_1758),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_2055),
.Y(n_2270)
);

BUFx6f_ASAP7_75t_L g2271 ( 
.A(n_1768),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_2062),
.Y(n_2272)
);

INVx3_ASAP7_75t_L g2273 ( 
.A(n_1768),
.Y(n_2273)
);

INVx1_ASAP7_75t_SL g2274 ( 
.A(n_1758),
.Y(n_2274)
);

INVx1_ASAP7_75t_L g2275 ( 
.A(n_2062),
.Y(n_2275)
);

BUFx6f_ASAP7_75t_L g2276 ( 
.A(n_1779),
.Y(n_2276)
);

INVxp67_ASAP7_75t_L g2277 ( 
.A(n_1832),
.Y(n_2277)
);

INVx2_ASAP7_75t_L g2278 ( 
.A(n_1908),
.Y(n_2278)
);

NOR2xp33_ASAP7_75t_L g2279 ( 
.A(n_1900),
.B(n_1677),
.Y(n_2279)
);

BUFx8_ASAP7_75t_L g2280 ( 
.A(n_1807),
.Y(n_2280)
);

NAND2xp5_ASAP7_75t_L g2281 ( 
.A(n_1737),
.B(n_1596),
.Y(n_2281)
);

XNOR2x1_ASAP7_75t_L g2282 ( 
.A(n_1798),
.B(n_1407),
.Y(n_2282)
);

HB1xp67_ASAP7_75t_L g2283 ( 
.A(n_1875),
.Y(n_2283)
);

INVx2_ASAP7_75t_L g2284 ( 
.A(n_1937),
.Y(n_2284)
);

BUFx6f_ASAP7_75t_L g2285 ( 
.A(n_1779),
.Y(n_2285)
);

BUFx2_ASAP7_75t_L g2286 ( 
.A(n_1726),
.Y(n_2286)
);

INVxp67_ASAP7_75t_L g2287 ( 
.A(n_1783),
.Y(n_2287)
);

NAND2x1_ASAP7_75t_L g2288 ( 
.A(n_1788),
.B(n_1220),
.Y(n_2288)
);

NAND2xp33_ASAP7_75t_L g2289 ( 
.A(n_1981),
.B(n_1999),
.Y(n_2289)
);

INVx3_ASAP7_75t_L g2290 ( 
.A(n_1779),
.Y(n_2290)
);

NAND2xp5_ASAP7_75t_L g2291 ( 
.A(n_1704),
.B(n_1718),
.Y(n_2291)
);

NAND2xp5_ASAP7_75t_L g2292 ( 
.A(n_1704),
.B(n_1619),
.Y(n_2292)
);

AND2x6_ASAP7_75t_L g2293 ( 
.A(n_1880),
.B(n_1120),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_L g2294 ( 
.A(n_1718),
.B(n_1619),
.Y(n_2294)
);

AND2x2_ASAP7_75t_L g2295 ( 
.A(n_1888),
.B(n_1626),
.Y(n_2295)
);

INVx1_ASAP7_75t_L g2296 ( 
.A(n_2062),
.Y(n_2296)
);

INVx2_ASAP7_75t_L g2297 ( 
.A(n_1937),
.Y(n_2297)
);

OA21x2_ASAP7_75t_L g2298 ( 
.A1(n_1894),
.A2(n_1688),
.B(n_1687),
.Y(n_2298)
);

NOR2xp33_ASAP7_75t_SL g2299 ( 
.A(n_1866),
.B(n_1607),
.Y(n_2299)
);

BUFx6f_ASAP7_75t_L g2300 ( 
.A(n_1780),
.Y(n_2300)
);

HB1xp67_ASAP7_75t_L g2301 ( 
.A(n_1875),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_2062),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_2010),
.Y(n_2303)
);

NAND2xp5_ASAP7_75t_L g2304 ( 
.A(n_1786),
.B(n_1626),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_2010),
.Y(n_2305)
);

INVx2_ASAP7_75t_L g2306 ( 
.A(n_1937),
.Y(n_2306)
);

HB1xp67_ASAP7_75t_L g2307 ( 
.A(n_1897),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_2043),
.Y(n_2308)
);

NAND2xp5_ASAP7_75t_L g2309 ( 
.A(n_1786),
.B(n_1628),
.Y(n_2309)
);

BUFx3_ASAP7_75t_L g2310 ( 
.A(n_1710),
.Y(n_2310)
);

AND2x2_ASAP7_75t_L g2311 ( 
.A(n_1898),
.B(n_1628),
.Y(n_2311)
);

INVx3_ASAP7_75t_L g2312 ( 
.A(n_1780),
.Y(n_2312)
);

AND2x4_ASAP7_75t_L g2313 ( 
.A(n_1897),
.B(n_1513),
.Y(n_2313)
);

NAND2x1p5_ASAP7_75t_L g2314 ( 
.A(n_2022),
.B(n_1423),
.Y(n_2314)
);

INVx2_ASAP7_75t_L g2315 ( 
.A(n_1951),
.Y(n_2315)
);

AND2x4_ASAP7_75t_L g2316 ( 
.A(n_1902),
.B(n_1517),
.Y(n_2316)
);

INVx2_ASAP7_75t_L g2317 ( 
.A(n_1951),
.Y(n_2317)
);

BUFx6f_ASAP7_75t_L g2318 ( 
.A(n_1780),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_2043),
.Y(n_2319)
);

INVxp67_ASAP7_75t_L g2320 ( 
.A(n_1783),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_1723),
.Y(n_2321)
);

INVxp33_ASAP7_75t_L g2322 ( 
.A(n_1784),
.Y(n_2322)
);

NAND2xp5_ASAP7_75t_L g2323 ( 
.A(n_1830),
.B(n_1630),
.Y(n_2323)
);

NAND2xp5_ASAP7_75t_SL g2324 ( 
.A(n_1830),
.B(n_1630),
.Y(n_2324)
);

AND2x4_ASAP7_75t_L g2325 ( 
.A(n_1902),
.B(n_1519),
.Y(n_2325)
);

OAI22xp33_ASAP7_75t_L g2326 ( 
.A1(n_1702),
.A2(n_1696),
.B1(n_1678),
.B2(n_1341),
.Y(n_2326)
);

OAI22xp5_ASAP7_75t_L g2327 ( 
.A1(n_1879),
.A2(n_1516),
.B1(n_1551),
.B2(n_1659),
.Y(n_2327)
);

INVx2_ASAP7_75t_L g2328 ( 
.A(n_1951),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_1728),
.Y(n_2329)
);

INVx1_ASAP7_75t_L g2330 ( 
.A(n_1744),
.Y(n_2330)
);

AND2x2_ASAP7_75t_L g2331 ( 
.A(n_1751),
.B(n_1659),
.Y(n_2331)
);

INVx2_ASAP7_75t_L g2332 ( 
.A(n_1952),
.Y(n_2332)
);

BUFx6f_ASAP7_75t_L g2333 ( 
.A(n_1787),
.Y(n_2333)
);

AND3x2_ASAP7_75t_L g2334 ( 
.A(n_1972),
.B(n_1072),
.C(n_1069),
.Y(n_2334)
);

INVx6_ASAP7_75t_L g2335 ( 
.A(n_2022),
.Y(n_2335)
);

BUFx3_ASAP7_75t_L g2336 ( 
.A(n_1906),
.Y(n_2336)
);

AND2x2_ASAP7_75t_L g2337 ( 
.A(n_1911),
.B(n_1665),
.Y(n_2337)
);

INVx1_ASAP7_75t_L g2338 ( 
.A(n_1770),
.Y(n_2338)
);

INVx2_ASAP7_75t_L g2339 ( 
.A(n_1952),
.Y(n_2339)
);

OA21x2_ASAP7_75t_L g2340 ( 
.A1(n_1944),
.A2(n_1684),
.B(n_1681),
.Y(n_2340)
);

NAND2xp5_ASAP7_75t_SL g2341 ( 
.A(n_1910),
.B(n_1665),
.Y(n_2341)
);

INVx2_ASAP7_75t_L g2342 ( 
.A(n_1952),
.Y(n_2342)
);

INVxp67_ASAP7_75t_L g2343 ( 
.A(n_1784),
.Y(n_2343)
);

OAI21x1_ASAP7_75t_L g2344 ( 
.A1(n_1947),
.A2(n_1690),
.B(n_1685),
.Y(n_2344)
);

INVx1_ASAP7_75t_L g2345 ( 
.A(n_1785),
.Y(n_2345)
);

AND2x2_ASAP7_75t_L g2346 ( 
.A(n_1955),
.B(n_1666),
.Y(n_2346)
);

INVx1_ASAP7_75t_L g2347 ( 
.A(n_1828),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_1860),
.Y(n_2348)
);

NAND2xp5_ASAP7_75t_L g2349 ( 
.A(n_1910),
.B(n_1666),
.Y(n_2349)
);

NOR2xp33_ASAP7_75t_L g2350 ( 
.A(n_1789),
.B(n_1692),
.Y(n_2350)
);

INVx2_ASAP7_75t_L g2351 ( 
.A(n_1954),
.Y(n_2351)
);

INVx2_ASAP7_75t_L g2352 ( 
.A(n_1954),
.Y(n_2352)
);

INVx2_ASAP7_75t_L g2353 ( 
.A(n_1954),
.Y(n_2353)
);

INVx2_ASAP7_75t_L g2354 ( 
.A(n_1957),
.Y(n_2354)
);

AND2x6_ASAP7_75t_L g2355 ( 
.A(n_1956),
.B(n_1120),
.Y(n_2355)
);

BUFx6f_ASAP7_75t_L g2356 ( 
.A(n_1787),
.Y(n_2356)
);

NAND2xp5_ASAP7_75t_L g2357 ( 
.A(n_1925),
.B(n_1521),
.Y(n_2357)
);

NAND2xp5_ASAP7_75t_L g2358 ( 
.A(n_1925),
.B(n_1522),
.Y(n_2358)
);

HB1xp67_ASAP7_75t_L g2359 ( 
.A(n_1906),
.Y(n_2359)
);

NAND2xp5_ASAP7_75t_L g2360 ( 
.A(n_1789),
.B(n_1524),
.Y(n_2360)
);

INVx2_ASAP7_75t_L g2361 ( 
.A(n_1957),
.Y(n_2361)
);

AND2x4_ASAP7_75t_L g2362 ( 
.A(n_1922),
.B(n_1526),
.Y(n_2362)
);

NOR2x1_ASAP7_75t_L g2363 ( 
.A(n_1719),
.B(n_1529),
.Y(n_2363)
);

NAND2xp33_ASAP7_75t_L g2364 ( 
.A(n_1981),
.B(n_1143),
.Y(n_2364)
);

INVx1_ASAP7_75t_L g2365 ( 
.A(n_1870),
.Y(n_2365)
);

INVx1_ASAP7_75t_SL g2366 ( 
.A(n_1767),
.Y(n_2366)
);

INVx2_ASAP7_75t_L g2367 ( 
.A(n_1957),
.Y(n_2367)
);

INVx1_ASAP7_75t_L g2368 ( 
.A(n_1884),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_1891),
.Y(n_2369)
);

INVx3_ASAP7_75t_L g2370 ( 
.A(n_1787),
.Y(n_2370)
);

INVx2_ASAP7_75t_L g2371 ( 
.A(n_1959),
.Y(n_2371)
);

NAND2xp5_ASAP7_75t_SL g2372 ( 
.A(n_1947),
.B(n_1143),
.Y(n_2372)
);

BUFx6f_ASAP7_75t_L g2373 ( 
.A(n_1791),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_2009),
.Y(n_2374)
);

NAND2xp5_ASAP7_75t_L g2375 ( 
.A(n_1796),
.B(n_1531),
.Y(n_2375)
);

AND2x2_ASAP7_75t_L g2376 ( 
.A(n_1966),
.B(n_1329),
.Y(n_2376)
);

INVx2_ASAP7_75t_L g2377 ( 
.A(n_1959),
.Y(n_2377)
);

HB1xp67_ASAP7_75t_L g2378 ( 
.A(n_1922),
.Y(n_2378)
);

INVx4_ASAP7_75t_L g2379 ( 
.A(n_2022),
.Y(n_2379)
);

NAND2xp5_ASAP7_75t_SL g2380 ( 
.A(n_2039),
.B(n_1186),
.Y(n_2380)
);

INVx1_ASAP7_75t_L g2381 ( 
.A(n_2037),
.Y(n_2381)
);

INVx1_ASAP7_75t_L g2382 ( 
.A(n_2038),
.Y(n_2382)
);

NAND2xp33_ASAP7_75t_L g2383 ( 
.A(n_1999),
.B(n_1186),
.Y(n_2383)
);

NAND2xp33_ASAP7_75t_SL g2384 ( 
.A(n_2057),
.B(n_1507),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_2049),
.Y(n_2385)
);

AND2x2_ASAP7_75t_L g2386 ( 
.A(n_1806),
.B(n_1329),
.Y(n_2386)
);

INVx2_ASAP7_75t_L g2387 ( 
.A(n_1959),
.Y(n_2387)
);

AND2x2_ASAP7_75t_L g2388 ( 
.A(n_1771),
.B(n_1341),
.Y(n_2388)
);

INVx3_ASAP7_75t_L g2389 ( 
.A(n_1791),
.Y(n_2389)
);

INVx1_ASAP7_75t_L g2390 ( 
.A(n_2061),
.Y(n_2390)
);

INVx2_ASAP7_75t_L g2391 ( 
.A(n_1960),
.Y(n_2391)
);

INVx1_ASAP7_75t_L g2392 ( 
.A(n_2059),
.Y(n_2392)
);

NAND2xp5_ASAP7_75t_SL g2393 ( 
.A(n_1725),
.B(n_1198),
.Y(n_2393)
);

INVx3_ASAP7_75t_L g2394 ( 
.A(n_1791),
.Y(n_2394)
);

NAND2xp5_ASAP7_75t_L g2395 ( 
.A(n_1796),
.B(n_1534),
.Y(n_2395)
);

INVx1_ASAP7_75t_L g2396 ( 
.A(n_1874),
.Y(n_2396)
);

INVx1_ASAP7_75t_L g2397 ( 
.A(n_1874),
.Y(n_2397)
);

NOR2xp33_ASAP7_75t_L g2398 ( 
.A(n_1797),
.B(n_1375),
.Y(n_2398)
);

INVx2_ASAP7_75t_L g2399 ( 
.A(n_1960),
.Y(n_2399)
);

INVx2_ASAP7_75t_L g2400 ( 
.A(n_1960),
.Y(n_2400)
);

NAND2x1p5_ASAP7_75t_L g2401 ( 
.A(n_2022),
.B(n_1680),
.Y(n_2401)
);

INVx4_ASAP7_75t_L g2402 ( 
.A(n_2026),
.Y(n_2402)
);

NAND2xp5_ASAP7_75t_L g2403 ( 
.A(n_1797),
.B(n_1799),
.Y(n_2403)
);

AND2x6_ASAP7_75t_L g2404 ( 
.A(n_1725),
.B(n_1198),
.Y(n_2404)
);

INVx1_ASAP7_75t_L g2405 ( 
.A(n_1874),
.Y(n_2405)
);

NAND2xp5_ASAP7_75t_L g2406 ( 
.A(n_1799),
.B(n_1536),
.Y(n_2406)
);

AND2x2_ASAP7_75t_L g2407 ( 
.A(n_1771),
.B(n_1375),
.Y(n_2407)
);

INVx2_ASAP7_75t_L g2408 ( 
.A(n_1961),
.Y(n_2408)
);

NAND2xp5_ASAP7_75t_L g2409 ( 
.A(n_1822),
.B(n_1539),
.Y(n_2409)
);

BUFx6f_ASAP7_75t_L g2410 ( 
.A(n_1812),
.Y(n_2410)
);

AND2x2_ASAP7_75t_L g2411 ( 
.A(n_1762),
.B(n_1395),
.Y(n_2411)
);

AND2x4_ASAP7_75t_L g2412 ( 
.A(n_1949),
.B(n_1541),
.Y(n_2412)
);

INVx2_ASAP7_75t_L g2413 ( 
.A(n_1961),
.Y(n_2413)
);

NAND2xp5_ASAP7_75t_L g2414 ( 
.A(n_1822),
.B(n_1544),
.Y(n_2414)
);

INVx2_ASAP7_75t_L g2415 ( 
.A(n_1961),
.Y(n_2415)
);

INVx3_ASAP7_75t_L g2416 ( 
.A(n_1812),
.Y(n_2416)
);

INVx3_ASAP7_75t_L g2417 ( 
.A(n_1812),
.Y(n_2417)
);

BUFx8_ASAP7_75t_L g2418 ( 
.A(n_1824),
.Y(n_2418)
);

NAND2xp5_ASAP7_75t_L g2419 ( 
.A(n_1837),
.B(n_1550),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_1878),
.Y(n_2420)
);

INVx1_ASAP7_75t_L g2421 ( 
.A(n_1878),
.Y(n_2421)
);

CKINVDCx5p33_ASAP7_75t_R g2422 ( 
.A(n_1767),
.Y(n_2422)
);

INVx2_ASAP7_75t_L g2423 ( 
.A(n_1983),
.Y(n_2423)
);

NAND2xp5_ASAP7_75t_SL g2424 ( 
.A(n_1727),
.B(n_1225),
.Y(n_2424)
);

BUFx8_ASAP7_75t_L g2425 ( 
.A(n_1838),
.Y(n_2425)
);

INVx1_ASAP7_75t_L g2426 ( 
.A(n_1878),
.Y(n_2426)
);

INVx1_ASAP7_75t_L g2427 ( 
.A(n_1885),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_1885),
.Y(n_2428)
);

OR2x6_ASAP7_75t_L g2429 ( 
.A(n_1792),
.B(n_1504),
.Y(n_2429)
);

INVx2_ASAP7_75t_L g2430 ( 
.A(n_1983),
.Y(n_2430)
);

NAND2xp5_ASAP7_75t_L g2431 ( 
.A(n_1837),
.B(n_1553),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_1885),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_1890),
.Y(n_2433)
);

INVx1_ASAP7_75t_L g2434 ( 
.A(n_1890),
.Y(n_2434)
);

BUFx6f_ASAP7_75t_L g2435 ( 
.A(n_1817),
.Y(n_2435)
);

BUFx3_ASAP7_75t_L g2436 ( 
.A(n_1949),
.Y(n_2436)
);

BUFx6f_ASAP7_75t_L g2437 ( 
.A(n_1817),
.Y(n_2437)
);

NOR2x1_ASAP7_75t_L g2438 ( 
.A(n_1719),
.B(n_1554),
.Y(n_2438)
);

HB1xp67_ASAP7_75t_L g2439 ( 
.A(n_1976),
.Y(n_2439)
);

AND2x4_ASAP7_75t_L g2440 ( 
.A(n_1976),
.B(n_1555),
.Y(n_2440)
);

NAND2xp5_ASAP7_75t_L g2441 ( 
.A(n_1841),
.B(n_1556),
.Y(n_2441)
);

INVx3_ASAP7_75t_L g2442 ( 
.A(n_1817),
.Y(n_2442)
);

INVx1_ASAP7_75t_L g2443 ( 
.A(n_1890),
.Y(n_2443)
);

BUFx6f_ASAP7_75t_L g2444 ( 
.A(n_1818),
.Y(n_2444)
);

INVx1_ASAP7_75t_L g2445 ( 
.A(n_1892),
.Y(n_2445)
);

BUFx8_ASAP7_75t_L g2446 ( 
.A(n_1754),
.Y(n_2446)
);

INVx1_ASAP7_75t_L g2447 ( 
.A(n_1983),
.Y(n_2447)
);

AND2x2_ASAP7_75t_L g2448 ( 
.A(n_1762),
.B(n_1395),
.Y(n_2448)
);

INVx1_ASAP7_75t_L g2449 ( 
.A(n_1987),
.Y(n_2449)
);

INVx1_ASAP7_75t_L g2450 ( 
.A(n_1987),
.Y(n_2450)
);

INVx1_ASAP7_75t_L g2451 ( 
.A(n_1987),
.Y(n_2451)
);

AND2x2_ASAP7_75t_L g2452 ( 
.A(n_1842),
.B(n_1403),
.Y(n_2452)
);

INVx2_ASAP7_75t_L g2453 ( 
.A(n_1820),
.Y(n_2453)
);

INVx2_ASAP7_75t_L g2454 ( 
.A(n_1820),
.Y(n_2454)
);

INVx4_ASAP7_75t_L g2455 ( 
.A(n_2026),
.Y(n_2455)
);

INVx1_ASAP7_75t_L g2456 ( 
.A(n_1775),
.Y(n_2456)
);

AND2x2_ASAP7_75t_L g2457 ( 
.A(n_1752),
.B(n_1403),
.Y(n_2457)
);

BUFx6f_ASAP7_75t_L g2458 ( 
.A(n_1818),
.Y(n_2458)
);

AND2x2_ASAP7_75t_L g2459 ( 
.A(n_1769),
.B(n_1404),
.Y(n_2459)
);

BUFx6f_ASAP7_75t_L g2460 ( 
.A(n_1818),
.Y(n_2460)
);

INVx1_ASAP7_75t_L g2461 ( 
.A(n_1775),
.Y(n_2461)
);

BUFx6f_ASAP7_75t_L g2462 ( 
.A(n_1810),
.Y(n_2462)
);

BUFx8_ASAP7_75t_L g2463 ( 
.A(n_1707),
.Y(n_2463)
);

INVx2_ASAP7_75t_L g2464 ( 
.A(n_1820),
.Y(n_2464)
);

INVx3_ASAP7_75t_L g2465 ( 
.A(n_1810),
.Y(n_2465)
);

OA21x2_ASAP7_75t_L g2466 ( 
.A1(n_1841),
.A2(n_1849),
.B(n_1958),
.Y(n_2466)
);

INVx3_ASAP7_75t_L g2467 ( 
.A(n_1810),
.Y(n_2467)
);

BUFx6f_ASAP7_75t_L g2468 ( 
.A(n_1810),
.Y(n_2468)
);

BUFx2_ASAP7_75t_L g2469 ( 
.A(n_1732),
.Y(n_2469)
);

INVx3_ASAP7_75t_L g2470 ( 
.A(n_1813),
.Y(n_2470)
);

INVx1_ASAP7_75t_L g2471 ( 
.A(n_1802),
.Y(n_2471)
);

INVxp67_ASAP7_75t_L g2472 ( 
.A(n_1803),
.Y(n_2472)
);

BUFx12f_ASAP7_75t_L g2473 ( 
.A(n_1941),
.Y(n_2473)
);

CKINVDCx20_ASAP7_75t_R g2474 ( 
.A(n_1781),
.Y(n_2474)
);

AND2x2_ASAP7_75t_L g2475 ( 
.A(n_1790),
.B(n_1833),
.Y(n_2475)
);

INVx1_ASAP7_75t_L g2476 ( 
.A(n_1802),
.Y(n_2476)
);

AND2x2_ASAP7_75t_L g2477 ( 
.A(n_1833),
.B(n_1404),
.Y(n_2477)
);

INVx3_ASAP7_75t_L g2478 ( 
.A(n_1813),
.Y(n_2478)
);

AND2x2_ASAP7_75t_L g2479 ( 
.A(n_1803),
.B(n_1411),
.Y(n_2479)
);

HB1xp67_ASAP7_75t_L g2480 ( 
.A(n_1997),
.Y(n_2480)
);

INVx1_ASAP7_75t_L g2481 ( 
.A(n_1826),
.Y(n_2481)
);

INVx2_ASAP7_75t_L g2482 ( 
.A(n_2065),
.Y(n_2482)
);

NOR2x1p5_ASAP7_75t_L g2483 ( 
.A(n_2473),
.B(n_1759),
.Y(n_2483)
);

INVx4_ASAP7_75t_L g2484 ( 
.A(n_2095),
.Y(n_2484)
);

BUFx6f_ASAP7_75t_L g2485 ( 
.A(n_2336),
.Y(n_2485)
);

AOI22xp5_ASAP7_75t_L g2486 ( 
.A1(n_2384),
.A2(n_1843),
.B1(n_1973),
.B2(n_1965),
.Y(n_2486)
);

INVx2_ASAP7_75t_SL g2487 ( 
.A(n_2376),
.Y(n_2487)
);

INVx2_ASAP7_75t_L g2488 ( 
.A(n_2065),
.Y(n_2488)
);

NAND2xp5_ASAP7_75t_SL g2489 ( 
.A(n_2291),
.B(n_1866),
.Y(n_2489)
);

INVx2_ASAP7_75t_L g2490 ( 
.A(n_2068),
.Y(n_2490)
);

INVx2_ASAP7_75t_L g2491 ( 
.A(n_2068),
.Y(n_2491)
);

INVx1_ASAP7_75t_L g2492 ( 
.A(n_2212),
.Y(n_2492)
);

INVx2_ASAP7_75t_L g2493 ( 
.A(n_2092),
.Y(n_2493)
);

INVx2_ASAP7_75t_L g2494 ( 
.A(n_2092),
.Y(n_2494)
);

NAND2xp5_ASAP7_75t_SL g2495 ( 
.A(n_2403),
.B(n_2002),
.Y(n_2495)
);

INVx3_ASAP7_75t_L g2496 ( 
.A(n_2218),
.Y(n_2496)
);

CKINVDCx5p33_ASAP7_75t_R g2497 ( 
.A(n_2167),
.Y(n_2497)
);

CKINVDCx5p33_ASAP7_75t_R g2498 ( 
.A(n_2167),
.Y(n_2498)
);

INVx8_ASAP7_75t_L g2499 ( 
.A(n_2293),
.Y(n_2499)
);

INVxp33_ASAP7_75t_L g2500 ( 
.A(n_2388),
.Y(n_2500)
);

NAND2xp5_ASAP7_75t_SL g2501 ( 
.A(n_2292),
.B(n_2002),
.Y(n_2501)
);

NOR2xp33_ASAP7_75t_L g2502 ( 
.A(n_2322),
.B(n_1735),
.Y(n_2502)
);

INVx2_ASAP7_75t_L g2503 ( 
.A(n_2093),
.Y(n_2503)
);

INVx2_ASAP7_75t_L g2504 ( 
.A(n_2093),
.Y(n_2504)
);

INVx1_ASAP7_75t_L g2505 ( 
.A(n_2212),
.Y(n_2505)
);

INVx1_ASAP7_75t_L g2506 ( 
.A(n_2220),
.Y(n_2506)
);

INVx2_ASAP7_75t_L g2507 ( 
.A(n_2098),
.Y(n_2507)
);

NOR2xp33_ASAP7_75t_L g2508 ( 
.A(n_2322),
.B(n_2192),
.Y(n_2508)
);

INVx2_ASAP7_75t_L g2509 ( 
.A(n_2098),
.Y(n_2509)
);

NOR2xp33_ASAP7_75t_L g2510 ( 
.A(n_2192),
.B(n_1829),
.Y(n_2510)
);

INVx2_ASAP7_75t_L g2511 ( 
.A(n_2112),
.Y(n_2511)
);

INVxp33_ASAP7_75t_SL g2512 ( 
.A(n_2299),
.Y(n_2512)
);

INVx3_ASAP7_75t_L g2513 ( 
.A(n_2218),
.Y(n_2513)
);

AO21x2_ASAP7_75t_L g2514 ( 
.A1(n_2372),
.A2(n_1849),
.B(n_1958),
.Y(n_2514)
);

INVx3_ASAP7_75t_L g2515 ( 
.A(n_2221),
.Y(n_2515)
);

INVx2_ASAP7_75t_L g2516 ( 
.A(n_2112),
.Y(n_2516)
);

INVx2_ASAP7_75t_L g2517 ( 
.A(n_2138),
.Y(n_2517)
);

INVx2_ASAP7_75t_SL g2518 ( 
.A(n_2171),
.Y(n_2518)
);

INVx6_ASAP7_75t_L g2519 ( 
.A(n_2103),
.Y(n_2519)
);

INVx1_ASAP7_75t_L g2520 ( 
.A(n_2220),
.Y(n_2520)
);

INVx1_ASAP7_75t_L g2521 ( 
.A(n_2241),
.Y(n_2521)
);

INVx2_ASAP7_75t_L g2522 ( 
.A(n_2138),
.Y(n_2522)
);

INVx2_ASAP7_75t_L g2523 ( 
.A(n_2148),
.Y(n_2523)
);

INVx1_ASAP7_75t_L g2524 ( 
.A(n_2241),
.Y(n_2524)
);

INVx2_ASAP7_75t_L g2525 ( 
.A(n_2148),
.Y(n_2525)
);

NAND2xp5_ASAP7_75t_SL g2526 ( 
.A(n_2294),
.B(n_2019),
.Y(n_2526)
);

INVx3_ASAP7_75t_L g2527 ( 
.A(n_2221),
.Y(n_2527)
);

AND2x6_ASAP7_75t_L g2528 ( 
.A(n_2475),
.B(n_1727),
.Y(n_2528)
);

INVx2_ASAP7_75t_L g2529 ( 
.A(n_2152),
.Y(n_2529)
);

CKINVDCx6p67_ASAP7_75t_R g2530 ( 
.A(n_2269),
.Y(n_2530)
);

NAND2xp5_ASAP7_75t_SL g2531 ( 
.A(n_2304),
.B(n_1731),
.Y(n_2531)
);

BUFx6f_ASAP7_75t_L g2532 ( 
.A(n_2336),
.Y(n_2532)
);

INVx2_ASAP7_75t_L g2533 ( 
.A(n_2152),
.Y(n_2533)
);

INVx1_ASAP7_75t_L g2534 ( 
.A(n_2256),
.Y(n_2534)
);

INVx2_ASAP7_75t_L g2535 ( 
.A(n_2155),
.Y(n_2535)
);

AND2x2_ASAP7_75t_L g2536 ( 
.A(n_2398),
.B(n_1997),
.Y(n_2536)
);

INVx1_ASAP7_75t_L g2537 ( 
.A(n_2256),
.Y(n_2537)
);

INVx1_ASAP7_75t_L g2538 ( 
.A(n_2264),
.Y(n_2538)
);

INVx1_ASAP7_75t_L g2539 ( 
.A(n_2264),
.Y(n_2539)
);

NOR2xp33_ASAP7_75t_L g2540 ( 
.A(n_2214),
.B(n_1855),
.Y(n_2540)
);

NAND2xp33_ASAP7_75t_L g2541 ( 
.A(n_2404),
.B(n_1788),
.Y(n_2541)
);

INVx2_ASAP7_75t_L g2542 ( 
.A(n_2155),
.Y(n_2542)
);

INVx1_ASAP7_75t_L g2543 ( 
.A(n_2283),
.Y(n_2543)
);

INVx1_ASAP7_75t_L g2544 ( 
.A(n_2283),
.Y(n_2544)
);

BUFx6f_ASAP7_75t_L g2545 ( 
.A(n_2436),
.Y(n_2545)
);

INVx2_ASAP7_75t_L g2546 ( 
.A(n_2161),
.Y(n_2546)
);

INVx3_ASAP7_75t_L g2547 ( 
.A(n_2222),
.Y(n_2547)
);

INVx2_ASAP7_75t_L g2548 ( 
.A(n_2161),
.Y(n_2548)
);

INVx1_ASAP7_75t_L g2549 ( 
.A(n_2301),
.Y(n_2549)
);

INVx1_ASAP7_75t_L g2550 ( 
.A(n_2301),
.Y(n_2550)
);

INVx3_ASAP7_75t_L g2551 ( 
.A(n_2222),
.Y(n_2551)
);

NAND2xp5_ASAP7_75t_SL g2552 ( 
.A(n_2309),
.B(n_1844),
.Y(n_2552)
);

INVx1_ASAP7_75t_L g2553 ( 
.A(n_2307),
.Y(n_2553)
);

INVx1_ASAP7_75t_L g2554 ( 
.A(n_2307),
.Y(n_2554)
);

INVx1_ASAP7_75t_L g2555 ( 
.A(n_2359),
.Y(n_2555)
);

NAND2xp5_ASAP7_75t_L g2556 ( 
.A(n_2398),
.B(n_1733),
.Y(n_2556)
);

NAND2xp5_ASAP7_75t_L g2557 ( 
.A(n_2350),
.B(n_1733),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_2359),
.Y(n_2558)
);

INVx2_ASAP7_75t_L g2559 ( 
.A(n_2166),
.Y(n_2559)
);

OR2x2_ASAP7_75t_L g2560 ( 
.A(n_2066),
.B(n_1452),
.Y(n_2560)
);

INVx2_ASAP7_75t_L g2561 ( 
.A(n_2166),
.Y(n_2561)
);

INVx2_ASAP7_75t_L g2562 ( 
.A(n_2177),
.Y(n_2562)
);

INVx1_ASAP7_75t_L g2563 ( 
.A(n_2378),
.Y(n_2563)
);

INVx3_ASAP7_75t_L g2564 ( 
.A(n_2224),
.Y(n_2564)
);

BUFx6f_ASAP7_75t_SL g2565 ( 
.A(n_2429),
.Y(n_2565)
);

NAND2xp5_ASAP7_75t_SL g2566 ( 
.A(n_2323),
.B(n_1862),
.Y(n_2566)
);

INVx2_ASAP7_75t_L g2567 ( 
.A(n_2177),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_2378),
.Y(n_2568)
);

INVx3_ASAP7_75t_L g2569 ( 
.A(n_2224),
.Y(n_2569)
);

INVx2_ASAP7_75t_L g2570 ( 
.A(n_2184),
.Y(n_2570)
);

INVx2_ASAP7_75t_L g2571 ( 
.A(n_2184),
.Y(n_2571)
);

NAND2xp5_ASAP7_75t_L g2572 ( 
.A(n_2350),
.B(n_1742),
.Y(n_2572)
);

NOR2xp33_ASAP7_75t_L g2573 ( 
.A(n_2214),
.B(n_1915),
.Y(n_2573)
);

NAND3xp33_ASAP7_75t_L g2574 ( 
.A(n_2132),
.B(n_1919),
.C(n_1876),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_2439),
.Y(n_2575)
);

NAND3xp33_ASAP7_75t_L g2576 ( 
.A(n_2132),
.B(n_1919),
.C(n_1876),
.Y(n_2576)
);

INVx1_ASAP7_75t_L g2577 ( 
.A(n_2439),
.Y(n_2577)
);

NOR2x1p5_ASAP7_75t_L g2578 ( 
.A(n_2473),
.B(n_1815),
.Y(n_2578)
);

INVx2_ASAP7_75t_L g2579 ( 
.A(n_2188),
.Y(n_2579)
);

INVx2_ASAP7_75t_L g2580 ( 
.A(n_2188),
.Y(n_2580)
);

INVx5_ASAP7_75t_L g2581 ( 
.A(n_2095),
.Y(n_2581)
);

INVx8_ASAP7_75t_L g2582 ( 
.A(n_2293),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_2436),
.Y(n_2583)
);

BUFx6f_ASAP7_75t_L g2584 ( 
.A(n_2064),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_2072),
.Y(n_2585)
);

NAND2xp5_ASAP7_75t_SL g2586 ( 
.A(n_2349),
.B(n_1917),
.Y(n_2586)
);

INVx2_ASAP7_75t_L g2587 ( 
.A(n_2202),
.Y(n_2587)
);

INVx3_ASAP7_75t_L g2588 ( 
.A(n_2227),
.Y(n_2588)
);

NAND2xp5_ASAP7_75t_L g2589 ( 
.A(n_2245),
.B(n_2067),
.Y(n_2589)
);

HB1xp67_ASAP7_75t_L g2590 ( 
.A(n_2071),
.Y(n_2590)
);

NAND2xp5_ASAP7_75t_SL g2591 ( 
.A(n_2357),
.B(n_1939),
.Y(n_2591)
);

INVx1_ASAP7_75t_L g2592 ( 
.A(n_2076),
.Y(n_2592)
);

INVx4_ASAP7_75t_L g2593 ( 
.A(n_2095),
.Y(n_2593)
);

AND2x2_ASAP7_75t_L g2594 ( 
.A(n_2411),
.B(n_2001),
.Y(n_2594)
);

AND2x2_ASAP7_75t_L g2595 ( 
.A(n_2448),
.B(n_2001),
.Y(n_2595)
);

NAND2xp5_ASAP7_75t_SL g2596 ( 
.A(n_2358),
.B(n_1765),
.Y(n_2596)
);

INVx2_ASAP7_75t_SL g2597 ( 
.A(n_2171),
.Y(n_2597)
);

INVx5_ASAP7_75t_L g2598 ( 
.A(n_2095),
.Y(n_2598)
);

NAND3xp33_ASAP7_75t_L g2599 ( 
.A(n_2189),
.B(n_1931),
.C(n_1927),
.Y(n_2599)
);

BUFx3_ASAP7_75t_L g2600 ( 
.A(n_2069),
.Y(n_2600)
);

NAND2xp5_ASAP7_75t_L g2601 ( 
.A(n_2077),
.B(n_1742),
.Y(n_2601)
);

BUFx10_ASAP7_75t_L g2602 ( 
.A(n_2189),
.Y(n_2602)
);

INVx1_ASAP7_75t_L g2603 ( 
.A(n_2079),
.Y(n_2603)
);

INVx2_ASAP7_75t_L g2604 ( 
.A(n_2202),
.Y(n_2604)
);

INVx2_ASAP7_75t_L g2605 ( 
.A(n_2204),
.Y(n_2605)
);

INVx3_ASAP7_75t_L g2606 ( 
.A(n_2227),
.Y(n_2606)
);

INVx3_ASAP7_75t_L g2607 ( 
.A(n_2236),
.Y(n_2607)
);

INVx1_ASAP7_75t_L g2608 ( 
.A(n_2085),
.Y(n_2608)
);

NAND2xp5_ASAP7_75t_L g2609 ( 
.A(n_2081),
.B(n_1747),
.Y(n_2609)
);

BUFx3_ASAP7_75t_L g2610 ( 
.A(n_2069),
.Y(n_2610)
);

INVx2_ASAP7_75t_SL g2611 ( 
.A(n_2074),
.Y(n_2611)
);

INVx4_ASAP7_75t_L g2612 ( 
.A(n_2462),
.Y(n_2612)
);

INVx1_ASAP7_75t_L g2613 ( 
.A(n_2089),
.Y(n_2613)
);

INVx1_ASAP7_75t_L g2614 ( 
.A(n_2091),
.Y(n_2614)
);

INVx2_ASAP7_75t_L g2615 ( 
.A(n_2204),
.Y(n_2615)
);

NAND2xp5_ASAP7_75t_L g2616 ( 
.A(n_2106),
.B(n_1747),
.Y(n_2616)
);

AND2x2_ASAP7_75t_L g2617 ( 
.A(n_2477),
.B(n_1750),
.Y(n_2617)
);

INVx1_ASAP7_75t_L g2618 ( 
.A(n_2094),
.Y(n_2618)
);

INVx3_ASAP7_75t_L g2619 ( 
.A(n_2236),
.Y(n_2619)
);

INVx2_ASAP7_75t_L g2620 ( 
.A(n_2207),
.Y(n_2620)
);

INVxp67_ASAP7_75t_L g2621 ( 
.A(n_2407),
.Y(n_2621)
);

INVx8_ASAP7_75t_L g2622 ( 
.A(n_2293),
.Y(n_2622)
);

BUFx2_ASAP7_75t_L g2623 ( 
.A(n_2066),
.Y(n_2623)
);

INVx1_ASAP7_75t_L g2624 ( 
.A(n_2108),
.Y(n_2624)
);

INVx3_ASAP7_75t_L g2625 ( 
.A(n_2237),
.Y(n_2625)
);

INVx2_ASAP7_75t_L g2626 ( 
.A(n_2207),
.Y(n_2626)
);

BUFx6f_ASAP7_75t_L g2627 ( 
.A(n_2064),
.Y(n_2627)
);

NAND3xp33_ASAP7_75t_L g2628 ( 
.A(n_2251),
.B(n_2279),
.C(n_2287),
.Y(n_2628)
);

NAND2xp5_ASAP7_75t_L g2629 ( 
.A(n_2127),
.B(n_1750),
.Y(n_2629)
);

INVx2_ASAP7_75t_L g2630 ( 
.A(n_2213),
.Y(n_2630)
);

INVx3_ASAP7_75t_L g2631 ( 
.A(n_2237),
.Y(n_2631)
);

NOR2xp33_ASAP7_75t_L g2632 ( 
.A(n_2266),
.B(n_1765),
.Y(n_2632)
);

INVx2_ASAP7_75t_L g2633 ( 
.A(n_2213),
.Y(n_2633)
);

NAND2xp5_ASAP7_75t_SL g2634 ( 
.A(n_2479),
.B(n_1850),
.Y(n_2634)
);

BUFx4f_ASAP7_75t_L g2635 ( 
.A(n_2097),
.Y(n_2635)
);

INVx3_ASAP7_75t_L g2636 ( 
.A(n_2240),
.Y(n_2636)
);

AO21x2_ASAP7_75t_L g2637 ( 
.A1(n_2372),
.A2(n_1995),
.B(n_1969),
.Y(n_2637)
);

NAND2xp5_ASAP7_75t_L g2638 ( 
.A(n_2134),
.B(n_1969),
.Y(n_2638)
);

INVx8_ASAP7_75t_L g2639 ( 
.A(n_2293),
.Y(n_2639)
);

INVxp33_ASAP7_75t_L g2640 ( 
.A(n_2105),
.Y(n_2640)
);

INVx1_ASAP7_75t_SL g2641 ( 
.A(n_2286),
.Y(n_2641)
);

BUFx3_ASAP7_75t_L g2642 ( 
.A(n_2103),
.Y(n_2642)
);

NAND2xp5_ASAP7_75t_SL g2643 ( 
.A(n_2266),
.B(n_1850),
.Y(n_2643)
);

INVx1_ASAP7_75t_L g2644 ( 
.A(n_2109),
.Y(n_2644)
);

INVx2_ASAP7_75t_SL g2645 ( 
.A(n_2386),
.Y(n_2645)
);

NAND3xp33_ASAP7_75t_L g2646 ( 
.A(n_2251),
.B(n_1931),
.C(n_1927),
.Y(n_2646)
);

INVx1_ASAP7_75t_L g2647 ( 
.A(n_2110),
.Y(n_2647)
);

INVx2_ASAP7_75t_SL g2648 ( 
.A(n_2131),
.Y(n_2648)
);

NAND2xp5_ASAP7_75t_L g2649 ( 
.A(n_2136),
.B(n_1995),
.Y(n_2649)
);

AND2x2_ASAP7_75t_L g2650 ( 
.A(n_2457),
.B(n_1701),
.Y(n_2650)
);

INVx2_ASAP7_75t_L g2651 ( 
.A(n_2165),
.Y(n_2651)
);

BUFx2_ASAP7_75t_L g2652 ( 
.A(n_2083),
.Y(n_2652)
);

INVx1_ASAP7_75t_L g2653 ( 
.A(n_2303),
.Y(n_2653)
);

INVx1_ASAP7_75t_L g2654 ( 
.A(n_2305),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_2308),
.Y(n_2655)
);

OR2x2_ASAP7_75t_L g2656 ( 
.A(n_2452),
.B(n_1463),
.Y(n_2656)
);

NOR2xp33_ASAP7_75t_L g2657 ( 
.A(n_2277),
.B(n_1963),
.Y(n_2657)
);

INVx2_ASAP7_75t_SL g2658 ( 
.A(n_2131),
.Y(n_2658)
);

INVx1_ASAP7_75t_L g2659 ( 
.A(n_2319),
.Y(n_2659)
);

INVx2_ASAP7_75t_L g2660 ( 
.A(n_2165),
.Y(n_2660)
);

NAND2xp5_ASAP7_75t_SL g2661 ( 
.A(n_2277),
.B(n_1843),
.Y(n_2661)
);

INVx2_ASAP7_75t_L g2662 ( 
.A(n_2165),
.Y(n_2662)
);

NAND2xp5_ASAP7_75t_L g2663 ( 
.A(n_2143),
.B(n_2015),
.Y(n_2663)
);

BUFx3_ASAP7_75t_L g2664 ( 
.A(n_2103),
.Y(n_2664)
);

NOR2xp33_ASAP7_75t_L g2665 ( 
.A(n_2287),
.B(n_1963),
.Y(n_2665)
);

AO21x2_ASAP7_75t_L g2666 ( 
.A1(n_2344),
.A2(n_2036),
.B(n_2015),
.Y(n_2666)
);

NAND2xp5_ASAP7_75t_SL g2667 ( 
.A(n_2320),
.B(n_1965),
.Y(n_2667)
);

BUFx6f_ASAP7_75t_L g2668 ( 
.A(n_2064),
.Y(n_2668)
);

INVx1_ASAP7_75t_L g2669 ( 
.A(n_2390),
.Y(n_2669)
);

NAND2xp5_ASAP7_75t_SL g2670 ( 
.A(n_2320),
.B(n_1973),
.Y(n_2670)
);

NAND3xp33_ASAP7_75t_L g2671 ( 
.A(n_2279),
.B(n_1994),
.C(n_1974),
.Y(n_2671)
);

INVx2_ASAP7_75t_L g2672 ( 
.A(n_2240),
.Y(n_2672)
);

INVx2_ASAP7_75t_L g2673 ( 
.A(n_2298),
.Y(n_2673)
);

BUFx3_ASAP7_75t_L g2674 ( 
.A(n_2149),
.Y(n_2674)
);

AOI22xp33_ASAP7_75t_L g2675 ( 
.A1(n_2298),
.A2(n_1701),
.B1(n_1753),
.B2(n_2052),
.Y(n_2675)
);

AND2x2_ASAP7_75t_L g2676 ( 
.A(n_2459),
.B(n_1753),
.Y(n_2676)
);

AOI22xp33_ASAP7_75t_L g2677 ( 
.A1(n_2298),
.A2(n_2060),
.B1(n_2052),
.B2(n_1994),
.Y(n_2677)
);

INVx3_ASAP7_75t_L g2678 ( 
.A(n_2453),
.Y(n_2678)
);

INVx3_ASAP7_75t_L g2679 ( 
.A(n_2453),
.Y(n_2679)
);

INVx3_ASAP7_75t_L g2680 ( 
.A(n_2454),
.Y(n_2680)
);

AND3x2_ASAP7_75t_L g2681 ( 
.A(n_2469),
.B(n_1734),
.C(n_1800),
.Y(n_2681)
);

INVx2_ASAP7_75t_SL g2682 ( 
.A(n_2176),
.Y(n_2682)
);

INVxp33_ASAP7_75t_L g2683 ( 
.A(n_2111),
.Y(n_2683)
);

INVx1_ASAP7_75t_L g2684 ( 
.A(n_2374),
.Y(n_2684)
);

INVx2_ASAP7_75t_L g2685 ( 
.A(n_2340),
.Y(n_2685)
);

INVx2_ASAP7_75t_L g2686 ( 
.A(n_2340),
.Y(n_2686)
);

INVx1_ASAP7_75t_L g2687 ( 
.A(n_2381),
.Y(n_2687)
);

INVx2_ASAP7_75t_L g2688 ( 
.A(n_2340),
.Y(n_2688)
);

AND2x2_ASAP7_75t_L g2689 ( 
.A(n_2480),
.B(n_1990),
.Y(n_2689)
);

INVx2_ASAP7_75t_L g2690 ( 
.A(n_2253),
.Y(n_2690)
);

AOI21x1_ASAP7_75t_L g2691 ( 
.A1(n_2146),
.A2(n_2185),
.B(n_2163),
.Y(n_2691)
);

AND2x4_ASAP7_75t_L g2692 ( 
.A(n_2113),
.B(n_2063),
.Y(n_2692)
);

INVx2_ASAP7_75t_L g2693 ( 
.A(n_2253),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_2382),
.Y(n_2694)
);

INVx2_ASAP7_75t_L g2695 ( 
.A(n_2255),
.Y(n_2695)
);

INVxp33_ASAP7_75t_SL g2696 ( 
.A(n_2422),
.Y(n_2696)
);

NAND2xp5_ASAP7_75t_L g2697 ( 
.A(n_2201),
.B(n_2036),
.Y(n_2697)
);

HB1xp67_ASAP7_75t_L g2698 ( 
.A(n_2083),
.Y(n_2698)
);

INVx3_ASAP7_75t_L g2699 ( 
.A(n_2454),
.Y(n_2699)
);

INVx2_ASAP7_75t_L g2700 ( 
.A(n_2255),
.Y(n_2700)
);

BUFx6f_ASAP7_75t_L g2701 ( 
.A(n_2064),
.Y(n_2701)
);

INVx2_ASAP7_75t_SL g2702 ( 
.A(n_2176),
.Y(n_2702)
);

INVx2_ASAP7_75t_SL g2703 ( 
.A(n_2205),
.Y(n_2703)
);

INVx2_ASAP7_75t_L g2704 ( 
.A(n_2257),
.Y(n_2704)
);

INVx3_ASAP7_75t_L g2705 ( 
.A(n_2464),
.Y(n_2705)
);

INVx2_ASAP7_75t_L g2706 ( 
.A(n_2257),
.Y(n_2706)
);

OR2x2_ASAP7_75t_L g2707 ( 
.A(n_2088),
.B(n_1478),
.Y(n_2707)
);

NOR2xp33_ASAP7_75t_L g2708 ( 
.A(n_2343),
.B(n_1974),
.Y(n_2708)
);

INVx2_ASAP7_75t_L g2709 ( 
.A(n_2263),
.Y(n_2709)
);

INVx1_ASAP7_75t_L g2710 ( 
.A(n_2385),
.Y(n_2710)
);

INVx1_ASAP7_75t_L g2711 ( 
.A(n_2480),
.Y(n_2711)
);

INVx2_ASAP7_75t_L g2712 ( 
.A(n_2263),
.Y(n_2712)
);

NAND2xp5_ASAP7_75t_L g2713 ( 
.A(n_2209),
.B(n_2042),
.Y(n_2713)
);

OR2x6_ASAP7_75t_L g2714 ( 
.A(n_2099),
.B(n_1864),
.Y(n_2714)
);

INVx2_ASAP7_75t_L g2715 ( 
.A(n_2265),
.Y(n_2715)
);

INVx1_ASAP7_75t_L g2716 ( 
.A(n_2082),
.Y(n_2716)
);

INVxp33_ASAP7_75t_L g2717 ( 
.A(n_2128),
.Y(n_2717)
);

INVx2_ASAP7_75t_L g2718 ( 
.A(n_2265),
.Y(n_2718)
);

INVx2_ASAP7_75t_L g2719 ( 
.A(n_2278),
.Y(n_2719)
);

INVx2_ASAP7_75t_SL g2720 ( 
.A(n_2205),
.Y(n_2720)
);

INVx1_ASAP7_75t_L g2721 ( 
.A(n_2082),
.Y(n_2721)
);

INVx2_ASAP7_75t_L g2722 ( 
.A(n_2278),
.Y(n_2722)
);

INVx5_ASAP7_75t_L g2723 ( 
.A(n_2404),
.Y(n_2723)
);

INVx11_ASAP7_75t_L g2724 ( 
.A(n_2118),
.Y(n_2724)
);

NAND2xp5_ASAP7_75t_L g2725 ( 
.A(n_2225),
.B(n_2042),
.Y(n_2725)
);

INVx2_ASAP7_75t_L g2726 ( 
.A(n_2284),
.Y(n_2726)
);

INVx2_ASAP7_75t_L g2727 ( 
.A(n_2284),
.Y(n_2727)
);

INVx2_ASAP7_75t_L g2728 ( 
.A(n_2297),
.Y(n_2728)
);

INVx1_ASAP7_75t_L g2729 ( 
.A(n_2082),
.Y(n_2729)
);

INVx2_ASAP7_75t_L g2730 ( 
.A(n_2297),
.Y(n_2730)
);

INVx2_ASAP7_75t_L g2731 ( 
.A(n_2306),
.Y(n_2731)
);

INVx1_ASAP7_75t_L g2732 ( 
.A(n_2321),
.Y(n_2732)
);

NOR2xp33_ASAP7_75t_L g2733 ( 
.A(n_2343),
.B(n_2006),
.Y(n_2733)
);

OAI22xp5_ASAP7_75t_L g2734 ( 
.A1(n_2472),
.A2(n_2040),
.B1(n_2060),
.B2(n_2006),
.Y(n_2734)
);

NAND2xp5_ASAP7_75t_SL g2735 ( 
.A(n_2472),
.B(n_2026),
.Y(n_2735)
);

INVx2_ASAP7_75t_L g2736 ( 
.A(n_2306),
.Y(n_2736)
);

INVx1_ASAP7_75t_L g2737 ( 
.A(n_2329),
.Y(n_2737)
);

AND3x2_ASAP7_75t_L g2738 ( 
.A(n_2088),
.B(n_1734),
.C(n_1808),
.Y(n_2738)
);

INVx1_ASAP7_75t_L g2739 ( 
.A(n_2330),
.Y(n_2739)
);

NAND2xp5_ASAP7_75t_L g2740 ( 
.A(n_2360),
.B(n_2045),
.Y(n_2740)
);

BUFx10_ASAP7_75t_L g2741 ( 
.A(n_2087),
.Y(n_2741)
);

INVx2_ASAP7_75t_L g2742 ( 
.A(n_2315),
.Y(n_2742)
);

CKINVDCx5p33_ASAP7_75t_R g2743 ( 
.A(n_2422),
.Y(n_2743)
);

NOR2xp33_ASAP7_75t_SL g2744 ( 
.A(n_2087),
.B(n_1886),
.Y(n_2744)
);

INVx3_ASAP7_75t_L g2745 ( 
.A(n_2464),
.Y(n_2745)
);

INVx1_ASAP7_75t_L g2746 ( 
.A(n_2338),
.Y(n_2746)
);

INVx2_ASAP7_75t_L g2747 ( 
.A(n_2315),
.Y(n_2747)
);

INVx2_ASAP7_75t_L g2748 ( 
.A(n_2317),
.Y(n_2748)
);

INVx1_ASAP7_75t_L g2749 ( 
.A(n_2345),
.Y(n_2749)
);

INVx2_ASAP7_75t_L g2750 ( 
.A(n_2317),
.Y(n_2750)
);

AND3x2_ASAP7_75t_L g2751 ( 
.A(n_2258),
.B(n_1943),
.C(n_1924),
.Y(n_2751)
);

INVx2_ASAP7_75t_L g2752 ( 
.A(n_2328),
.Y(n_2752)
);

INVx2_ASAP7_75t_L g2753 ( 
.A(n_2328),
.Y(n_2753)
);

NAND2xp5_ASAP7_75t_L g2754 ( 
.A(n_2375),
.B(n_2045),
.Y(n_2754)
);

INVxp67_ASAP7_75t_L g2755 ( 
.A(n_2162),
.Y(n_2755)
);

INVx1_ASAP7_75t_L g2756 ( 
.A(n_2347),
.Y(n_2756)
);

INVx2_ASAP7_75t_L g2757 ( 
.A(n_2332),
.Y(n_2757)
);

INVx4_ASAP7_75t_L g2758 ( 
.A(n_2462),
.Y(n_2758)
);

NAND2xp5_ASAP7_75t_L g2759 ( 
.A(n_2395),
.B(n_2040),
.Y(n_2759)
);

INVx1_ASAP7_75t_L g2760 ( 
.A(n_2348),
.Y(n_2760)
);

INVx2_ASAP7_75t_L g2761 ( 
.A(n_2332),
.Y(n_2761)
);

NOR2xp33_ASAP7_75t_L g2762 ( 
.A(n_2324),
.B(n_1882),
.Y(n_2762)
);

INVx2_ASAP7_75t_L g2763 ( 
.A(n_2339),
.Y(n_2763)
);

INVx3_ASAP7_75t_L g2764 ( 
.A(n_2339),
.Y(n_2764)
);

BUFx3_ASAP7_75t_L g2765 ( 
.A(n_2149),
.Y(n_2765)
);

INVx2_ASAP7_75t_L g2766 ( 
.A(n_2342),
.Y(n_2766)
);

INVx1_ASAP7_75t_L g2767 ( 
.A(n_2365),
.Y(n_2767)
);

INVxp67_ASAP7_75t_SL g2768 ( 
.A(n_2342),
.Y(n_2768)
);

INVx3_ASAP7_75t_L g2769 ( 
.A(n_2351),
.Y(n_2769)
);

INVx2_ASAP7_75t_L g2770 ( 
.A(n_2351),
.Y(n_2770)
);

NAND2xp5_ASAP7_75t_L g2771 ( 
.A(n_2406),
.B(n_2011),
.Y(n_2771)
);

NOR2xp33_ASAP7_75t_L g2772 ( 
.A(n_2324),
.B(n_1882),
.Y(n_2772)
);

NAND2xp5_ASAP7_75t_L g2773 ( 
.A(n_2466),
.B(n_2016),
.Y(n_2773)
);

BUFx2_ASAP7_75t_L g2774 ( 
.A(n_2203),
.Y(n_2774)
);

NAND3xp33_ASAP7_75t_L g2775 ( 
.A(n_2384),
.B(n_2031),
.C(n_1896),
.Y(n_2775)
);

NAND2xp5_ASAP7_75t_SL g2776 ( 
.A(n_2326),
.B(n_2026),
.Y(n_2776)
);

INVx2_ASAP7_75t_L g2777 ( 
.A(n_2352),
.Y(n_2777)
);

INVx2_ASAP7_75t_L g2778 ( 
.A(n_2352),
.Y(n_2778)
);

INVx2_ASAP7_75t_L g2779 ( 
.A(n_2353),
.Y(n_2779)
);

INVx2_ASAP7_75t_L g2780 ( 
.A(n_2353),
.Y(n_2780)
);

INVx2_ASAP7_75t_L g2781 ( 
.A(n_2354),
.Y(n_2781)
);

INVx2_ASAP7_75t_L g2782 ( 
.A(n_2354),
.Y(n_2782)
);

NOR2xp33_ASAP7_75t_L g2783 ( 
.A(n_2341),
.B(n_1889),
.Y(n_2783)
);

INVx1_ASAP7_75t_L g2784 ( 
.A(n_2368),
.Y(n_2784)
);

BUFx6f_ASAP7_75t_SL g2785 ( 
.A(n_2429),
.Y(n_2785)
);

BUFx10_ASAP7_75t_L g2786 ( 
.A(n_2107),
.Y(n_2786)
);

INVx1_ASAP7_75t_L g2787 ( 
.A(n_2369),
.Y(n_2787)
);

INVx1_ASAP7_75t_L g2788 ( 
.A(n_2114),
.Y(n_2788)
);

INVx2_ASAP7_75t_L g2789 ( 
.A(n_2361),
.Y(n_2789)
);

INVx2_ASAP7_75t_L g2790 ( 
.A(n_2361),
.Y(n_2790)
);

INVx1_ASAP7_75t_L g2791 ( 
.A(n_2116),
.Y(n_2791)
);

NAND2xp5_ASAP7_75t_L g2792 ( 
.A(n_2466),
.B(n_1999),
.Y(n_2792)
);

BUFx3_ASAP7_75t_L g2793 ( 
.A(n_2149),
.Y(n_2793)
);

BUFx6f_ASAP7_75t_L g2794 ( 
.A(n_2070),
.Y(n_2794)
);

NAND2xp5_ASAP7_75t_L g2795 ( 
.A(n_2466),
.B(n_1999),
.Y(n_2795)
);

BUFx6f_ASAP7_75t_L g2796 ( 
.A(n_2070),
.Y(n_2796)
);

INVx1_ASAP7_75t_L g2797 ( 
.A(n_2117),
.Y(n_2797)
);

INVx2_ASAP7_75t_SL g2798 ( 
.A(n_2107),
.Y(n_2798)
);

INVx2_ASAP7_75t_L g2799 ( 
.A(n_2367),
.Y(n_2799)
);

NAND2xp5_ASAP7_75t_L g2800 ( 
.A(n_2409),
.B(n_1999),
.Y(n_2800)
);

NAND2xp5_ASAP7_75t_SL g2801 ( 
.A(n_2326),
.B(n_1988),
.Y(n_2801)
);

INVx2_ASAP7_75t_SL g2802 ( 
.A(n_2115),
.Y(n_2802)
);

NAND2xp5_ASAP7_75t_SL g2803 ( 
.A(n_2341),
.B(n_1998),
.Y(n_2803)
);

INVx1_ASAP7_75t_L g2804 ( 
.A(n_2119),
.Y(n_2804)
);

NOR2xp33_ASAP7_75t_L g2805 ( 
.A(n_2268),
.B(n_1889),
.Y(n_2805)
);

INVx2_ASAP7_75t_L g2806 ( 
.A(n_2367),
.Y(n_2806)
);

INVx3_ASAP7_75t_L g2807 ( 
.A(n_2371),
.Y(n_2807)
);

INVx1_ASAP7_75t_L g2808 ( 
.A(n_2124),
.Y(n_2808)
);

BUFx2_ASAP7_75t_L g2809 ( 
.A(n_2229),
.Y(n_2809)
);

INVx1_ASAP7_75t_L g2810 ( 
.A(n_2125),
.Y(n_2810)
);

BUFx6f_ASAP7_75t_L g2811 ( 
.A(n_2070),
.Y(n_2811)
);

INVx1_ASAP7_75t_L g2812 ( 
.A(n_2126),
.Y(n_2812)
);

NAND2xp5_ASAP7_75t_SL g2813 ( 
.A(n_2331),
.B(n_1896),
.Y(n_2813)
);

INVx3_ASAP7_75t_L g2814 ( 
.A(n_2371),
.Y(n_2814)
);

INVx3_ASAP7_75t_L g2815 ( 
.A(n_2377),
.Y(n_2815)
);

NAND2xp5_ASAP7_75t_L g2816 ( 
.A(n_2414),
.B(n_2014),
.Y(n_2816)
);

INVx1_ASAP7_75t_L g2817 ( 
.A(n_2130),
.Y(n_2817)
);

OA22x2_ASAP7_75t_L g2818 ( 
.A1(n_2182),
.A2(n_1920),
.B1(n_1953),
.B2(n_1916),
.Y(n_2818)
);

INVx2_ASAP7_75t_L g2819 ( 
.A(n_2377),
.Y(n_2819)
);

NOR2xp33_ASAP7_75t_L g2820 ( 
.A(n_2281),
.B(n_1916),
.Y(n_2820)
);

NAND2xp5_ASAP7_75t_L g2821 ( 
.A(n_2419),
.B(n_2014),
.Y(n_2821)
);

INVx1_ASAP7_75t_L g2822 ( 
.A(n_2135),
.Y(n_2822)
);

NAND2xp5_ASAP7_75t_SL g2823 ( 
.A(n_2295),
.B(n_1920),
.Y(n_2823)
);

INVx2_ASAP7_75t_L g2824 ( 
.A(n_2387),
.Y(n_2824)
);

NAND2xp5_ASAP7_75t_SL g2825 ( 
.A(n_2311),
.B(n_2337),
.Y(n_2825)
);

INVx2_ASAP7_75t_SL g2826 ( 
.A(n_2115),
.Y(n_2826)
);

INVx2_ASAP7_75t_L g2827 ( 
.A(n_2387),
.Y(n_2827)
);

BUFx6f_ASAP7_75t_SL g2828 ( 
.A(n_2429),
.Y(n_2828)
);

BUFx10_ASAP7_75t_L g2829 ( 
.A(n_2140),
.Y(n_2829)
);

INVx1_ASAP7_75t_L g2830 ( 
.A(n_2362),
.Y(n_2830)
);

INVx1_ASAP7_75t_L g2831 ( 
.A(n_2362),
.Y(n_2831)
);

BUFx6f_ASAP7_75t_SL g2832 ( 
.A(n_2099),
.Y(n_2832)
);

INVx2_ASAP7_75t_L g2833 ( 
.A(n_2391),
.Y(n_2833)
);

INVx3_ASAP7_75t_L g2834 ( 
.A(n_2391),
.Y(n_2834)
);

INVx2_ASAP7_75t_SL g2835 ( 
.A(n_2140),
.Y(n_2835)
);

NAND2xp5_ASAP7_75t_SL g2836 ( 
.A(n_2346),
.B(n_1953),
.Y(n_2836)
);

INVx2_ASAP7_75t_L g2837 ( 
.A(n_2399),
.Y(n_2837)
);

NAND2xp5_ASAP7_75t_SL g2838 ( 
.A(n_2431),
.B(n_2008),
.Y(n_2838)
);

CKINVDCx5p33_ASAP7_75t_R g2839 ( 
.A(n_2269),
.Y(n_2839)
);

OAI22xp33_ASAP7_75t_L g2840 ( 
.A1(n_2243),
.A2(n_2032),
.B1(n_2008),
.B2(n_1639),
.Y(n_2840)
);

INVx2_ASAP7_75t_L g2841 ( 
.A(n_2399),
.Y(n_2841)
);

BUFx2_ASAP7_75t_L g2842 ( 
.A(n_2175),
.Y(n_2842)
);

INVx1_ASAP7_75t_L g2843 ( 
.A(n_2362),
.Y(n_2843)
);

AND2x2_ASAP7_75t_L g2844 ( 
.A(n_2090),
.B(n_2032),
.Y(n_2844)
);

AOI22xp5_ASAP7_75t_L g2845 ( 
.A1(n_2097),
.A2(n_1907),
.B1(n_1914),
.B2(n_1901),
.Y(n_2845)
);

INVx2_ASAP7_75t_L g2846 ( 
.A(n_2400),
.Y(n_2846)
);

INVxp67_ASAP7_75t_SL g2847 ( 
.A(n_2400),
.Y(n_2847)
);

INVx2_ASAP7_75t_SL g2848 ( 
.A(n_2208),
.Y(n_2848)
);

INVxp33_ASAP7_75t_L g2849 ( 
.A(n_2282),
.Y(n_2849)
);

NAND2xp5_ASAP7_75t_SL g2850 ( 
.A(n_2441),
.B(n_1732),
.Y(n_2850)
);

NOR2xp33_ASAP7_75t_L g2851 ( 
.A(n_2249),
.B(n_1634),
.Y(n_2851)
);

BUFx6f_ASAP7_75t_L g2852 ( 
.A(n_2070),
.Y(n_2852)
);

BUFx6f_ASAP7_75t_L g2853 ( 
.A(n_2075),
.Y(n_2853)
);

INVx1_ASAP7_75t_L g2854 ( 
.A(n_2151),
.Y(n_2854)
);

INVx1_ASAP7_75t_L g2855 ( 
.A(n_2090),
.Y(n_2855)
);

NAND2xp5_ASAP7_75t_L g2856 ( 
.A(n_2244),
.B(n_2248),
.Y(n_2856)
);

INVx1_ASAP7_75t_L g2857 ( 
.A(n_2090),
.Y(n_2857)
);

INVx1_ASAP7_75t_L g2858 ( 
.A(n_2313),
.Y(n_2858)
);

NAND2xp5_ASAP7_75t_SL g2859 ( 
.A(n_2215),
.B(n_1873),
.Y(n_2859)
);

NOR2xp33_ASAP7_75t_L g2860 ( 
.A(n_2226),
.B(n_1873),
.Y(n_2860)
);

INVxp67_ASAP7_75t_L g2861 ( 
.A(n_2198),
.Y(n_2861)
);

NOR2xp33_ASAP7_75t_L g2862 ( 
.A(n_2226),
.B(n_1979),
.Y(n_2862)
);

AO22x2_ASAP7_75t_L g2863 ( 
.A1(n_2282),
.A2(n_1075),
.B1(n_1079),
.B2(n_1072),
.Y(n_2863)
);

INVx2_ASAP7_75t_L g2864 ( 
.A(n_2408),
.Y(n_2864)
);

AOI22xp33_ASAP7_75t_L g2865 ( 
.A1(n_2244),
.A2(n_2014),
.B1(n_1788),
.B2(n_1811),
.Y(n_2865)
);

INVx2_ASAP7_75t_L g2866 ( 
.A(n_2408),
.Y(n_2866)
);

INVx3_ASAP7_75t_L g2867 ( 
.A(n_2413),
.Y(n_2867)
);

INVx2_ASAP7_75t_L g2868 ( 
.A(n_2413),
.Y(n_2868)
);

BUFx6f_ASAP7_75t_L g2869 ( 
.A(n_2075),
.Y(n_2869)
);

INVx5_ASAP7_75t_L g2870 ( 
.A(n_2404),
.Y(n_2870)
);

INVx2_ASAP7_75t_L g2871 ( 
.A(n_2415),
.Y(n_2871)
);

NAND2xp5_ASAP7_75t_L g2872 ( 
.A(n_2244),
.B(n_2014),
.Y(n_2872)
);

INVx3_ASAP7_75t_L g2873 ( 
.A(n_2415),
.Y(n_2873)
);

INVx1_ASAP7_75t_L g2874 ( 
.A(n_2313),
.Y(n_2874)
);

AO21x2_ASAP7_75t_L g2875 ( 
.A1(n_2272),
.A2(n_2044),
.B(n_2029),
.Y(n_2875)
);

INVx1_ASAP7_75t_L g2876 ( 
.A(n_2316),
.Y(n_2876)
);

INVx1_ASAP7_75t_L g2877 ( 
.A(n_2316),
.Y(n_2877)
);

NAND2xp5_ASAP7_75t_L g2878 ( 
.A(n_2097),
.B(n_2014),
.Y(n_2878)
);

INVx2_ASAP7_75t_L g2879 ( 
.A(n_2423),
.Y(n_2879)
);

INVx2_ASAP7_75t_L g2880 ( 
.A(n_2423),
.Y(n_2880)
);

NOR2xp33_ASAP7_75t_L g2881 ( 
.A(n_2157),
.B(n_1979),
.Y(n_2881)
);

INVx2_ASAP7_75t_L g2882 ( 
.A(n_2430),
.Y(n_2882)
);

NOR2xp33_ASAP7_75t_L g2883 ( 
.A(n_2210),
.B(n_1991),
.Y(n_2883)
);

INVx1_ASAP7_75t_L g2884 ( 
.A(n_2325),
.Y(n_2884)
);

NAND2xp5_ASAP7_75t_L g2885 ( 
.A(n_2097),
.B(n_1826),
.Y(n_2885)
);

INVx2_ASAP7_75t_L g2886 ( 
.A(n_2430),
.Y(n_2886)
);

BUFx6f_ASAP7_75t_L g2887 ( 
.A(n_2075),
.Y(n_2887)
);

OAI22xp33_ASAP7_75t_L g2888 ( 
.A1(n_2099),
.A2(n_1933),
.B1(n_1942),
.B2(n_1936),
.Y(n_2888)
);

INVx1_ASAP7_75t_L g2889 ( 
.A(n_2325),
.Y(n_2889)
);

NAND2xp5_ASAP7_75t_SL g2890 ( 
.A(n_2198),
.B(n_1991),
.Y(n_2890)
);

NAND2xp5_ASAP7_75t_L g2891 ( 
.A(n_2097),
.B(n_1826),
.Y(n_2891)
);

INVx1_ASAP7_75t_L g2892 ( 
.A(n_2412),
.Y(n_2892)
);

NAND2xp5_ASAP7_75t_L g2893 ( 
.A(n_2137),
.B(n_1834),
.Y(n_2893)
);

INVxp67_ASAP7_75t_SL g2894 ( 
.A(n_2462),
.Y(n_2894)
);

NOR2xp33_ASAP7_75t_L g2895 ( 
.A(n_2101),
.B(n_2051),
.Y(n_2895)
);

INVx1_ASAP7_75t_L g2896 ( 
.A(n_2412),
.Y(n_2896)
);

INVx2_ASAP7_75t_L g2897 ( 
.A(n_2141),
.Y(n_2897)
);

NAND2xp5_ASAP7_75t_SL g2898 ( 
.A(n_2275),
.B(n_1819),
.Y(n_2898)
);

NAND2xp5_ASAP7_75t_L g2899 ( 
.A(n_2144),
.B(n_1834),
.Y(n_2899)
);

INVx1_ASAP7_75t_L g2900 ( 
.A(n_2440),
.Y(n_2900)
);

INVx2_ASAP7_75t_L g2901 ( 
.A(n_2150),
.Y(n_2901)
);

OR2x6_ASAP7_75t_L g2902 ( 
.A(n_2156),
.B(n_1977),
.Y(n_2902)
);

OR2x2_ASAP7_75t_L g2903 ( 
.A(n_2392),
.B(n_834),
.Y(n_2903)
);

INVx2_ASAP7_75t_L g2904 ( 
.A(n_2445),
.Y(n_2904)
);

INVx1_ASAP7_75t_L g2905 ( 
.A(n_2440),
.Y(n_2905)
);

INVx1_ASAP7_75t_L g2906 ( 
.A(n_2208),
.Y(n_2906)
);

NOR2xp33_ASAP7_75t_L g2907 ( 
.A(n_2101),
.B(n_2035),
.Y(n_2907)
);

BUFx6f_ASAP7_75t_L g2908 ( 
.A(n_2075),
.Y(n_2908)
);

AOI21x1_ASAP7_75t_L g2909 ( 
.A1(n_2296),
.A2(n_2044),
.B(n_2029),
.Y(n_2909)
);

INVx1_ASAP7_75t_L g2910 ( 
.A(n_2233),
.Y(n_2910)
);

NAND2xp5_ASAP7_75t_L g2911 ( 
.A(n_2355),
.B(n_1834),
.Y(n_2911)
);

NAND2xp5_ASAP7_75t_SL g2912 ( 
.A(n_2302),
.B(n_1819),
.Y(n_2912)
);

NOR2xp33_ASAP7_75t_L g2913 ( 
.A(n_2657),
.B(n_2200),
.Y(n_2913)
);

NOR2xp33_ASAP7_75t_L g2914 ( 
.A(n_2665),
.B(n_1367),
.Y(n_2914)
);

AND2x2_ASAP7_75t_L g2915 ( 
.A(n_2536),
.B(n_2183),
.Y(n_2915)
);

XOR2xp5_ASAP7_75t_L g2916 ( 
.A(n_2849),
.B(n_2474),
.Y(n_2916)
);

INVx1_ASAP7_75t_L g2917 ( 
.A(n_2482),
.Y(n_2917)
);

INVx1_ASAP7_75t_L g2918 ( 
.A(n_2482),
.Y(n_2918)
);

INVx1_ASAP7_75t_L g2919 ( 
.A(n_2488),
.Y(n_2919)
);

INVx1_ASAP7_75t_L g2920 ( 
.A(n_2488),
.Y(n_2920)
);

INVx1_ASAP7_75t_SL g2921 ( 
.A(n_2652),
.Y(n_2921)
);

INVx1_ASAP7_75t_L g2922 ( 
.A(n_2490),
.Y(n_2922)
);

AND2x2_ASAP7_75t_L g2923 ( 
.A(n_2536),
.B(n_2183),
.Y(n_2923)
);

INVx1_ASAP7_75t_L g2924 ( 
.A(n_2490),
.Y(n_2924)
);

INVx1_ASAP7_75t_L g2925 ( 
.A(n_2491),
.Y(n_2925)
);

INVx1_ASAP7_75t_L g2926 ( 
.A(n_2491),
.Y(n_2926)
);

XNOR2xp5_ASAP7_75t_L g2927 ( 
.A(n_2849),
.B(n_2474),
.Y(n_2927)
);

INVx1_ASAP7_75t_L g2928 ( 
.A(n_2493),
.Y(n_2928)
);

INVx2_ASAP7_75t_L g2929 ( 
.A(n_2493),
.Y(n_2929)
);

CKINVDCx20_ASAP7_75t_R g2930 ( 
.A(n_2530),
.Y(n_2930)
);

INVx1_ASAP7_75t_L g2931 ( 
.A(n_2494),
.Y(n_2931)
);

INVx1_ASAP7_75t_L g2932 ( 
.A(n_2494),
.Y(n_2932)
);

XOR2x2_ASAP7_75t_L g2933 ( 
.A(n_2574),
.B(n_2182),
.Y(n_2933)
);

NOR2xp67_ASAP7_75t_L g2934 ( 
.A(n_2895),
.B(n_1711),
.Y(n_2934)
);

INVxp67_ASAP7_75t_SL g2935 ( 
.A(n_2584),
.Y(n_2935)
);

INVx1_ASAP7_75t_L g2936 ( 
.A(n_2503),
.Y(n_2936)
);

INVx1_ASAP7_75t_L g2937 ( 
.A(n_2503),
.Y(n_2937)
);

INVx1_ASAP7_75t_L g2938 ( 
.A(n_2504),
.Y(n_2938)
);

NOR2xp33_ASAP7_75t_L g2939 ( 
.A(n_2708),
.B(n_1367),
.Y(n_2939)
);

INVx2_ASAP7_75t_SL g2940 ( 
.A(n_2590),
.Y(n_2940)
);

INVx1_ASAP7_75t_L g2941 ( 
.A(n_2504),
.Y(n_2941)
);

INVx1_ASAP7_75t_L g2942 ( 
.A(n_2507),
.Y(n_2942)
);

CKINVDCx20_ASAP7_75t_R g2943 ( 
.A(n_2530),
.Y(n_2943)
);

AND2x4_ASAP7_75t_L g2944 ( 
.A(n_2642),
.B(n_2310),
.Y(n_2944)
);

NAND2xp5_ASAP7_75t_L g2945 ( 
.A(n_2589),
.B(n_2404),
.Y(n_2945)
);

NOR2xp33_ASAP7_75t_L g2946 ( 
.A(n_2733),
.B(n_1373),
.Y(n_2946)
);

XOR2xp5_ASAP7_75t_L g2947 ( 
.A(n_2696),
.B(n_1373),
.Y(n_2947)
);

INVx1_ASAP7_75t_L g2948 ( 
.A(n_2507),
.Y(n_2948)
);

CKINVDCx20_ASAP7_75t_R g2949 ( 
.A(n_2839),
.Y(n_2949)
);

INVx1_ASAP7_75t_L g2950 ( 
.A(n_2509),
.Y(n_2950)
);

AND2x2_ASAP7_75t_L g2951 ( 
.A(n_2594),
.B(n_2310),
.Y(n_2951)
);

CKINVDCx16_ASAP7_75t_R g2952 ( 
.A(n_2744),
.Y(n_2952)
);

AND2x4_ASAP7_75t_L g2953 ( 
.A(n_2642),
.B(n_2233),
.Y(n_2953)
);

AOI21x1_ASAP7_75t_L g2954 ( 
.A1(n_2872),
.A2(n_2288),
.B(n_2481),
.Y(n_2954)
);

INVxp33_ASAP7_75t_SL g2955 ( 
.A(n_2497),
.Y(n_2955)
);

NOR2xp33_ASAP7_75t_L g2956 ( 
.A(n_2628),
.B(n_2219),
.Y(n_2956)
);

CKINVDCx20_ASAP7_75t_R g2957 ( 
.A(n_2839),
.Y(n_2957)
);

XOR2xp5_ASAP7_75t_L g2958 ( 
.A(n_2696),
.B(n_1380),
.Y(n_2958)
);

INVx1_ASAP7_75t_L g2959 ( 
.A(n_2509),
.Y(n_2959)
);

INVx1_ASAP7_75t_L g2960 ( 
.A(n_2511),
.Y(n_2960)
);

NOR2xp33_ASAP7_75t_L g2961 ( 
.A(n_2508),
.B(n_2219),
.Y(n_2961)
);

NOR2xp33_ASAP7_75t_L g2962 ( 
.A(n_2661),
.B(n_2230),
.Y(n_2962)
);

INVx2_ASAP7_75t_L g2963 ( 
.A(n_2511),
.Y(n_2963)
);

NOR2xp33_ASAP7_75t_L g2964 ( 
.A(n_2661),
.B(n_2230),
.Y(n_2964)
);

INVx1_ASAP7_75t_L g2965 ( 
.A(n_2516),
.Y(n_2965)
);

NAND2xp5_ASAP7_75t_SL g2966 ( 
.A(n_2557),
.B(n_2363),
.Y(n_2966)
);

NOR2xp33_ASAP7_75t_L g2967 ( 
.A(n_2667),
.B(n_2380),
.Y(n_2967)
);

NOR2xp33_ASAP7_75t_L g2968 ( 
.A(n_2667),
.B(n_2380),
.Y(n_2968)
);

INVx1_ASAP7_75t_L g2969 ( 
.A(n_2516),
.Y(n_2969)
);

INVx1_ASAP7_75t_L g2970 ( 
.A(n_2517),
.Y(n_2970)
);

INVx2_ASAP7_75t_SL g2971 ( 
.A(n_2698),
.Y(n_2971)
);

INVx1_ASAP7_75t_L g2972 ( 
.A(n_2517),
.Y(n_2972)
);

INVx1_ASAP7_75t_L g2973 ( 
.A(n_2522),
.Y(n_2973)
);

NOR2xp33_ASAP7_75t_L g2974 ( 
.A(n_2510),
.B(n_1380),
.Y(n_2974)
);

INVx1_ASAP7_75t_SL g2975 ( 
.A(n_2641),
.Y(n_2975)
);

CKINVDCx5p33_ASAP7_75t_R g2976 ( 
.A(n_2497),
.Y(n_2976)
);

INVx2_ASAP7_75t_L g2977 ( 
.A(n_2522),
.Y(n_2977)
);

INVx1_ASAP7_75t_L g2978 ( 
.A(n_2523),
.Y(n_2978)
);

INVx1_ASAP7_75t_L g2979 ( 
.A(n_2523),
.Y(n_2979)
);

INVx1_ASAP7_75t_L g2980 ( 
.A(n_2525),
.Y(n_2980)
);

INVxp33_ASAP7_75t_L g2981 ( 
.A(n_2707),
.Y(n_2981)
);

CKINVDCx20_ASAP7_75t_R g2982 ( 
.A(n_2498),
.Y(n_2982)
);

NOR2xp33_ASAP7_75t_L g2983 ( 
.A(n_2540),
.B(n_1381),
.Y(n_2983)
);

INVx1_ASAP7_75t_L g2984 ( 
.A(n_2525),
.Y(n_2984)
);

INVx1_ASAP7_75t_L g2985 ( 
.A(n_2529),
.Y(n_2985)
);

NOR2xp33_ASAP7_75t_L g2986 ( 
.A(n_2573),
.B(n_1381),
.Y(n_2986)
);

INVx1_ASAP7_75t_L g2987 ( 
.A(n_2529),
.Y(n_2987)
);

INVx2_ASAP7_75t_L g2988 ( 
.A(n_2533),
.Y(n_2988)
);

AND2x6_ASAP7_75t_L g2989 ( 
.A(n_2651),
.B(n_2438),
.Y(n_2989)
);

INVx1_ASAP7_75t_L g2990 ( 
.A(n_2533),
.Y(n_2990)
);

INVx1_ASAP7_75t_L g2991 ( 
.A(n_2535),
.Y(n_2991)
);

AND2x2_ASAP7_75t_L g2992 ( 
.A(n_2594),
.B(n_2235),
.Y(n_2992)
);

INVx1_ASAP7_75t_L g2993 ( 
.A(n_2535),
.Y(n_2993)
);

OR2x6_ASAP7_75t_L g2994 ( 
.A(n_2902),
.B(n_2714),
.Y(n_2994)
);

NAND2xp5_ASAP7_75t_L g2995 ( 
.A(n_2638),
.B(n_2404),
.Y(n_2995)
);

INVxp33_ASAP7_75t_L g2996 ( 
.A(n_2707),
.Y(n_2996)
);

AND2x2_ASAP7_75t_L g2997 ( 
.A(n_2595),
.B(n_2617),
.Y(n_2997)
);

INVx1_ASAP7_75t_L g2998 ( 
.A(n_2542),
.Y(n_2998)
);

CKINVDCx20_ASAP7_75t_R g2999 ( 
.A(n_2498),
.Y(n_2999)
);

AOI21xp5_ASAP7_75t_L g3000 ( 
.A1(n_2856),
.A2(n_2289),
.B(n_2364),
.Y(n_3000)
);

HB1xp67_ASAP7_75t_L g3001 ( 
.A(n_2842),
.Y(n_3001)
);

OR2x2_ASAP7_75t_L g3002 ( 
.A(n_2656),
.B(n_2123),
.Y(n_3002)
);

AND2x2_ASAP7_75t_L g3003 ( 
.A(n_2595),
.B(n_2235),
.Y(n_3003)
);

AND2x6_ASAP7_75t_L g3004 ( 
.A(n_2651),
.B(n_2252),
.Y(n_3004)
);

INVx1_ASAP7_75t_L g3005 ( 
.A(n_2542),
.Y(n_3005)
);

NAND2xp5_ASAP7_75t_L g3006 ( 
.A(n_2649),
.B(n_2663),
.Y(n_3006)
);

INVx1_ASAP7_75t_L g3007 ( 
.A(n_2546),
.Y(n_3007)
);

INVx1_ASAP7_75t_L g3008 ( 
.A(n_2546),
.Y(n_3008)
);

HB1xp67_ASAP7_75t_L g3009 ( 
.A(n_2648),
.Y(n_3009)
);

NAND2xp33_ASAP7_75t_R g3010 ( 
.A(n_2512),
.B(n_2232),
.Y(n_3010)
);

INVx2_ASAP7_75t_L g3011 ( 
.A(n_2548),
.Y(n_3011)
);

XOR2xp5_ASAP7_75t_L g3012 ( 
.A(n_2743),
.B(n_1433),
.Y(n_3012)
);

NOR2xp67_ASAP7_75t_L g3013 ( 
.A(n_2907),
.B(n_2327),
.Y(n_3013)
);

INVx1_ASAP7_75t_L g3014 ( 
.A(n_2548),
.Y(n_3014)
);

INVx1_ASAP7_75t_L g3015 ( 
.A(n_2559),
.Y(n_3015)
);

INVxp33_ASAP7_75t_L g3016 ( 
.A(n_2560),
.Y(n_3016)
);

NOR2xp33_ASAP7_75t_L g3017 ( 
.A(n_2576),
.B(n_1433),
.Y(n_3017)
);

INVx1_ASAP7_75t_L g3018 ( 
.A(n_2559),
.Y(n_3018)
);

INVx1_ASAP7_75t_L g3019 ( 
.A(n_2561),
.Y(n_3019)
);

AND2x2_ASAP7_75t_L g3020 ( 
.A(n_2617),
.B(n_2650),
.Y(n_3020)
);

BUFx6f_ASAP7_75t_SL g3021 ( 
.A(n_2902),
.Y(n_3021)
);

INVxp67_ASAP7_75t_SL g3022 ( 
.A(n_2584),
.Y(n_3022)
);

INVx1_ASAP7_75t_L g3023 ( 
.A(n_2561),
.Y(n_3023)
);

INVx1_ASAP7_75t_SL g3024 ( 
.A(n_2623),
.Y(n_3024)
);

INVxp33_ASAP7_75t_L g3025 ( 
.A(n_2560),
.Y(n_3025)
);

INVx1_ASAP7_75t_L g3026 ( 
.A(n_2562),
.Y(n_3026)
);

INVx1_ASAP7_75t_L g3027 ( 
.A(n_2562),
.Y(n_3027)
);

INVx1_ASAP7_75t_L g3028 ( 
.A(n_2567),
.Y(n_3028)
);

AND2x4_ASAP7_75t_L g3029 ( 
.A(n_2664),
.B(n_2252),
.Y(n_3029)
);

INVx1_ASAP7_75t_L g3030 ( 
.A(n_2567),
.Y(n_3030)
);

INVx1_ASAP7_75t_L g3031 ( 
.A(n_2570),
.Y(n_3031)
);

AND2x2_ASAP7_75t_L g3032 ( 
.A(n_2650),
.B(n_2086),
.Y(n_3032)
);

NOR2xp33_ASAP7_75t_SL g3033 ( 
.A(n_2599),
.B(n_2232),
.Y(n_3033)
);

NOR2xp33_ASAP7_75t_L g3034 ( 
.A(n_2670),
.B(n_2334),
.Y(n_3034)
);

INVx1_ASAP7_75t_L g3035 ( 
.A(n_2570),
.Y(n_3035)
);

INVx1_ASAP7_75t_L g3036 ( 
.A(n_2571),
.Y(n_3036)
);

INVx1_ASAP7_75t_L g3037 ( 
.A(n_2571),
.Y(n_3037)
);

INVx1_ASAP7_75t_L g3038 ( 
.A(n_2579),
.Y(n_3038)
);

INVxp67_ASAP7_75t_L g3039 ( 
.A(n_2656),
.Y(n_3039)
);

XNOR2xp5_ASAP7_75t_L g3040 ( 
.A(n_2743),
.B(n_2274),
.Y(n_3040)
);

INVx1_ASAP7_75t_L g3041 ( 
.A(n_2579),
.Y(n_3041)
);

AND2x2_ASAP7_75t_L g3042 ( 
.A(n_2676),
.B(n_2393),
.Y(n_3042)
);

INVx4_ASAP7_75t_SL g3043 ( 
.A(n_2528),
.Y(n_3043)
);

INVx1_ASAP7_75t_L g3044 ( 
.A(n_2580),
.Y(n_3044)
);

NAND2xp5_ASAP7_75t_L g3045 ( 
.A(n_2697),
.B(n_2293),
.Y(n_3045)
);

INVx1_ASAP7_75t_L g3046 ( 
.A(n_2580),
.Y(n_3046)
);

OR2x2_ASAP7_75t_L g3047 ( 
.A(n_2759),
.B(n_2366),
.Y(n_3047)
);

INVx2_ASAP7_75t_L g3048 ( 
.A(n_2587),
.Y(n_3048)
);

INVx2_ASAP7_75t_L g3049 ( 
.A(n_2587),
.Y(n_3049)
);

INVxp33_ASAP7_75t_L g3050 ( 
.A(n_2903),
.Y(n_3050)
);

INVx2_ASAP7_75t_L g3051 ( 
.A(n_2604),
.Y(n_3051)
);

INVx2_ASAP7_75t_L g3052 ( 
.A(n_2604),
.Y(n_3052)
);

NAND2xp33_ASAP7_75t_R g3053 ( 
.A(n_2512),
.B(n_2334),
.Y(n_3053)
);

AND2x2_ASAP7_75t_L g3054 ( 
.A(n_2676),
.B(n_2393),
.Y(n_3054)
);

INVx1_ASAP7_75t_L g3055 ( 
.A(n_2605),
.Y(n_3055)
);

INVx1_ASAP7_75t_L g3056 ( 
.A(n_2605),
.Y(n_3056)
);

INVx2_ASAP7_75t_SL g3057 ( 
.A(n_2648),
.Y(n_3057)
);

INVx1_ASAP7_75t_L g3058 ( 
.A(n_2615),
.Y(n_3058)
);

INVxp33_ASAP7_75t_L g3059 ( 
.A(n_2903),
.Y(n_3059)
);

NAND2xp5_ASAP7_75t_L g3060 ( 
.A(n_2713),
.B(n_2355),
.Y(n_3060)
);

BUFx5_ASAP7_75t_L g3061 ( 
.A(n_2528),
.Y(n_3061)
);

INVx1_ASAP7_75t_L g3062 ( 
.A(n_2615),
.Y(n_3062)
);

BUFx6f_ASAP7_75t_L g3063 ( 
.A(n_2485),
.Y(n_3063)
);

OR2x6_ASAP7_75t_L g3064 ( 
.A(n_2902),
.B(n_2156),
.Y(n_3064)
);

BUFx6f_ASAP7_75t_L g3065 ( 
.A(n_2485),
.Y(n_3065)
);

INVx2_ASAP7_75t_L g3066 ( 
.A(n_2620),
.Y(n_3066)
);

CKINVDCx20_ASAP7_75t_R g3067 ( 
.A(n_2774),
.Y(n_3067)
);

NAND2xp5_ASAP7_75t_L g3068 ( 
.A(n_2725),
.B(n_2355),
.Y(n_3068)
);

INVx1_ASAP7_75t_L g3069 ( 
.A(n_2620),
.Y(n_3069)
);

NOR2xp33_ASAP7_75t_L g3070 ( 
.A(n_2646),
.B(n_1448),
.Y(n_3070)
);

INVx1_ASAP7_75t_L g3071 ( 
.A(n_2626),
.Y(n_3071)
);

INVx1_ASAP7_75t_L g3072 ( 
.A(n_2626),
.Y(n_3072)
);

INVx1_ASAP7_75t_L g3073 ( 
.A(n_2630),
.Y(n_3073)
);

NOR2xp33_ASAP7_75t_L g3074 ( 
.A(n_2671),
.B(n_2632),
.Y(n_3074)
);

AND2x4_ASAP7_75t_L g3075 ( 
.A(n_2664),
.B(n_2154),
.Y(n_3075)
);

INVx1_ASAP7_75t_L g3076 ( 
.A(n_2630),
.Y(n_3076)
);

INVx1_ASAP7_75t_L g3077 ( 
.A(n_2633),
.Y(n_3077)
);

OR2x6_ASAP7_75t_L g3078 ( 
.A(n_2902),
.B(n_2156),
.Y(n_3078)
);

NOR2xp33_ASAP7_75t_L g3079 ( 
.A(n_2502),
.B(n_1448),
.Y(n_3079)
);

AND2x2_ASAP7_75t_L g3080 ( 
.A(n_2500),
.B(n_2424),
.Y(n_3080)
);

INVx1_ASAP7_75t_L g3081 ( 
.A(n_2633),
.Y(n_3081)
);

INVx1_ASAP7_75t_L g3082 ( 
.A(n_2585),
.Y(n_3082)
);

INVx1_ASAP7_75t_L g3083 ( 
.A(n_2592),
.Y(n_3083)
);

XOR2xp5_ASAP7_75t_L g3084 ( 
.A(n_2486),
.B(n_1462),
.Y(n_3084)
);

NAND2xp5_ASAP7_75t_SL g3085 ( 
.A(n_2572),
.B(n_2314),
.Y(n_3085)
);

INVx1_ASAP7_75t_L g3086 ( 
.A(n_2603),
.Y(n_3086)
);

INVx2_ASAP7_75t_L g3087 ( 
.A(n_2672),
.Y(n_3087)
);

NOR2xp33_ASAP7_75t_SL g3088 ( 
.A(n_2762),
.B(n_2355),
.Y(n_3088)
);

NOR2xp33_ASAP7_75t_L g3089 ( 
.A(n_2670),
.B(n_2424),
.Y(n_3089)
);

CKINVDCx5p33_ASAP7_75t_R g3090 ( 
.A(n_2724),
.Y(n_3090)
);

AND2x2_ASAP7_75t_SL g3091 ( 
.A(n_2851),
.B(n_2122),
.Y(n_3091)
);

AND2x2_ASAP7_75t_L g3092 ( 
.A(n_2500),
.B(n_2621),
.Y(n_3092)
);

AND2x2_ASAP7_75t_L g3093 ( 
.A(n_2689),
.B(n_1411),
.Y(n_3093)
);

INVx1_ASAP7_75t_L g3094 ( 
.A(n_2608),
.Y(n_3094)
);

AND2x2_ASAP7_75t_L g3095 ( 
.A(n_2689),
.B(n_1483),
.Y(n_3095)
);

NOR2xp67_ASAP7_75t_L g3096 ( 
.A(n_2881),
.B(n_2158),
.Y(n_3096)
);

BUFx8_ASAP7_75t_L g3097 ( 
.A(n_2565),
.Y(n_3097)
);

XOR2x2_ASAP7_75t_L g3098 ( 
.A(n_2734),
.B(n_1781),
.Y(n_3098)
);

NOR2xp33_ASAP7_75t_L g3099 ( 
.A(n_2640),
.B(n_2160),
.Y(n_3099)
);

INVx1_ASAP7_75t_L g3100 ( 
.A(n_2613),
.Y(n_3100)
);

INVxp67_ASAP7_75t_SL g3101 ( 
.A(n_2584),
.Y(n_3101)
);

INVx1_ASAP7_75t_L g3102 ( 
.A(n_2614),
.Y(n_3102)
);

INVx1_ASAP7_75t_L g3103 ( 
.A(n_2618),
.Y(n_3103)
);

INVx1_ASAP7_75t_L g3104 ( 
.A(n_2624),
.Y(n_3104)
);

INVx1_ASAP7_75t_L g3105 ( 
.A(n_2644),
.Y(n_3105)
);

NAND2xp5_ASAP7_75t_L g3106 ( 
.A(n_2740),
.B(n_2355),
.Y(n_3106)
);

INVx1_ASAP7_75t_L g3107 ( 
.A(n_2647),
.Y(n_3107)
);

INVx1_ASAP7_75t_L g3108 ( 
.A(n_2732),
.Y(n_3108)
);

AND2x4_ASAP7_75t_L g3109 ( 
.A(n_2674),
.B(n_2164),
.Y(n_3109)
);

INVx1_ASAP7_75t_L g3110 ( 
.A(n_2737),
.Y(n_3110)
);

INVx1_ASAP7_75t_L g3111 ( 
.A(n_2739),
.Y(n_3111)
);

INVx1_ASAP7_75t_L g3112 ( 
.A(n_2746),
.Y(n_3112)
);

BUFx12f_ASAP7_75t_L g3113 ( 
.A(n_2483),
.Y(n_3113)
);

AND2x2_ASAP7_75t_L g3114 ( 
.A(n_2658),
.B(n_1483),
.Y(n_3114)
);

INVx2_ASAP7_75t_L g3115 ( 
.A(n_2672),
.Y(n_3115)
);

INVx1_ASAP7_75t_L g3116 ( 
.A(n_2749),
.Y(n_3116)
);

INVx1_ASAP7_75t_L g3117 ( 
.A(n_2756),
.Y(n_3117)
);

INVx2_ASAP7_75t_L g3118 ( 
.A(n_2690),
.Y(n_3118)
);

INVx1_ASAP7_75t_L g3119 ( 
.A(n_2760),
.Y(n_3119)
);

AND2x6_ASAP7_75t_L g3120 ( 
.A(n_2660),
.B(n_1075),
.Y(n_3120)
);

NOR2xp33_ASAP7_75t_L g3121 ( 
.A(n_2805),
.B(n_1462),
.Y(n_3121)
);

AND2x2_ASAP7_75t_L g3122 ( 
.A(n_2658),
.B(n_1494),
.Y(n_3122)
);

OR2x2_ASAP7_75t_L g3123 ( 
.A(n_2645),
.B(n_2611),
.Y(n_3123)
);

XOR2xp5_ASAP7_75t_L g3124 ( 
.A(n_2845),
.B(n_1511),
.Y(n_3124)
);

XOR2xp5_ASAP7_75t_L g3125 ( 
.A(n_2640),
.B(n_1511),
.Y(n_3125)
);

INVx2_ASAP7_75t_L g3126 ( 
.A(n_2690),
.Y(n_3126)
);

INVx1_ASAP7_75t_L g3127 ( 
.A(n_2767),
.Y(n_3127)
);

INVx1_ASAP7_75t_L g3128 ( 
.A(n_2784),
.Y(n_3128)
);

NAND2xp5_ASAP7_75t_L g3129 ( 
.A(n_2754),
.B(n_2447),
.Y(n_3129)
);

NAND2xp5_ASAP7_75t_L g3130 ( 
.A(n_2556),
.B(n_2449),
.Y(n_3130)
);

INVx1_ASAP7_75t_L g3131 ( 
.A(n_2787),
.Y(n_3131)
);

INVx1_ASAP7_75t_L g3132 ( 
.A(n_2492),
.Y(n_3132)
);

AND2x2_ASAP7_75t_L g3133 ( 
.A(n_2844),
.B(n_1494),
.Y(n_3133)
);

NOR2xp33_ASAP7_75t_L g3134 ( 
.A(n_2820),
.B(n_1520),
.Y(n_3134)
);

INVx1_ASAP7_75t_L g3135 ( 
.A(n_2505),
.Y(n_3135)
);

XOR2xp5_ASAP7_75t_L g3136 ( 
.A(n_2683),
.B(n_1520),
.Y(n_3136)
);

INVx1_ASAP7_75t_L g3137 ( 
.A(n_2506),
.Y(n_3137)
);

BUFx5_ASAP7_75t_L g3138 ( 
.A(n_2528),
.Y(n_3138)
);

CKINVDCx5p33_ASAP7_75t_R g3139 ( 
.A(n_2724),
.Y(n_3139)
);

INVx1_ASAP7_75t_L g3140 ( 
.A(n_2520),
.Y(n_3140)
);

AND2x2_ASAP7_75t_L g3141 ( 
.A(n_2844),
.B(n_1495),
.Y(n_3141)
);

INVx2_ASAP7_75t_L g3142 ( 
.A(n_2693),
.Y(n_3142)
);

INVx4_ASAP7_75t_L g3143 ( 
.A(n_2485),
.Y(n_3143)
);

INVx1_ASAP7_75t_L g3144 ( 
.A(n_2521),
.Y(n_3144)
);

INVx1_ASAP7_75t_L g3145 ( 
.A(n_2524),
.Y(n_3145)
);

INVxp33_ASAP7_75t_L g3146 ( 
.A(n_2813),
.Y(n_3146)
);

INVx1_ASAP7_75t_L g3147 ( 
.A(n_2534),
.Y(n_3147)
);

INVx1_ASAP7_75t_L g3148 ( 
.A(n_2537),
.Y(n_3148)
);

INVx1_ASAP7_75t_L g3149 ( 
.A(n_2538),
.Y(n_3149)
);

AND2x2_ASAP7_75t_L g3150 ( 
.A(n_2645),
.B(n_1495),
.Y(n_3150)
);

INVx1_ASAP7_75t_L g3151 ( 
.A(n_2539),
.Y(n_3151)
);

XOR2xp5_ASAP7_75t_L g3152 ( 
.A(n_2683),
.B(n_1535),
.Y(n_3152)
);

INVxp33_ASAP7_75t_L g3153 ( 
.A(n_2813),
.Y(n_3153)
);

INVx1_ASAP7_75t_L g3154 ( 
.A(n_2543),
.Y(n_3154)
);

HB1xp67_ASAP7_75t_L g3155 ( 
.A(n_2611),
.Y(n_3155)
);

XNOR2xp5_ASAP7_75t_SL g3156 ( 
.A(n_2681),
.B(n_1868),
.Y(n_3156)
);

INVx1_ASAP7_75t_L g3157 ( 
.A(n_2544),
.Y(n_3157)
);

INVx1_ASAP7_75t_L g3158 ( 
.A(n_2549),
.Y(n_3158)
);

INVx1_ASAP7_75t_L g3159 ( 
.A(n_2550),
.Y(n_3159)
);

BUFx6f_ASAP7_75t_SL g3160 ( 
.A(n_2714),
.Y(n_3160)
);

HB1xp67_ASAP7_75t_L g3161 ( 
.A(n_2755),
.Y(n_3161)
);

INVx1_ASAP7_75t_L g3162 ( 
.A(n_2553),
.Y(n_3162)
);

NOR2xp33_ASAP7_75t_L g3163 ( 
.A(n_2717),
.B(n_2170),
.Y(n_3163)
);

AND2x2_ASAP7_75t_L g3164 ( 
.A(n_2717),
.B(n_1502),
.Y(n_3164)
);

XOR2xp5_ASAP7_75t_L g3165 ( 
.A(n_2809),
.B(n_1535),
.Y(n_3165)
);

AND2x2_ASAP7_75t_SL g3166 ( 
.A(n_2860),
.B(n_2122),
.Y(n_3166)
);

AND2x4_ASAP7_75t_L g3167 ( 
.A(n_2674),
.B(n_2173),
.Y(n_3167)
);

INVx1_ASAP7_75t_L g3168 ( 
.A(n_2554),
.Y(n_3168)
);

AND2x2_ASAP7_75t_L g3169 ( 
.A(n_2487),
.B(n_1502),
.Y(n_3169)
);

INVx1_ASAP7_75t_L g3170 ( 
.A(n_2555),
.Y(n_3170)
);

INVx1_ASAP7_75t_L g3171 ( 
.A(n_2558),
.Y(n_3171)
);

XOR2xp5_ASAP7_75t_L g3172 ( 
.A(n_2775),
.B(n_1540),
.Y(n_3172)
);

INVx1_ASAP7_75t_L g3173 ( 
.A(n_2563),
.Y(n_3173)
);

AND2x2_ASAP7_75t_L g3174 ( 
.A(n_2487),
.B(n_1506),
.Y(n_3174)
);

AND2x4_ASAP7_75t_L g3175 ( 
.A(n_2765),
.B(n_2174),
.Y(n_3175)
);

INVx1_ASAP7_75t_L g3176 ( 
.A(n_2568),
.Y(n_3176)
);

INVx1_ASAP7_75t_L g3177 ( 
.A(n_2575),
.Y(n_3177)
);

CKINVDCx20_ASAP7_75t_R g3178 ( 
.A(n_2586),
.Y(n_3178)
);

HB1xp67_ASAP7_75t_L g3179 ( 
.A(n_2711),
.Y(n_3179)
);

INVx1_ASAP7_75t_L g3180 ( 
.A(n_2577),
.Y(n_3180)
);

INVx1_ASAP7_75t_L g3181 ( 
.A(n_2854),
.Y(n_3181)
);

INVx2_ASAP7_75t_L g3182 ( 
.A(n_2693),
.Y(n_3182)
);

INVxp33_ASAP7_75t_L g3183 ( 
.A(n_2836),
.Y(n_3183)
);

INVx1_ASAP7_75t_L g3184 ( 
.A(n_2897),
.Y(n_3184)
);

INVxp33_ASAP7_75t_L g3185 ( 
.A(n_2836),
.Y(n_3185)
);

BUFx6f_ASAP7_75t_L g3186 ( 
.A(n_2485),
.Y(n_3186)
);

INVx1_ASAP7_75t_L g3187 ( 
.A(n_2897),
.Y(n_3187)
);

INVx1_ASAP7_75t_L g3188 ( 
.A(n_2901),
.Y(n_3188)
);

INVx1_ASAP7_75t_L g3189 ( 
.A(n_2901),
.Y(n_3189)
);

AND2x2_ASAP7_75t_L g3190 ( 
.A(n_2771),
.B(n_1506),
.Y(n_3190)
);

INVx2_ASAP7_75t_L g3191 ( 
.A(n_2695),
.Y(n_3191)
);

CKINVDCx20_ASAP7_75t_R g3192 ( 
.A(n_2586),
.Y(n_3192)
);

AOI21xp5_ASAP7_75t_L g3193 ( 
.A1(n_2792),
.A2(n_2289),
.B(n_2364),
.Y(n_3193)
);

INVx1_ASAP7_75t_L g3194 ( 
.A(n_2904),
.Y(n_3194)
);

INVx1_ASAP7_75t_L g3195 ( 
.A(n_2904),
.Y(n_3195)
);

INVx1_ASAP7_75t_L g3196 ( 
.A(n_2716),
.Y(n_3196)
);

INVx1_ASAP7_75t_L g3197 ( 
.A(n_2721),
.Y(n_3197)
);

INVx2_ASAP7_75t_L g3198 ( 
.A(n_2695),
.Y(n_3198)
);

INVx1_ASAP7_75t_L g3199 ( 
.A(n_2729),
.Y(n_3199)
);

INVx1_ASAP7_75t_L g3200 ( 
.A(n_2788),
.Y(n_3200)
);

INVx2_ASAP7_75t_SL g3201 ( 
.A(n_2692),
.Y(n_3201)
);

AND2x2_ASAP7_75t_L g3202 ( 
.A(n_2601),
.B(n_1576),
.Y(n_3202)
);

NAND2xp33_ASAP7_75t_SL g3203 ( 
.A(n_2859),
.B(n_1253),
.Y(n_3203)
);

XNOR2x1_ASAP7_75t_L g3204 ( 
.A(n_2863),
.B(n_887),
.Y(n_3204)
);

INVx1_ASAP7_75t_L g3205 ( 
.A(n_2791),
.Y(n_3205)
);

OR2x2_ASAP7_75t_L g3206 ( 
.A(n_2801),
.B(n_2314),
.Y(n_3206)
);

INVx1_ASAP7_75t_L g3207 ( 
.A(n_2797),
.Y(n_3207)
);

AND2x2_ASAP7_75t_L g3208 ( 
.A(n_2609),
.B(n_1576),
.Y(n_3208)
);

XOR2xp5_ASAP7_75t_L g3209 ( 
.A(n_2825),
.B(n_1540),
.Y(n_3209)
);

INVx1_ASAP7_75t_L g3210 ( 
.A(n_2804),
.Y(n_3210)
);

INVx1_ASAP7_75t_L g3211 ( 
.A(n_2808),
.Y(n_3211)
);

INVx1_ASAP7_75t_L g3212 ( 
.A(n_2810),
.Y(n_3212)
);

INVx1_ASAP7_75t_L g3213 ( 
.A(n_2812),
.Y(n_3213)
);

XOR2xp5_ASAP7_75t_L g3214 ( 
.A(n_2825),
.B(n_1558),
.Y(n_3214)
);

INVx1_ASAP7_75t_L g3215 ( 
.A(n_2817),
.Y(n_3215)
);

NOR2xp33_ASAP7_75t_L g3216 ( 
.A(n_2495),
.B(n_2178),
.Y(n_3216)
);

INVx1_ASAP7_75t_L g3217 ( 
.A(n_2822),
.Y(n_3217)
);

INVx1_ASAP7_75t_L g3218 ( 
.A(n_2700),
.Y(n_3218)
);

INVx1_ASAP7_75t_L g3219 ( 
.A(n_2700),
.Y(n_3219)
);

INVx1_ASAP7_75t_L g3220 ( 
.A(n_2704),
.Y(n_3220)
);

INVx4_ASAP7_75t_SL g3221 ( 
.A(n_2528),
.Y(n_3221)
);

INVx2_ASAP7_75t_L g3222 ( 
.A(n_2704),
.Y(n_3222)
);

INVx1_ASAP7_75t_L g3223 ( 
.A(n_2706),
.Y(n_3223)
);

INVx1_ASAP7_75t_L g3224 ( 
.A(n_2706),
.Y(n_3224)
);

HB1xp67_ASAP7_75t_L g3225 ( 
.A(n_2861),
.Y(n_3225)
);

INVx1_ASAP7_75t_L g3226 ( 
.A(n_2709),
.Y(n_3226)
);

AND2x4_ASAP7_75t_L g3227 ( 
.A(n_2765),
.B(n_2180),
.Y(n_3227)
);

INVx1_ASAP7_75t_L g3228 ( 
.A(n_2709),
.Y(n_3228)
);

INVx1_ASAP7_75t_L g3229 ( 
.A(n_2712),
.Y(n_3229)
);

CKINVDCx5p33_ASAP7_75t_R g3230 ( 
.A(n_2565),
.Y(n_3230)
);

INVx1_ASAP7_75t_L g3231 ( 
.A(n_2712),
.Y(n_3231)
);

INVx1_ASAP7_75t_L g3232 ( 
.A(n_2715),
.Y(n_3232)
);

OAI21xp5_ASAP7_75t_L g3233 ( 
.A1(n_2673),
.A2(n_2168),
.B(n_2159),
.Y(n_3233)
);

BUFx2_ASAP7_75t_L g3234 ( 
.A(n_2518),
.Y(n_3234)
);

INVx1_ASAP7_75t_L g3235 ( 
.A(n_2715),
.Y(n_3235)
);

INVx1_ASAP7_75t_L g3236 ( 
.A(n_2718),
.Y(n_3236)
);

INVx1_ASAP7_75t_L g3237 ( 
.A(n_2718),
.Y(n_3237)
);

INVxp67_ASAP7_75t_SL g3238 ( 
.A(n_2584),
.Y(n_3238)
);

INVx1_ASAP7_75t_L g3239 ( 
.A(n_2719),
.Y(n_3239)
);

NOR2xp33_ASAP7_75t_L g3240 ( 
.A(n_2772),
.B(n_1558),
.Y(n_3240)
);

INVx1_ASAP7_75t_L g3241 ( 
.A(n_2719),
.Y(n_3241)
);

INVxp33_ASAP7_75t_L g3242 ( 
.A(n_2823),
.Y(n_3242)
);

INVx1_ASAP7_75t_L g3243 ( 
.A(n_2722),
.Y(n_3243)
);

INVx1_ASAP7_75t_L g3244 ( 
.A(n_2722),
.Y(n_3244)
);

INVx1_ASAP7_75t_L g3245 ( 
.A(n_2726),
.Y(n_3245)
);

INVx2_ASAP7_75t_L g3246 ( 
.A(n_2726),
.Y(n_3246)
);

BUFx5_ASAP7_75t_L g3247 ( 
.A(n_2528),
.Y(n_3247)
);

INVx2_ASAP7_75t_L g3248 ( 
.A(n_2727),
.Y(n_3248)
);

NAND2xp5_ASAP7_75t_L g3249 ( 
.A(n_2637),
.B(n_2450),
.Y(n_3249)
);

XOR2xp5_ASAP7_75t_L g3250 ( 
.A(n_2634),
.B(n_1595),
.Y(n_3250)
);

BUFx6f_ASAP7_75t_L g3251 ( 
.A(n_2532),
.Y(n_3251)
);

INVx1_ASAP7_75t_L g3252 ( 
.A(n_2727),
.Y(n_3252)
);

CKINVDCx20_ASAP7_75t_R g3253 ( 
.A(n_2602),
.Y(n_3253)
);

INVx1_ASAP7_75t_L g3254 ( 
.A(n_2728),
.Y(n_3254)
);

XNOR2xp5_ASAP7_75t_L g3255 ( 
.A(n_2751),
.B(n_1595),
.Y(n_3255)
);

NOR2xp33_ASAP7_75t_L g3256 ( 
.A(n_2783),
.B(n_1638),
.Y(n_3256)
);

XNOR2xp5_ASAP7_75t_L g3257 ( 
.A(n_2738),
.B(n_1638),
.Y(n_3257)
);

INVx1_ASAP7_75t_L g3258 ( 
.A(n_2728),
.Y(n_3258)
);

INVx1_ASAP7_75t_L g3259 ( 
.A(n_2730),
.Y(n_3259)
);

INVx1_ASAP7_75t_L g3260 ( 
.A(n_2730),
.Y(n_3260)
);

INVx1_ASAP7_75t_L g3261 ( 
.A(n_2731),
.Y(n_3261)
);

NOR2xp33_ASAP7_75t_L g3262 ( 
.A(n_2495),
.B(n_1641),
.Y(n_3262)
);

NOR2xp33_ASAP7_75t_L g3263 ( 
.A(n_2801),
.B(n_2181),
.Y(n_3263)
);

NAND2xp5_ASAP7_75t_L g3264 ( 
.A(n_2637),
.B(n_2451),
.Y(n_3264)
);

INVx1_ASAP7_75t_L g3265 ( 
.A(n_2731),
.Y(n_3265)
);

INVx1_ASAP7_75t_L g3266 ( 
.A(n_2736),
.Y(n_3266)
);

NOR2xp33_ASAP7_75t_L g3267 ( 
.A(n_2838),
.B(n_2187),
.Y(n_3267)
);

AND2x2_ASAP7_75t_L g3268 ( 
.A(n_2616),
.B(n_1621),
.Y(n_3268)
);

BUFx3_ASAP7_75t_L g3269 ( 
.A(n_2519),
.Y(n_3269)
);

INVx1_ASAP7_75t_L g3270 ( 
.A(n_2736),
.Y(n_3270)
);

CKINVDCx5p33_ASAP7_75t_R g3271 ( 
.A(n_2565),
.Y(n_3271)
);

INVx1_ASAP7_75t_L g3272 ( 
.A(n_2742),
.Y(n_3272)
);

INVx1_ASAP7_75t_L g3273 ( 
.A(n_2742),
.Y(n_3273)
);

CKINVDCx5p33_ASAP7_75t_R g3274 ( 
.A(n_2785),
.Y(n_3274)
);

AND2x2_ASAP7_75t_L g3275 ( 
.A(n_2629),
.B(n_1621),
.Y(n_3275)
);

INVx1_ASAP7_75t_L g3276 ( 
.A(n_2747),
.Y(n_3276)
);

XOR2xp5_ASAP7_75t_L g3277 ( 
.A(n_2634),
.B(n_1641),
.Y(n_3277)
);

INVxp33_ASAP7_75t_L g3278 ( 
.A(n_2823),
.Y(n_3278)
);

NAND2xp5_ASAP7_75t_L g3279 ( 
.A(n_2637),
.B(n_2691),
.Y(n_3279)
);

INVxp33_ASAP7_75t_L g3280 ( 
.A(n_2838),
.Y(n_3280)
);

INVx1_ASAP7_75t_L g3281 ( 
.A(n_2747),
.Y(n_3281)
);

OR2x2_ASAP7_75t_L g3282 ( 
.A(n_2489),
.B(n_2191),
.Y(n_3282)
);

AND2x2_ASAP7_75t_L g3283 ( 
.A(n_2682),
.B(n_1678),
.Y(n_3283)
);

BUFx8_ASAP7_75t_L g3284 ( 
.A(n_2785),
.Y(n_3284)
);

INVx2_ASAP7_75t_L g3285 ( 
.A(n_2748),
.Y(n_3285)
);

INVx1_ASAP7_75t_L g3286 ( 
.A(n_2748),
.Y(n_3286)
);

INVx1_ASAP7_75t_L g3287 ( 
.A(n_2750),
.Y(n_3287)
);

INVx2_ASAP7_75t_L g3288 ( 
.A(n_2750),
.Y(n_3288)
);

INVx2_ASAP7_75t_L g3289 ( 
.A(n_2752),
.Y(n_3289)
);

INVx2_ASAP7_75t_L g3290 ( 
.A(n_2752),
.Y(n_3290)
);

INVx1_ASAP7_75t_L g3291 ( 
.A(n_2753),
.Y(n_3291)
);

INVx1_ASAP7_75t_L g3292 ( 
.A(n_2753),
.Y(n_3292)
);

INVx1_ASAP7_75t_L g3293 ( 
.A(n_2757),
.Y(n_3293)
);

NAND2xp5_ASAP7_75t_L g3294 ( 
.A(n_2773),
.B(n_2159),
.Y(n_3294)
);

CKINVDCx16_ASAP7_75t_R g3295 ( 
.A(n_2785),
.Y(n_3295)
);

INVx1_ASAP7_75t_L g3296 ( 
.A(n_2757),
.Y(n_3296)
);

INVx1_ASAP7_75t_L g3297 ( 
.A(n_2761),
.Y(n_3297)
);

INVxp33_ASAP7_75t_SL g3298 ( 
.A(n_2862),
.Y(n_3298)
);

INVxp33_ASAP7_75t_L g3299 ( 
.A(n_2863),
.Y(n_3299)
);

INVx2_ASAP7_75t_L g3300 ( 
.A(n_2761),
.Y(n_3300)
);

INVx1_ASAP7_75t_L g3301 ( 
.A(n_2763),
.Y(n_3301)
);

AOI21xp5_ASAP7_75t_L g3302 ( 
.A1(n_2795),
.A2(n_2383),
.B(n_2168),
.Y(n_3302)
);

INVx2_ASAP7_75t_L g3303 ( 
.A(n_2763),
.Y(n_3303)
);

CKINVDCx20_ASAP7_75t_R g3304 ( 
.A(n_2602),
.Y(n_3304)
);

INVx1_ASAP7_75t_L g3305 ( 
.A(n_2766),
.Y(n_3305)
);

INVx1_ASAP7_75t_L g3306 ( 
.A(n_2766),
.Y(n_3306)
);

INVx1_ASAP7_75t_L g3307 ( 
.A(n_2770),
.Y(n_3307)
);

INVx1_ASAP7_75t_L g3308 ( 
.A(n_2770),
.Y(n_3308)
);

NAND2xp5_ASAP7_75t_L g3309 ( 
.A(n_2875),
.B(n_2193),
.Y(n_3309)
);

INVx1_ASAP7_75t_L g3310 ( 
.A(n_2777),
.Y(n_3310)
);

AND2x4_ASAP7_75t_L g3311 ( 
.A(n_2793),
.B(n_2194),
.Y(n_3311)
);

INVx1_ASAP7_75t_L g3312 ( 
.A(n_2777),
.Y(n_3312)
);

INVx1_ASAP7_75t_SL g3313 ( 
.A(n_2741),
.Y(n_3313)
);

XOR2xp5_ASAP7_75t_L g3314 ( 
.A(n_2526),
.B(n_1651),
.Y(n_3314)
);

INVx1_ASAP7_75t_L g3315 ( 
.A(n_2778),
.Y(n_3315)
);

INVxp33_ASAP7_75t_SL g3316 ( 
.A(n_2883),
.Y(n_3316)
);

NOR2xp33_ASAP7_75t_L g3317 ( 
.A(n_2602),
.B(n_2195),
.Y(n_3317)
);

INVx1_ASAP7_75t_L g3318 ( 
.A(n_2778),
.Y(n_3318)
);

INVx2_ASAP7_75t_L g3319 ( 
.A(n_2779),
.Y(n_3319)
);

BUFx3_ASAP7_75t_L g3320 ( 
.A(n_2519),
.Y(n_3320)
);

NOR2xp33_ASAP7_75t_L g3321 ( 
.A(n_2489),
.B(n_2197),
.Y(n_3321)
);

INVx2_ASAP7_75t_L g3322 ( 
.A(n_2779),
.Y(n_3322)
);

INVx1_ASAP7_75t_L g3323 ( 
.A(n_2780),
.Y(n_3323)
);

NAND2xp5_ASAP7_75t_L g3324 ( 
.A(n_2875),
.B(n_2206),
.Y(n_3324)
);

INVx1_ASAP7_75t_L g3325 ( 
.A(n_2780),
.Y(n_3325)
);

INVx1_ASAP7_75t_SL g3326 ( 
.A(n_2741),
.Y(n_3326)
);

BUFx6f_ASAP7_75t_L g3327 ( 
.A(n_2532),
.Y(n_3327)
);

INVx1_ASAP7_75t_L g3328 ( 
.A(n_2781),
.Y(n_3328)
);

NOR2xp33_ASAP7_75t_L g3329 ( 
.A(n_2643),
.B(n_1651),
.Y(n_3329)
);

INVx1_ASAP7_75t_L g3330 ( 
.A(n_2781),
.Y(n_3330)
);

AND2x2_ASAP7_75t_L g3331 ( 
.A(n_2682),
.B(n_1696),
.Y(n_3331)
);

INVxp67_ASAP7_75t_SL g3332 ( 
.A(n_2627),
.Y(n_3332)
);

XOR2xp5_ASAP7_75t_L g3333 ( 
.A(n_2526),
.B(n_2401),
.Y(n_3333)
);

BUFx6f_ASAP7_75t_L g3334 ( 
.A(n_2532),
.Y(n_3334)
);

NOR2xp33_ASAP7_75t_L g3335 ( 
.A(n_2643),
.B(n_1868),
.Y(n_3335)
);

INVx1_ASAP7_75t_L g3336 ( 
.A(n_2782),
.Y(n_3336)
);

INVx1_ASAP7_75t_L g3337 ( 
.A(n_2782),
.Y(n_3337)
);

INVx2_ASAP7_75t_L g3338 ( 
.A(n_2789),
.Y(n_3338)
);

INVx8_ASAP7_75t_L g3339 ( 
.A(n_2528),
.Y(n_3339)
);

INVx1_ASAP7_75t_L g3340 ( 
.A(n_2789),
.Y(n_3340)
);

NAND2xp33_ASAP7_75t_R g3341 ( 
.A(n_2692),
.B(n_1895),
.Y(n_3341)
);

INVx1_ASAP7_75t_L g3342 ( 
.A(n_2790),
.Y(n_3342)
);

INVx1_ASAP7_75t_L g3343 ( 
.A(n_2790),
.Y(n_3343)
);

AND2x2_ASAP7_75t_L g3344 ( 
.A(n_2702),
.B(n_2004),
.Y(n_3344)
);

INVx1_ASAP7_75t_L g3345 ( 
.A(n_2799),
.Y(n_3345)
);

XOR2xp5_ASAP7_75t_L g3346 ( 
.A(n_2818),
.B(n_2401),
.Y(n_3346)
);

INVx2_ASAP7_75t_L g3347 ( 
.A(n_2799),
.Y(n_3347)
);

INVx2_ASAP7_75t_L g3348 ( 
.A(n_3087),
.Y(n_3348)
);

NAND2xp5_ASAP7_75t_L g3349 ( 
.A(n_3006),
.B(n_2677),
.Y(n_3349)
);

NAND2xp5_ASAP7_75t_SL g3350 ( 
.A(n_3006),
.B(n_2741),
.Y(n_3350)
);

INVx2_ASAP7_75t_L g3351 ( 
.A(n_3115),
.Y(n_3351)
);

INVx2_ASAP7_75t_L g3352 ( 
.A(n_3118),
.Y(n_3352)
);

INVx4_ASAP7_75t_L g3353 ( 
.A(n_3063),
.Y(n_3353)
);

NAND2xp5_ASAP7_75t_SL g3354 ( 
.A(n_2961),
.B(n_2532),
.Y(n_3354)
);

NAND2xp5_ASAP7_75t_L g3355 ( 
.A(n_3020),
.B(n_2675),
.Y(n_3355)
);

NAND2xp5_ASAP7_75t_SL g3356 ( 
.A(n_2961),
.B(n_2545),
.Y(n_3356)
);

BUFx12f_ASAP7_75t_L g3357 ( 
.A(n_3097),
.Y(n_3357)
);

NAND2xp5_ASAP7_75t_L g3358 ( 
.A(n_3074),
.B(n_2875),
.Y(n_3358)
);

INVx2_ASAP7_75t_L g3359 ( 
.A(n_3126),
.Y(n_3359)
);

NAND2xp5_ASAP7_75t_L g3360 ( 
.A(n_3129),
.B(n_2514),
.Y(n_3360)
);

OAI221xp5_ASAP7_75t_L g3361 ( 
.A1(n_3240),
.A2(n_2803),
.B1(n_2501),
.B2(n_2703),
.C(n_2720),
.Y(n_3361)
);

NAND2x1_ASAP7_75t_L g3362 ( 
.A(n_3143),
.B(n_2612),
.Y(n_3362)
);

OAI221xp5_ASAP7_75t_L g3363 ( 
.A1(n_3256),
.A2(n_2803),
.B1(n_2501),
.B2(n_2703),
.C(n_2720),
.Y(n_3363)
);

NAND2xp5_ASAP7_75t_SL g3364 ( 
.A(n_3091),
.B(n_2545),
.Y(n_3364)
);

INVx8_ASAP7_75t_L g3365 ( 
.A(n_3064),
.Y(n_3365)
);

NAND2xp5_ASAP7_75t_L g3366 ( 
.A(n_3129),
.B(n_2514),
.Y(n_3366)
);

AOI22xp5_ASAP7_75t_L g3367 ( 
.A1(n_2956),
.A2(n_2552),
.B1(n_2566),
.B2(n_2531),
.Y(n_3367)
);

INVx2_ASAP7_75t_L g3368 ( 
.A(n_3142),
.Y(n_3368)
);

INVxp33_ASAP7_75t_L g3369 ( 
.A(n_3165),
.Y(n_3369)
);

NOR2xp33_ASAP7_75t_L g3370 ( 
.A(n_2913),
.B(n_2840),
.Y(n_3370)
);

INVx1_ASAP7_75t_L g3371 ( 
.A(n_3082),
.Y(n_3371)
);

NOR2xp33_ASAP7_75t_R g3372 ( 
.A(n_2976),
.B(n_3341),
.Y(n_3372)
);

NAND2xp5_ASAP7_75t_L g3373 ( 
.A(n_3042),
.B(n_2514),
.Y(n_3373)
);

AND2x4_ASAP7_75t_L g3374 ( 
.A(n_2944),
.B(n_2793),
.Y(n_3374)
);

NAND2xp5_ASAP7_75t_L g3375 ( 
.A(n_3054),
.B(n_2660),
.Y(n_3375)
);

NOR2xp33_ASAP7_75t_L g3376 ( 
.A(n_2913),
.B(n_2591),
.Y(n_3376)
);

NAND2xp5_ASAP7_75t_L g3377 ( 
.A(n_3190),
.B(n_2662),
.Y(n_3377)
);

NAND2xp5_ASAP7_75t_SL g3378 ( 
.A(n_3013),
.B(n_2545),
.Y(n_3378)
);

NAND2xp5_ASAP7_75t_L g3379 ( 
.A(n_2967),
.B(n_2662),
.Y(n_3379)
);

INVx4_ASAP7_75t_L g3380 ( 
.A(n_3063),
.Y(n_3380)
);

NAND2xp5_ASAP7_75t_L g3381 ( 
.A(n_2967),
.B(n_2673),
.Y(n_3381)
);

INVx1_ASAP7_75t_L g3382 ( 
.A(n_3083),
.Y(n_3382)
);

AOI22xp33_ASAP7_75t_L g3383 ( 
.A1(n_2997),
.A2(n_2818),
.B1(n_2776),
.B2(n_2830),
.Y(n_3383)
);

NAND2xp5_ASAP7_75t_L g3384 ( 
.A(n_2968),
.B(n_2685),
.Y(n_3384)
);

INVxp67_ASAP7_75t_L g3385 ( 
.A(n_2975),
.Y(n_3385)
);

NAND2xp5_ASAP7_75t_SL g3386 ( 
.A(n_2956),
.B(n_2962),
.Y(n_3386)
);

NAND2xp5_ASAP7_75t_SL g3387 ( 
.A(n_2962),
.B(n_2545),
.Y(n_3387)
);

AOI22xp33_ASAP7_75t_L g3388 ( 
.A1(n_3032),
.A2(n_2776),
.B1(n_2843),
.B2(n_2831),
.Y(n_3388)
);

INVx1_ASAP7_75t_L g3389 ( 
.A(n_3086),
.Y(n_3389)
);

AND2x2_ASAP7_75t_L g3390 ( 
.A(n_3133),
.B(n_2702),
.Y(n_3390)
);

AND2x4_ASAP7_75t_L g3391 ( 
.A(n_2944),
.B(n_2600),
.Y(n_3391)
);

OR2x2_ASAP7_75t_L g3392 ( 
.A(n_3039),
.B(n_2518),
.Y(n_3392)
);

NAND2xp5_ASAP7_75t_SL g3393 ( 
.A(n_2964),
.B(n_2597),
.Y(n_3393)
);

NOR2xp33_ASAP7_75t_L g3394 ( 
.A(n_2914),
.B(n_2591),
.Y(n_3394)
);

AOI22xp5_ASAP7_75t_L g3395 ( 
.A1(n_2964),
.A2(n_2531),
.B1(n_2566),
.B2(n_2552),
.Y(n_3395)
);

NAND2xp5_ASAP7_75t_L g3396 ( 
.A(n_2968),
.B(n_2685),
.Y(n_3396)
);

INVx1_ASAP7_75t_L g3397 ( 
.A(n_3094),
.Y(n_3397)
);

NAND2xp5_ASAP7_75t_L g3398 ( 
.A(n_3202),
.B(n_2686),
.Y(n_3398)
);

NOR2xp33_ASAP7_75t_L g3399 ( 
.A(n_2939),
.B(n_1895),
.Y(n_3399)
);

AOI22xp5_ASAP7_75t_L g3400 ( 
.A1(n_3262),
.A2(n_2597),
.B1(n_2596),
.B2(n_2798),
.Y(n_3400)
);

INVx1_ASAP7_75t_L g3401 ( 
.A(n_3100),
.Y(n_3401)
);

NAND2xp5_ASAP7_75t_SL g3402 ( 
.A(n_2915),
.B(n_2798),
.Y(n_3402)
);

NAND2xp5_ASAP7_75t_SL g3403 ( 
.A(n_2923),
.B(n_2802),
.Y(n_3403)
);

NAND2xp5_ASAP7_75t_L g3404 ( 
.A(n_3208),
.B(n_2596),
.Y(n_3404)
);

NAND2xp5_ASAP7_75t_L g3405 ( 
.A(n_3268),
.B(n_2583),
.Y(n_3405)
);

NOR2xp33_ASAP7_75t_L g3406 ( 
.A(n_2946),
.B(n_1985),
.Y(n_3406)
);

NAND2xp5_ASAP7_75t_L g3407 ( 
.A(n_3275),
.B(n_2855),
.Y(n_3407)
);

BUFx3_ASAP7_75t_L g3408 ( 
.A(n_3067),
.Y(n_3408)
);

NAND2xp5_ASAP7_75t_L g3409 ( 
.A(n_3089),
.B(n_2857),
.Y(n_3409)
);

NAND2xp5_ASAP7_75t_SL g3410 ( 
.A(n_2951),
.B(n_2802),
.Y(n_3410)
);

NOR2xp33_ASAP7_75t_L g3411 ( 
.A(n_3121),
.B(n_1985),
.Y(n_3411)
);

INVxp67_ASAP7_75t_SL g3412 ( 
.A(n_2935),
.Y(n_3412)
);

INVx2_ASAP7_75t_L g3413 ( 
.A(n_3182),
.Y(n_3413)
);

NAND2xp5_ASAP7_75t_L g3414 ( 
.A(n_3089),
.B(n_2735),
.Y(n_3414)
);

NAND2xp5_ASAP7_75t_L g3415 ( 
.A(n_3093),
.B(n_2735),
.Y(n_3415)
);

INVx1_ASAP7_75t_L g3416 ( 
.A(n_3102),
.Y(n_3416)
);

INVx1_ASAP7_75t_L g3417 ( 
.A(n_3103),
.Y(n_3417)
);

INVx1_ASAP7_75t_L g3418 ( 
.A(n_3104),
.Y(n_3418)
);

NAND2xp5_ASAP7_75t_SL g3419 ( 
.A(n_3206),
.B(n_2826),
.Y(n_3419)
);

AOI22xp33_ASAP7_75t_L g3420 ( 
.A1(n_3033),
.A2(n_2692),
.B1(n_2654),
.B2(n_2655),
.Y(n_3420)
);

INVx5_ASAP7_75t_L g3421 ( 
.A(n_3339),
.Y(n_3421)
);

BUFx12f_ASAP7_75t_L g3422 ( 
.A(n_3097),
.Y(n_3422)
);

AND2x6_ASAP7_75t_SL g3423 ( 
.A(n_3079),
.B(n_2714),
.Y(n_3423)
);

A2O1A1Ixp33_ASAP7_75t_L g3424 ( 
.A1(n_3034),
.A2(n_2635),
.B(n_2816),
.C(n_2800),
.Y(n_3424)
);

NAND2xp5_ASAP7_75t_L g3425 ( 
.A(n_3095),
.B(n_2653),
.Y(n_3425)
);

AND2x4_ASAP7_75t_L g3426 ( 
.A(n_3269),
.B(n_2600),
.Y(n_3426)
);

AOI21xp5_ASAP7_75t_L g3427 ( 
.A1(n_2945),
.A2(n_2635),
.B(n_2723),
.Y(n_3427)
);

INVx2_ASAP7_75t_L g3428 ( 
.A(n_3191),
.Y(n_3428)
);

NOR2x1p5_ASAP7_75t_L g3429 ( 
.A(n_3090),
.B(n_2610),
.Y(n_3429)
);

NOR2xp33_ASAP7_75t_SL g3430 ( 
.A(n_2955),
.B(n_1992),
.Y(n_3430)
);

NAND2xp5_ASAP7_75t_L g3431 ( 
.A(n_3141),
.B(n_2659),
.Y(n_3431)
);

NOR2xp33_ASAP7_75t_L g3432 ( 
.A(n_3134),
.B(n_1992),
.Y(n_3432)
);

INVx1_ASAP7_75t_L g3433 ( 
.A(n_3105),
.Y(n_3433)
);

NOR2xp33_ASAP7_75t_L g3434 ( 
.A(n_3016),
.B(n_1996),
.Y(n_3434)
);

INVx2_ASAP7_75t_L g3435 ( 
.A(n_3198),
.Y(n_3435)
);

NAND2xp5_ASAP7_75t_L g3436 ( 
.A(n_3263),
.B(n_2610),
.Y(n_3436)
);

INVxp67_ASAP7_75t_L g3437 ( 
.A(n_2975),
.Y(n_3437)
);

NOR2xp33_ASAP7_75t_L g3438 ( 
.A(n_3025),
.B(n_1996),
.Y(n_3438)
);

INVx3_ASAP7_75t_L g3439 ( 
.A(n_3063),
.Y(n_3439)
);

AND2x2_ASAP7_75t_SL g3440 ( 
.A(n_2974),
.B(n_2635),
.Y(n_3440)
);

INVx1_ASAP7_75t_L g3441 ( 
.A(n_3107),
.Y(n_3441)
);

INVx3_ASAP7_75t_L g3442 ( 
.A(n_3065),
.Y(n_3442)
);

AND2x4_ASAP7_75t_L g3443 ( 
.A(n_3320),
.B(n_2826),
.Y(n_3443)
);

AO221x1_ASAP7_75t_L g3444 ( 
.A1(n_3039),
.A2(n_2888),
.B1(n_2863),
.B2(n_2680),
.C(n_2699),
.Y(n_3444)
);

INVx2_ASAP7_75t_L g3445 ( 
.A(n_3222),
.Y(n_3445)
);

NOR2xp33_ASAP7_75t_L g3446 ( 
.A(n_3298),
.B(n_3047),
.Y(n_3446)
);

INVx2_ASAP7_75t_L g3447 ( 
.A(n_3246),
.Y(n_3447)
);

INVx2_ASAP7_75t_L g3448 ( 
.A(n_3248),
.Y(n_3448)
);

NAND2xp5_ASAP7_75t_SL g3449 ( 
.A(n_3057),
.B(n_2835),
.Y(n_3449)
);

INVx2_ASAP7_75t_L g3450 ( 
.A(n_3285),
.Y(n_3450)
);

AND2x2_ASAP7_75t_L g3451 ( 
.A(n_3114),
.B(n_2848),
.Y(n_3451)
);

CKINVDCx11_ASAP7_75t_R g3452 ( 
.A(n_2949),
.Y(n_3452)
);

NAND2xp5_ASAP7_75t_L g3453 ( 
.A(n_3263),
.B(n_2848),
.Y(n_3453)
);

NOR2xp33_ASAP7_75t_L g3454 ( 
.A(n_3050),
.B(n_2023),
.Y(n_3454)
);

NAND2xp5_ASAP7_75t_L g3455 ( 
.A(n_3164),
.B(n_2669),
.Y(n_3455)
);

INVx1_ASAP7_75t_L g3456 ( 
.A(n_3108),
.Y(n_3456)
);

NOR2xp67_ASAP7_75t_L g3457 ( 
.A(n_2940),
.B(n_2859),
.Y(n_3457)
);

INVx2_ASAP7_75t_L g3458 ( 
.A(n_3288),
.Y(n_3458)
);

NAND2xp33_ASAP7_75t_L g3459 ( 
.A(n_3061),
.B(n_2499),
.Y(n_3459)
);

INVx2_ASAP7_75t_SL g3460 ( 
.A(n_2921),
.Y(n_3460)
);

AND2x2_ASAP7_75t_L g3461 ( 
.A(n_3122),
.B(n_2835),
.Y(n_3461)
);

INVx3_ASAP7_75t_L g3462 ( 
.A(n_3065),
.Y(n_3462)
);

INVx1_ASAP7_75t_L g3463 ( 
.A(n_3110),
.Y(n_3463)
);

NAND2xp5_ASAP7_75t_L g3464 ( 
.A(n_3150),
.B(n_2684),
.Y(n_3464)
);

NOR2xp33_ASAP7_75t_L g3465 ( 
.A(n_3059),
.B(n_2023),
.Y(n_3465)
);

AND2x2_ASAP7_75t_L g3466 ( 
.A(n_3169),
.B(n_2858),
.Y(n_3466)
);

NAND2xp5_ASAP7_75t_L g3467 ( 
.A(n_3174),
.B(n_3080),
.Y(n_3467)
);

NAND2xp5_ASAP7_75t_SL g3468 ( 
.A(n_2952),
.B(n_2786),
.Y(n_3468)
);

NOR2xp33_ASAP7_75t_L g3469 ( 
.A(n_2981),
.B(n_2996),
.Y(n_3469)
);

OR2x6_ASAP7_75t_L g3470 ( 
.A(n_3064),
.B(n_2714),
.Y(n_3470)
);

NOR2xp33_ASAP7_75t_L g3471 ( 
.A(n_2983),
.B(n_2034),
.Y(n_3471)
);

INVx2_ASAP7_75t_L g3472 ( 
.A(n_3289),
.Y(n_3472)
);

INVx2_ASAP7_75t_L g3473 ( 
.A(n_3290),
.Y(n_3473)
);

NAND2xp5_ASAP7_75t_L g3474 ( 
.A(n_3034),
.B(n_2687),
.Y(n_3474)
);

INVx1_ASAP7_75t_L g3475 ( 
.A(n_3111),
.Y(n_3475)
);

AOI22xp33_ASAP7_75t_L g3476 ( 
.A1(n_3033),
.A2(n_2694),
.B1(n_2710),
.B2(n_2900),
.Y(n_3476)
);

INVx2_ASAP7_75t_L g3477 ( 
.A(n_3300),
.Y(n_3477)
);

NAND2xp5_ASAP7_75t_L g3478 ( 
.A(n_3130),
.B(n_2874),
.Y(n_3478)
);

INVx1_ASAP7_75t_L g3479 ( 
.A(n_3112),
.Y(n_3479)
);

INVx8_ASAP7_75t_L g3480 ( 
.A(n_3064),
.Y(n_3480)
);

INVx1_ASAP7_75t_L g3481 ( 
.A(n_3116),
.Y(n_3481)
);

NAND2xp5_ASAP7_75t_L g3482 ( 
.A(n_3130),
.B(n_2876),
.Y(n_3482)
);

AND2x2_ASAP7_75t_L g3483 ( 
.A(n_3283),
.B(n_2877),
.Y(n_3483)
);

NAND2xp5_ASAP7_75t_L g3484 ( 
.A(n_3225),
.B(n_2686),
.Y(n_3484)
);

A2O1A1Ixp33_ASAP7_75t_L g3485 ( 
.A1(n_3216),
.A2(n_2821),
.B(n_2890),
.C(n_2889),
.Y(n_3485)
);

AOI22xp5_ASAP7_75t_L g3486 ( 
.A1(n_3017),
.A2(n_2884),
.B1(n_2896),
.B2(n_2892),
.Y(n_3486)
);

INVx1_ASAP7_75t_L g3487 ( 
.A(n_3117),
.Y(n_3487)
);

NAND2xp5_ASAP7_75t_L g3488 ( 
.A(n_3225),
.B(n_2688),
.Y(n_3488)
);

NAND2xp5_ASAP7_75t_L g3489 ( 
.A(n_3216),
.B(n_2688),
.Y(n_3489)
);

INVx3_ASAP7_75t_L g3490 ( 
.A(n_3065),
.Y(n_3490)
);

INVx2_ASAP7_75t_L g3491 ( 
.A(n_3303),
.Y(n_3491)
);

INVx2_ASAP7_75t_L g3492 ( 
.A(n_3319),
.Y(n_3492)
);

INVx3_ASAP7_75t_L g3493 ( 
.A(n_3186),
.Y(n_3493)
);

AND2x2_ASAP7_75t_L g3494 ( 
.A(n_3331),
.B(n_2905),
.Y(n_3494)
);

AO221x1_ASAP7_75t_L g3495 ( 
.A1(n_3186),
.A2(n_2680),
.B1(n_2699),
.B2(n_2679),
.C(n_2678),
.Y(n_3495)
);

NAND2xp5_ASAP7_75t_SL g3496 ( 
.A(n_3024),
.B(n_2786),
.Y(n_3496)
);

NAND2xp5_ASAP7_75t_SL g3497 ( 
.A(n_3024),
.B(n_2786),
.Y(n_3497)
);

NOR2xp67_ASAP7_75t_L g3498 ( 
.A(n_2934),
.B(n_2890),
.Y(n_3498)
);

NAND2xp5_ASAP7_75t_L g3499 ( 
.A(n_3045),
.B(n_2909),
.Y(n_3499)
);

INVx2_ASAP7_75t_SL g3500 ( 
.A(n_2921),
.Y(n_3500)
);

NAND2xp5_ASAP7_75t_L g3501 ( 
.A(n_3045),
.B(n_2806),
.Y(n_3501)
);

HB1xp67_ASAP7_75t_L g3502 ( 
.A(n_3001),
.Y(n_3502)
);

NAND2xp33_ASAP7_75t_L g3503 ( 
.A(n_3061),
.B(n_2499),
.Y(n_3503)
);

NAND2xp5_ASAP7_75t_L g3504 ( 
.A(n_2995),
.B(n_2806),
.Y(n_3504)
);

NOR2xp67_ASAP7_75t_L g3505 ( 
.A(n_3139),
.B(n_2850),
.Y(n_3505)
);

NAND2xp5_ASAP7_75t_L g3506 ( 
.A(n_2995),
.B(n_2819),
.Y(n_3506)
);

NAND2xp5_ASAP7_75t_L g3507 ( 
.A(n_3060),
.B(n_2819),
.Y(n_3507)
);

NAND2xp5_ASAP7_75t_L g3508 ( 
.A(n_3060),
.B(n_2824),
.Y(n_3508)
);

NAND2xp5_ASAP7_75t_L g3509 ( 
.A(n_3068),
.B(n_2824),
.Y(n_3509)
);

NOR2xp33_ASAP7_75t_L g3510 ( 
.A(n_2986),
.B(n_2034),
.Y(n_3510)
);

INVx1_ASAP7_75t_L g3511 ( 
.A(n_3119),
.Y(n_3511)
);

NAND2xp5_ASAP7_75t_L g3512 ( 
.A(n_3068),
.B(n_2827),
.Y(n_3512)
);

NAND2xp33_ASAP7_75t_L g3513 ( 
.A(n_3061),
.B(n_2499),
.Y(n_3513)
);

NAND2xp5_ASAP7_75t_L g3514 ( 
.A(n_3106),
.B(n_2827),
.Y(n_3514)
);

INVx2_ASAP7_75t_L g3515 ( 
.A(n_3322),
.Y(n_3515)
);

NOR2xp33_ASAP7_75t_L g3516 ( 
.A(n_3316),
.B(n_2850),
.Y(n_3516)
);

INVx3_ASAP7_75t_L g3517 ( 
.A(n_3186),
.Y(n_3517)
);

AOI22xp5_ASAP7_75t_L g3518 ( 
.A1(n_3070),
.A2(n_2906),
.B1(n_2910),
.B2(n_2519),
.Y(n_3518)
);

INVx1_ASAP7_75t_L g3519 ( 
.A(n_3127),
.Y(n_3519)
);

NAND2xp5_ASAP7_75t_SL g3520 ( 
.A(n_3123),
.B(n_2829),
.Y(n_3520)
);

NAND2xp5_ASAP7_75t_SL g3521 ( 
.A(n_3280),
.B(n_2829),
.Y(n_3521)
);

NOR2xp67_ASAP7_75t_L g3522 ( 
.A(n_3002),
.B(n_2893),
.Y(n_3522)
);

INVx2_ASAP7_75t_L g3523 ( 
.A(n_3338),
.Y(n_3523)
);

OR2x6_ASAP7_75t_L g3524 ( 
.A(n_3078),
.B(n_2578),
.Y(n_3524)
);

NOR2xp33_ASAP7_75t_L g3525 ( 
.A(n_3146),
.B(n_3153),
.Y(n_3525)
);

NOR2xp67_ASAP7_75t_SL g3526 ( 
.A(n_3251),
.B(n_2723),
.Y(n_3526)
);

NAND2xp5_ASAP7_75t_L g3527 ( 
.A(n_3106),
.B(n_2833),
.Y(n_3527)
);

NOR2xp33_ASAP7_75t_L g3528 ( 
.A(n_3183),
.B(n_2832),
.Y(n_3528)
);

NOR2xp33_ASAP7_75t_L g3529 ( 
.A(n_3185),
.B(n_2832),
.Y(n_3529)
);

NOR3xp33_ASAP7_75t_L g3530 ( 
.A(n_3203),
.B(n_1142),
.C(n_2056),
.Y(n_3530)
);

INVx1_ASAP7_75t_L g3531 ( 
.A(n_3128),
.Y(n_3531)
);

BUFx3_ASAP7_75t_L g3532 ( 
.A(n_2982),
.Y(n_3532)
);

NOR2xp33_ASAP7_75t_SL g3533 ( 
.A(n_2999),
.B(n_2463),
.Y(n_3533)
);

INVx1_ASAP7_75t_L g3534 ( 
.A(n_3131),
.Y(n_3534)
);

NAND2xp5_ASAP7_75t_L g3535 ( 
.A(n_3267),
.B(n_2768),
.Y(n_3535)
);

NAND2xp5_ASAP7_75t_L g3536 ( 
.A(n_3267),
.B(n_2847),
.Y(n_3536)
);

NAND2xp5_ASAP7_75t_L g3537 ( 
.A(n_3099),
.B(n_3163),
.Y(n_3537)
);

INVx2_ASAP7_75t_L g3538 ( 
.A(n_3347),
.Y(n_3538)
);

NAND2xp5_ASAP7_75t_SL g3539 ( 
.A(n_3166),
.B(n_2829),
.Y(n_3539)
);

NAND2xp5_ASAP7_75t_L g3540 ( 
.A(n_3099),
.B(n_2833),
.Y(n_3540)
);

NAND2xp5_ASAP7_75t_SL g3541 ( 
.A(n_2992),
.B(n_2723),
.Y(n_3541)
);

NAND2xp5_ASAP7_75t_SL g3542 ( 
.A(n_3003),
.B(n_2723),
.Y(n_3542)
);

NOR2xp33_ASAP7_75t_L g3543 ( 
.A(n_3242),
.B(n_3278),
.Y(n_3543)
);

NAND2xp33_ASAP7_75t_L g3544 ( 
.A(n_3061),
.B(n_2499),
.Y(n_3544)
);

INVx4_ASAP7_75t_L g3545 ( 
.A(n_3251),
.Y(n_3545)
);

BUFx6f_ASAP7_75t_SL g3546 ( 
.A(n_2994),
.Y(n_3546)
);

NOR2xp33_ASAP7_75t_L g3547 ( 
.A(n_3313),
.B(n_3326),
.Y(n_3547)
);

INVx2_ASAP7_75t_SL g3548 ( 
.A(n_2971),
.Y(n_3548)
);

INVx1_ASAP7_75t_L g3549 ( 
.A(n_3181),
.Y(n_3549)
);

NAND2xp5_ASAP7_75t_L g3550 ( 
.A(n_3163),
.B(n_2837),
.Y(n_3550)
);

INVx1_ASAP7_75t_L g3551 ( 
.A(n_2917),
.Y(n_3551)
);

NAND2xp5_ASAP7_75t_SL g3552 ( 
.A(n_3313),
.B(n_2723),
.Y(n_3552)
);

INVx2_ASAP7_75t_L g3553 ( 
.A(n_2929),
.Y(n_3553)
);

INVx2_ASAP7_75t_SL g3554 ( 
.A(n_3009),
.Y(n_3554)
);

INVx2_ASAP7_75t_L g3555 ( 
.A(n_2963),
.Y(n_3555)
);

NOR2xp33_ASAP7_75t_L g3556 ( 
.A(n_3326),
.B(n_3001),
.Y(n_3556)
);

INVx2_ASAP7_75t_L g3557 ( 
.A(n_2977),
.Y(n_3557)
);

AOI22xp5_ASAP7_75t_L g3558 ( 
.A1(n_3178),
.A2(n_2832),
.B1(n_2216),
.B2(n_2217),
.Y(n_3558)
);

NAND2xp5_ASAP7_75t_L g3559 ( 
.A(n_2945),
.B(n_2837),
.Y(n_3559)
);

NAND2xp5_ASAP7_75t_L g3560 ( 
.A(n_3321),
.B(n_3309),
.Y(n_3560)
);

INVxp67_ASAP7_75t_L g3561 ( 
.A(n_3161),
.Y(n_3561)
);

NAND2xp5_ASAP7_75t_L g3562 ( 
.A(n_3321),
.B(n_2841),
.Y(n_3562)
);

NAND2xp5_ASAP7_75t_L g3563 ( 
.A(n_3309),
.B(n_2841),
.Y(n_3563)
);

INVx2_ASAP7_75t_SL g3564 ( 
.A(n_3009),
.Y(n_3564)
);

INVx2_ASAP7_75t_L g3565 ( 
.A(n_2988),
.Y(n_3565)
);

INVx2_ASAP7_75t_SL g3566 ( 
.A(n_3179),
.Y(n_3566)
);

INVxp67_ASAP7_75t_L g3567 ( 
.A(n_3161),
.Y(n_3567)
);

CKINVDCx14_ASAP7_75t_R g3568 ( 
.A(n_3156),
.Y(n_3568)
);

NAND2xp5_ASAP7_75t_SL g3569 ( 
.A(n_3092),
.B(n_2870),
.Y(n_3569)
);

INVx1_ASAP7_75t_L g3570 ( 
.A(n_2918),
.Y(n_3570)
);

NAND2xp5_ASAP7_75t_L g3571 ( 
.A(n_3324),
.B(n_2846),
.Y(n_3571)
);

NAND2xp5_ASAP7_75t_L g3572 ( 
.A(n_3324),
.B(n_2846),
.Y(n_3572)
);

NAND2xp5_ASAP7_75t_L g3573 ( 
.A(n_3184),
.B(n_2864),
.Y(n_3573)
);

AND2x4_ASAP7_75t_L g3574 ( 
.A(n_2953),
.B(n_2864),
.Y(n_3574)
);

NOR2xp67_ASAP7_75t_L g3575 ( 
.A(n_3040),
.B(n_3096),
.Y(n_3575)
);

NAND2xp5_ASAP7_75t_L g3576 ( 
.A(n_3187),
.B(n_2866),
.Y(n_3576)
);

INVx2_ASAP7_75t_L g3577 ( 
.A(n_3011),
.Y(n_3577)
);

NAND2xp5_ASAP7_75t_L g3578 ( 
.A(n_3188),
.B(n_2866),
.Y(n_3578)
);

NAND2xp5_ASAP7_75t_L g3579 ( 
.A(n_3189),
.B(n_2868),
.Y(n_3579)
);

NOR3xp33_ASAP7_75t_L g3580 ( 
.A(n_3329),
.B(n_2056),
.C(n_908),
.Y(n_3580)
);

INVx1_ASAP7_75t_L g3581 ( 
.A(n_2919),
.Y(n_3581)
);

AOI22xp5_ASAP7_75t_L g3582 ( 
.A1(n_3192),
.A2(n_2223),
.B1(n_2228),
.B2(n_2211),
.Y(n_3582)
);

NOR2xp67_ASAP7_75t_L g3583 ( 
.A(n_3132),
.B(n_2899),
.Y(n_3583)
);

NAND2xp5_ASAP7_75t_SL g3584 ( 
.A(n_3155),
.B(n_3201),
.Y(n_3584)
);

NAND2xp5_ASAP7_75t_L g3585 ( 
.A(n_3194),
.B(n_2868),
.Y(n_3585)
);

NAND2xp5_ASAP7_75t_L g3586 ( 
.A(n_3195),
.B(n_2871),
.Y(n_3586)
);

NAND2xp5_ASAP7_75t_SL g3587 ( 
.A(n_3155),
.B(n_2870),
.Y(n_3587)
);

NAND2xp5_ASAP7_75t_L g3588 ( 
.A(n_3196),
.B(n_2871),
.Y(n_3588)
);

NAND2xp5_ASAP7_75t_SL g3589 ( 
.A(n_3234),
.B(n_2870),
.Y(n_3589)
);

AO22x1_ASAP7_75t_L g3590 ( 
.A1(n_3299),
.A2(n_2446),
.B1(n_2020),
.B2(n_2280),
.Y(n_3590)
);

INVx2_ASAP7_75t_L g3591 ( 
.A(n_3048),
.Y(n_3591)
);

OAI22xp33_ASAP7_75t_L g3592 ( 
.A1(n_3010),
.A2(n_2870),
.B1(n_2622),
.B2(n_2639),
.Y(n_3592)
);

NAND2xp5_ASAP7_75t_L g3593 ( 
.A(n_3197),
.B(n_2879),
.Y(n_3593)
);

INVx2_ASAP7_75t_L g3594 ( 
.A(n_3049),
.Y(n_3594)
);

NOR2xp33_ASAP7_75t_L g3595 ( 
.A(n_3125),
.B(n_2446),
.Y(n_3595)
);

NAND2xp5_ASAP7_75t_L g3596 ( 
.A(n_3199),
.B(n_2879),
.Y(n_3596)
);

OAI21xp5_ASAP7_75t_L g3597 ( 
.A1(n_3294),
.A2(n_3000),
.B(n_3193),
.Y(n_3597)
);

NAND2xp5_ASAP7_75t_L g3598 ( 
.A(n_3317),
.B(n_3282),
.Y(n_3598)
);

BUFx2_ASAP7_75t_L g3599 ( 
.A(n_2957),
.Y(n_3599)
);

AOI22xp33_ASAP7_75t_SL g3600 ( 
.A1(n_3088),
.A2(n_2828),
.B1(n_2622),
.B2(n_2639),
.Y(n_3600)
);

INVx2_ASAP7_75t_SL g3601 ( 
.A(n_3179),
.Y(n_3601)
);

INVx2_ASAP7_75t_L g3602 ( 
.A(n_3051),
.Y(n_3602)
);

OAI22xp5_ASAP7_75t_L g3603 ( 
.A1(n_3294),
.A2(n_2865),
.B1(n_2870),
.B2(n_2622),
.Y(n_3603)
);

INVx2_ASAP7_75t_L g3604 ( 
.A(n_3052),
.Y(n_3604)
);

NOR2xp33_ASAP7_75t_L g3605 ( 
.A(n_3136),
.B(n_2828),
.Y(n_3605)
);

NAND2xp5_ASAP7_75t_L g3606 ( 
.A(n_3317),
.B(n_2880),
.Y(n_3606)
);

A2O1A1Ixp33_ASAP7_75t_L g3607 ( 
.A1(n_3088),
.A2(n_3233),
.B(n_3302),
.C(n_3200),
.Y(n_3607)
);

NAND2xp5_ASAP7_75t_L g3608 ( 
.A(n_3205),
.B(n_2880),
.Y(n_3608)
);

NAND2xp5_ASAP7_75t_L g3609 ( 
.A(n_2920),
.B(n_2882),
.Y(n_3609)
);

INVxp67_ASAP7_75t_SL g3610 ( 
.A(n_2935),
.Y(n_3610)
);

NAND2xp5_ASAP7_75t_L g3611 ( 
.A(n_2922),
.B(n_2882),
.Y(n_3611)
);

OAI22xp5_ASAP7_75t_L g3612 ( 
.A1(n_3346),
.A2(n_3084),
.B1(n_3233),
.B2(n_3210),
.Y(n_3612)
);

NAND2xp5_ASAP7_75t_SL g3613 ( 
.A(n_3251),
.B(n_2627),
.Y(n_3613)
);

INVx2_ASAP7_75t_L g3614 ( 
.A(n_3066),
.Y(n_3614)
);

INVx2_ASAP7_75t_L g3615 ( 
.A(n_3218),
.Y(n_3615)
);

O2A1O1Ixp33_ASAP7_75t_L g3616 ( 
.A1(n_2966),
.A2(n_2234),
.B(n_2238),
.C(n_2231),
.Y(n_3616)
);

INVx1_ASAP7_75t_L g3617 ( 
.A(n_2924),
.Y(n_3617)
);

NAND2xp33_ASAP7_75t_SL g3618 ( 
.A(n_3053),
.B(n_2828),
.Y(n_3618)
);

INVx1_ASAP7_75t_L g3619 ( 
.A(n_2925),
.Y(n_3619)
);

NOR2xp33_ASAP7_75t_L g3620 ( 
.A(n_3152),
.B(n_2678),
.Y(n_3620)
);

NAND2xp5_ASAP7_75t_L g3621 ( 
.A(n_2926),
.B(n_2886),
.Y(n_3621)
);

OAI221xp5_ASAP7_75t_L g3622 ( 
.A1(n_3172),
.A2(n_1011),
.B1(n_1041),
.B2(n_986),
.C(n_893),
.Y(n_3622)
);

AND2x2_ASAP7_75t_L g3623 ( 
.A(n_3344),
.B(n_3135),
.Y(n_3623)
);

NAND2xp5_ASAP7_75t_SL g3624 ( 
.A(n_3327),
.B(n_2627),
.Y(n_3624)
);

NOR2xp33_ASAP7_75t_L g3625 ( 
.A(n_3209),
.B(n_2678),
.Y(n_3625)
);

NAND2xp5_ASAP7_75t_SL g3626 ( 
.A(n_3327),
.B(n_2627),
.Y(n_3626)
);

AND2x2_ASAP7_75t_L g3627 ( 
.A(n_3137),
.B(n_2004),
.Y(n_3627)
);

INVx2_ASAP7_75t_L g3628 ( 
.A(n_3219),
.Y(n_3628)
);

INVx1_ASAP7_75t_L g3629 ( 
.A(n_2928),
.Y(n_3629)
);

CKINVDCx11_ASAP7_75t_R g3630 ( 
.A(n_3113),
.Y(n_3630)
);

INVx2_ASAP7_75t_SL g3631 ( 
.A(n_3140),
.Y(n_3631)
);

AND2x4_ASAP7_75t_L g3632 ( 
.A(n_2953),
.B(n_3029),
.Y(n_3632)
);

INVx1_ASAP7_75t_L g3633 ( 
.A(n_2931),
.Y(n_3633)
);

INVx2_ASAP7_75t_L g3634 ( 
.A(n_3220),
.Y(n_3634)
);

AND2x4_ASAP7_75t_L g3635 ( 
.A(n_3029),
.B(n_2886),
.Y(n_3635)
);

INVx8_ASAP7_75t_L g3636 ( 
.A(n_3078),
.Y(n_3636)
);

NAND2xp5_ASAP7_75t_L g3637 ( 
.A(n_2932),
.B(n_2496),
.Y(n_3637)
);

OR2x2_ASAP7_75t_L g3638 ( 
.A(n_3214),
.B(n_2898),
.Y(n_3638)
);

INVx1_ASAP7_75t_L g3639 ( 
.A(n_2936),
.Y(n_3639)
);

INVx1_ASAP7_75t_L g3640 ( 
.A(n_2937),
.Y(n_3640)
);

NAND2xp5_ASAP7_75t_L g3641 ( 
.A(n_2938),
.B(n_2941),
.Y(n_3641)
);

NOR2xp33_ASAP7_75t_L g3642 ( 
.A(n_3250),
.B(n_2679),
.Y(n_3642)
);

INVxp67_ASAP7_75t_SL g3643 ( 
.A(n_3022),
.Y(n_3643)
);

AOI22xp5_ASAP7_75t_L g3644 ( 
.A1(n_2933),
.A2(n_2242),
.B1(n_2246),
.B2(n_2239),
.Y(n_3644)
);

BUFx2_ASAP7_75t_L g3645 ( 
.A(n_3078),
.Y(n_3645)
);

NOR2xp33_ASAP7_75t_L g3646 ( 
.A(n_3277),
.B(n_2679),
.Y(n_3646)
);

NAND2xp5_ASAP7_75t_L g3647 ( 
.A(n_2942),
.B(n_2496),
.Y(n_3647)
);

NOR2xp33_ASAP7_75t_L g3648 ( 
.A(n_3314),
.B(n_2680),
.Y(n_3648)
);

NAND2xp5_ASAP7_75t_SL g3649 ( 
.A(n_3327),
.B(n_2668),
.Y(n_3649)
);

OR2x6_ASAP7_75t_L g3650 ( 
.A(n_2994),
.B(n_2582),
.Y(n_3650)
);

INVx2_ASAP7_75t_L g3651 ( 
.A(n_3223),
.Y(n_3651)
);

NAND2xp5_ASAP7_75t_L g3652 ( 
.A(n_3207),
.B(n_2699),
.Y(n_3652)
);

INVx2_ASAP7_75t_L g3653 ( 
.A(n_3224),
.Y(n_3653)
);

INVx2_ASAP7_75t_L g3654 ( 
.A(n_3226),
.Y(n_3654)
);

NAND2xp5_ASAP7_75t_SL g3655 ( 
.A(n_3334),
.B(n_2668),
.Y(n_3655)
);

NAND2xp5_ASAP7_75t_L g3656 ( 
.A(n_3211),
.B(n_2705),
.Y(n_3656)
);

NAND2xp5_ASAP7_75t_L g3657 ( 
.A(n_3212),
.B(n_3213),
.Y(n_3657)
);

NOR2xp33_ASAP7_75t_L g3658 ( 
.A(n_3335),
.B(n_2705),
.Y(n_3658)
);

NAND2xp5_ASAP7_75t_L g3659 ( 
.A(n_3215),
.B(n_2705),
.Y(n_3659)
);

INVx2_ASAP7_75t_L g3660 ( 
.A(n_3228),
.Y(n_3660)
);

OAI21xp5_ASAP7_75t_L g3661 ( 
.A1(n_3000),
.A2(n_2878),
.B(n_2541),
.Y(n_3661)
);

INVx1_ASAP7_75t_L g3662 ( 
.A(n_2948),
.Y(n_3662)
);

INVx2_ASAP7_75t_SL g3663 ( 
.A(n_3144),
.Y(n_3663)
);

NAND2xp5_ASAP7_75t_L g3664 ( 
.A(n_3217),
.B(n_2745),
.Y(n_3664)
);

NAND2xp5_ASAP7_75t_L g3665 ( 
.A(n_2950),
.B(n_2496),
.Y(n_3665)
);

INVx2_ASAP7_75t_L g3666 ( 
.A(n_3229),
.Y(n_3666)
);

OR2x6_ASAP7_75t_L g3667 ( 
.A(n_2994),
.B(n_2582),
.Y(n_3667)
);

NAND2xp5_ASAP7_75t_SL g3668 ( 
.A(n_3334),
.B(n_2668),
.Y(n_3668)
);

INVx1_ASAP7_75t_L g3669 ( 
.A(n_2959),
.Y(n_3669)
);

NOR2xp33_ASAP7_75t_L g3670 ( 
.A(n_3257),
.B(n_2745),
.Y(n_3670)
);

INVx2_ASAP7_75t_L g3671 ( 
.A(n_3231),
.Y(n_3671)
);

NOR2xp33_ASAP7_75t_L g3672 ( 
.A(n_3333),
.B(n_2745),
.Y(n_3672)
);

OAI22xp33_ASAP7_75t_L g3673 ( 
.A1(n_3145),
.A2(n_2622),
.B1(n_2639),
.B2(n_2582),
.Y(n_3673)
);

INVx1_ASAP7_75t_L g3674 ( 
.A(n_2960),
.Y(n_3674)
);

AOI21xp5_ASAP7_75t_L g3675 ( 
.A1(n_3302),
.A2(n_2639),
.B(n_2582),
.Y(n_3675)
);

NAND3xp33_ASAP7_75t_SL g3676 ( 
.A(n_3012),
.B(n_1165),
.C(n_1154),
.Y(n_3676)
);

AND2x2_ASAP7_75t_L g3677 ( 
.A(n_3147),
.B(n_2007),
.Y(n_3677)
);

NAND2xp5_ASAP7_75t_SL g3678 ( 
.A(n_3334),
.B(n_2668),
.Y(n_3678)
);

INVxp67_ASAP7_75t_SL g3679 ( 
.A(n_3022),
.Y(n_3679)
);

AND2x2_ASAP7_75t_L g3680 ( 
.A(n_3148),
.B(n_2007),
.Y(n_3680)
);

NAND2xp5_ASAP7_75t_SL g3681 ( 
.A(n_3143),
.B(n_2701),
.Y(n_3681)
);

INVx1_ASAP7_75t_L g3682 ( 
.A(n_2965),
.Y(n_3682)
);

NAND3xp33_ASAP7_75t_L g3683 ( 
.A(n_3204),
.B(n_3151),
.C(n_3149),
.Y(n_3683)
);

AOI21xp5_ASAP7_75t_L g3684 ( 
.A1(n_3279),
.A2(n_2758),
.B(n_2612),
.Y(n_3684)
);

NAND2xp5_ASAP7_75t_L g3685 ( 
.A(n_3085),
.B(n_2764),
.Y(n_3685)
);

NOR2xp33_ASAP7_75t_L g3686 ( 
.A(n_2947),
.B(n_2764),
.Y(n_3686)
);

NAND2xp5_ASAP7_75t_L g3687 ( 
.A(n_3101),
.B(n_3238),
.Y(n_3687)
);

INVx2_ASAP7_75t_SL g3688 ( 
.A(n_3154),
.Y(n_3688)
);

INVx1_ASAP7_75t_L g3689 ( 
.A(n_2969),
.Y(n_3689)
);

NAND2xp5_ASAP7_75t_SL g3690 ( 
.A(n_3157),
.B(n_2701),
.Y(n_3690)
);

INVx1_ASAP7_75t_L g3691 ( 
.A(n_2970),
.Y(n_3691)
);

INVx2_ASAP7_75t_L g3692 ( 
.A(n_3232),
.Y(n_3692)
);

NAND2xp5_ASAP7_75t_SL g3693 ( 
.A(n_3158),
.B(n_2701),
.Y(n_3693)
);

NAND2xp5_ASAP7_75t_L g3694 ( 
.A(n_3101),
.B(n_2764),
.Y(n_3694)
);

INVx2_ASAP7_75t_L g3695 ( 
.A(n_3235),
.Y(n_3695)
);

NOR2xp33_ASAP7_75t_L g3696 ( 
.A(n_2958),
.B(n_2769),
.Y(n_3696)
);

INVx4_ASAP7_75t_L g3697 ( 
.A(n_3339),
.Y(n_3697)
);

NAND2xp5_ASAP7_75t_L g3698 ( 
.A(n_3238),
.B(n_3332),
.Y(n_3698)
);

INVxp67_ASAP7_75t_L g3699 ( 
.A(n_3159),
.Y(n_3699)
);

INVx3_ASAP7_75t_L g3700 ( 
.A(n_3004),
.Y(n_3700)
);

NAND2xp5_ASAP7_75t_SL g3701 ( 
.A(n_3162),
.B(n_2701),
.Y(n_3701)
);

NOR2xp33_ASAP7_75t_L g3702 ( 
.A(n_3168),
.B(n_2769),
.Y(n_3702)
);

INVx1_ASAP7_75t_L g3703 ( 
.A(n_2972),
.Y(n_3703)
);

AND2x2_ASAP7_75t_L g3704 ( 
.A(n_3170),
.B(n_2058),
.Y(n_3704)
);

INVxp67_ASAP7_75t_SL g3705 ( 
.A(n_3332),
.Y(n_3705)
);

NAND2xp5_ASAP7_75t_L g3706 ( 
.A(n_3171),
.B(n_2769),
.Y(n_3706)
);

A2O1A1Ixp33_ASAP7_75t_L g3707 ( 
.A1(n_3193),
.A2(n_2885),
.B(n_2891),
.C(n_2541),
.Y(n_3707)
);

AND2x2_ASAP7_75t_L g3708 ( 
.A(n_3173),
.B(n_2058),
.Y(n_3708)
);

HB1xp67_ASAP7_75t_L g3709 ( 
.A(n_3176),
.Y(n_3709)
);

BUFx6f_ASAP7_75t_L g3710 ( 
.A(n_3075),
.Y(n_3710)
);

NAND2xp5_ASAP7_75t_L g3711 ( 
.A(n_3177),
.B(n_2807),
.Y(n_3711)
);

INVxp67_ASAP7_75t_L g3712 ( 
.A(n_3180),
.Y(n_3712)
);

NAND2xp5_ASAP7_75t_SL g3713 ( 
.A(n_3075),
.B(n_2794),
.Y(n_3713)
);

AND2x2_ASAP7_75t_L g3714 ( 
.A(n_3109),
.B(n_3167),
.Y(n_3714)
);

NAND2xp5_ASAP7_75t_L g3715 ( 
.A(n_2973),
.B(n_2807),
.Y(n_3715)
);

NAND2xp5_ASAP7_75t_L g3716 ( 
.A(n_2978),
.B(n_2513),
.Y(n_3716)
);

AND2x4_ASAP7_75t_L g3717 ( 
.A(n_3109),
.B(n_2898),
.Y(n_3717)
);

HB1xp67_ASAP7_75t_L g3718 ( 
.A(n_3167),
.Y(n_3718)
);

INVx1_ASAP7_75t_L g3719 ( 
.A(n_2979),
.Y(n_3719)
);

INVxp67_ASAP7_75t_L g3720 ( 
.A(n_2916),
.Y(n_3720)
);

BUFx6f_ASAP7_75t_L g3721 ( 
.A(n_3175),
.Y(n_3721)
);

NAND2xp5_ASAP7_75t_L g3722 ( 
.A(n_2980),
.B(n_2984),
.Y(n_3722)
);

INVx1_ASAP7_75t_L g3723 ( 
.A(n_2985),
.Y(n_3723)
);

NAND2xp5_ASAP7_75t_L g3724 ( 
.A(n_2987),
.B(n_2513),
.Y(n_3724)
);

INVx2_ASAP7_75t_L g3725 ( 
.A(n_3236),
.Y(n_3725)
);

INVx3_ASAP7_75t_L g3726 ( 
.A(n_3004),
.Y(n_3726)
);

INVx2_ASAP7_75t_SL g3727 ( 
.A(n_3175),
.Y(n_3727)
);

INVx2_ASAP7_75t_SL g3728 ( 
.A(n_3227),
.Y(n_3728)
);

AND2x2_ASAP7_75t_L g3729 ( 
.A(n_3227),
.B(n_3311),
.Y(n_3729)
);

NAND2xp5_ASAP7_75t_L g3730 ( 
.A(n_2990),
.B(n_2513),
.Y(n_3730)
);

AND2x6_ASAP7_75t_L g3731 ( 
.A(n_3279),
.B(n_2911),
.Y(n_3731)
);

NOR2xp33_ASAP7_75t_L g3732 ( 
.A(n_3253),
.B(n_2807),
.Y(n_3732)
);

NAND2xp5_ASAP7_75t_L g3733 ( 
.A(n_2991),
.B(n_2515),
.Y(n_3733)
);

NAND2xp5_ASAP7_75t_SL g3734 ( 
.A(n_3311),
.B(n_2794),
.Y(n_3734)
);

NAND2xp5_ASAP7_75t_L g3735 ( 
.A(n_2993),
.B(n_2515),
.Y(n_3735)
);

OAI22xp5_ASAP7_75t_L g3736 ( 
.A1(n_2998),
.A2(n_2894),
.B1(n_1094),
.B2(n_1098),
.Y(n_3736)
);

NAND2xp5_ASAP7_75t_SL g3737 ( 
.A(n_3061),
.B(n_2794),
.Y(n_3737)
);

AOI22xp5_ASAP7_75t_SL g3738 ( 
.A1(n_3124),
.A2(n_1189),
.B1(n_1177),
.B2(n_880),
.Y(n_3738)
);

AOI22xp33_ASAP7_75t_L g3739 ( 
.A1(n_3120),
.A2(n_2666),
.B1(n_2247),
.B2(n_2259),
.Y(n_3739)
);

NAND2xp5_ASAP7_75t_SL g3740 ( 
.A(n_3138),
.B(n_2794),
.Y(n_3740)
);

CKINVDCx5p33_ASAP7_75t_R g3741 ( 
.A(n_2930),
.Y(n_3741)
);

NOR2xp33_ASAP7_75t_L g3742 ( 
.A(n_3304),
.B(n_2814),
.Y(n_3742)
);

INVx1_ASAP7_75t_L g3743 ( 
.A(n_3005),
.Y(n_3743)
);

NAND2xp5_ASAP7_75t_L g3744 ( 
.A(n_3007),
.B(n_3008),
.Y(n_3744)
);

NAND2xp5_ASAP7_75t_SL g3745 ( 
.A(n_3138),
.B(n_2796),
.Y(n_3745)
);

AOI22xp33_ASAP7_75t_L g3746 ( 
.A1(n_3120),
.A2(n_2666),
.B1(n_2250),
.B2(n_2270),
.Y(n_3746)
);

INVx2_ASAP7_75t_L g3747 ( 
.A(n_3237),
.Y(n_3747)
);

NAND3xp33_ASAP7_75t_L g3748 ( 
.A(n_3255),
.B(n_2020),
.C(n_2118),
.Y(n_3748)
);

NOR2xp33_ASAP7_75t_L g3749 ( 
.A(n_2927),
.B(n_3249),
.Y(n_3749)
);

INVxp67_ASAP7_75t_L g3750 ( 
.A(n_3021),
.Y(n_3750)
);

INVx1_ASAP7_75t_L g3751 ( 
.A(n_3014),
.Y(n_3751)
);

AOI22xp5_ASAP7_75t_L g3752 ( 
.A1(n_3394),
.A2(n_3098),
.B1(n_2943),
.B2(n_3230),
.Y(n_3752)
);

O2A1O1Ixp33_ASAP7_75t_L g3753 ( 
.A1(n_3370),
.A2(n_2260),
.B(n_1528),
.C(n_1632),
.Y(n_3753)
);

O2A1O1Ixp33_ASAP7_75t_SL g3754 ( 
.A1(n_3485),
.A2(n_3264),
.B(n_3249),
.C(n_3015),
.Y(n_3754)
);

AND2x2_ASAP7_75t_L g3755 ( 
.A(n_3749),
.B(n_2063),
.Y(n_3755)
);

AOI21xp5_ASAP7_75t_L g3756 ( 
.A1(n_3459),
.A2(n_3513),
.B(n_3503),
.Y(n_3756)
);

A2O1A1Ixp33_ASAP7_75t_L g3757 ( 
.A1(n_3376),
.A2(n_3339),
.B(n_3019),
.C(n_3023),
.Y(n_3757)
);

O2A1O1Ixp33_ASAP7_75t_L g3758 ( 
.A1(n_3386),
.A2(n_1636),
.B(n_1682),
.C(n_1525),
.Y(n_3758)
);

NAND2x1p5_ASAP7_75t_L g3759 ( 
.A(n_3421),
.B(n_3018),
.Y(n_3759)
);

NAND2xp5_ASAP7_75t_L g3760 ( 
.A(n_3537),
.B(n_2989),
.Y(n_3760)
);

CKINVDCx20_ASAP7_75t_R g3761 ( 
.A(n_3452),
.Y(n_3761)
);

BUFx2_ASAP7_75t_L g3762 ( 
.A(n_3385),
.Y(n_3762)
);

AOI21x1_ASAP7_75t_L g3763 ( 
.A1(n_3354),
.A2(n_3356),
.B(n_3350),
.Y(n_3763)
);

NOR2xp33_ASAP7_75t_R g3764 ( 
.A(n_3741),
.B(n_3271),
.Y(n_3764)
);

AOI21xp5_ASAP7_75t_L g3765 ( 
.A1(n_3544),
.A2(n_2758),
.B(n_2612),
.Y(n_3765)
);

AOI21xp5_ASAP7_75t_L g3766 ( 
.A1(n_3535),
.A2(n_2758),
.B(n_3264),
.Y(n_3766)
);

AOI21xp5_ASAP7_75t_L g3767 ( 
.A1(n_3536),
.A2(n_2593),
.B(n_2484),
.Y(n_3767)
);

NAND2xp5_ASAP7_75t_L g3768 ( 
.A(n_3467),
.B(n_2989),
.Y(n_3768)
);

NAND2xp5_ASAP7_75t_L g3769 ( 
.A(n_3598),
.B(n_2989),
.Y(n_3769)
);

OAI21xp5_ASAP7_75t_L g3770 ( 
.A1(n_3349),
.A2(n_2989),
.B(n_3026),
.Y(n_3770)
);

NAND2xp5_ASAP7_75t_SL g3771 ( 
.A(n_3460),
.B(n_3295),
.Y(n_3771)
);

HB1xp67_ASAP7_75t_L g3772 ( 
.A(n_3502),
.Y(n_3772)
);

OAI21xp5_ASAP7_75t_L g3773 ( 
.A1(n_3367),
.A2(n_3028),
.B(n_3027),
.Y(n_3773)
);

A2O1A1Ixp33_ASAP7_75t_L g3774 ( 
.A1(n_3395),
.A2(n_3031),
.B(n_3035),
.C(n_3030),
.Y(n_3774)
);

AOI21xp33_ASAP7_75t_L g3775 ( 
.A1(n_3469),
.A2(n_3404),
.B(n_3612),
.Y(n_3775)
);

NAND2xp5_ASAP7_75t_SL g3776 ( 
.A(n_3500),
.B(n_3274),
.Y(n_3776)
);

NAND2xp5_ASAP7_75t_L g3777 ( 
.A(n_3478),
.B(n_3036),
.Y(n_3777)
);

AOI21xp5_ASAP7_75t_L g3778 ( 
.A1(n_3607),
.A2(n_2593),
.B(n_2484),
.Y(n_3778)
);

BUFx3_ASAP7_75t_L g3779 ( 
.A(n_3408),
.Y(n_3779)
);

AOI21xp33_ASAP7_75t_L g3780 ( 
.A1(n_3612),
.A2(n_3038),
.B(n_3037),
.Y(n_3780)
);

NAND2xp5_ASAP7_75t_SL g3781 ( 
.A(n_3446),
.B(n_3284),
.Y(n_3781)
);

NOR2xp33_ASAP7_75t_L g3782 ( 
.A(n_3437),
.B(n_3021),
.Y(n_3782)
);

AND2x2_ASAP7_75t_L g3783 ( 
.A(n_3625),
.B(n_1686),
.Y(n_3783)
);

BUFx2_ASAP7_75t_L g3784 ( 
.A(n_3548),
.Y(n_3784)
);

NAND2xp5_ASAP7_75t_L g3785 ( 
.A(n_3482),
.B(n_3041),
.Y(n_3785)
);

OAI21xp5_ASAP7_75t_L g3786 ( 
.A1(n_3424),
.A2(n_3120),
.B(n_3046),
.Y(n_3786)
);

NAND2xp5_ASAP7_75t_SL g3787 ( 
.A(n_3525),
.B(n_3543),
.Y(n_3787)
);

O2A1O1Ixp33_ASAP7_75t_L g3788 ( 
.A1(n_3361),
.A2(n_1094),
.B(n_1098),
.C(n_1079),
.Y(n_3788)
);

AOI22xp33_ASAP7_75t_L g3789 ( 
.A1(n_3580),
.A2(n_3004),
.B1(n_3120),
.B2(n_3160),
.Y(n_3789)
);

BUFx3_ASAP7_75t_L g3790 ( 
.A(n_3599),
.Y(n_3790)
);

AND2x2_ASAP7_75t_L g3791 ( 
.A(n_3466),
.B(n_3044),
.Y(n_3791)
);

NOR2xp67_ASAP7_75t_L g3792 ( 
.A(n_3720),
.B(n_3055),
.Y(n_3792)
);

INVx11_ASAP7_75t_L g3793 ( 
.A(n_3357),
.Y(n_3793)
);

OAI21xp5_ASAP7_75t_L g3794 ( 
.A1(n_3358),
.A2(n_3058),
.B(n_3056),
.Y(n_3794)
);

NAND2xp5_ASAP7_75t_L g3795 ( 
.A(n_3414),
.B(n_3062),
.Y(n_3795)
);

NAND2xp5_ASAP7_75t_L g3796 ( 
.A(n_3560),
.B(n_3069),
.Y(n_3796)
);

NAND2xp5_ASAP7_75t_L g3797 ( 
.A(n_3560),
.B(n_3071),
.Y(n_3797)
);

INVxp67_ASAP7_75t_L g3798 ( 
.A(n_3556),
.Y(n_3798)
);

INVx1_ASAP7_75t_L g3799 ( 
.A(n_3371),
.Y(n_3799)
);

NAND2xp5_ASAP7_75t_L g3800 ( 
.A(n_3455),
.B(n_3474),
.Y(n_3800)
);

CKINVDCx6p67_ASAP7_75t_R g3801 ( 
.A(n_3630),
.Y(n_3801)
);

NAND2xp33_ASAP7_75t_L g3802 ( 
.A(n_3421),
.B(n_3138),
.Y(n_3802)
);

INVx1_ASAP7_75t_L g3803 ( 
.A(n_3382),
.Y(n_3803)
);

NAND2xp5_ASAP7_75t_L g3804 ( 
.A(n_3451),
.B(n_3461),
.Y(n_3804)
);

AOI21xp5_ASAP7_75t_L g3805 ( 
.A1(n_3675),
.A2(n_2593),
.B(n_2484),
.Y(n_3805)
);

INVx2_ASAP7_75t_L g3806 ( 
.A(n_3615),
.Y(n_3806)
);

AOI21xp5_ASAP7_75t_L g3807 ( 
.A1(n_3597),
.A2(n_2811),
.B(n_2796),
.Y(n_3807)
);

NAND2xp5_ASAP7_75t_SL g3808 ( 
.A(n_3522),
.B(n_3284),
.Y(n_3808)
);

NAND2xp5_ASAP7_75t_L g3809 ( 
.A(n_3390),
.B(n_3072),
.Y(n_3809)
);

AOI21xp5_ASAP7_75t_L g3810 ( 
.A1(n_3597),
.A2(n_2811),
.B(n_2796),
.Y(n_3810)
);

O2A1O1Ixp33_ASAP7_75t_L g3811 ( 
.A1(n_3363),
.A2(n_1101),
.B(n_1103),
.C(n_1099),
.Y(n_3811)
);

INVx1_ASAP7_75t_L g3812 ( 
.A(n_3389),
.Y(n_3812)
);

AOI21xp5_ASAP7_75t_L g3813 ( 
.A1(n_3427),
.A2(n_2811),
.B(n_2796),
.Y(n_3813)
);

BUFx3_ASAP7_75t_L g3814 ( 
.A(n_3532),
.Y(n_3814)
);

BUFx3_ASAP7_75t_L g3815 ( 
.A(n_3422),
.Y(n_3815)
);

OAI21xp5_ASAP7_75t_L g3816 ( 
.A1(n_3358),
.A2(n_3076),
.B(n_3073),
.Y(n_3816)
);

AND2x2_ASAP7_75t_L g3817 ( 
.A(n_3648),
.B(n_3077),
.Y(n_3817)
);

AOI21xp5_ASAP7_75t_L g3818 ( 
.A1(n_3360),
.A2(n_3366),
.B(n_3603),
.Y(n_3818)
);

AOI22xp33_ASAP7_75t_L g3819 ( 
.A1(n_3530),
.A2(n_3004),
.B1(n_3160),
.B2(n_3081),
.Y(n_3819)
);

INVx2_ASAP7_75t_L g3820 ( 
.A(n_3628),
.Y(n_3820)
);

O2A1O1Ixp33_ASAP7_75t_L g3821 ( 
.A1(n_3622),
.A2(n_1101),
.B(n_1103),
.C(n_1099),
.Y(n_3821)
);

AOI21xp5_ASAP7_75t_L g3822 ( 
.A1(n_3360),
.A2(n_2852),
.B(n_2811),
.Y(n_3822)
);

AOI21xp5_ASAP7_75t_L g3823 ( 
.A1(n_3366),
.A2(n_2853),
.B(n_2852),
.Y(n_3823)
);

NOR2xp33_ASAP7_75t_L g3824 ( 
.A(n_3642),
.B(n_3239),
.Y(n_3824)
);

NAND2xp5_ASAP7_75t_SL g3825 ( 
.A(n_3683),
.B(n_3138),
.Y(n_3825)
);

AND2x4_ASAP7_75t_L g3826 ( 
.A(n_3632),
.B(n_3043),
.Y(n_3826)
);

AOI22xp5_ASAP7_75t_L g3827 ( 
.A1(n_3411),
.A2(n_3247),
.B1(n_3138),
.B2(n_2418),
.Y(n_3827)
);

AOI21xp5_ASAP7_75t_L g3828 ( 
.A1(n_3603),
.A2(n_2853),
.B(n_2852),
.Y(n_3828)
);

NAND2xp5_ASAP7_75t_L g3829 ( 
.A(n_3453),
.B(n_3623),
.Y(n_3829)
);

NAND2xp5_ASAP7_75t_L g3830 ( 
.A(n_3407),
.B(n_3241),
.Y(n_3830)
);

INVx1_ASAP7_75t_L g3831 ( 
.A(n_3397),
.Y(n_3831)
);

INVx2_ASAP7_75t_L g3832 ( 
.A(n_3634),
.Y(n_3832)
);

AOI21xp5_ASAP7_75t_L g3833 ( 
.A1(n_3684),
.A2(n_2853),
.B(n_2852),
.Y(n_3833)
);

NAND2xp5_ASAP7_75t_L g3834 ( 
.A(n_3464),
.B(n_3243),
.Y(n_3834)
);

NOR2xp33_ASAP7_75t_L g3835 ( 
.A(n_3646),
.B(n_3244),
.Y(n_3835)
);

AOI21xp5_ASAP7_75t_L g3836 ( 
.A1(n_3499),
.A2(n_2869),
.B(n_2853),
.Y(n_3836)
);

AO21x1_ASAP7_75t_L g3837 ( 
.A1(n_3387),
.A2(n_3252),
.B(n_3245),
.Y(n_3837)
);

NAND2xp5_ASAP7_75t_SL g3838 ( 
.A(n_3547),
.B(n_3247),
.Y(n_3838)
);

OAI21xp5_ASAP7_75t_L g3839 ( 
.A1(n_3707),
.A2(n_3258),
.B(n_3254),
.Y(n_3839)
);

OAI22xp5_ASAP7_75t_L g3840 ( 
.A1(n_3440),
.A2(n_3260),
.B1(n_3261),
.B2(n_3259),
.Y(n_3840)
);

INVx2_ASAP7_75t_L g3841 ( 
.A(n_3651),
.Y(n_3841)
);

BUFx4f_ASAP7_75t_L g3842 ( 
.A(n_3365),
.Y(n_3842)
);

AOI21xp5_ASAP7_75t_L g3843 ( 
.A1(n_3499),
.A2(n_2887),
.B(n_2869),
.Y(n_3843)
);

NOR2xp33_ASAP7_75t_L g3844 ( 
.A(n_3620),
.B(n_3265),
.Y(n_3844)
);

NAND2xp5_ASAP7_75t_SL g3845 ( 
.A(n_3575),
.B(n_3247),
.Y(n_3845)
);

NAND2xp5_ASAP7_75t_SL g3846 ( 
.A(n_3516),
.B(n_3566),
.Y(n_3846)
);

O2A1O1Ixp33_ASAP7_75t_L g3847 ( 
.A1(n_3676),
.A2(n_1115),
.B(n_1133),
.C(n_1107),
.Y(n_3847)
);

NAND2xp5_ASAP7_75t_L g3848 ( 
.A(n_3415),
.B(n_3266),
.Y(n_3848)
);

AOI21xp5_ASAP7_75t_L g3849 ( 
.A1(n_3489),
.A2(n_2887),
.B(n_2869),
.Y(n_3849)
);

AOI21xp5_ASAP7_75t_L g3850 ( 
.A1(n_3489),
.A2(n_2887),
.B(n_2869),
.Y(n_3850)
);

INVx2_ASAP7_75t_L g3851 ( 
.A(n_3653),
.Y(n_3851)
);

NAND2xp5_ASAP7_75t_SL g3852 ( 
.A(n_3601),
.B(n_3400),
.Y(n_3852)
);

NOR2xp33_ASAP7_75t_L g3853 ( 
.A(n_3638),
.B(n_3270),
.Y(n_3853)
);

OR2x6_ASAP7_75t_SL g3854 ( 
.A(n_3748),
.B(n_2280),
.Y(n_3854)
);

AOI21xp5_ASAP7_75t_L g3855 ( 
.A1(n_3378),
.A2(n_2908),
.B(n_2887),
.Y(n_3855)
);

NAND2xp5_ASAP7_75t_L g3856 ( 
.A(n_3405),
.B(n_3272),
.Y(n_3856)
);

NAND2xp5_ASAP7_75t_L g3857 ( 
.A(n_3425),
.B(n_3273),
.Y(n_3857)
);

NOR3xp33_ASAP7_75t_L g3858 ( 
.A(n_3432),
.B(n_2000),
.C(n_1115),
.Y(n_3858)
);

NOR2xp33_ASAP7_75t_L g3859 ( 
.A(n_3686),
.B(n_3276),
.Y(n_3859)
);

AOI22xp33_ASAP7_75t_L g3860 ( 
.A1(n_3444),
.A2(n_2666),
.B1(n_3286),
.B2(n_3281),
.Y(n_3860)
);

NAND2x1_ASAP7_75t_L g3861 ( 
.A(n_3526),
.B(n_3697),
.Y(n_3861)
);

A2O1A1Ixp33_ASAP7_75t_L g3862 ( 
.A1(n_3658),
.A2(n_3291),
.B(n_3292),
.C(n_3287),
.Y(n_3862)
);

NAND2xp5_ASAP7_75t_L g3863 ( 
.A(n_3377),
.B(n_3293),
.Y(n_3863)
);

AOI21xp5_ASAP7_75t_L g3864 ( 
.A1(n_3592),
.A2(n_2908),
.B(n_2598),
.Y(n_3864)
);

NAND2xp5_ASAP7_75t_L g3865 ( 
.A(n_3377),
.B(n_3296),
.Y(n_3865)
);

AOI21xp5_ASAP7_75t_L g3866 ( 
.A1(n_3379),
.A2(n_2908),
.B(n_2598),
.Y(n_3866)
);

OAI21xp5_ASAP7_75t_L g3867 ( 
.A1(n_3355),
.A2(n_3301),
.B(n_3297),
.Y(n_3867)
);

AOI21xp5_ASAP7_75t_L g3868 ( 
.A1(n_3379),
.A2(n_2908),
.B(n_2598),
.Y(n_3868)
);

NAND2xp5_ASAP7_75t_L g3869 ( 
.A(n_3409),
.B(n_3305),
.Y(n_3869)
);

INVx1_ASAP7_75t_L g3870 ( 
.A(n_3401),
.Y(n_3870)
);

AOI21xp5_ASAP7_75t_L g3871 ( 
.A1(n_3381),
.A2(n_2598),
.B(n_2581),
.Y(n_3871)
);

AOI21xp5_ASAP7_75t_L g3872 ( 
.A1(n_3381),
.A2(n_3396),
.B(n_3384),
.Y(n_3872)
);

AOI21xp5_ASAP7_75t_L g3873 ( 
.A1(n_3384),
.A2(n_2598),
.B(n_2581),
.Y(n_3873)
);

INVx1_ASAP7_75t_L g3874 ( 
.A(n_3416),
.Y(n_3874)
);

AOI21xp5_ASAP7_75t_L g3875 ( 
.A1(n_3396),
.A2(n_2581),
.B(n_3306),
.Y(n_3875)
);

AOI21xp5_ASAP7_75t_L g3876 ( 
.A1(n_3661),
.A2(n_2581),
.B(n_3307),
.Y(n_3876)
);

INVx1_ASAP7_75t_L g3877 ( 
.A(n_3417),
.Y(n_3877)
);

AOI21xp5_ASAP7_75t_L g3878 ( 
.A1(n_3661),
.A2(n_2581),
.B(n_3308),
.Y(n_3878)
);

NAND3xp33_ASAP7_75t_L g3879 ( 
.A(n_3738),
.B(n_2463),
.C(n_2425),
.Y(n_3879)
);

NAND2xp5_ASAP7_75t_SL g3880 ( 
.A(n_3561),
.B(n_3247),
.Y(n_3880)
);

INVx1_ASAP7_75t_L g3881 ( 
.A(n_3418),
.Y(n_3881)
);

NAND2xp5_ASAP7_75t_L g3882 ( 
.A(n_3431),
.B(n_3310),
.Y(n_3882)
);

NAND2x1p5_ASAP7_75t_L g3883 ( 
.A(n_3421),
.B(n_3312),
.Y(n_3883)
);

AOI21xp5_ASAP7_75t_L g3884 ( 
.A1(n_3563),
.A2(n_3318),
.B(n_3315),
.Y(n_3884)
);

NAND2xp5_ASAP7_75t_SL g3885 ( 
.A(n_3567),
.B(n_3247),
.Y(n_3885)
);

NAND2xp5_ASAP7_75t_L g3886 ( 
.A(n_3483),
.B(n_3323),
.Y(n_3886)
);

NOR2xp33_ASAP7_75t_L g3887 ( 
.A(n_3696),
.B(n_3325),
.Y(n_3887)
);

NAND2xp5_ASAP7_75t_L g3888 ( 
.A(n_3494),
.B(n_3328),
.Y(n_3888)
);

NOR3xp33_ASAP7_75t_L g3889 ( 
.A(n_3399),
.B(n_1133),
.C(n_1107),
.Y(n_3889)
);

OAI22xp5_ASAP7_75t_L g3890 ( 
.A1(n_3420),
.A2(n_3336),
.B1(n_3337),
.B2(n_3330),
.Y(n_3890)
);

O2A1O1Ixp33_ASAP7_75t_L g3891 ( 
.A1(n_3393),
.A2(n_1138),
.B(n_1145),
.C(n_1134),
.Y(n_3891)
);

AOI33xp33_ASAP7_75t_L g3892 ( 
.A1(n_3383),
.A2(n_1563),
.A3(n_1560),
.B1(n_1564),
.B2(n_1561),
.B3(n_1559),
.Y(n_3892)
);

AOI21xp5_ASAP7_75t_L g3893 ( 
.A1(n_3563),
.A2(n_3342),
.B(n_3340),
.Y(n_3893)
);

AOI21xp5_ASAP7_75t_L g3894 ( 
.A1(n_3571),
.A2(n_3345),
.B(n_3343),
.Y(n_3894)
);

NAND2xp5_ASAP7_75t_L g3895 ( 
.A(n_3398),
.B(n_2814),
.Y(n_3895)
);

NAND2xp33_ASAP7_75t_L g3896 ( 
.A(n_3421),
.B(n_2814),
.Y(n_3896)
);

AND2x4_ASAP7_75t_L g3897 ( 
.A(n_3632),
.B(n_3043),
.Y(n_3897)
);

AOI22xp5_ASAP7_75t_L g3898 ( 
.A1(n_3406),
.A2(n_2425),
.B1(n_2418),
.B2(n_3043),
.Y(n_3898)
);

BUFx6f_ASAP7_75t_L g3899 ( 
.A(n_3365),
.Y(n_3899)
);

NAND2xp5_ASAP7_75t_L g3900 ( 
.A(n_3398),
.B(n_3355),
.Y(n_3900)
);

AOI21xp5_ASAP7_75t_L g3901 ( 
.A1(n_3571),
.A2(n_3572),
.B(n_3673),
.Y(n_3901)
);

AOI21xp5_ASAP7_75t_L g3902 ( 
.A1(n_3572),
.A2(n_2383),
.B(n_2515),
.Y(n_3902)
);

BUFx3_ASAP7_75t_L g3903 ( 
.A(n_3374),
.Y(n_3903)
);

AOI21xp5_ASAP7_75t_L g3904 ( 
.A1(n_3687),
.A2(n_2547),
.B(n_2527),
.Y(n_3904)
);

OAI21xp5_ASAP7_75t_L g3905 ( 
.A1(n_3373),
.A2(n_3559),
.B(n_3506),
.Y(n_3905)
);

AOI21xp5_ASAP7_75t_L g3906 ( 
.A1(n_3698),
.A2(n_2547),
.B(n_2527),
.Y(n_3906)
);

NAND2xp5_ASAP7_75t_L g3907 ( 
.A(n_3436),
.B(n_3657),
.Y(n_3907)
);

AOI21xp5_ASAP7_75t_L g3908 ( 
.A1(n_3373),
.A2(n_2547),
.B(n_2527),
.Y(n_3908)
);

NAND2xp5_ASAP7_75t_L g3909 ( 
.A(n_3375),
.B(n_2815),
.Y(n_3909)
);

AOI21xp5_ASAP7_75t_L g3910 ( 
.A1(n_3559),
.A2(n_2564),
.B(n_2551),
.Y(n_3910)
);

INVx1_ASAP7_75t_L g3911 ( 
.A(n_3433),
.Y(n_3911)
);

AOI21xp5_ASAP7_75t_L g3912 ( 
.A1(n_3501),
.A2(n_2564),
.B(n_2551),
.Y(n_3912)
);

AOI21xp5_ASAP7_75t_L g3913 ( 
.A1(n_3501),
.A2(n_2564),
.B(n_2551),
.Y(n_3913)
);

AND2x4_ASAP7_75t_L g3914 ( 
.A(n_3374),
.B(n_3221),
.Y(n_3914)
);

AOI21xp5_ASAP7_75t_L g3915 ( 
.A1(n_3507),
.A2(n_2588),
.B(n_2569),
.Y(n_3915)
);

AOI22xp5_ASAP7_75t_L g3916 ( 
.A1(n_3471),
.A2(n_3221),
.B1(n_2912),
.B2(n_2396),
.Y(n_3916)
);

AOI21x1_ASAP7_75t_L g3917 ( 
.A1(n_3562),
.A2(n_2954),
.B(n_2405),
.Y(n_3917)
);

INVx3_ASAP7_75t_L g3918 ( 
.A(n_3697),
.Y(n_3918)
);

INVx3_ASAP7_75t_L g3919 ( 
.A(n_3650),
.Y(n_3919)
);

INVx2_ASAP7_75t_L g3920 ( 
.A(n_3654),
.Y(n_3920)
);

CKINVDCx10_ASAP7_75t_R g3921 ( 
.A(n_3546),
.Y(n_3921)
);

INVx3_ASAP7_75t_L g3922 ( 
.A(n_3650),
.Y(n_3922)
);

NAND2xp5_ASAP7_75t_L g3923 ( 
.A(n_3375),
.B(n_2815),
.Y(n_3923)
);

OAI21x1_ASAP7_75t_L g3924 ( 
.A1(n_3504),
.A2(n_2588),
.B(n_2569),
.Y(n_3924)
);

OAI22xp5_ASAP7_75t_L g3925 ( 
.A1(n_3388),
.A2(n_2834),
.B1(n_2867),
.B2(n_2815),
.Y(n_3925)
);

NAND2xp5_ASAP7_75t_L g3926 ( 
.A(n_3441),
.B(n_2834),
.Y(n_3926)
);

AOI21x1_ASAP7_75t_L g3927 ( 
.A1(n_3562),
.A2(n_2420),
.B(n_2397),
.Y(n_3927)
);

INVx2_ASAP7_75t_SL g3928 ( 
.A(n_3365),
.Y(n_3928)
);

NAND2xp5_ASAP7_75t_L g3929 ( 
.A(n_3456),
.B(n_2834),
.Y(n_3929)
);

INVx1_ASAP7_75t_L g3930 ( 
.A(n_3463),
.Y(n_3930)
);

AOI22xp33_ASAP7_75t_L g3931 ( 
.A1(n_3670),
.A2(n_2912),
.B1(n_2873),
.B2(n_2867),
.Y(n_3931)
);

NOR2xp33_ASAP7_75t_L g3932 ( 
.A(n_3369),
.B(n_2867),
.Y(n_3932)
);

NOR2xp33_ASAP7_75t_L g3933 ( 
.A(n_3672),
.B(n_2873),
.Y(n_3933)
);

HB1xp67_ASAP7_75t_L g3934 ( 
.A(n_3554),
.Y(n_3934)
);

NAND2xp5_ASAP7_75t_L g3935 ( 
.A(n_3475),
.B(n_2873),
.Y(n_3935)
);

OAI21xp5_ASAP7_75t_L g3936 ( 
.A1(n_3364),
.A2(n_2631),
.B(n_2625),
.Y(n_3936)
);

NOR2xp33_ASAP7_75t_L g3937 ( 
.A(n_3510),
.B(n_2569),
.Y(n_3937)
);

AND2x4_ASAP7_75t_L g3938 ( 
.A(n_3714),
.B(n_3221),
.Y(n_3938)
);

INVx2_ASAP7_75t_SL g3939 ( 
.A(n_3480),
.Y(n_3939)
);

INVx1_ASAP7_75t_L g3940 ( 
.A(n_3479),
.Y(n_3940)
);

AND2x4_ASAP7_75t_L g3941 ( 
.A(n_3729),
.B(n_2588),
.Y(n_3941)
);

NAND2xp5_ASAP7_75t_L g3942 ( 
.A(n_3481),
.B(n_2606),
.Y(n_3942)
);

AOI22xp33_ASAP7_75t_L g3943 ( 
.A1(n_3618),
.A2(n_2607),
.B1(n_2619),
.B2(n_2606),
.Y(n_3943)
);

AOI22xp33_ASAP7_75t_L g3944 ( 
.A1(n_3539),
.A2(n_2607),
.B1(n_2619),
.B2(n_2606),
.Y(n_3944)
);

AOI21xp5_ASAP7_75t_L g3945 ( 
.A1(n_3507),
.A2(n_2619),
.B(n_2607),
.Y(n_3945)
);

AOI21xp5_ASAP7_75t_L g3946 ( 
.A1(n_3508),
.A2(n_2631),
.B(n_2625),
.Y(n_3946)
);

HB1xp67_ASAP7_75t_L g3947 ( 
.A(n_3564),
.Y(n_3947)
);

AOI222xp33_ASAP7_75t_L g3948 ( 
.A1(n_3699),
.A2(n_1146),
.B1(n_1138),
.B2(n_1148),
.C1(n_1145),
.C2(n_1134),
.Y(n_3948)
);

NAND2xp5_ASAP7_75t_L g3949 ( 
.A(n_3487),
.B(n_2625),
.Y(n_3949)
);

OAI21xp33_ASAP7_75t_L g3950 ( 
.A1(n_3486),
.A2(n_881),
.B(n_879),
.Y(n_3950)
);

INVx2_ASAP7_75t_L g3951 ( 
.A(n_3660),
.Y(n_3951)
);

INVx2_ASAP7_75t_SL g3952 ( 
.A(n_3480),
.Y(n_3952)
);

NAND2xp5_ASAP7_75t_L g3953 ( 
.A(n_3511),
.B(n_2631),
.Y(n_3953)
);

OAI21xp33_ASAP7_75t_L g3954 ( 
.A1(n_3644),
.A2(n_888),
.B(n_885),
.Y(n_3954)
);

OAI321xp33_ASAP7_75t_L g3955 ( 
.A1(n_3476),
.A2(n_1156),
.A3(n_1148),
.B1(n_1160),
.B2(n_1149),
.C(n_1146),
.Y(n_3955)
);

INVx1_ASAP7_75t_L g3956 ( 
.A(n_3519),
.Y(n_3956)
);

O2A1O1Ixp33_ASAP7_75t_L g3957 ( 
.A1(n_3419),
.A2(n_1156),
.B(n_1160),
.C(n_1149),
.Y(n_3957)
);

AOI21xp5_ASAP7_75t_L g3958 ( 
.A1(n_3508),
.A2(n_2636),
.B(n_2468),
.Y(n_3958)
);

AOI21xp5_ASAP7_75t_L g3959 ( 
.A1(n_3509),
.A2(n_2636),
.B(n_2468),
.Y(n_3959)
);

NOR2xp67_ASAP7_75t_L g3960 ( 
.A(n_3712),
.B(n_2636),
.Y(n_3960)
);

AOI22xp5_ASAP7_75t_L g3961 ( 
.A1(n_3434),
.A2(n_2421),
.B1(n_2427),
.B2(n_2426),
.Y(n_3961)
);

AOI21xp5_ASAP7_75t_L g3962 ( 
.A1(n_3509),
.A2(n_2468),
.B(n_2462),
.Y(n_3962)
);

AOI21xp5_ASAP7_75t_L g3963 ( 
.A1(n_3512),
.A2(n_2468),
.B(n_2402),
.Y(n_3963)
);

NAND2xp5_ASAP7_75t_L g3964 ( 
.A(n_3531),
.B(n_1945),
.Y(n_3964)
);

OAI21xp5_ASAP7_75t_L g3965 ( 
.A1(n_3504),
.A2(n_3506),
.B(n_3512),
.Y(n_3965)
);

NAND2xp5_ASAP7_75t_L g3966 ( 
.A(n_3534),
.B(n_1948),
.Y(n_3966)
);

NAND2xp5_ASAP7_75t_L g3967 ( 
.A(n_3549),
.B(n_1970),
.Y(n_3967)
);

NAND2xp5_ASAP7_75t_L g3968 ( 
.A(n_3484),
.B(n_3488),
.Y(n_3968)
);

INVx1_ASAP7_75t_L g3969 ( 
.A(n_3551),
.Y(n_3969)
);

CKINVDCx20_ASAP7_75t_R g3970 ( 
.A(n_3372),
.Y(n_3970)
);

NAND2xp5_ASAP7_75t_L g3971 ( 
.A(n_3484),
.B(n_2456),
.Y(n_3971)
);

A2O1A1Ixp33_ASAP7_75t_L g3972 ( 
.A1(n_3498),
.A2(n_2471),
.B(n_2476),
.C(n_2461),
.Y(n_3972)
);

NAND2xp5_ASAP7_75t_L g3973 ( 
.A(n_3488),
.B(n_1883),
.Y(n_3973)
);

INVx2_ASAP7_75t_L g3974 ( 
.A(n_3666),
.Y(n_3974)
);

O2A1O1Ixp5_ASAP7_75t_L g3975 ( 
.A1(n_3552),
.A2(n_2432),
.B(n_2433),
.C(n_2428),
.Y(n_3975)
);

INVx1_ASAP7_75t_L g3976 ( 
.A(n_3570),
.Y(n_3976)
);

NOR3xp33_ASAP7_75t_L g3977 ( 
.A(n_3454),
.B(n_1172),
.C(n_1170),
.Y(n_3977)
);

OAI21xp33_ASAP7_75t_L g3978 ( 
.A1(n_3582),
.A2(n_3709),
.B(n_3677),
.Y(n_3978)
);

AOI21xp5_ASAP7_75t_L g3979 ( 
.A1(n_3514),
.A2(n_2402),
.B(n_2379),
.Y(n_3979)
);

NAND2xp5_ASAP7_75t_L g3980 ( 
.A(n_3540),
.B(n_1883),
.Y(n_3980)
);

NAND2xp5_ASAP7_75t_L g3981 ( 
.A(n_3550),
.B(n_1904),
.Y(n_3981)
);

OAI321xp33_ASAP7_75t_L g3982 ( 
.A1(n_3736),
.A2(n_1185),
.A3(n_1172),
.B1(n_1190),
.B2(n_1181),
.C(n_1170),
.Y(n_3982)
);

INVx3_ASAP7_75t_L g3983 ( 
.A(n_3650),
.Y(n_3983)
);

INVx1_ASAP7_75t_SL g3984 ( 
.A(n_3392),
.Y(n_3984)
);

NOR2xp33_ASAP7_75t_L g3985 ( 
.A(n_3438),
.B(n_2434),
.Y(n_3985)
);

NAND2xp5_ASAP7_75t_L g3986 ( 
.A(n_3412),
.B(n_1904),
.Y(n_3986)
);

OAI22xp5_ASAP7_75t_L g3987 ( 
.A1(n_3610),
.A2(n_2335),
.B1(n_2455),
.B2(n_2379),
.Y(n_3987)
);

INVx1_ASAP7_75t_L g3988 ( 
.A(n_3581),
.Y(n_3988)
);

INVx2_ASAP7_75t_L g3989 ( 
.A(n_3671),
.Y(n_3989)
);

AOI21xp5_ASAP7_75t_L g3990 ( 
.A1(n_3514),
.A2(n_2455),
.B(n_2169),
.Y(n_3990)
);

NOR2xp33_ASAP7_75t_L g3991 ( 
.A(n_3465),
.B(n_2443),
.Y(n_3991)
);

NAND2xp5_ASAP7_75t_SL g3992 ( 
.A(n_3391),
.B(n_889),
.Y(n_3992)
);

A2O1A1Ixp33_ASAP7_75t_L g3993 ( 
.A1(n_3583),
.A2(n_1185),
.B(n_1190),
.C(n_1181),
.Y(n_3993)
);

AOI21xp5_ASAP7_75t_L g3994 ( 
.A1(n_3527),
.A2(n_2190),
.B(n_2084),
.Y(n_3994)
);

AOI21xp5_ASAP7_75t_L g3995 ( 
.A1(n_3527),
.A2(n_2190),
.B(n_2084),
.Y(n_3995)
);

NOR2xp33_ASAP7_75t_L g3996 ( 
.A(n_3631),
.B(n_890),
.Y(n_3996)
);

AOI21xp5_ASAP7_75t_L g3997 ( 
.A1(n_3643),
.A2(n_3705),
.B(n_3679),
.Y(n_3997)
);

INVx1_ASAP7_75t_L g3998 ( 
.A(n_3617),
.Y(n_3998)
);

AOI21xp5_ASAP7_75t_L g3999 ( 
.A1(n_3606),
.A2(n_2145),
.B(n_2102),
.Y(n_3999)
);

NAND2xp5_ASAP7_75t_L g4000 ( 
.A(n_3663),
.B(n_1934),
.Y(n_4000)
);

NAND2xp5_ASAP7_75t_L g4001 ( 
.A(n_3688),
.B(n_1934),
.Y(n_4001)
);

NAND2xp5_ASAP7_75t_SL g4002 ( 
.A(n_3391),
.B(n_891),
.Y(n_4002)
);

O2A1O1Ixp33_ASAP7_75t_SL g4003 ( 
.A1(n_3737),
.A2(n_1201),
.B(n_1202),
.C(n_1195),
.Y(n_4003)
);

AOI21xp5_ASAP7_75t_L g4004 ( 
.A1(n_3740),
.A2(n_2254),
.B(n_2153),
.Y(n_4004)
);

AO21x1_ASAP7_75t_L g4005 ( 
.A1(n_3569),
.A2(n_1201),
.B(n_1195),
.Y(n_4005)
);

AOI21xp5_ASAP7_75t_L g4006 ( 
.A1(n_3745),
.A2(n_2129),
.B(n_2080),
.Y(n_4006)
);

INVx3_ASAP7_75t_L g4007 ( 
.A(n_3667),
.Y(n_4007)
);

OAI21xp33_ASAP7_75t_L g4008 ( 
.A1(n_3627),
.A2(n_3704),
.B(n_3680),
.Y(n_4008)
);

AOI21xp5_ASAP7_75t_L g4009 ( 
.A1(n_3694),
.A2(n_2129),
.B(n_2080),
.Y(n_4009)
);

INVx2_ASAP7_75t_L g4010 ( 
.A(n_3692),
.Y(n_4010)
);

AOI21xp5_ASAP7_75t_L g4011 ( 
.A1(n_3541),
.A2(n_2129),
.B(n_2080),
.Y(n_4011)
);

AOI21xp5_ASAP7_75t_L g4012 ( 
.A1(n_3542),
.A2(n_2129),
.B(n_2080),
.Y(n_4012)
);

AOI21xp5_ASAP7_75t_L g4013 ( 
.A1(n_3685),
.A2(n_2139),
.B(n_2084),
.Y(n_4013)
);

BUFx2_ASAP7_75t_L g4014 ( 
.A(n_3645),
.Y(n_4014)
);

AOI21xp5_ASAP7_75t_L g4015 ( 
.A1(n_3587),
.A2(n_2139),
.B(n_2084),
.Y(n_4015)
);

NAND2xp5_ASAP7_75t_L g4016 ( 
.A(n_3708),
.B(n_1980),
.Y(n_4016)
);

NAND2xp5_ASAP7_75t_L g4017 ( 
.A(n_3727),
.B(n_1980),
.Y(n_4017)
);

AOI21xp5_ASAP7_75t_L g4018 ( 
.A1(n_3600),
.A2(n_2196),
.B(n_2145),
.Y(n_4018)
);

INVx1_ASAP7_75t_L g4019 ( 
.A(n_3619),
.Y(n_4019)
);

AOI21xp5_ASAP7_75t_L g4020 ( 
.A1(n_3589),
.A2(n_2196),
.B(n_2145),
.Y(n_4020)
);

O2A1O1Ixp33_ASAP7_75t_L g4021 ( 
.A1(n_3402),
.A2(n_1205),
.B(n_1207),
.C(n_1202),
.Y(n_4021)
);

OAI21xp5_ASAP7_75t_L g4022 ( 
.A1(n_3739),
.A2(n_2467),
.B(n_2465),
.Y(n_4022)
);

OAI21xp5_ASAP7_75t_L g4023 ( 
.A1(n_3746),
.A2(n_2467),
.B(n_2465),
.Y(n_4023)
);

AOI21x1_ASAP7_75t_L g4024 ( 
.A1(n_3573),
.A2(n_1569),
.B(n_1568),
.Y(n_4024)
);

NAND2xp5_ASAP7_75t_L g4025 ( 
.A(n_3728),
.B(n_3403),
.Y(n_4025)
);

AOI21xp33_ASAP7_75t_L g4026 ( 
.A1(n_3528),
.A2(n_895),
.B(n_892),
.Y(n_4026)
);

NAND2xp5_ASAP7_75t_SL g4027 ( 
.A(n_3710),
.B(n_897),
.Y(n_4027)
);

NAND2xp5_ASAP7_75t_SL g4028 ( 
.A(n_3710),
.B(n_899),
.Y(n_4028)
);

INVx2_ASAP7_75t_L g4029 ( 
.A(n_3695),
.Y(n_4029)
);

AOI21xp5_ASAP7_75t_L g4030 ( 
.A1(n_3641),
.A2(n_2190),
.B(n_2096),
.Y(n_4030)
);

NAND2xp5_ASAP7_75t_SL g4031 ( 
.A(n_3710),
.B(n_903),
.Y(n_4031)
);

OAI22xp5_ASAP7_75t_L g4032 ( 
.A1(n_3667),
.A2(n_2335),
.B1(n_2078),
.B2(n_2100),
.Y(n_4032)
);

AND2x4_ASAP7_75t_L g4033 ( 
.A(n_3429),
.B(n_2073),
.Y(n_4033)
);

NAND2xp5_ASAP7_75t_L g4034 ( 
.A(n_3718),
.B(n_2073),
.Y(n_4034)
);

AOI21xp5_ASAP7_75t_L g4035 ( 
.A1(n_3641),
.A2(n_2285),
.B(n_2102),
.Y(n_4035)
);

AOI22xp5_ASAP7_75t_L g4036 ( 
.A1(n_3529),
.A2(n_2335),
.B1(n_905),
.B2(n_907),
.Y(n_4036)
);

AOI21xp5_ASAP7_75t_L g4037 ( 
.A1(n_3722),
.A2(n_2300),
.B(n_2169),
.Y(n_4037)
);

AOI21xp5_ASAP7_75t_L g4038 ( 
.A1(n_3722),
.A2(n_2300),
.B(n_2169),
.Y(n_4038)
);

OAI22xp5_ASAP7_75t_L g4039 ( 
.A1(n_3798),
.A2(n_3558),
.B1(n_3742),
.B2(n_3732),
.Y(n_4039)
);

NAND2xp5_ASAP7_75t_L g4040 ( 
.A(n_3800),
.B(n_3426),
.Y(n_4040)
);

INVx4_ASAP7_75t_L g4041 ( 
.A(n_3842),
.Y(n_4041)
);

NAND2xp5_ASAP7_75t_L g4042 ( 
.A(n_3783),
.B(n_3426),
.Y(n_4042)
);

INVx2_ASAP7_75t_SL g4043 ( 
.A(n_3921),
.Y(n_4043)
);

INVx2_ASAP7_75t_L g4044 ( 
.A(n_3806),
.Y(n_4044)
);

INVx11_ASAP7_75t_L g4045 ( 
.A(n_3793),
.Y(n_4045)
);

OAI21xp33_ASAP7_75t_L g4046 ( 
.A1(n_3889),
.A2(n_3430),
.B(n_3518),
.Y(n_4046)
);

OAI21xp5_ASAP7_75t_L g4047 ( 
.A1(n_3775),
.A2(n_3457),
.B(n_3410),
.Y(n_4047)
);

NAND2xp5_ASAP7_75t_L g4048 ( 
.A(n_3829),
.B(n_3443),
.Y(n_4048)
);

NAND2xp5_ASAP7_75t_L g4049 ( 
.A(n_3907),
.B(n_3443),
.Y(n_4049)
);

NAND2xp5_ASAP7_75t_L g4050 ( 
.A(n_3859),
.B(n_3584),
.Y(n_4050)
);

AO22x1_ASAP7_75t_L g4051 ( 
.A1(n_3824),
.A2(n_3595),
.B1(n_3605),
.B2(n_3750),
.Y(n_4051)
);

AOI22xp33_ASAP7_75t_L g4052 ( 
.A1(n_3977),
.A2(n_3546),
.B1(n_3521),
.B2(n_3505),
.Y(n_4052)
);

O2A1O1Ixp33_ASAP7_75t_L g4053 ( 
.A1(n_3821),
.A2(n_3468),
.B(n_3520),
.C(n_3497),
.Y(n_4053)
);

HB1xp67_ASAP7_75t_L g4054 ( 
.A(n_3762),
.Y(n_4054)
);

OR2x2_ASAP7_75t_L g4055 ( 
.A(n_3984),
.B(n_3496),
.Y(n_4055)
);

AOI21xp5_ASAP7_75t_L g4056 ( 
.A1(n_3756),
.A2(n_3667),
.B(n_3495),
.Y(n_4056)
);

NAND2xp5_ASAP7_75t_SL g4057 ( 
.A(n_3844),
.B(n_3533),
.Y(n_4057)
);

NOR3xp33_ASAP7_75t_L g4058 ( 
.A(n_4008),
.B(n_3590),
.C(n_3568),
.Y(n_4058)
);

AOI21xp5_ASAP7_75t_L g4059 ( 
.A1(n_3802),
.A2(n_3744),
.B(n_3576),
.Y(n_4059)
);

AOI21xp5_ASAP7_75t_L g4060 ( 
.A1(n_3765),
.A2(n_3744),
.B(n_3576),
.Y(n_4060)
);

O2A1O1Ixp5_ASAP7_75t_L g4061 ( 
.A1(n_3825),
.A2(n_3690),
.B(n_3701),
.C(n_3693),
.Y(n_4061)
);

OR2x6_ASAP7_75t_SL g4062 ( 
.A(n_3879),
.B(n_3736),
.Y(n_4062)
);

NAND2xp5_ASAP7_75t_L g4063 ( 
.A(n_3887),
.B(n_3574),
.Y(n_4063)
);

BUFx2_ASAP7_75t_L g4064 ( 
.A(n_3784),
.Y(n_4064)
);

NAND2xp5_ASAP7_75t_L g4065 ( 
.A(n_3835),
.B(n_3574),
.Y(n_4065)
);

NOR2xp33_ASAP7_75t_R g4066 ( 
.A(n_3761),
.B(n_3480),
.Y(n_4066)
);

NAND2xp5_ASAP7_75t_L g4067 ( 
.A(n_3817),
.B(n_3635),
.Y(n_4067)
);

INVx1_ASAP7_75t_L g4068 ( 
.A(n_3799),
.Y(n_4068)
);

O2A1O1Ixp33_ASAP7_75t_L g4069 ( 
.A1(n_3788),
.A2(n_3449),
.B(n_1207),
.C(n_1210),
.Y(n_4069)
);

NAND2xp5_ASAP7_75t_L g4070 ( 
.A(n_3755),
.B(n_3635),
.Y(n_4070)
);

NOR2xp33_ASAP7_75t_L g4071 ( 
.A(n_3787),
.B(n_3721),
.Y(n_4071)
);

INVx1_ASAP7_75t_L g4072 ( 
.A(n_3803),
.Y(n_4072)
);

AOI21xp5_ASAP7_75t_L g4073 ( 
.A1(n_3896),
.A2(n_3578),
.B(n_3573),
.Y(n_4073)
);

HB1xp67_ASAP7_75t_L g4074 ( 
.A(n_3772),
.Y(n_4074)
);

CKINVDCx20_ASAP7_75t_R g4075 ( 
.A(n_3970),
.Y(n_4075)
);

HB1xp67_ASAP7_75t_L g4076 ( 
.A(n_3934),
.Y(n_4076)
);

AOI22xp33_ASAP7_75t_L g4077 ( 
.A1(n_3978),
.A2(n_3717),
.B1(n_3470),
.B2(n_3636),
.Y(n_4077)
);

NOR2xp33_ASAP7_75t_SL g4078 ( 
.A(n_3801),
.B(n_3636),
.Y(n_4078)
);

OAI22xp5_ASAP7_75t_L g4079 ( 
.A1(n_3846),
.A2(n_3470),
.B1(n_3636),
.B2(n_3702),
.Y(n_4079)
);

NAND2xp5_ASAP7_75t_SL g4080 ( 
.A(n_3792),
.B(n_3721),
.Y(n_4080)
);

NAND2xp5_ASAP7_75t_SL g4081 ( 
.A(n_3853),
.B(n_3721),
.Y(n_4081)
);

NAND2xp5_ASAP7_75t_L g4082 ( 
.A(n_3804),
.B(n_3717),
.Y(n_4082)
);

OAI22xp5_ASAP7_75t_L g4083 ( 
.A1(n_3752),
.A2(n_3470),
.B1(n_3711),
.B2(n_3706),
.Y(n_4083)
);

BUFx12f_ASAP7_75t_L g4084 ( 
.A(n_3899),
.Y(n_4084)
);

OAI22xp5_ASAP7_75t_L g4085 ( 
.A1(n_3933),
.A2(n_3961),
.B1(n_3827),
.B2(n_3819),
.Y(n_4085)
);

NAND2xp5_ASAP7_75t_SL g4086 ( 
.A(n_3985),
.B(n_3725),
.Y(n_4086)
);

INVx2_ASAP7_75t_L g4087 ( 
.A(n_3820),
.Y(n_4087)
);

OAI22xp5_ASAP7_75t_L g4088 ( 
.A1(n_3984),
.A2(n_3524),
.B1(n_3633),
.B2(n_3629),
.Y(n_4088)
);

OR2x2_ASAP7_75t_L g4089 ( 
.A(n_3809),
.B(n_3747),
.Y(n_4089)
);

OAI21xp33_ASAP7_75t_SL g4090 ( 
.A1(n_3892),
.A2(n_3734),
.B(n_3713),
.Y(n_4090)
);

AOI21xp5_ASAP7_75t_L g4091 ( 
.A1(n_3901),
.A2(n_3579),
.B(n_3578),
.Y(n_4091)
);

OAI21xp5_ASAP7_75t_L g4092 ( 
.A1(n_3811),
.A2(n_3616),
.B(n_3731),
.Y(n_4092)
);

NAND2xp5_ASAP7_75t_SL g4093 ( 
.A(n_3991),
.B(n_3639),
.Y(n_4093)
);

NOR2xp33_ASAP7_75t_L g4094 ( 
.A(n_3932),
.B(n_3423),
.Y(n_4094)
);

OR2x6_ASAP7_75t_L g4095 ( 
.A(n_3899),
.B(n_3524),
.Y(n_4095)
);

AND2x4_ASAP7_75t_L g4096 ( 
.A(n_3826),
.B(n_3353),
.Y(n_4096)
);

INVx4_ASAP7_75t_L g4097 ( 
.A(n_3842),
.Y(n_4097)
);

OR2x6_ASAP7_75t_L g4098 ( 
.A(n_3899),
.B(n_3524),
.Y(n_4098)
);

NAND2xp5_ASAP7_75t_L g4099 ( 
.A(n_3857),
.B(n_3640),
.Y(n_4099)
);

NAND2xp5_ASAP7_75t_SL g4100 ( 
.A(n_3937),
.B(n_3662),
.Y(n_4100)
);

INVx1_ASAP7_75t_L g4101 ( 
.A(n_3812),
.Y(n_4101)
);

AOI21xp5_ASAP7_75t_L g4102 ( 
.A1(n_3766),
.A2(n_3585),
.B(n_3579),
.Y(n_4102)
);

NAND2xp5_ASAP7_75t_L g4103 ( 
.A(n_3882),
.B(n_3791),
.Y(n_4103)
);

INVx3_ASAP7_75t_SL g4104 ( 
.A(n_3771),
.Y(n_4104)
);

BUFx3_ASAP7_75t_L g4105 ( 
.A(n_3779),
.Y(n_4105)
);

INVx1_ASAP7_75t_L g4106 ( 
.A(n_3831),
.Y(n_4106)
);

NOR2xp33_ASAP7_75t_L g4107 ( 
.A(n_4026),
.B(n_3790),
.Y(n_4107)
);

NOR2xp33_ASAP7_75t_SL g4108 ( 
.A(n_3782),
.B(n_3353),
.Y(n_4108)
);

HB1xp67_ASAP7_75t_L g4109 ( 
.A(n_3947),
.Y(n_4109)
);

NAND2xp5_ASAP7_75t_SL g4110 ( 
.A(n_3834),
.B(n_3669),
.Y(n_4110)
);

NOR3xp33_ASAP7_75t_L g4111 ( 
.A(n_3992),
.B(n_1575),
.C(n_1574),
.Y(n_4111)
);

INVx2_ASAP7_75t_L g4112 ( 
.A(n_3832),
.Y(n_4112)
);

CKINVDCx5p33_ASAP7_75t_R g4113 ( 
.A(n_3764),
.Y(n_4113)
);

NAND2x1p5_ASAP7_75t_L g4114 ( 
.A(n_3918),
.B(n_3380),
.Y(n_4114)
);

AOI21xp5_ASAP7_75t_L g4115 ( 
.A1(n_3754),
.A2(n_3586),
.B(n_3585),
.Y(n_4115)
);

AOI21xp5_ASAP7_75t_L g4116 ( 
.A1(n_3872),
.A2(n_3586),
.B(n_3362),
.Y(n_4116)
);

INVxp67_ASAP7_75t_L g4117 ( 
.A(n_4014),
.Y(n_4117)
);

O2A1O1Ixp33_ASAP7_75t_SL g4118 ( 
.A1(n_3757),
.A2(n_3613),
.B(n_3626),
.C(n_3624),
.Y(n_4118)
);

NOR2xp67_ASAP7_75t_L g4119 ( 
.A(n_3928),
.B(n_3439),
.Y(n_4119)
);

BUFx6f_ASAP7_75t_L g4120 ( 
.A(n_3903),
.Y(n_4120)
);

NAND2xp5_ASAP7_75t_SL g4121 ( 
.A(n_3886),
.B(n_3674),
.Y(n_4121)
);

NAND2xp5_ASAP7_75t_L g4122 ( 
.A(n_3856),
.B(n_3888),
.Y(n_4122)
);

OR2x6_ASAP7_75t_SL g4123 ( 
.A(n_3768),
.B(n_904),
.Y(n_4123)
);

AOI21xp5_ASAP7_75t_L g4124 ( 
.A1(n_3807),
.A2(n_3611),
.B(n_3609),
.Y(n_4124)
);

NAND2xp5_ASAP7_75t_L g4125 ( 
.A(n_3830),
.B(n_3682),
.Y(n_4125)
);

AOI21xp5_ASAP7_75t_L g4126 ( 
.A1(n_3810),
.A2(n_3611),
.B(n_3609),
.Y(n_4126)
);

NAND2xp5_ASAP7_75t_L g4127 ( 
.A(n_3848),
.B(n_3689),
.Y(n_4127)
);

OAI21xp5_ASAP7_75t_L g4128 ( 
.A1(n_3862),
.A2(n_3753),
.B(n_3760),
.Y(n_4128)
);

O2A1O1Ixp33_ASAP7_75t_SL g4129 ( 
.A1(n_3845),
.A2(n_3649),
.B(n_3668),
.C(n_3655),
.Y(n_4129)
);

NOR2xp67_ASAP7_75t_SL g4130 ( 
.A(n_3982),
.B(n_3700),
.Y(n_4130)
);

OAI22xp5_ASAP7_75t_L g4131 ( 
.A1(n_3789),
.A2(n_3691),
.B1(n_3703),
.B2(n_3719),
.Y(n_4131)
);

NOR2xp33_ASAP7_75t_L g4132 ( 
.A(n_3814),
.B(n_3348),
.Y(n_4132)
);

OR2x6_ASAP7_75t_SL g4133 ( 
.A(n_3769),
.B(n_909),
.Y(n_4133)
);

AOI21xp5_ASAP7_75t_L g4134 ( 
.A1(n_3818),
.A2(n_3621),
.B(n_3637),
.Y(n_4134)
);

NAND2xp5_ASAP7_75t_L g4135 ( 
.A(n_3900),
.B(n_3723),
.Y(n_4135)
);

AOI21xp5_ASAP7_75t_L g4136 ( 
.A1(n_3997),
.A2(n_3621),
.B(n_3637),
.Y(n_4136)
);

OAI21xp33_ASAP7_75t_L g4137 ( 
.A1(n_3954),
.A2(n_913),
.B(n_911),
.Y(n_4137)
);

A2O1A1Ixp33_ASAP7_75t_L g4138 ( 
.A1(n_3780),
.A2(n_3758),
.B(n_3858),
.C(n_3950),
.Y(n_4138)
);

AND2x4_ASAP7_75t_L g4139 ( 
.A(n_3826),
.B(n_3380),
.Y(n_4139)
);

NOR2xp67_ASAP7_75t_L g4140 ( 
.A(n_3939),
.B(n_3439),
.Y(n_4140)
);

OAI22xp5_ASAP7_75t_L g4141 ( 
.A1(n_3916),
.A2(n_3743),
.B1(n_3751),
.B2(n_3608),
.Y(n_4141)
);

AOI21xp5_ASAP7_75t_L g4142 ( 
.A1(n_3794),
.A2(n_3647),
.B(n_3665),
.Y(n_4142)
);

BUFx6f_ASAP7_75t_L g4143 ( 
.A(n_3914),
.Y(n_4143)
);

INVx1_ASAP7_75t_L g4144 ( 
.A(n_3870),
.Y(n_4144)
);

NAND2xp5_ASAP7_75t_L g4145 ( 
.A(n_3777),
.B(n_3351),
.Y(n_4145)
);

NOR2xp33_ASAP7_75t_L g4146 ( 
.A(n_3781),
.B(n_3352),
.Y(n_4146)
);

O2A1O1Ixp33_ASAP7_75t_L g4147 ( 
.A1(n_3847),
.A2(n_1210),
.B(n_1211),
.C(n_1205),
.Y(n_4147)
);

AO21x1_ASAP7_75t_L g4148 ( 
.A1(n_3840),
.A2(n_3678),
.B(n_3681),
.Y(n_4148)
);

OAI22xp5_ASAP7_75t_L g4149 ( 
.A1(n_3785),
.A2(n_3656),
.B1(n_3659),
.B2(n_3652),
.Y(n_4149)
);

BUFx2_ASAP7_75t_L g4150 ( 
.A(n_3941),
.Y(n_4150)
);

NAND2xp5_ASAP7_75t_SL g4151 ( 
.A(n_3941),
.B(n_3664),
.Y(n_4151)
);

AO32x1_ASAP7_75t_L g4152 ( 
.A1(n_3890),
.A2(n_1227),
.A3(n_1232),
.B1(n_1216),
.B2(n_1211),
.Y(n_4152)
);

INVx4_ASAP7_75t_L g4153 ( 
.A(n_3918),
.Y(n_4153)
);

NOR2xp67_ASAP7_75t_L g4154 ( 
.A(n_3952),
.B(n_3442),
.Y(n_4154)
);

INVx2_ASAP7_75t_L g4155 ( 
.A(n_3841),
.Y(n_4155)
);

O2A1O1Ixp33_ASAP7_75t_L g4156 ( 
.A1(n_3852),
.A2(n_1227),
.B(n_1232),
.C(n_1216),
.Y(n_4156)
);

A2O1A1Ixp33_ASAP7_75t_L g4157 ( 
.A1(n_3955),
.A2(n_3726),
.B(n_3700),
.C(n_3593),
.Y(n_4157)
);

INVx1_ASAP7_75t_L g4158 ( 
.A(n_3874),
.Y(n_4158)
);

NAND2xp5_ASAP7_75t_L g4159 ( 
.A(n_3795),
.B(n_3359),
.Y(n_4159)
);

INVx2_ASAP7_75t_L g4160 ( 
.A(n_3851),
.Y(n_4160)
);

BUFx6f_ASAP7_75t_L g4161 ( 
.A(n_3914),
.Y(n_4161)
);

INVx4_ASAP7_75t_L g4162 ( 
.A(n_3897),
.Y(n_4162)
);

NAND2xp5_ASAP7_75t_SL g4163 ( 
.A(n_4025),
.B(n_3588),
.Y(n_4163)
);

AOI21xp5_ASAP7_75t_L g4164 ( 
.A1(n_3794),
.A2(n_3665),
.B(n_3647),
.Y(n_4164)
);

A2O1A1Ixp33_ASAP7_75t_L g4165 ( 
.A1(n_3955),
.A2(n_3726),
.B(n_3596),
.C(n_3413),
.Y(n_4165)
);

INVx1_ASAP7_75t_L g4166 ( 
.A(n_3877),
.Y(n_4166)
);

NAND3xp33_ASAP7_75t_L g4167 ( 
.A(n_3948),
.B(n_918),
.C(n_917),
.Y(n_4167)
);

AOI21xp5_ASAP7_75t_L g4168 ( 
.A1(n_3816),
.A2(n_3724),
.B(n_3716),
.Y(n_4168)
);

O2A1O1Ixp5_ASAP7_75t_L g4169 ( 
.A1(n_3786),
.A2(n_3716),
.B(n_3730),
.C(n_3724),
.Y(n_4169)
);

BUFx6f_ASAP7_75t_L g4170 ( 
.A(n_3897),
.Y(n_4170)
);

NAND2xp5_ASAP7_75t_L g4171 ( 
.A(n_3996),
.B(n_3368),
.Y(n_4171)
);

O2A1O1Ixp33_ASAP7_75t_L g4172 ( 
.A1(n_3993),
.A2(n_1236),
.B(n_1238),
.C(n_1237),
.Y(n_4172)
);

AND2x2_ASAP7_75t_L g4173 ( 
.A(n_3938),
.B(n_3428),
.Y(n_4173)
);

NOR3xp33_ASAP7_75t_L g4174 ( 
.A(n_4002),
.B(n_1580),
.C(n_1579),
.Y(n_4174)
);

INVx1_ASAP7_75t_L g4175 ( 
.A(n_3881),
.Y(n_4175)
);

AOI21xp5_ASAP7_75t_L g4176 ( 
.A1(n_3816),
.A2(n_3733),
.B(n_3730),
.Y(n_4176)
);

OAI21xp5_ASAP7_75t_L g4177 ( 
.A1(n_3770),
.A2(n_3731),
.B(n_3715),
.Y(n_4177)
);

A2O1A1Ixp33_ASAP7_75t_L g4178 ( 
.A1(n_3891),
.A2(n_3445),
.B(n_3447),
.C(n_3435),
.Y(n_4178)
);

INVx1_ASAP7_75t_SL g4179 ( 
.A(n_3776),
.Y(n_4179)
);

OAI22xp5_ASAP7_75t_L g4180 ( 
.A1(n_3796),
.A2(n_3591),
.B1(n_3594),
.B2(n_3577),
.Y(n_4180)
);

AND2x2_ASAP7_75t_L g4181 ( 
.A(n_3938),
.B(n_3448),
.Y(n_4181)
);

AND2x2_ASAP7_75t_L g4182 ( 
.A(n_3920),
.B(n_3450),
.Y(n_4182)
);

O2A1O1Ixp33_ASAP7_75t_L g4183 ( 
.A1(n_3808),
.A2(n_3948),
.B(n_4028),
.C(n_4027),
.Y(n_4183)
);

NAND2x1p5_ASAP7_75t_L g4184 ( 
.A(n_3861),
.B(n_3545),
.Y(n_4184)
);

O2A1O1Ixp33_ASAP7_75t_SL g4185 ( 
.A1(n_3880),
.A2(n_3885),
.B(n_3838),
.C(n_3797),
.Y(n_4185)
);

O2A1O1Ixp33_ASAP7_75t_L g4186 ( 
.A1(n_4031),
.A2(n_1236),
.B(n_1238),
.C(n_1237),
.Y(n_4186)
);

HB1xp67_ASAP7_75t_L g4187 ( 
.A(n_3911),
.Y(n_4187)
);

AOI21x1_ASAP7_75t_L g4188 ( 
.A1(n_3917),
.A2(n_3735),
.B(n_3733),
.Y(n_4188)
);

INVx1_ASAP7_75t_L g4189 ( 
.A(n_3930),
.Y(n_4189)
);

NAND2xp5_ASAP7_75t_L g4190 ( 
.A(n_3968),
.B(n_3458),
.Y(n_4190)
);

OA22x2_ASAP7_75t_L g4191 ( 
.A1(n_3898),
.A2(n_924),
.B1(n_925),
.B2(n_919),
.Y(n_4191)
);

HB1xp67_ASAP7_75t_L g4192 ( 
.A(n_3940),
.Y(n_4192)
);

NAND2xp5_ASAP7_75t_SL g4193 ( 
.A(n_3960),
.B(n_3472),
.Y(n_4193)
);

NAND2xp5_ASAP7_75t_L g4194 ( 
.A(n_3869),
.B(n_3951),
.Y(n_4194)
);

AOI21xp5_ASAP7_75t_L g4195 ( 
.A1(n_3767),
.A2(n_3878),
.B(n_3876),
.Y(n_4195)
);

INVx3_ASAP7_75t_L g4196 ( 
.A(n_3919),
.Y(n_4196)
);

HB1xp67_ASAP7_75t_L g4197 ( 
.A(n_3956),
.Y(n_4197)
);

INVxp67_ASAP7_75t_L g4198 ( 
.A(n_3974),
.Y(n_4198)
);

INVx1_ASAP7_75t_SL g4199 ( 
.A(n_4034),
.Y(n_4199)
);

AOI22xp33_ASAP7_75t_L g4200 ( 
.A1(n_4005),
.A2(n_3731),
.B1(n_3477),
.B2(n_3491),
.Y(n_4200)
);

AOI21xp5_ASAP7_75t_L g4201 ( 
.A1(n_3833),
.A2(n_3965),
.B(n_3905),
.Y(n_4201)
);

OAI22xp5_ASAP7_75t_L g4202 ( 
.A1(n_4036),
.A2(n_3555),
.B1(n_3557),
.B2(n_3553),
.Y(n_4202)
);

NOR2xp33_ASAP7_75t_L g4203 ( 
.A(n_4000),
.B(n_3473),
.Y(n_4203)
);

NAND2xp5_ASAP7_75t_L g4204 ( 
.A(n_3989),
.B(n_3492),
.Y(n_4204)
);

INVx2_ASAP7_75t_L g4205 ( 
.A(n_4010),
.Y(n_4205)
);

INVx4_ASAP7_75t_L g4206 ( 
.A(n_3919),
.Y(n_4206)
);

AOI21xp5_ASAP7_75t_L g4207 ( 
.A1(n_3965),
.A2(n_3735),
.B(n_3545),
.Y(n_4207)
);

AOI21xp5_ASAP7_75t_L g4208 ( 
.A1(n_3905),
.A2(n_3523),
.B(n_3515),
.Y(n_4208)
);

NAND2xp5_ASAP7_75t_L g4209 ( 
.A(n_4029),
.B(n_3538),
.Y(n_4209)
);

NAND2xp5_ASAP7_75t_SL g4210 ( 
.A(n_4016),
.B(n_3565),
.Y(n_4210)
);

AOI21xp5_ASAP7_75t_L g4211 ( 
.A1(n_3822),
.A2(n_3604),
.B(n_3602),
.Y(n_4211)
);

NOR2xp33_ASAP7_75t_L g4212 ( 
.A(n_4001),
.B(n_3614),
.Y(n_4212)
);

NOR2xp67_ASAP7_75t_SL g4213 ( 
.A(n_3982),
.B(n_3442),
.Y(n_4213)
);

NOR2xp33_ASAP7_75t_L g4214 ( 
.A(n_4017),
.B(n_3964),
.Y(n_4214)
);

BUFx2_ASAP7_75t_L g4215 ( 
.A(n_4033),
.Y(n_4215)
);

OAI22xp5_ASAP7_75t_L g4216 ( 
.A1(n_3931),
.A2(n_3490),
.B1(n_3493),
.B2(n_3462),
.Y(n_4216)
);

AOI21xp5_ASAP7_75t_L g4217 ( 
.A1(n_3823),
.A2(n_3731),
.B(n_3490),
.Y(n_4217)
);

NOR2xp33_ASAP7_75t_L g4218 ( 
.A(n_3966),
.B(n_3462),
.Y(n_4218)
);

AOI22xp5_ASAP7_75t_L g4219 ( 
.A1(n_3922),
.A2(n_3731),
.B1(n_929),
.B2(n_933),
.Y(n_4219)
);

BUFx6f_ASAP7_75t_L g4220 ( 
.A(n_3922),
.Y(n_4220)
);

A2O1A1Ixp33_ASAP7_75t_L g4221 ( 
.A1(n_3786),
.A2(n_3517),
.B(n_3493),
.C(n_1249),
.Y(n_4221)
);

OAI22x1_ASAP7_75t_L g4222 ( 
.A1(n_3983),
.A2(n_1249),
.B1(n_1254),
.B2(n_3517),
.Y(n_4222)
);

NAND2xp5_ASAP7_75t_L g4223 ( 
.A(n_3969),
.B(n_928),
.Y(n_4223)
);

INVx2_ASAP7_75t_L g4224 ( 
.A(n_3976),
.Y(n_4224)
);

O2A1O1Ixp33_ASAP7_75t_L g4225 ( 
.A1(n_3957),
.A2(n_4021),
.B(n_4003),
.C(n_3972),
.Y(n_4225)
);

INVx5_ASAP7_75t_L g4226 ( 
.A(n_3983),
.Y(n_4226)
);

NAND2xp5_ASAP7_75t_L g4227 ( 
.A(n_3988),
.B(n_3998),
.Y(n_4227)
);

A2O1A1Ixp33_ASAP7_75t_L g4228 ( 
.A1(n_3867),
.A2(n_1254),
.B(n_1225),
.C(n_940),
.Y(n_4228)
);

INVx3_ASAP7_75t_L g4229 ( 
.A(n_4007),
.Y(n_4229)
);

CKINVDCx5p33_ASAP7_75t_R g4230 ( 
.A(n_3815),
.Y(n_4230)
);

NOR2xp67_ASAP7_75t_L g4231 ( 
.A(n_4033),
.B(n_2078),
.Y(n_4231)
);

CKINVDCx20_ASAP7_75t_R g4232 ( 
.A(n_4007),
.Y(n_4232)
);

NAND2xp5_ASAP7_75t_L g4233 ( 
.A(n_4019),
.B(n_935),
.Y(n_4233)
);

INVx2_ASAP7_75t_L g4234 ( 
.A(n_3942),
.Y(n_4234)
);

NAND2xp5_ASAP7_75t_L g4235 ( 
.A(n_3980),
.B(n_942),
.Y(n_4235)
);

AOI21x1_ASAP7_75t_L g4236 ( 
.A1(n_3927),
.A2(n_1583),
.B(n_1581),
.Y(n_4236)
);

INVx1_ASAP7_75t_L g4237 ( 
.A(n_3967),
.Y(n_4237)
);

O2A1O1Ixp33_ASAP7_75t_L g4238 ( 
.A1(n_3774),
.A2(n_1587),
.B(n_1593),
.C(n_1584),
.Y(n_4238)
);

INVx1_ASAP7_75t_L g4239 ( 
.A(n_3926),
.Y(n_4239)
);

NAND2xp5_ASAP7_75t_L g4240 ( 
.A(n_3981),
.B(n_943),
.Y(n_4240)
);

AOI21xp5_ASAP7_75t_L g4241 ( 
.A1(n_3884),
.A2(n_2102),
.B(n_2096),
.Y(n_4241)
);

AOI21xp5_ASAP7_75t_L g4242 ( 
.A1(n_3893),
.A2(n_2102),
.B(n_2096),
.Y(n_4242)
);

OAI22xp5_ASAP7_75t_L g4243 ( 
.A1(n_3860),
.A2(n_3943),
.B1(n_3944),
.B2(n_3863),
.Y(n_4243)
);

OAI21xp5_ASAP7_75t_L g4244 ( 
.A1(n_3867),
.A2(n_2120),
.B(n_2100),
.Y(n_4244)
);

AND2x2_ASAP7_75t_L g4245 ( 
.A(n_3973),
.B(n_1597),
.Y(n_4245)
);

INVx2_ASAP7_75t_L g4246 ( 
.A(n_3949),
.Y(n_4246)
);

AOI21xp5_ASAP7_75t_L g4247 ( 
.A1(n_3894),
.A2(n_2104),
.B(n_2096),
.Y(n_4247)
);

AND2x4_ASAP7_75t_L g4248 ( 
.A(n_3929),
.B(n_2186),
.Y(n_4248)
);

NAND2xp5_ASAP7_75t_SL g4249 ( 
.A(n_3773),
.B(n_3865),
.Y(n_4249)
);

NAND2xp5_ASAP7_75t_L g4250 ( 
.A(n_3971),
.B(n_945),
.Y(n_4250)
);

AOI21xp5_ASAP7_75t_L g4251 ( 
.A1(n_3778),
.A2(n_2121),
.B(n_2104),
.Y(n_4251)
);

BUFx4f_ASAP7_75t_L g4252 ( 
.A(n_3759),
.Y(n_4252)
);

NOR3xp33_ASAP7_75t_L g4253 ( 
.A(n_3763),
.B(n_1599),
.C(n_1598),
.Y(n_4253)
);

NAND2xp5_ASAP7_75t_L g4254 ( 
.A(n_3986),
.B(n_949),
.Y(n_4254)
);

INVx2_ASAP7_75t_SL g4255 ( 
.A(n_3759),
.Y(n_4255)
);

NAND2xp5_ASAP7_75t_L g4256 ( 
.A(n_3935),
.B(n_951),
.Y(n_4256)
);

AOI22xp5_ASAP7_75t_L g4257 ( 
.A1(n_4032),
.A2(n_953),
.B1(n_955),
.B2(n_952),
.Y(n_4257)
);

AOI21xp5_ASAP7_75t_L g4258 ( 
.A1(n_3864),
.A2(n_2121),
.B(n_2104),
.Y(n_4258)
);

INVx1_ASAP7_75t_L g4259 ( 
.A(n_3953),
.Y(n_4259)
);

NOR2xp33_ASAP7_75t_SL g4260 ( 
.A(n_3883),
.B(n_957),
.Y(n_4260)
);

BUFx6f_ASAP7_75t_L g4261 ( 
.A(n_3883),
.Y(n_4261)
);

AOI21xp5_ASAP7_75t_L g4262 ( 
.A1(n_3836),
.A2(n_2121),
.B(n_2104),
.Y(n_4262)
);

AOI21xp5_ASAP7_75t_L g4263 ( 
.A1(n_3843),
.A2(n_2139),
.B(n_2121),
.Y(n_4263)
);

NOR2x1_ASAP7_75t_L g4264 ( 
.A(n_3839),
.B(n_2120),
.Y(n_4264)
);

NOR2xp33_ASAP7_75t_L g4265 ( 
.A(n_3854),
.B(n_959),
.Y(n_4265)
);

INVx1_ASAP7_75t_L g4266 ( 
.A(n_3837),
.Y(n_4266)
);

INVx3_ASAP7_75t_L g4267 ( 
.A(n_4024),
.Y(n_4267)
);

NAND2xp5_ASAP7_75t_L g4268 ( 
.A(n_3909),
.B(n_961),
.Y(n_4268)
);

CKINVDCx20_ASAP7_75t_R g4269 ( 
.A(n_3839),
.Y(n_4269)
);

AND2x2_ASAP7_75t_L g4270 ( 
.A(n_3936),
.B(n_1604),
.Y(n_4270)
);

BUFx3_ASAP7_75t_L g4271 ( 
.A(n_3923),
.Y(n_4271)
);

NOR2xp33_ASAP7_75t_L g4272 ( 
.A(n_3895),
.B(n_962),
.Y(n_4272)
);

OAI22xp5_ASAP7_75t_L g4273 ( 
.A1(n_3828),
.A2(n_968),
.B1(n_970),
.B2(n_965),
.Y(n_4273)
);

NOR2xp33_ASAP7_75t_L g4274 ( 
.A(n_3979),
.B(n_972),
.Y(n_4274)
);

AOI21xp5_ASAP7_75t_L g4275 ( 
.A1(n_3805),
.A2(n_2145),
.B(n_2139),
.Y(n_4275)
);

OAI21x1_ASAP7_75t_L g4276 ( 
.A1(n_3924),
.A2(n_2478),
.B(n_2470),
.Y(n_4276)
);

INVx2_ASAP7_75t_L g4277 ( 
.A(n_3975),
.Y(n_4277)
);

AOI21xp5_ASAP7_75t_L g4278 ( 
.A1(n_3813),
.A2(n_2169),
.B(n_2153),
.Y(n_4278)
);

NAND2xp5_ASAP7_75t_L g4279 ( 
.A(n_3849),
.B(n_973),
.Y(n_4279)
);

BUFx6f_ASAP7_75t_L g4280 ( 
.A(n_4020),
.Y(n_4280)
);

BUFx4f_ASAP7_75t_L g4281 ( 
.A(n_4018),
.Y(n_4281)
);

A2O1A1Ixp33_ASAP7_75t_L g4282 ( 
.A1(n_3875),
.A2(n_977),
.B(n_979),
.C(n_975),
.Y(n_4282)
);

A2O1A1Ixp33_ASAP7_75t_L g4283 ( 
.A1(n_4030),
.A2(n_983),
.B(n_985),
.C(n_981),
.Y(n_4283)
);

NAND2xp5_ASAP7_75t_L g4284 ( 
.A(n_3850),
.B(n_988),
.Y(n_4284)
);

NAND2xp5_ASAP7_75t_L g4285 ( 
.A(n_3902),
.B(n_991),
.Y(n_4285)
);

AND2x2_ASAP7_75t_L g4286 ( 
.A(n_4022),
.B(n_1605),
.Y(n_4286)
);

AND2x2_ASAP7_75t_L g4287 ( 
.A(n_4022),
.B(n_1606),
.Y(n_4287)
);

NAND2xp5_ASAP7_75t_L g4288 ( 
.A(n_3904),
.B(n_992),
.Y(n_4288)
);

INVx1_ASAP7_75t_SL g4289 ( 
.A(n_3855),
.Y(n_4289)
);

AOI21xp5_ASAP7_75t_L g4290 ( 
.A1(n_3962),
.A2(n_2172),
.B(n_2153),
.Y(n_4290)
);

NAND2xp5_ASAP7_75t_L g4291 ( 
.A(n_3906),
.B(n_994),
.Y(n_4291)
);

OR2x2_ASAP7_75t_SL g4292 ( 
.A(n_4023),
.B(n_1609),
.Y(n_4292)
);

NAND2x1p5_ASAP7_75t_L g4293 ( 
.A(n_3866),
.B(n_2133),
.Y(n_4293)
);

NOR2x1_ASAP7_75t_L g4294 ( 
.A(n_3987),
.B(n_2133),
.Y(n_4294)
);

NAND2xp5_ASAP7_75t_L g4295 ( 
.A(n_3908),
.B(n_1000),
.Y(n_4295)
);

NAND2xp5_ASAP7_75t_SL g4296 ( 
.A(n_3925),
.B(n_1003),
.Y(n_4296)
);

NAND2xp5_ASAP7_75t_L g4297 ( 
.A(n_3910),
.B(n_1004),
.Y(n_4297)
);

AND2x2_ASAP7_75t_SL g4298 ( 
.A(n_4035),
.B(n_1610),
.Y(n_4298)
);

NOR2xp67_ASAP7_75t_L g4299 ( 
.A(n_4011),
.B(n_2142),
.Y(n_4299)
);

AOI21xp5_ASAP7_75t_L g4300 ( 
.A1(n_3994),
.A2(n_2172),
.B(n_2153),
.Y(n_4300)
);

INVx1_ASAP7_75t_L g4301 ( 
.A(n_3912),
.Y(n_4301)
);

BUFx2_ASAP7_75t_R g4302 ( 
.A(n_4113),
.Y(n_4302)
);

OAI21xp5_ASAP7_75t_L g4303 ( 
.A1(n_4138),
.A2(n_4038),
.B(n_4037),
.Y(n_4303)
);

OAI21xp5_ASAP7_75t_L g4304 ( 
.A1(n_4274),
.A2(n_3990),
.B(n_3963),
.Y(n_4304)
);

AOI21xp5_ASAP7_75t_SL g4305 ( 
.A1(n_4183),
.A2(n_4023),
.B(n_3868),
.Y(n_4305)
);

OAI21x1_ASAP7_75t_L g4306 ( 
.A1(n_4195),
.A2(n_3999),
.B(n_3995),
.Y(n_4306)
);

A2O1A1Ixp33_ASAP7_75t_L g4307 ( 
.A1(n_4046),
.A2(n_4009),
.B(n_4013),
.C(n_3959),
.Y(n_4307)
);

INVx1_ASAP7_75t_L g4308 ( 
.A(n_4187),
.Y(n_4308)
);

AOI21xp5_ASAP7_75t_L g4309 ( 
.A1(n_4201),
.A2(n_3958),
.B(n_3873),
.Y(n_4309)
);

NAND2xp5_ASAP7_75t_L g4310 ( 
.A(n_4122),
.B(n_1014),
.Y(n_4310)
);

NAND2xp5_ASAP7_75t_L g4311 ( 
.A(n_4040),
.B(n_1015),
.Y(n_4311)
);

NAND2xp5_ASAP7_75t_SL g4312 ( 
.A(n_4050),
.B(n_4012),
.Y(n_4312)
);

OR2x2_ASAP7_75t_L g4313 ( 
.A(n_4055),
.B(n_1611),
.Y(n_4313)
);

NAND2xp5_ASAP7_75t_L g4314 ( 
.A(n_4049),
.B(n_1017),
.Y(n_4314)
);

NAND2xp5_ASAP7_75t_L g4315 ( 
.A(n_4103),
.B(n_4063),
.Y(n_4315)
);

HB1xp67_ASAP7_75t_L g4316 ( 
.A(n_4074),
.Y(n_4316)
);

OAI211xp5_ASAP7_75t_SL g4317 ( 
.A1(n_4057),
.A2(n_1616),
.B(n_1618),
.C(n_1613),
.Y(n_4317)
);

NAND2xp5_ASAP7_75t_SL g4318 ( 
.A(n_4047),
.B(n_4015),
.Y(n_4318)
);

OAI21x1_ASAP7_75t_L g4319 ( 
.A1(n_4276),
.A2(n_3915),
.B(n_3913),
.Y(n_4319)
);

NAND2x1p5_ASAP7_75t_L g4320 ( 
.A(n_4041),
.B(n_4004),
.Y(n_4320)
);

NAND2xp5_ASAP7_75t_L g4321 ( 
.A(n_4065),
.B(n_1019),
.Y(n_4321)
);

OAI21xp5_ASAP7_75t_L g4322 ( 
.A1(n_4128),
.A2(n_3871),
.B(n_3945),
.Y(n_4322)
);

NAND2xp5_ASAP7_75t_L g4323 ( 
.A(n_4048),
.B(n_1020),
.Y(n_4323)
);

AOI21xp5_ASAP7_75t_L g4324 ( 
.A1(n_4059),
.A2(n_3946),
.B(n_4006),
.Y(n_4324)
);

NAND2x1_ASAP7_75t_L g4325 ( 
.A(n_4267),
.B(n_2470),
.Y(n_4325)
);

OAI21x1_ASAP7_75t_L g4326 ( 
.A1(n_4217),
.A2(n_4116),
.B(n_4251),
.Y(n_4326)
);

INVx2_ASAP7_75t_L g4327 ( 
.A(n_4224),
.Y(n_4327)
);

AO31x2_ASAP7_75t_L g4328 ( 
.A1(n_4148),
.A2(n_1622),
.A3(n_1624),
.B(n_1620),
.Y(n_4328)
);

AOI21xp5_ASAP7_75t_L g4329 ( 
.A1(n_4060),
.A2(n_2478),
.B(n_2179),
.Y(n_4329)
);

NOR2x1_ASAP7_75t_SL g4330 ( 
.A(n_4249),
.B(n_1625),
.Y(n_4330)
);

AOI21xp5_ASAP7_75t_L g4331 ( 
.A1(n_4091),
.A2(n_2179),
.B(n_2172),
.Y(n_4331)
);

INVx2_ASAP7_75t_L g4332 ( 
.A(n_4044),
.Y(n_4332)
);

A2O1A1Ixp33_ASAP7_75t_L g4333 ( 
.A1(n_4053),
.A2(n_1633),
.B(n_1635),
.C(n_1631),
.Y(n_4333)
);

AOI21xp5_ASAP7_75t_L g4334 ( 
.A1(n_4134),
.A2(n_2179),
.B(n_2172),
.Y(n_4334)
);

CKINVDCx6p67_ASAP7_75t_R g4335 ( 
.A(n_4075),
.Y(n_4335)
);

AO31x2_ASAP7_75t_L g4336 ( 
.A1(n_4266),
.A2(n_1642),
.A3(n_1643),
.B(n_1637),
.Y(n_4336)
);

NAND2xp5_ASAP7_75t_SL g4337 ( 
.A(n_4107),
.B(n_1644),
.Y(n_4337)
);

INVxp67_ASAP7_75t_L g4338 ( 
.A(n_4054),
.Y(n_4338)
);

INVx2_ASAP7_75t_SL g4339 ( 
.A(n_4045),
.Y(n_4339)
);

BUFx4f_ASAP7_75t_L g4340 ( 
.A(n_4043),
.Y(n_4340)
);

OAI21x1_ASAP7_75t_L g4341 ( 
.A1(n_4236),
.A2(n_2147),
.B(n_2142),
.Y(n_4341)
);

AO31x2_ASAP7_75t_L g4342 ( 
.A1(n_4056),
.A2(n_1648),
.A3(n_1649),
.B(n_1646),
.Y(n_4342)
);

OAI22xp5_ASAP7_75t_L g4343 ( 
.A1(n_4269),
.A2(n_1023),
.B1(n_1026),
.B2(n_1022),
.Y(n_4343)
);

OAI21x1_ASAP7_75t_L g4344 ( 
.A1(n_4275),
.A2(n_2186),
.B(n_2147),
.Y(n_4344)
);

NOR2x1_ASAP7_75t_SL g4345 ( 
.A(n_4277),
.B(n_1652),
.Y(n_4345)
);

OAI21xp5_ASAP7_75t_SL g4346 ( 
.A1(n_4167),
.A2(n_1655),
.B(n_1654),
.Y(n_4346)
);

NAND2xp5_ASAP7_75t_L g4347 ( 
.A(n_4194),
.B(n_1031),
.Y(n_4347)
);

AND2x2_ASAP7_75t_L g4348 ( 
.A(n_4150),
.B(n_1656),
.Y(n_4348)
);

NAND2xp5_ASAP7_75t_L g4349 ( 
.A(n_4237),
.B(n_1037),
.Y(n_4349)
);

OR2x2_ASAP7_75t_L g4350 ( 
.A(n_4192),
.B(n_1657),
.Y(n_4350)
);

AND2x2_ASAP7_75t_L g4351 ( 
.A(n_4067),
.B(n_1658),
.Y(n_4351)
);

AO31x2_ASAP7_75t_L g4352 ( 
.A1(n_4301),
.A2(n_1661),
.A3(n_1662),
.B(n_1660),
.Y(n_4352)
);

NAND2xp5_ASAP7_75t_L g4353 ( 
.A(n_4082),
.B(n_1039),
.Y(n_4353)
);

INVx5_ASAP7_75t_L g4354 ( 
.A(n_4041),
.Y(n_4354)
);

OAI22xp5_ASAP7_75t_L g4355 ( 
.A1(n_4077),
.A2(n_4052),
.B1(n_4179),
.B2(n_4062),
.Y(n_4355)
);

NAND2xp5_ASAP7_75t_L g4356 ( 
.A(n_4089),
.B(n_1042),
.Y(n_4356)
);

AND2x2_ASAP7_75t_L g4357 ( 
.A(n_4199),
.B(n_1663),
.Y(n_4357)
);

NAND2xp5_ASAP7_75t_L g4358 ( 
.A(n_4135),
.B(n_1044),
.Y(n_4358)
);

OAI21x1_ASAP7_75t_L g4359 ( 
.A1(n_4102),
.A2(n_2261),
.B(n_2199),
.Y(n_4359)
);

INVx4_ASAP7_75t_L g4360 ( 
.A(n_4084),
.Y(n_4360)
);

OAI22xp5_ASAP7_75t_L g4361 ( 
.A1(n_4104),
.A2(n_1047),
.B1(n_1050),
.B2(n_1045),
.Y(n_4361)
);

OAI21xp5_ASAP7_75t_L g4362 ( 
.A1(n_4228),
.A2(n_1668),
.B(n_1664),
.Y(n_4362)
);

NAND2xp5_ASAP7_75t_L g4363 ( 
.A(n_4127),
.B(n_1057),
.Y(n_4363)
);

NAND2xp5_ASAP7_75t_L g4364 ( 
.A(n_4099),
.B(n_1058),
.Y(n_4364)
);

OAI22xp5_ASAP7_75t_L g4365 ( 
.A1(n_4039),
.A2(n_4094),
.B1(n_4042),
.B2(n_4070),
.Y(n_4365)
);

AOI21xp5_ASAP7_75t_L g4366 ( 
.A1(n_4281),
.A2(n_2190),
.B(n_2179),
.Y(n_4366)
);

OAI21xp5_ASAP7_75t_L g4367 ( 
.A1(n_4085),
.A2(n_1671),
.B(n_1669),
.Y(n_4367)
);

BUFx8_ASAP7_75t_SL g4368 ( 
.A(n_4230),
.Y(n_4368)
);

BUFx6f_ASAP7_75t_L g4369 ( 
.A(n_4143),
.Y(n_4369)
);

AOI21xp5_ASAP7_75t_L g4370 ( 
.A1(n_4281),
.A2(n_4073),
.B(n_4142),
.Y(n_4370)
);

AO31x2_ASAP7_75t_L g4371 ( 
.A1(n_4115),
.A2(n_1675),
.A3(n_1676),
.B(n_1672),
.Y(n_4371)
);

NAND2xp5_ASAP7_75t_L g4372 ( 
.A(n_4125),
.B(n_1061),
.Y(n_4372)
);

NAND2xp5_ASAP7_75t_SL g4373 ( 
.A(n_4058),
.B(n_1679),
.Y(n_4373)
);

AOI21xp5_ASAP7_75t_L g4374 ( 
.A1(n_4164),
.A2(n_2254),
.B(n_2196),
.Y(n_4374)
);

OAI21xp33_ASAP7_75t_L g4375 ( 
.A1(n_4137),
.A2(n_1066),
.B(n_1065),
.Y(n_4375)
);

AOI21xp5_ASAP7_75t_L g4376 ( 
.A1(n_4168),
.A2(n_2254),
.B(n_2196),
.Y(n_4376)
);

AOI22xp5_ASAP7_75t_L g4377 ( 
.A1(n_4191),
.A2(n_1077),
.B1(n_1078),
.B2(n_1076),
.Y(n_4377)
);

OAI21x1_ASAP7_75t_L g4378 ( 
.A1(n_4124),
.A2(n_2261),
.B(n_2199),
.Y(n_4378)
);

OAI21xp5_ASAP7_75t_L g4379 ( 
.A1(n_4282),
.A2(n_1698),
.B(n_1693),
.Y(n_4379)
);

INVx3_ASAP7_75t_L g4380 ( 
.A(n_4105),
.Y(n_4380)
);

OAI22xp5_ASAP7_75t_L g4381 ( 
.A1(n_4146),
.A2(n_1083),
.B1(n_1084),
.B2(n_1080),
.Y(n_4381)
);

AOI21xp5_ASAP7_75t_L g4382 ( 
.A1(n_4176),
.A2(n_2267),
.B(n_2254),
.Y(n_4382)
);

OAI21x1_ASAP7_75t_L g4383 ( 
.A1(n_4126),
.A2(n_2273),
.B(n_2262),
.Y(n_4383)
);

NAND2xp5_ASAP7_75t_L g4384 ( 
.A(n_4214),
.B(n_1085),
.Y(n_4384)
);

AO31x2_ASAP7_75t_L g4385 ( 
.A1(n_4221),
.A2(n_1700),
.A3(n_1968),
.B(n_1811),
.Y(n_4385)
);

AOI221x1_ASAP7_75t_L g4386 ( 
.A1(n_4092),
.A2(n_2290),
.B1(n_2312),
.B2(n_2273),
.C(n_2262),
.Y(n_4386)
);

NAND2xp5_ASAP7_75t_L g4387 ( 
.A(n_4190),
.B(n_1086),
.Y(n_4387)
);

INVx1_ASAP7_75t_L g4388 ( 
.A(n_4197),
.Y(n_4388)
);

INVxp67_ASAP7_75t_SL g4389 ( 
.A(n_4271),
.Y(n_4389)
);

NAND3xp33_ASAP7_75t_L g4390 ( 
.A(n_4147),
.B(n_1088),
.C(n_1087),
.Y(n_4390)
);

AND2x2_ASAP7_75t_L g4391 ( 
.A(n_4071),
.B(n_600),
.Y(n_4391)
);

AOI21xp5_ASAP7_75t_L g4392 ( 
.A1(n_4136),
.A2(n_2271),
.B(n_2267),
.Y(n_4392)
);

OA21x2_ASAP7_75t_L g4393 ( 
.A1(n_4169),
.A2(n_1093),
.B(n_1089),
.Y(n_4393)
);

OAI21x1_ASAP7_75t_L g4394 ( 
.A1(n_4290),
.A2(n_2312),
.B(n_2290),
.Y(n_4394)
);

OAI21xp5_ASAP7_75t_L g4395 ( 
.A1(n_4285),
.A2(n_1096),
.B(n_1095),
.Y(n_4395)
);

INVx3_ASAP7_75t_L g4396 ( 
.A(n_4097),
.Y(n_4396)
);

BUFx6f_ASAP7_75t_L g4397 ( 
.A(n_4143),
.Y(n_4397)
);

O2A1O1Ixp5_ASAP7_75t_L g4398 ( 
.A1(n_4130),
.A2(n_2389),
.B(n_2394),
.C(n_2370),
.Y(n_4398)
);

AO31x2_ASAP7_75t_L g4399 ( 
.A1(n_4207),
.A2(n_1968),
.A3(n_1811),
.B(n_1788),
.Y(n_4399)
);

AND2x4_ASAP7_75t_L g4400 ( 
.A(n_4232),
.B(n_2370),
.Y(n_4400)
);

OAI21x1_ASAP7_75t_L g4401 ( 
.A1(n_4300),
.A2(n_2394),
.B(n_2389),
.Y(n_4401)
);

INVx1_ASAP7_75t_L g4402 ( 
.A(n_4068),
.Y(n_4402)
);

OAI21xp5_ASAP7_75t_L g4403 ( 
.A1(n_4295),
.A2(n_1104),
.B(n_1100),
.Y(n_4403)
);

AOI21xp5_ASAP7_75t_L g4404 ( 
.A1(n_4118),
.A2(n_2271),
.B(n_2267),
.Y(n_4404)
);

NAND2xp5_ASAP7_75t_L g4405 ( 
.A(n_4159),
.B(n_1109),
.Y(n_4405)
);

OA21x2_ASAP7_75t_L g4406 ( 
.A1(n_4177),
.A2(n_1111),
.B(n_1110),
.Y(n_4406)
);

OAI21x1_ASAP7_75t_L g4407 ( 
.A1(n_4241),
.A2(n_2417),
.B(n_2416),
.Y(n_4407)
);

OAI21x1_ASAP7_75t_L g4408 ( 
.A1(n_4242),
.A2(n_2417),
.B(n_2416),
.Y(n_4408)
);

OAI21x1_ASAP7_75t_L g4409 ( 
.A1(n_4247),
.A2(n_2442),
.B(n_1848),
.Y(n_4409)
);

AOI21xp5_ASAP7_75t_L g4410 ( 
.A1(n_4185),
.A2(n_2271),
.B(n_2267),
.Y(n_4410)
);

AND2x2_ASAP7_75t_L g4411 ( 
.A(n_4173),
.B(n_4181),
.Y(n_4411)
);

NAND2xp5_ASAP7_75t_SL g4412 ( 
.A(n_4108),
.B(n_1114),
.Y(n_4412)
);

AOI21xp5_ASAP7_75t_L g4413 ( 
.A1(n_4252),
.A2(n_2276),
.B(n_2271),
.Y(n_4413)
);

OAI21x1_ASAP7_75t_L g4414 ( 
.A1(n_4188),
.A2(n_2442),
.B(n_1848),
.Y(n_4414)
);

INVx1_ASAP7_75t_L g4415 ( 
.A(n_4072),
.Y(n_4415)
);

OAI21x1_ASAP7_75t_L g4416 ( 
.A1(n_4211),
.A2(n_1863),
.B(n_1835),
.Y(n_4416)
);

OAI21xp5_ASAP7_75t_L g4417 ( 
.A1(n_4272),
.A2(n_1117),
.B(n_1116),
.Y(n_4417)
);

OAI21x1_ASAP7_75t_L g4418 ( 
.A1(n_4278),
.A2(n_1863),
.B(n_1835),
.Y(n_4418)
);

AOI31xp67_ASAP7_75t_L g4419 ( 
.A1(n_4100),
.A2(n_1968),
.A3(n_1839),
.B(n_1852),
.Y(n_4419)
);

OAI21x1_ASAP7_75t_L g4420 ( 
.A1(n_4208),
.A2(n_1851),
.B(n_1839),
.Y(n_4420)
);

AOI21xp33_ASAP7_75t_L g4421 ( 
.A1(n_4288),
.A2(n_4291),
.B(n_4284),
.Y(n_4421)
);

OAI21x1_ASAP7_75t_L g4422 ( 
.A1(n_4262),
.A2(n_4263),
.B(n_4267),
.Y(n_4422)
);

OAI21xp5_ASAP7_75t_L g4423 ( 
.A1(n_4279),
.A2(n_1123),
.B(n_1121),
.Y(n_4423)
);

OAI21x1_ASAP7_75t_L g4424 ( 
.A1(n_4258),
.A2(n_1851),
.B(n_1839),
.Y(n_4424)
);

OAI21x1_ASAP7_75t_L g4425 ( 
.A1(n_4293),
.A2(n_1852),
.B(n_1851),
.Y(n_4425)
);

OA22x2_ASAP7_75t_L g4426 ( 
.A1(n_4222),
.A2(n_1127),
.B1(n_1128),
.B2(n_1126),
.Y(n_4426)
);

BUFx2_ASAP7_75t_L g4427 ( 
.A(n_4064),
.Y(n_4427)
);

OAI21x1_ASAP7_75t_L g4428 ( 
.A1(n_4264),
.A2(n_1854),
.B(n_1852),
.Y(n_4428)
);

OAI21x1_ASAP7_75t_SL g4429 ( 
.A1(n_4088),
.A2(n_4),
.B(n_5),
.Y(n_4429)
);

AOI21xp5_ASAP7_75t_L g4430 ( 
.A1(n_4252),
.A2(n_2285),
.B(n_2276),
.Y(n_4430)
);

NOR2x1p5_ASAP7_75t_L g4431 ( 
.A(n_4097),
.B(n_1129),
.Y(n_4431)
);

INVx2_ASAP7_75t_L g4432 ( 
.A(n_4087),
.Y(n_4432)
);

A2O1A1Ixp33_ASAP7_75t_L g4433 ( 
.A1(n_4225),
.A2(n_1163),
.B(n_1193),
.C(n_1141),
.Y(n_4433)
);

NAND2xp5_ASAP7_75t_L g4434 ( 
.A(n_4145),
.B(n_1130),
.Y(n_4434)
);

OA21x2_ASAP7_75t_L g4435 ( 
.A1(n_4061),
.A2(n_1135),
.B(n_1131),
.Y(n_4435)
);

NOR2xp33_ASAP7_75t_L g4436 ( 
.A(n_4051),
.B(n_4132),
.Y(n_4436)
);

OAI21x1_ASAP7_75t_L g4437 ( 
.A1(n_4294),
.A2(n_1857),
.B(n_1854),
.Y(n_4437)
);

INVx3_ASAP7_75t_L g4438 ( 
.A(n_4120),
.Y(n_4438)
);

NAND2xp5_ASAP7_75t_SL g4439 ( 
.A(n_4079),
.B(n_4086),
.Y(n_4439)
);

CKINVDCx5p33_ASAP7_75t_R g4440 ( 
.A(n_4066),
.Y(n_4440)
);

NAND2xp5_ASAP7_75t_L g4441 ( 
.A(n_4110),
.B(n_1137),
.Y(n_4441)
);

AOI21x1_ASAP7_75t_L g4442 ( 
.A1(n_4299),
.A2(n_2285),
.B(n_2276),
.Y(n_4442)
);

INVx2_ASAP7_75t_L g4443 ( 
.A(n_4112),
.Y(n_4443)
);

NOR2xp67_ASAP7_75t_L g4444 ( 
.A(n_4198),
.B(n_4171),
.Y(n_4444)
);

AO31x2_ASAP7_75t_L g4445 ( 
.A1(n_4243),
.A2(n_1968),
.A3(n_1811),
.B(n_605),
.Y(n_4445)
);

OAI21x1_ASAP7_75t_L g4446 ( 
.A1(n_4244),
.A2(n_1857),
.B(n_1854),
.Y(n_4446)
);

OAI21x1_ASAP7_75t_L g4447 ( 
.A1(n_4200),
.A2(n_1861),
.B(n_1857),
.Y(n_4447)
);

OR2x6_ASAP7_75t_L g4448 ( 
.A(n_4095),
.B(n_1861),
.Y(n_4448)
);

INVx2_ASAP7_75t_SL g4449 ( 
.A(n_4120),
.Y(n_4449)
);

OAI21xp5_ASAP7_75t_L g4450 ( 
.A1(n_4297),
.A2(n_1140),
.B(n_1139),
.Y(n_4450)
);

OAI21x1_ASAP7_75t_L g4451 ( 
.A1(n_4196),
.A2(n_4229),
.B(n_4149),
.Y(n_4451)
);

NAND3xp33_ASAP7_75t_SL g4452 ( 
.A(n_4265),
.B(n_1150),
.C(n_1147),
.Y(n_4452)
);

NAND2xp5_ASAP7_75t_L g4453 ( 
.A(n_4163),
.B(n_1155),
.Y(n_4453)
);

OAI21x1_ASAP7_75t_L g4454 ( 
.A1(n_4196),
.A2(n_1871),
.B(n_1861),
.Y(n_4454)
);

NAND2xp5_ASAP7_75t_L g4455 ( 
.A(n_4121),
.B(n_1157),
.Y(n_4455)
);

OAI21xp5_ASAP7_75t_L g4456 ( 
.A1(n_4283),
.A2(n_1159),
.B(n_1158),
.Y(n_4456)
);

AO31x2_ASAP7_75t_L g4457 ( 
.A1(n_4157),
.A2(n_1968),
.A3(n_1811),
.B(n_607),
.Y(n_4457)
);

AOI21xp5_ASAP7_75t_L g4458 ( 
.A1(n_4093),
.A2(n_2285),
.B(n_2276),
.Y(n_4458)
);

CKINVDCx5p33_ASAP7_75t_R g4459 ( 
.A(n_4076),
.Y(n_4459)
);

NAND2xp5_ASAP7_75t_L g4460 ( 
.A(n_4081),
.B(n_1162),
.Y(n_4460)
);

OAI21x1_ASAP7_75t_L g4461 ( 
.A1(n_4229),
.A2(n_4210),
.B(n_4141),
.Y(n_4461)
);

AOI22xp5_ASAP7_75t_L g4462 ( 
.A1(n_4083),
.A2(n_1169),
.B1(n_1173),
.B2(n_1167),
.Y(n_4462)
);

BUFx6f_ASAP7_75t_L g4463 ( 
.A(n_4143),
.Y(n_4463)
);

INVx3_ASAP7_75t_SL g4464 ( 
.A(n_4120),
.Y(n_4464)
);

HB1xp67_ASAP7_75t_L g4465 ( 
.A(n_4109),
.Y(n_4465)
);

NOR2xp33_ASAP7_75t_SL g4466 ( 
.A(n_4162),
.B(n_1175),
.Y(n_4466)
);

AOI21xp5_ASAP7_75t_L g4467 ( 
.A1(n_4129),
.A2(n_2318),
.B(n_2300),
.Y(n_4467)
);

AOI21xp5_ASAP7_75t_L g4468 ( 
.A1(n_4298),
.A2(n_2318),
.B(n_2300),
.Y(n_4468)
);

NOR2x1_ASAP7_75t_SL g4469 ( 
.A(n_4226),
.B(n_4261),
.Y(n_4469)
);

OAI22xp5_ASAP7_75t_L g4470 ( 
.A1(n_4292),
.A2(n_1179),
.B1(n_1187),
.B2(n_1176),
.Y(n_4470)
);

NAND2xp5_ASAP7_75t_SL g4471 ( 
.A(n_4260),
.B(n_1194),
.Y(n_4471)
);

NAND3xp33_ASAP7_75t_L g4472 ( 
.A(n_4273),
.B(n_1209),
.C(n_1204),
.Y(n_4472)
);

OA22x2_ASAP7_75t_L g4473 ( 
.A1(n_4080),
.A2(n_1215),
.B1(n_1218),
.B2(n_1213),
.Y(n_4473)
);

AOI211x1_ASAP7_75t_L g4474 ( 
.A1(n_4227),
.A2(n_1222),
.B(n_1223),
.C(n_1219),
.Y(n_4474)
);

INVx3_ASAP7_75t_L g4475 ( 
.A(n_4161),
.Y(n_4475)
);

AOI21xp5_ASAP7_75t_L g4476 ( 
.A1(n_4289),
.A2(n_2333),
.B(n_2318),
.Y(n_4476)
);

O2A1O1Ixp5_ASAP7_75t_SL g4477 ( 
.A1(n_4101),
.A2(n_1228),
.B(n_1229),
.C(n_1226),
.Y(n_4477)
);

A2O1A1Ixp33_ASAP7_75t_L g4478 ( 
.A1(n_4069),
.A2(n_1251),
.B(n_1233),
.C(n_1240),
.Y(n_4478)
);

INVx2_ASAP7_75t_L g4479 ( 
.A(n_4155),
.Y(n_4479)
);

AOI21xp5_ASAP7_75t_L g4480 ( 
.A1(n_4151),
.A2(n_2333),
.B(n_2318),
.Y(n_4480)
);

BUFx6f_ASAP7_75t_L g4481 ( 
.A(n_4161),
.Y(n_4481)
);

INVx8_ASAP7_75t_L g4482 ( 
.A(n_4095),
.Y(n_4482)
);

AND2x4_ASAP7_75t_L g4483 ( 
.A(n_4226),
.B(n_602),
.Y(n_4483)
);

AOI21xp5_ASAP7_75t_L g4484 ( 
.A1(n_4286),
.A2(n_2356),
.B(n_2333),
.Y(n_4484)
);

AO22x2_ASAP7_75t_L g4485 ( 
.A1(n_4131),
.A2(n_8),
.B1(n_6),
.B2(n_7),
.Y(n_4485)
);

NAND2xp5_ASAP7_75t_L g4486 ( 
.A(n_4239),
.B(n_1234),
.Y(n_4486)
);

NOR2xp33_ASAP7_75t_L g4487 ( 
.A(n_4117),
.B(n_1242),
.Y(n_4487)
);

AOI21xp5_ASAP7_75t_SL g4488 ( 
.A1(n_4178),
.A2(n_1244),
.B(n_1243),
.Y(n_4488)
);

NAND2xp5_ASAP7_75t_L g4489 ( 
.A(n_4259),
.B(n_1248),
.Y(n_4489)
);

AOI21xp5_ASAP7_75t_L g4490 ( 
.A1(n_4287),
.A2(n_2356),
.B(n_2333),
.Y(n_4490)
);

NOR2xp33_ASAP7_75t_L g4491 ( 
.A(n_4133),
.B(n_4123),
.Y(n_4491)
);

OAI22xp5_ASAP7_75t_L g4492 ( 
.A1(n_4098),
.A2(n_1252),
.B1(n_1250),
.B2(n_2356),
.Y(n_4492)
);

INVx3_ASAP7_75t_L g4493 ( 
.A(n_4161),
.Y(n_4493)
);

AOI21xp5_ASAP7_75t_L g4494 ( 
.A1(n_4165),
.A2(n_2373),
.B(n_2356),
.Y(n_4494)
);

O2A1O1Ixp5_ASAP7_75t_L g4495 ( 
.A1(n_4213),
.A2(n_10),
.B(n_6),
.C(n_9),
.Y(n_4495)
);

NAND2xp5_ASAP7_75t_SL g4496 ( 
.A(n_4220),
.B(n_1871),
.Y(n_4496)
);

AOI21xp5_ASAP7_75t_L g4497 ( 
.A1(n_4152),
.A2(n_2410),
.B(n_2373),
.Y(n_4497)
);

AOI21x1_ASAP7_75t_L g4498 ( 
.A1(n_4270),
.A2(n_2410),
.B(n_2373),
.Y(n_4498)
);

AND2x2_ASAP7_75t_L g4499 ( 
.A(n_4182),
.B(n_4160),
.Y(n_4499)
);

AOI22xp5_ASAP7_75t_L g4500 ( 
.A1(n_4111),
.A2(n_2041),
.B1(n_2047),
.B2(n_2027),
.Y(n_4500)
);

AO31x2_ASAP7_75t_L g4501 ( 
.A1(n_4206),
.A2(n_610),
.A3(n_612),
.B(n_608),
.Y(n_4501)
);

NAND2xp5_ASAP7_75t_L g4502 ( 
.A(n_4245),
.B(n_9),
.Y(n_4502)
);

CKINVDCx5p33_ASAP7_75t_R g4503 ( 
.A(n_4215),
.Y(n_4503)
);

NAND2xp5_ASAP7_75t_L g4504 ( 
.A(n_4205),
.B(n_10),
.Y(n_4504)
);

OAI21x1_ASAP7_75t_SL g4505 ( 
.A1(n_4206),
.A2(n_11),
.B(n_12),
.Y(n_4505)
);

OAI21xp5_ASAP7_75t_L g4506 ( 
.A1(n_4090),
.A2(n_2041),
.B(n_2027),
.Y(n_4506)
);

OAI21x1_ASAP7_75t_L g4507 ( 
.A1(n_4234),
.A2(n_1872),
.B(n_1871),
.Y(n_4507)
);

AOI21xp33_ASAP7_75t_L g4508 ( 
.A1(n_4296),
.A2(n_1872),
.B(n_2373),
.Y(n_4508)
);

OAI21x1_ASAP7_75t_L g4509 ( 
.A1(n_4246),
.A2(n_1872),
.B(n_2410),
.Y(n_4509)
);

AOI221x1_ASAP7_75t_L g4510 ( 
.A1(n_4253),
.A2(n_2437),
.B1(n_2444),
.B2(n_2435),
.C(n_2410),
.Y(n_4510)
);

INVx2_ASAP7_75t_L g4511 ( 
.A(n_4106),
.Y(n_4511)
);

OAI21xp5_ASAP7_75t_L g4512 ( 
.A1(n_4250),
.A2(n_2041),
.B(n_2027),
.Y(n_4512)
);

HB1xp67_ASAP7_75t_L g4513 ( 
.A(n_4144),
.Y(n_4513)
);

AOI221x1_ASAP7_75t_L g4514 ( 
.A1(n_4216),
.A2(n_2444),
.B1(n_2458),
.B2(n_2437),
.C(n_2435),
.Y(n_4514)
);

AOI22xp5_ASAP7_75t_L g4515 ( 
.A1(n_4174),
.A2(n_2041),
.B1(n_2047),
.B2(n_2027),
.Y(n_4515)
);

NAND2xp5_ASAP7_75t_L g4516 ( 
.A(n_4268),
.B(n_13),
.Y(n_4516)
);

OAI21xp5_ASAP7_75t_L g4517 ( 
.A1(n_4235),
.A2(n_4240),
.B(n_4254),
.Y(n_4517)
);

INVx1_ASAP7_75t_L g4518 ( 
.A(n_4158),
.Y(n_4518)
);

INVx2_ASAP7_75t_L g4519 ( 
.A(n_4166),
.Y(n_4519)
);

OAI21x1_ASAP7_75t_L g4520 ( 
.A1(n_4180),
.A2(n_2437),
.B(n_2435),
.Y(n_4520)
);

INVx1_ASAP7_75t_L g4521 ( 
.A(n_4175),
.Y(n_4521)
);

NOR2xp33_ASAP7_75t_SL g4522 ( 
.A(n_4162),
.B(n_2047),
.Y(n_4522)
);

OA21x2_ASAP7_75t_L g4523 ( 
.A1(n_4189),
.A2(n_2437),
.B(n_2435),
.Y(n_4523)
);

AOI21xp5_ASAP7_75t_L g4524 ( 
.A1(n_4152),
.A2(n_2458),
.B(n_2444),
.Y(n_4524)
);

INVx1_ASAP7_75t_L g4525 ( 
.A(n_4204),
.Y(n_4525)
);

NAND2x1p5_ASAP7_75t_L g4526 ( 
.A(n_4153),
.B(n_2444),
.Y(n_4526)
);

BUFx3_ASAP7_75t_L g4527 ( 
.A(n_4170),
.Y(n_4527)
);

INVx3_ASAP7_75t_L g4528 ( 
.A(n_4170),
.Y(n_4528)
);

INVx1_ASAP7_75t_L g4529 ( 
.A(n_4209),
.Y(n_4529)
);

OAI21x1_ASAP7_75t_L g4530 ( 
.A1(n_4238),
.A2(n_2460),
.B(n_2458),
.Y(n_4530)
);

NAND2xp5_ASAP7_75t_L g4531 ( 
.A(n_4203),
.B(n_15),
.Y(n_4531)
);

OAI21x1_ASAP7_75t_L g4532 ( 
.A1(n_4193),
.A2(n_4202),
.B(n_4219),
.Y(n_4532)
);

OAI21x1_ASAP7_75t_L g4533 ( 
.A1(n_4184),
.A2(n_4156),
.B(n_4172),
.Y(n_4533)
);

OAI21x1_ASAP7_75t_L g4534 ( 
.A1(n_4114),
.A2(n_2460),
.B(n_2458),
.Y(n_4534)
);

BUFx2_ASAP7_75t_L g4535 ( 
.A(n_4098),
.Y(n_4535)
);

OAI21x1_ASAP7_75t_L g4536 ( 
.A1(n_4186),
.A2(n_2460),
.B(n_615),
.Y(n_4536)
);

OAI21x1_ASAP7_75t_L g4537 ( 
.A1(n_4218),
.A2(n_2460),
.B(n_617),
.Y(n_4537)
);

INVx4_ASAP7_75t_L g4538 ( 
.A(n_4170),
.Y(n_4538)
);

INVx3_ASAP7_75t_L g4539 ( 
.A(n_4220),
.Y(n_4539)
);

AND2x2_ASAP7_75t_L g4540 ( 
.A(n_4212),
.B(n_613),
.Y(n_4540)
);

OA22x2_ASAP7_75t_L g4541 ( 
.A1(n_4257),
.A2(n_19),
.B1(n_16),
.B2(n_18),
.Y(n_4541)
);

INVx2_ASAP7_75t_L g4542 ( 
.A(n_4220),
.Y(n_4542)
);

INVx6_ASAP7_75t_L g4543 ( 
.A(n_4096),
.Y(n_4543)
);

NAND2xp5_ASAP7_75t_L g4544 ( 
.A(n_4256),
.B(n_16),
.Y(n_4544)
);

OR2x6_ASAP7_75t_L g4545 ( 
.A(n_4261),
.B(n_4153),
.Y(n_4545)
);

NAND2xp5_ASAP7_75t_L g4546 ( 
.A(n_4223),
.B(n_19),
.Y(n_4546)
);

BUFx3_ASAP7_75t_L g4547 ( 
.A(n_4096),
.Y(n_4547)
);

NAND2xp5_ASAP7_75t_L g4548 ( 
.A(n_4233),
.B(n_20),
.Y(n_4548)
);

OAI21xp33_ASAP7_75t_L g4549 ( 
.A1(n_4078),
.A2(n_21),
.B(n_22),
.Y(n_4549)
);

OAI21x1_ASAP7_75t_L g4550 ( 
.A1(n_4280),
.A2(n_620),
.B(n_618),
.Y(n_4550)
);

NAND2xp5_ASAP7_75t_L g4551 ( 
.A(n_4139),
.B(n_22),
.Y(n_4551)
);

OAI21x1_ASAP7_75t_L g4552 ( 
.A1(n_4280),
.A2(n_4154),
.B(n_4140),
.Y(n_4552)
);

AO32x2_ASAP7_75t_L g4553 ( 
.A1(n_4255),
.A2(n_26),
.A3(n_23),
.B1(n_25),
.B2(n_27),
.Y(n_4553)
);

A2O1A1Ixp33_ASAP7_75t_L g4554 ( 
.A1(n_4231),
.A2(n_28),
.B(n_23),
.C(n_27),
.Y(n_4554)
);

NAND2xp5_ASAP7_75t_L g4555 ( 
.A(n_4139),
.B(n_28),
.Y(n_4555)
);

BUFx2_ASAP7_75t_L g4556 ( 
.A(n_4261),
.Y(n_4556)
);

INVx1_ASAP7_75t_L g4557 ( 
.A(n_4226),
.Y(n_4557)
);

CKINVDCx5p33_ASAP7_75t_R g4558 ( 
.A(n_4368),
.Y(n_4558)
);

NAND2xp5_ASAP7_75t_L g4559 ( 
.A(n_4315),
.B(n_4248),
.Y(n_4559)
);

OAI22xp5_ASAP7_75t_L g4560 ( 
.A1(n_4436),
.A2(n_4119),
.B1(n_4248),
.B2(n_4280),
.Y(n_4560)
);

NAND2xp5_ASAP7_75t_L g4561 ( 
.A(n_4316),
.B(n_4389),
.Y(n_4561)
);

INVx1_ASAP7_75t_SL g4562 ( 
.A(n_4459),
.Y(n_4562)
);

AND2x2_ASAP7_75t_L g4563 ( 
.A(n_4411),
.B(n_29),
.Y(n_4563)
);

BUFx3_ASAP7_75t_L g4564 ( 
.A(n_4380),
.Y(n_4564)
);

INVx3_ASAP7_75t_L g4565 ( 
.A(n_4482),
.Y(n_4565)
);

CKINVDCx5p33_ASAP7_75t_R g4566 ( 
.A(n_4335),
.Y(n_4566)
);

BUFx2_ASAP7_75t_L g4567 ( 
.A(n_4535),
.Y(n_4567)
);

AOI21xp5_ASAP7_75t_L g4568 ( 
.A1(n_4370),
.A2(n_4152),
.B(n_1836),
.Y(n_4568)
);

BUFx3_ASAP7_75t_L g4569 ( 
.A(n_4464),
.Y(n_4569)
);

AND2x2_ASAP7_75t_L g4570 ( 
.A(n_4308),
.B(n_30),
.Y(n_4570)
);

NOR2xp33_ASAP7_75t_SL g4571 ( 
.A(n_4302),
.B(n_1819),
.Y(n_4571)
);

AND2x2_ASAP7_75t_L g4572 ( 
.A(n_4388),
.B(n_30),
.Y(n_4572)
);

AND2x2_ASAP7_75t_L g4573 ( 
.A(n_4499),
.B(n_31),
.Y(n_4573)
);

BUFx2_ASAP7_75t_L g4574 ( 
.A(n_4556),
.Y(n_4574)
);

NAND2xp5_ASAP7_75t_SL g4575 ( 
.A(n_4444),
.B(n_2047),
.Y(n_4575)
);

OAI21xp33_ASAP7_75t_L g4576 ( 
.A1(n_4549),
.A2(n_32),
.B(n_34),
.Y(n_4576)
);

AND2x2_ASAP7_75t_L g4577 ( 
.A(n_4513),
.B(n_32),
.Y(n_4577)
);

OAI22xp5_ASAP7_75t_SL g4578 ( 
.A1(n_4491),
.A2(n_36),
.B1(n_34),
.B2(n_35),
.Y(n_4578)
);

AND2x4_ASAP7_75t_L g4579 ( 
.A(n_4511),
.B(n_624),
.Y(n_4579)
);

AOI21xp5_ASAP7_75t_L g4580 ( 
.A1(n_4304),
.A2(n_1836),
.B(n_1819),
.Y(n_4580)
);

AND2x2_ASAP7_75t_L g4581 ( 
.A(n_4519),
.B(n_37),
.Y(n_4581)
);

OR2x2_ASAP7_75t_L g4582 ( 
.A(n_4465),
.B(n_4402),
.Y(n_4582)
);

NAND2xp5_ASAP7_75t_L g4583 ( 
.A(n_4525),
.B(n_37),
.Y(n_4583)
);

CKINVDCx5p33_ASAP7_75t_R g4584 ( 
.A(n_4440),
.Y(n_4584)
);

BUFx2_ASAP7_75t_L g4585 ( 
.A(n_4427),
.Y(n_4585)
);

AOI22xp5_ASAP7_75t_L g4586 ( 
.A1(n_4355),
.A2(n_1926),
.B1(n_1928),
.B2(n_1881),
.Y(n_4586)
);

NAND2xp5_ASAP7_75t_L g4587 ( 
.A(n_4529),
.B(n_38),
.Y(n_4587)
);

INVx2_ASAP7_75t_SL g4588 ( 
.A(n_4503),
.Y(n_4588)
);

INVx2_ASAP7_75t_SL g4589 ( 
.A(n_4438),
.Y(n_4589)
);

AND2x4_ASAP7_75t_L g4590 ( 
.A(n_4415),
.B(n_625),
.Y(n_4590)
);

BUFx2_ASAP7_75t_L g4591 ( 
.A(n_4482),
.Y(n_4591)
);

INVx2_ASAP7_75t_L g4592 ( 
.A(n_4327),
.Y(n_4592)
);

AOI21xp5_ASAP7_75t_L g4593 ( 
.A1(n_4305),
.A2(n_1840),
.B(n_1836),
.Y(n_4593)
);

OAI21xp33_ASAP7_75t_L g4594 ( 
.A1(n_4462),
.A2(n_39),
.B(n_40),
.Y(n_4594)
);

INVx1_ASAP7_75t_SL g4595 ( 
.A(n_4357),
.Y(n_4595)
);

AND2x2_ASAP7_75t_L g4596 ( 
.A(n_4518),
.B(n_39),
.Y(n_4596)
);

INVx1_ASAP7_75t_L g4597 ( 
.A(n_4521),
.Y(n_4597)
);

NAND2xp5_ASAP7_75t_L g4598 ( 
.A(n_4338),
.B(n_40),
.Y(n_4598)
);

NOR2xp33_ASAP7_75t_L g4599 ( 
.A(n_4365),
.B(n_41),
.Y(n_4599)
);

NAND2xp5_ASAP7_75t_SL g4600 ( 
.A(n_4421),
.B(n_1836),
.Y(n_4600)
);

BUFx6f_ASAP7_75t_L g4601 ( 
.A(n_4369),
.Y(n_4601)
);

OAI21xp5_ASAP7_75t_L g4602 ( 
.A1(n_4433),
.A2(n_4367),
.B(n_4472),
.Y(n_4602)
);

CKINVDCx20_ASAP7_75t_R g4603 ( 
.A(n_4340),
.Y(n_4603)
);

AOI21xp5_ASAP7_75t_L g4604 ( 
.A1(n_4488),
.A2(n_4512),
.B(n_4322),
.Y(n_4604)
);

NOR2x1_ASAP7_75t_SL g4605 ( 
.A(n_4545),
.B(n_1840),
.Y(n_4605)
);

INVx2_ASAP7_75t_SL g4606 ( 
.A(n_4449),
.Y(n_4606)
);

NOR2xp33_ASAP7_75t_SL g4607 ( 
.A(n_4360),
.B(n_1840),
.Y(n_4607)
);

INVx3_ASAP7_75t_R g4608 ( 
.A(n_4313),
.Y(n_4608)
);

INVx1_ASAP7_75t_L g4609 ( 
.A(n_4336),
.Y(n_4609)
);

OR2x2_ASAP7_75t_L g4610 ( 
.A(n_4350),
.B(n_42),
.Y(n_4610)
);

BUFx2_ASAP7_75t_L g4611 ( 
.A(n_4557),
.Y(n_4611)
);

A2O1A1Ixp33_ASAP7_75t_L g4612 ( 
.A1(n_4495),
.A2(n_45),
.B(n_42),
.C(n_43),
.Y(n_4612)
);

AOI21xp5_ASAP7_75t_L g4613 ( 
.A1(n_4303),
.A2(n_1840),
.B(n_1813),
.Y(n_4613)
);

INVx1_ASAP7_75t_SL g4614 ( 
.A(n_4400),
.Y(n_4614)
);

NAND2xp5_ASAP7_75t_SL g4615 ( 
.A(n_4439),
.B(n_1881),
.Y(n_4615)
);

NAND2xp5_ASAP7_75t_L g4616 ( 
.A(n_4332),
.B(n_43),
.Y(n_4616)
);

AND2x2_ASAP7_75t_L g4617 ( 
.A(n_4542),
.B(n_45),
.Y(n_4617)
);

INVx2_ASAP7_75t_SL g4618 ( 
.A(n_4543),
.Y(n_4618)
);

INVx1_ASAP7_75t_L g4619 ( 
.A(n_4336),
.Y(n_4619)
);

INVx4_ASAP7_75t_L g4620 ( 
.A(n_4354),
.Y(n_4620)
);

OAI22xp5_ASAP7_75t_L g4621 ( 
.A1(n_4377),
.A2(n_48),
.B1(n_46),
.B2(n_47),
.Y(n_4621)
);

INVx3_ASAP7_75t_L g4622 ( 
.A(n_4545),
.Y(n_4622)
);

NOR2xp33_ASAP7_75t_R g4623 ( 
.A(n_4339),
.B(n_626),
.Y(n_4623)
);

OAI21xp33_ASAP7_75t_L g4624 ( 
.A1(n_4417),
.A2(n_4554),
.B(n_4541),
.Y(n_4624)
);

NAND2xp5_ASAP7_75t_L g4625 ( 
.A(n_4432),
.B(n_46),
.Y(n_4625)
);

AOI22xp5_ASAP7_75t_L g4626 ( 
.A1(n_4452),
.A2(n_1881),
.B1(n_1928),
.B2(n_1926),
.Y(n_4626)
);

CKINVDCx20_ASAP7_75t_R g4627 ( 
.A(n_4547),
.Y(n_4627)
);

BUFx6f_ASAP7_75t_L g4628 ( 
.A(n_4369),
.Y(n_4628)
);

NAND2xp5_ASAP7_75t_SL g4629 ( 
.A(n_4517),
.B(n_1881),
.Y(n_4629)
);

AOI22xp33_ASAP7_75t_L g4630 ( 
.A1(n_4426),
.A2(n_1926),
.B1(n_1950),
.B2(n_1928),
.Y(n_4630)
);

CKINVDCx20_ASAP7_75t_R g4631 ( 
.A(n_4543),
.Y(n_4631)
);

INVx1_ASAP7_75t_L g4632 ( 
.A(n_4336),
.Y(n_4632)
);

CKINVDCx11_ASAP7_75t_R g4633 ( 
.A(n_4360),
.Y(n_4633)
);

INVx1_ASAP7_75t_SL g4634 ( 
.A(n_4400),
.Y(n_4634)
);

INVx2_ASAP7_75t_SL g4635 ( 
.A(n_4369),
.Y(n_4635)
);

AND2x2_ASAP7_75t_L g4636 ( 
.A(n_4443),
.B(n_47),
.Y(n_4636)
);

INVx1_ASAP7_75t_L g4637 ( 
.A(n_4479),
.Y(n_4637)
);

AND2x4_ASAP7_75t_L g4638 ( 
.A(n_4451),
.B(n_627),
.Y(n_4638)
);

INVx2_ASAP7_75t_SL g4639 ( 
.A(n_4397),
.Y(n_4639)
);

BUFx12f_ASAP7_75t_L g4640 ( 
.A(n_4431),
.Y(n_4640)
);

AND2x4_ASAP7_75t_L g4641 ( 
.A(n_4469),
.B(n_4396),
.Y(n_4641)
);

AND2x2_ASAP7_75t_L g4642 ( 
.A(n_4351),
.B(n_48),
.Y(n_4642)
);

INVx1_ASAP7_75t_L g4643 ( 
.A(n_4352),
.Y(n_4643)
);

INVx4_ASAP7_75t_L g4644 ( 
.A(n_4354),
.Y(n_4644)
);

AOI21xp5_ASAP7_75t_L g4645 ( 
.A1(n_4410),
.A2(n_1813),
.B(n_1926),
.Y(n_4645)
);

INVx1_ASAP7_75t_L g4646 ( 
.A(n_4352),
.Y(n_4646)
);

BUFx3_ASAP7_75t_L g4647 ( 
.A(n_4527),
.Y(n_4647)
);

BUFx6f_ASAP7_75t_L g4648 ( 
.A(n_4397),
.Y(n_4648)
);

CKINVDCx5p33_ASAP7_75t_R g4649 ( 
.A(n_4397),
.Y(n_4649)
);

INVx1_ASAP7_75t_SL g4650 ( 
.A(n_4348),
.Y(n_4650)
);

INVxp67_ASAP7_75t_SL g4651 ( 
.A(n_4461),
.Y(n_4651)
);

AND2x2_ASAP7_75t_L g4652 ( 
.A(n_4391),
.B(n_49),
.Y(n_4652)
);

AND2x2_ASAP7_75t_SL g4653 ( 
.A(n_4406),
.B(n_49),
.Y(n_4653)
);

AND2x2_ASAP7_75t_L g4654 ( 
.A(n_4539),
.B(n_50),
.Y(n_4654)
);

INVx1_ASAP7_75t_L g4655 ( 
.A(n_4352),
.Y(n_4655)
);

INVx1_ASAP7_75t_L g4656 ( 
.A(n_4553),
.Y(n_4656)
);

NAND2xp5_ASAP7_75t_L g4657 ( 
.A(n_4353),
.B(n_51),
.Y(n_4657)
);

INVx2_ASAP7_75t_L g4658 ( 
.A(n_4463),
.Y(n_4658)
);

NAND2xp5_ASAP7_75t_L g4659 ( 
.A(n_4314),
.B(n_51),
.Y(n_4659)
);

OAI22xp5_ASAP7_75t_L g4660 ( 
.A1(n_4474),
.A2(n_4473),
.B1(n_4384),
.B2(n_4531),
.Y(n_4660)
);

INVx2_ASAP7_75t_L g4661 ( 
.A(n_4463),
.Y(n_4661)
);

NOR2x1_ASAP7_75t_SL g4662 ( 
.A(n_4318),
.B(n_1928),
.Y(n_4662)
);

AND2x4_ASAP7_75t_L g4663 ( 
.A(n_4354),
.B(n_628),
.Y(n_4663)
);

INVxp67_ASAP7_75t_L g4664 ( 
.A(n_4487),
.Y(n_4664)
);

INVx1_ASAP7_75t_L g4665 ( 
.A(n_4553),
.Y(n_4665)
);

NAND2xp5_ASAP7_75t_L g4666 ( 
.A(n_4323),
.B(n_53),
.Y(n_4666)
);

AND2x2_ASAP7_75t_L g4667 ( 
.A(n_4540),
.B(n_53),
.Y(n_4667)
);

BUFx6f_ASAP7_75t_L g4668 ( 
.A(n_4463),
.Y(n_4668)
);

INVx2_ASAP7_75t_L g4669 ( 
.A(n_4481),
.Y(n_4669)
);

NAND2xp5_ASAP7_75t_L g4670 ( 
.A(n_4311),
.B(n_54),
.Y(n_4670)
);

AND2x4_ASAP7_75t_SL g4671 ( 
.A(n_4538),
.B(n_633),
.Y(n_4671)
);

A2O1A1Ixp33_ASAP7_75t_L g4672 ( 
.A1(n_4375),
.A2(n_56),
.B(n_54),
.C(n_55),
.Y(n_4672)
);

CKINVDCx5p33_ASAP7_75t_R g4673 ( 
.A(n_4481),
.Y(n_4673)
);

AND2x4_ASAP7_75t_L g4674 ( 
.A(n_4538),
.B(n_638),
.Y(n_4674)
);

BUFx6f_ASAP7_75t_L g4675 ( 
.A(n_4481),
.Y(n_4675)
);

INVx1_ASAP7_75t_L g4676 ( 
.A(n_4553),
.Y(n_4676)
);

INVx2_ASAP7_75t_L g4677 ( 
.A(n_4504),
.Y(n_4677)
);

NAND2xp5_ASAP7_75t_L g4678 ( 
.A(n_4321),
.B(n_55),
.Y(n_4678)
);

AND2x2_ASAP7_75t_L g4679 ( 
.A(n_4551),
.B(n_56),
.Y(n_4679)
);

INVx2_ASAP7_75t_SL g4680 ( 
.A(n_4475),
.Y(n_4680)
);

NAND3xp33_ASAP7_75t_L g4681 ( 
.A(n_4395),
.B(n_1962),
.C(n_1950),
.Y(n_4681)
);

INVx2_ASAP7_75t_L g4682 ( 
.A(n_4371),
.Y(n_4682)
);

BUFx3_ASAP7_75t_L g4683 ( 
.A(n_4493),
.Y(n_4683)
);

OAI21xp5_ASAP7_75t_L g4684 ( 
.A1(n_4477),
.A2(n_1962),
.B(n_1950),
.Y(n_4684)
);

INVx2_ASAP7_75t_L g4685 ( 
.A(n_4371),
.Y(n_4685)
);

NAND2xp5_ASAP7_75t_L g4686 ( 
.A(n_4358),
.B(n_4387),
.Y(n_4686)
);

OAI21x1_ASAP7_75t_L g4687 ( 
.A1(n_4326),
.A2(n_642),
.B(n_640),
.Y(n_4687)
);

NAND2xp5_ASAP7_75t_L g4688 ( 
.A(n_4310),
.B(n_4356),
.Y(n_4688)
);

INVx1_ASAP7_75t_L g4689 ( 
.A(n_4371),
.Y(n_4689)
);

BUFx3_ASAP7_75t_L g4690 ( 
.A(n_4528),
.Y(n_4690)
);

AND2x2_ASAP7_75t_L g4691 ( 
.A(n_4555),
.B(n_57),
.Y(n_4691)
);

AND2x2_ASAP7_75t_L g4692 ( 
.A(n_4406),
.B(n_57),
.Y(n_4692)
);

AND2x4_ASAP7_75t_L g4693 ( 
.A(n_4552),
.B(n_647),
.Y(n_4693)
);

INVx1_ASAP7_75t_L g4694 ( 
.A(n_4485),
.Y(n_4694)
);

AND2x2_ASAP7_75t_L g4695 ( 
.A(n_4502),
.B(n_58),
.Y(n_4695)
);

HB1xp67_ASAP7_75t_L g4696 ( 
.A(n_4342),
.Y(n_4696)
);

CKINVDCx20_ASAP7_75t_R g4697 ( 
.A(n_4337),
.Y(n_4697)
);

A2O1A1Ixp33_ASAP7_75t_SL g4698 ( 
.A1(n_4423),
.A2(n_62),
.B(n_58),
.C(n_60),
.Y(n_4698)
);

AOI21xp5_ASAP7_75t_L g4699 ( 
.A1(n_4404),
.A2(n_1962),
.B(n_1950),
.Y(n_4699)
);

A2O1A1Ixp33_ASAP7_75t_L g4700 ( 
.A1(n_4390),
.A2(n_66),
.B(n_62),
.C(n_64),
.Y(n_4700)
);

A2O1A1Ixp33_ASAP7_75t_L g4701 ( 
.A1(n_4478),
.A2(n_68),
.B(n_64),
.C(n_67),
.Y(n_4701)
);

BUFx3_ASAP7_75t_L g4702 ( 
.A(n_4483),
.Y(n_4702)
);

AND2x4_ASAP7_75t_L g4703 ( 
.A(n_4448),
.B(n_653),
.Y(n_4703)
);

INVxp67_ASAP7_75t_SL g4704 ( 
.A(n_4312),
.Y(n_4704)
);

INVx3_ASAP7_75t_L g4705 ( 
.A(n_4483),
.Y(n_4705)
);

INVx2_ASAP7_75t_L g4706 ( 
.A(n_4509),
.Y(n_4706)
);

INVx1_ASAP7_75t_L g4707 ( 
.A(n_4485),
.Y(n_4707)
);

INVx2_ASAP7_75t_L g4708 ( 
.A(n_4342),
.Y(n_4708)
);

BUFx2_ASAP7_75t_SL g4709 ( 
.A(n_4413),
.Y(n_4709)
);

INVx5_ASAP7_75t_L g4710 ( 
.A(n_4448),
.Y(n_4710)
);

NAND2xp5_ASAP7_75t_L g4711 ( 
.A(n_4405),
.B(n_67),
.Y(n_4711)
);

BUFx3_ASAP7_75t_L g4712 ( 
.A(n_4526),
.Y(n_4712)
);

CKINVDCx5p33_ASAP7_75t_R g4713 ( 
.A(n_4546),
.Y(n_4713)
);

INVx4_ASAP7_75t_L g4714 ( 
.A(n_4320),
.Y(n_4714)
);

AOI21xp5_ASAP7_75t_L g4715 ( 
.A1(n_4309),
.A2(n_1975),
.B(n_1962),
.Y(n_4715)
);

AND2x2_ASAP7_75t_L g4716 ( 
.A(n_4342),
.B(n_68),
.Y(n_4716)
);

INVx1_ASAP7_75t_L g4717 ( 
.A(n_4328),
.Y(n_4717)
);

NAND2xp5_ASAP7_75t_L g4718 ( 
.A(n_4434),
.B(n_69),
.Y(n_4718)
);

NAND2x1p5_ASAP7_75t_L g4719 ( 
.A(n_4496),
.B(n_1975),
.Y(n_4719)
);

AOI21xp5_ASAP7_75t_L g4720 ( 
.A1(n_4324),
.A2(n_1982),
.B(n_1975),
.Y(n_4720)
);

OR2x6_ASAP7_75t_L g4721 ( 
.A(n_4430),
.B(n_654),
.Y(n_4721)
);

HB1xp67_ASAP7_75t_L g4722 ( 
.A(n_4532),
.Y(n_4722)
);

NOR2xp33_ASAP7_75t_L g4723 ( 
.A(n_4516),
.B(n_69),
.Y(n_4723)
);

INVx2_ASAP7_75t_SL g4724 ( 
.A(n_4548),
.Y(n_4724)
);

AND2x2_ASAP7_75t_L g4725 ( 
.A(n_4330),
.B(n_4328),
.Y(n_4725)
);

INVx4_ASAP7_75t_L g4726 ( 
.A(n_4435),
.Y(n_4726)
);

INVx2_ASAP7_75t_L g4727 ( 
.A(n_4422),
.Y(n_4727)
);

AOI21xp5_ASAP7_75t_L g4728 ( 
.A1(n_4514),
.A2(n_1982),
.B(n_1975),
.Y(n_4728)
);

BUFx3_ASAP7_75t_L g4729 ( 
.A(n_4544),
.Y(n_4729)
);

OR2x6_ASAP7_75t_L g4730 ( 
.A(n_4480),
.B(n_655),
.Y(n_4730)
);

INVx1_ASAP7_75t_SL g4731 ( 
.A(n_4412),
.Y(n_4731)
);

NAND3xp33_ASAP7_75t_L g4732 ( 
.A(n_4403),
.B(n_1984),
.C(n_1982),
.Y(n_4732)
);

OR2x2_ASAP7_75t_L g4733 ( 
.A(n_4453),
.B(n_70),
.Y(n_4733)
);

AND2x2_ASAP7_75t_L g4734 ( 
.A(n_4328),
.B(n_71),
.Y(n_4734)
);

INVxp67_ASAP7_75t_SL g4735 ( 
.A(n_4345),
.Y(n_4735)
);

AOI21xp5_ASAP7_75t_L g4736 ( 
.A1(n_4514),
.A2(n_1984),
.B(n_1982),
.Y(n_4736)
);

NAND2xp5_ASAP7_75t_L g4737 ( 
.A(n_4363),
.B(n_72),
.Y(n_4737)
);

INVx1_ASAP7_75t_L g4738 ( 
.A(n_4501),
.Y(n_4738)
);

AOI21xp5_ASAP7_75t_L g4739 ( 
.A1(n_4366),
.A2(n_1986),
.B(n_1984),
.Y(n_4739)
);

AND2x4_ASAP7_75t_L g4740 ( 
.A(n_4501),
.B(n_663),
.Y(n_4740)
);

O2A1O1Ixp5_ASAP7_75t_L g4741 ( 
.A1(n_4506),
.A2(n_75),
.B(n_73),
.C(n_74),
.Y(n_4741)
);

OR2x6_ASAP7_75t_L g4742 ( 
.A(n_4537),
.B(n_666),
.Y(n_4742)
);

AND2x4_ASAP7_75t_L g4743 ( 
.A(n_4501),
.B(n_668),
.Y(n_4743)
);

INVx2_ASAP7_75t_L g4744 ( 
.A(n_4393),
.Y(n_4744)
);

NOR3xp33_ASAP7_75t_L g4745 ( 
.A(n_4471),
.B(n_4343),
.C(n_4450),
.Y(n_4745)
);

INVx2_ASAP7_75t_L g4746 ( 
.A(n_4393),
.Y(n_4746)
);

INVx2_ASAP7_75t_L g4747 ( 
.A(n_4523),
.Y(n_4747)
);

A2O1A1Ixp33_ASAP7_75t_L g4748 ( 
.A1(n_4456),
.A2(n_77),
.B(n_73),
.C(n_75),
.Y(n_4748)
);

INVx6_ASAP7_75t_L g4749 ( 
.A(n_4466),
.Y(n_4749)
);

NOR2x1_ASAP7_75t_SL g4750 ( 
.A(n_4498),
.B(n_4442),
.Y(n_4750)
);

AND2x2_ASAP7_75t_L g4751 ( 
.A(n_4460),
.B(n_78),
.Y(n_4751)
);

AOI21xp33_ASAP7_75t_SL g4752 ( 
.A1(n_4361),
.A2(n_78),
.B(n_79),
.Y(n_4752)
);

INVx1_ASAP7_75t_L g4753 ( 
.A(n_4523),
.Y(n_4753)
);

A2O1A1Ixp33_ASAP7_75t_L g4754 ( 
.A1(n_4346),
.A2(n_83),
.B(n_80),
.C(n_82),
.Y(n_4754)
);

NAND2xp5_ASAP7_75t_L g4755 ( 
.A(n_4364),
.B(n_83),
.Y(n_4755)
);

AND2x4_ASAP7_75t_L g4756 ( 
.A(n_4550),
.B(n_671),
.Y(n_4756)
);

INVx1_ASAP7_75t_L g4757 ( 
.A(n_4325),
.Y(n_4757)
);

CKINVDCx8_ASAP7_75t_R g4758 ( 
.A(n_4435),
.Y(n_4758)
);

NOR2xp33_ASAP7_75t_SL g4759 ( 
.A(n_4522),
.B(n_1984),
.Y(n_4759)
);

OR2x2_ASAP7_75t_L g4760 ( 
.A(n_4441),
.B(n_84),
.Y(n_4760)
);

CKINVDCx5p33_ASAP7_75t_R g4761 ( 
.A(n_4349),
.Y(n_4761)
);

INVx1_ASAP7_75t_L g4762 ( 
.A(n_4325),
.Y(n_4762)
);

INVx2_ASAP7_75t_L g4763 ( 
.A(n_4507),
.Y(n_4763)
);

INVx3_ASAP7_75t_SL g4764 ( 
.A(n_4373),
.Y(n_4764)
);

INVx3_ASAP7_75t_L g4765 ( 
.A(n_4534),
.Y(n_4765)
);

INVx2_ASAP7_75t_L g4766 ( 
.A(n_4378),
.Y(n_4766)
);

BUFx3_ASAP7_75t_L g4767 ( 
.A(n_4486),
.Y(n_4767)
);

OAI21xp33_ASAP7_75t_L g4768 ( 
.A1(n_4470),
.A2(n_84),
.B(n_86),
.Y(n_4768)
);

NOR2xp33_ASAP7_75t_L g4769 ( 
.A(n_4347),
.B(n_86),
.Y(n_4769)
);

AND2x4_ASAP7_75t_L g4770 ( 
.A(n_4520),
.B(n_674),
.Y(n_4770)
);

AOI22xp5_ASAP7_75t_L g4771 ( 
.A1(n_4492),
.A2(n_1986),
.B1(n_2003),
.B2(n_1993),
.Y(n_4771)
);

OAI22xp33_ASAP7_75t_L g4772 ( 
.A1(n_4455),
.A2(n_89),
.B1(n_87),
.B2(n_88),
.Y(n_4772)
);

INVx2_ASAP7_75t_L g4773 ( 
.A(n_4383),
.Y(n_4773)
);

INVx8_ASAP7_75t_L g4774 ( 
.A(n_4505),
.Y(n_4774)
);

BUFx2_ASAP7_75t_L g4775 ( 
.A(n_4428),
.Y(n_4775)
);

INVx1_ASAP7_75t_L g4776 ( 
.A(n_4306),
.Y(n_4776)
);

NOR2xp33_ASAP7_75t_L g4777 ( 
.A(n_4372),
.B(n_88),
.Y(n_4777)
);

INVx6_ASAP7_75t_L g4778 ( 
.A(n_4429),
.Y(n_4778)
);

AND2x2_ASAP7_75t_L g4779 ( 
.A(n_4489),
.B(n_91),
.Y(n_4779)
);

INVx1_ASAP7_75t_L g4780 ( 
.A(n_4414),
.Y(n_4780)
);

INVx1_ASAP7_75t_L g4781 ( 
.A(n_4447),
.Y(n_4781)
);

NOR2x1_ASAP7_75t_L g4782 ( 
.A(n_4458),
.B(n_91),
.Y(n_4782)
);

AND2x2_ASAP7_75t_L g4783 ( 
.A(n_4445),
.B(n_95),
.Y(n_4783)
);

INVx2_ASAP7_75t_L g4784 ( 
.A(n_4359),
.Y(n_4784)
);

INVx3_ASAP7_75t_L g4785 ( 
.A(n_4425),
.Y(n_4785)
);

INVx2_ASAP7_75t_L g4786 ( 
.A(n_4407),
.Y(n_4786)
);

OAI22xp5_ASAP7_75t_L g4787 ( 
.A1(n_4381),
.A2(n_98),
.B1(n_96),
.B2(n_97),
.Y(n_4787)
);

OAI22xp5_ASAP7_75t_L g4788 ( 
.A1(n_4333),
.A2(n_100),
.B1(n_98),
.B2(n_99),
.Y(n_4788)
);

OAI22xp5_ASAP7_75t_L g4789 ( 
.A1(n_4500),
.A2(n_102),
.B1(n_99),
.B2(n_101),
.Y(n_4789)
);

NOR2xp33_ASAP7_75t_L g4790 ( 
.A(n_4317),
.B(n_102),
.Y(n_4790)
);

BUFx6f_ASAP7_75t_L g4791 ( 
.A(n_4533),
.Y(n_4791)
);

AOI21xp5_ASAP7_75t_L g4792 ( 
.A1(n_4467),
.A2(n_1993),
.B(n_1986),
.Y(n_4792)
);

INVx4_ASAP7_75t_L g4793 ( 
.A(n_4508),
.Y(n_4793)
);

AND2x2_ASAP7_75t_L g4794 ( 
.A(n_4445),
.B(n_103),
.Y(n_4794)
);

BUFx6f_ASAP7_75t_L g4795 ( 
.A(n_4454),
.Y(n_4795)
);

AOI22xp5_ASAP7_75t_L g4796 ( 
.A1(n_4362),
.A2(n_4379),
.B1(n_4515),
.B2(n_4536),
.Y(n_4796)
);

BUFx2_ASAP7_75t_L g4797 ( 
.A(n_4445),
.Y(n_4797)
);

AOI21xp5_ASAP7_75t_L g4798 ( 
.A1(n_4510),
.A2(n_4392),
.B(n_4331),
.Y(n_4798)
);

NAND2xp5_ASAP7_75t_L g4799 ( 
.A(n_4307),
.B(n_103),
.Y(n_4799)
);

INVx1_ASAP7_75t_L g4800 ( 
.A(n_4319),
.Y(n_4800)
);

HB1xp67_ASAP7_75t_L g4801 ( 
.A(n_4457),
.Y(n_4801)
);

AOI22xp5_ASAP7_75t_L g4802 ( 
.A1(n_4468),
.A2(n_4494),
.B1(n_4490),
.B2(n_4484),
.Y(n_4802)
);

BUFx3_ASAP7_75t_L g4803 ( 
.A(n_4437),
.Y(n_4803)
);

OR2x2_ASAP7_75t_L g4804 ( 
.A(n_4457),
.B(n_4374),
.Y(n_4804)
);

INVx1_ASAP7_75t_L g4805 ( 
.A(n_4420),
.Y(n_4805)
);

NAND2xp5_ASAP7_75t_L g4806 ( 
.A(n_4386),
.B(n_104),
.Y(n_4806)
);

AO31x2_ASAP7_75t_L g4807 ( 
.A1(n_4386),
.A2(n_106),
.A3(n_104),
.B(n_105),
.Y(n_4807)
);

NAND2xp5_ASAP7_75t_L g4808 ( 
.A(n_4476),
.B(n_107),
.Y(n_4808)
);

INVx2_ASAP7_75t_L g4809 ( 
.A(n_4582),
.Y(n_4809)
);

BUFx3_ASAP7_75t_L g4810 ( 
.A(n_4603),
.Y(n_4810)
);

INVx1_ASAP7_75t_L g4811 ( 
.A(n_4597),
.Y(n_4811)
);

OAI22xp5_ASAP7_75t_L g4812 ( 
.A1(n_4748),
.A2(n_4382),
.B1(n_4376),
.B2(n_4497),
.Y(n_4812)
);

AOI21xp33_ASAP7_75t_L g4813 ( 
.A1(n_4653),
.A2(n_4398),
.B(n_4530),
.Y(n_4813)
);

BUFx10_ASAP7_75t_L g4814 ( 
.A(n_4749),
.Y(n_4814)
);

INVx1_ASAP7_75t_L g4815 ( 
.A(n_4637),
.Y(n_4815)
);

NAND2x1_ASAP7_75t_L g4816 ( 
.A(n_4714),
.B(n_4334),
.Y(n_4816)
);

BUFx12f_ASAP7_75t_L g4817 ( 
.A(n_4633),
.Y(n_4817)
);

BUFx3_ASAP7_75t_L g4818 ( 
.A(n_4569),
.Y(n_4818)
);

INVx6_ASAP7_75t_L g4819 ( 
.A(n_4640),
.Y(n_4819)
);

AOI22xp5_ASAP7_75t_SL g4820 ( 
.A1(n_4599),
.A2(n_4329),
.B1(n_4524),
.B2(n_110),
.Y(n_4820)
);

AOI22xp33_ASAP7_75t_SL g4821 ( 
.A1(n_4602),
.A2(n_4446),
.B1(n_4424),
.B2(n_4341),
.Y(n_4821)
);

AOI22xp33_ASAP7_75t_SL g4822 ( 
.A1(n_4578),
.A2(n_4408),
.B1(n_4394),
.B2(n_4401),
.Y(n_4822)
);

BUFx6f_ASAP7_75t_L g4823 ( 
.A(n_4601),
.Y(n_4823)
);

CKINVDCx11_ASAP7_75t_R g4824 ( 
.A(n_4631),
.Y(n_4824)
);

AND2x2_ASAP7_75t_L g4825 ( 
.A(n_4585),
.B(n_4567),
.Y(n_4825)
);

INVx1_ASAP7_75t_L g4826 ( 
.A(n_4592),
.Y(n_4826)
);

INVx1_ASAP7_75t_L g4827 ( 
.A(n_4611),
.Y(n_4827)
);

CKINVDCx20_ASAP7_75t_R g4828 ( 
.A(n_4558),
.Y(n_4828)
);

INVx1_ASAP7_75t_L g4829 ( 
.A(n_4561),
.Y(n_4829)
);

INVx6_ASAP7_75t_L g4830 ( 
.A(n_4749),
.Y(n_4830)
);

INVx4_ASAP7_75t_L g4831 ( 
.A(n_4710),
.Y(n_4831)
);

NAND2xp5_ASAP7_75t_L g4832 ( 
.A(n_4704),
.B(n_4457),
.Y(n_4832)
);

INVx1_ASAP7_75t_L g4833 ( 
.A(n_4694),
.Y(n_4833)
);

BUFx2_ASAP7_75t_SL g4834 ( 
.A(n_4627),
.Y(n_4834)
);

OAI22xp33_ASAP7_75t_SL g4835 ( 
.A1(n_4758),
.A2(n_111),
.B1(n_107),
.B2(n_109),
.Y(n_4835)
);

INVx2_ASAP7_75t_L g4836 ( 
.A(n_4574),
.Y(n_4836)
);

INVx1_ASAP7_75t_SL g4837 ( 
.A(n_4595),
.Y(n_4837)
);

INVx6_ASAP7_75t_L g4838 ( 
.A(n_4564),
.Y(n_4838)
);

INVx1_ASAP7_75t_L g4839 ( 
.A(n_4707),
.Y(n_4839)
);

AND2x2_ASAP7_75t_L g4840 ( 
.A(n_4650),
.B(n_4344),
.Y(n_4840)
);

OAI22xp5_ASAP7_75t_L g4841 ( 
.A1(n_4764),
.A2(n_4510),
.B1(n_4385),
.B2(n_4399),
.Y(n_4841)
);

INVx6_ASAP7_75t_L g4842 ( 
.A(n_4601),
.Y(n_4842)
);

AOI22xp33_ASAP7_75t_L g4843 ( 
.A1(n_4745),
.A2(n_4624),
.B1(n_4594),
.B2(n_4576),
.Y(n_4843)
);

AND2x2_ASAP7_75t_L g4844 ( 
.A(n_4614),
.B(n_4385),
.Y(n_4844)
);

INVx1_ASAP7_75t_SL g4845 ( 
.A(n_4562),
.Y(n_4845)
);

AOI22xp33_ASAP7_75t_L g4846 ( 
.A1(n_4768),
.A2(n_4409),
.B1(n_4418),
.B2(n_4416),
.Y(n_4846)
);

BUFx2_ASAP7_75t_L g4847 ( 
.A(n_4622),
.Y(n_4847)
);

AOI22xp33_ASAP7_75t_L g4848 ( 
.A1(n_4799),
.A2(n_1993),
.B1(n_2003),
.B2(n_1986),
.Y(n_4848)
);

AOI22xp33_ASAP7_75t_L g4849 ( 
.A1(n_4767),
.A2(n_2003),
.B1(n_1993),
.B2(n_113),
.Y(n_4849)
);

INVx1_ASAP7_75t_L g4850 ( 
.A(n_4609),
.Y(n_4850)
);

INVx1_ASAP7_75t_L g4851 ( 
.A(n_4619),
.Y(n_4851)
);

INVx1_ASAP7_75t_L g4852 ( 
.A(n_4632),
.Y(n_4852)
);

BUFx3_ASAP7_75t_L g4853 ( 
.A(n_4588),
.Y(n_4853)
);

BUFx12f_ASAP7_75t_L g4854 ( 
.A(n_4584),
.Y(n_4854)
);

INVx2_ASAP7_75t_L g4855 ( 
.A(n_4658),
.Y(n_4855)
);

INVx2_ASAP7_75t_SL g4856 ( 
.A(n_4647),
.Y(n_4856)
);

OAI22xp5_ASAP7_75t_L g4857 ( 
.A1(n_4754),
.A2(n_4697),
.B1(n_4672),
.B2(n_4701),
.Y(n_4857)
);

AOI22xp33_ASAP7_75t_L g4858 ( 
.A1(n_4604),
.A2(n_2003),
.B1(n_113),
.B2(n_109),
.Y(n_4858)
);

AOI22xp33_ASAP7_75t_SL g4859 ( 
.A1(n_4783),
.A2(n_116),
.B1(n_112),
.B2(n_115),
.Y(n_4859)
);

BUFx12f_ASAP7_75t_L g4860 ( 
.A(n_4566),
.Y(n_4860)
);

AOI22xp33_ASAP7_75t_L g4861 ( 
.A1(n_4778),
.A2(n_117),
.B1(n_115),
.B2(n_116),
.Y(n_4861)
);

OAI22xp33_ASAP7_75t_L g4862 ( 
.A1(n_4796),
.A2(n_4721),
.B1(n_4586),
.B2(n_4730),
.Y(n_4862)
);

INVx1_ASAP7_75t_L g4863 ( 
.A(n_4738),
.Y(n_4863)
);

INVx2_ASAP7_75t_L g4864 ( 
.A(n_4661),
.Y(n_4864)
);

BUFx6f_ASAP7_75t_L g4865 ( 
.A(n_4601),
.Y(n_4865)
);

AOI22xp33_ASAP7_75t_L g4866 ( 
.A1(n_4778),
.A2(n_124),
.B1(n_121),
.B2(n_123),
.Y(n_4866)
);

INVx4_ASAP7_75t_L g4867 ( 
.A(n_4710),
.Y(n_4867)
);

INVx1_ASAP7_75t_L g4868 ( 
.A(n_4643),
.Y(n_4868)
);

INVx1_ASAP7_75t_L g4869 ( 
.A(n_4722),
.Y(n_4869)
);

INVx3_ASAP7_75t_L g4870 ( 
.A(n_4622),
.Y(n_4870)
);

AOI22xp33_ASAP7_75t_L g4871 ( 
.A1(n_4621),
.A2(n_124),
.B1(n_121),
.B2(n_123),
.Y(n_4871)
);

BUFx4_ASAP7_75t_R g4872 ( 
.A(n_4702),
.Y(n_4872)
);

NAND2x1p5_ASAP7_75t_L g4873 ( 
.A(n_4710),
.B(n_4419),
.Y(n_4873)
);

INVx2_ASAP7_75t_L g4874 ( 
.A(n_4669),
.Y(n_4874)
);

INVx1_ASAP7_75t_L g4875 ( 
.A(n_4646),
.Y(n_4875)
);

AOI22xp5_ASAP7_75t_L g4876 ( 
.A1(n_4788),
.A2(n_4385),
.B1(n_4399),
.B2(n_127),
.Y(n_4876)
);

BUFx2_ASAP7_75t_L g4877 ( 
.A(n_4641),
.Y(n_4877)
);

OAI22xp5_ASAP7_75t_L g4878 ( 
.A1(n_4761),
.A2(n_4700),
.B1(n_4612),
.B2(n_4630),
.Y(n_4878)
);

BUFx3_ASAP7_75t_L g4879 ( 
.A(n_4591),
.Y(n_4879)
);

INVx2_ASAP7_75t_L g4880 ( 
.A(n_4747),
.Y(n_4880)
);

INVx1_ASAP7_75t_L g4881 ( 
.A(n_4655),
.Y(n_4881)
);

AOI22xp33_ASAP7_75t_SL g4882 ( 
.A1(n_4794),
.A2(n_128),
.B1(n_125),
.B2(n_126),
.Y(n_4882)
);

AOI22xp5_ASAP7_75t_L g4883 ( 
.A1(n_4660),
.A2(n_4399),
.B1(n_130),
.B2(n_126),
.Y(n_4883)
);

INVx2_ASAP7_75t_L g4884 ( 
.A(n_4677),
.Y(n_4884)
);

HB1xp67_ASAP7_75t_L g4885 ( 
.A(n_4801),
.Y(n_4885)
);

INVx1_ASAP7_75t_L g4886 ( 
.A(n_4656),
.Y(n_4886)
);

AOI22xp33_ASAP7_75t_SL g4887 ( 
.A1(n_4692),
.A2(n_132),
.B1(n_129),
.B2(n_131),
.Y(n_4887)
);

AOI22xp33_ASAP7_75t_SL g4888 ( 
.A1(n_4774),
.A2(n_132),
.B1(n_129),
.B2(n_131),
.Y(n_4888)
);

BUFx4f_ASAP7_75t_SL g4889 ( 
.A(n_4565),
.Y(n_4889)
);

AND2x2_ASAP7_75t_L g4890 ( 
.A(n_4634),
.B(n_133),
.Y(n_4890)
);

NAND2xp5_ASAP7_75t_L g4891 ( 
.A(n_4559),
.B(n_134),
.Y(n_4891)
);

INVx1_ASAP7_75t_L g4892 ( 
.A(n_4665),
.Y(n_4892)
);

BUFx4_ASAP7_75t_SL g4893 ( 
.A(n_4649),
.Y(n_4893)
);

INVx2_ASAP7_75t_L g4894 ( 
.A(n_4753),
.Y(n_4894)
);

OAI22xp33_ASAP7_75t_L g4895 ( 
.A1(n_4721),
.A2(n_137),
.B1(n_135),
.B2(n_136),
.Y(n_4895)
);

INVx1_ASAP7_75t_L g4896 ( 
.A(n_4676),
.Y(n_4896)
);

INVx1_ASAP7_75t_L g4897 ( 
.A(n_4689),
.Y(n_4897)
);

INVx2_ASAP7_75t_L g4898 ( 
.A(n_4727),
.Y(n_4898)
);

BUFx10_ASAP7_75t_L g4899 ( 
.A(n_4769),
.Y(n_4899)
);

AOI22xp33_ASAP7_75t_L g4900 ( 
.A1(n_4729),
.A2(n_139),
.B1(n_135),
.B2(n_137),
.Y(n_4900)
);

INVx1_ASAP7_75t_L g4901 ( 
.A(n_4717),
.Y(n_4901)
);

NAND2xp5_ASAP7_75t_L g4902 ( 
.A(n_4724),
.B(n_139),
.Y(n_4902)
);

BUFx3_ASAP7_75t_L g4903 ( 
.A(n_4673),
.Y(n_4903)
);

INVx1_ASAP7_75t_SL g4904 ( 
.A(n_4731),
.Y(n_4904)
);

NAND2xp5_ASAP7_75t_L g4905 ( 
.A(n_4686),
.B(n_140),
.Y(n_4905)
);

AOI22xp33_ASAP7_75t_L g4906 ( 
.A1(n_4774),
.A2(n_143),
.B1(n_141),
.B2(n_142),
.Y(n_4906)
);

AOI22xp33_ASAP7_75t_L g4907 ( 
.A1(n_4777),
.A2(n_145),
.B1(n_142),
.B2(n_144),
.Y(n_4907)
);

NAND2x1p5_ASAP7_75t_L g4908 ( 
.A(n_4714),
.B(n_1867),
.Y(n_4908)
);

INVx2_ASAP7_75t_L g4909 ( 
.A(n_4744),
.Y(n_4909)
);

AOI22xp33_ASAP7_75t_L g4910 ( 
.A1(n_4723),
.A2(n_147),
.B1(n_145),
.B2(n_146),
.Y(n_4910)
);

INVx6_ASAP7_75t_L g4911 ( 
.A(n_4628),
.Y(n_4911)
);

INVx1_ASAP7_75t_SL g4912 ( 
.A(n_4683),
.Y(n_4912)
);

AOI22xp33_ASAP7_75t_SL g4913 ( 
.A1(n_4790),
.A2(n_151),
.B1(n_148),
.B2(n_149),
.Y(n_4913)
);

NAND2xp5_ASAP7_75t_L g4914 ( 
.A(n_4688),
.B(n_152),
.Y(n_4914)
);

INVx6_ASAP7_75t_L g4915 ( 
.A(n_4628),
.Y(n_4915)
);

INVx1_ASAP7_75t_L g4916 ( 
.A(n_4696),
.Y(n_4916)
);

INVx2_ASAP7_75t_L g4917 ( 
.A(n_4746),
.Y(n_4917)
);

AOI22xp33_ASAP7_75t_L g4918 ( 
.A1(n_4600),
.A2(n_154),
.B1(n_152),
.B2(n_153),
.Y(n_4918)
);

AOI22xp33_ASAP7_75t_L g4919 ( 
.A1(n_4772),
.A2(n_157),
.B1(n_155),
.B2(n_156),
.Y(n_4919)
);

AOI22xp33_ASAP7_75t_L g4920 ( 
.A1(n_4716),
.A2(n_158),
.B1(n_155),
.B2(n_157),
.Y(n_4920)
);

INVx6_ASAP7_75t_L g4921 ( 
.A(n_4628),
.Y(n_4921)
);

AOI22xp33_ASAP7_75t_SL g4922 ( 
.A1(n_4740),
.A2(n_160),
.B1(n_158),
.B2(n_159),
.Y(n_4922)
);

BUFx4f_ASAP7_75t_SL g4923 ( 
.A(n_4565),
.Y(n_4923)
);

OAI21xp5_ASAP7_75t_L g4924 ( 
.A1(n_4741),
.A2(n_159),
.B(n_161),
.Y(n_4924)
);

INVx2_ASAP7_75t_L g4925 ( 
.A(n_4706),
.Y(n_4925)
);

CKINVDCx20_ASAP7_75t_R g4926 ( 
.A(n_4608),
.Y(n_4926)
);

INVx4_ASAP7_75t_L g4927 ( 
.A(n_4648),
.Y(n_4927)
);

INVx2_ASAP7_75t_SL g4928 ( 
.A(n_4648),
.Y(n_4928)
);

INVx1_ASAP7_75t_L g4929 ( 
.A(n_4651),
.Y(n_4929)
);

CKINVDCx6p67_ASAP7_75t_R g4930 ( 
.A(n_4690),
.Y(n_4930)
);

OAI22x1_ASAP7_75t_L g4931 ( 
.A1(n_4713),
.A2(n_165),
.B1(n_163),
.B2(n_164),
.Y(n_4931)
);

INVx2_ASAP7_75t_L g4932 ( 
.A(n_4765),
.Y(n_4932)
);

INVx1_ASAP7_75t_L g4933 ( 
.A(n_4682),
.Y(n_4933)
);

INVx2_ASAP7_75t_SL g4934 ( 
.A(n_4648),
.Y(n_4934)
);

BUFx12f_ASAP7_75t_L g4935 ( 
.A(n_4610),
.Y(n_4935)
);

BUFx2_ASAP7_75t_SL g4936 ( 
.A(n_4606),
.Y(n_4936)
);

CKINVDCx6p67_ASAP7_75t_R g4937 ( 
.A(n_4642),
.Y(n_4937)
);

INVx1_ASAP7_75t_L g4938 ( 
.A(n_4685),
.Y(n_4938)
);

INVxp67_ASAP7_75t_SL g4939 ( 
.A(n_4797),
.Y(n_4939)
);

OAI22xp33_ASAP7_75t_L g4940 ( 
.A1(n_4730),
.A2(n_171),
.B1(n_167),
.B2(n_169),
.Y(n_4940)
);

BUFx6f_ASAP7_75t_L g4941 ( 
.A(n_4668),
.Y(n_4941)
);

OAI22xp5_ASAP7_75t_SL g4942 ( 
.A1(n_4664),
.A2(n_172),
.B1(n_167),
.B2(n_169),
.Y(n_4942)
);

OAI22xp33_ASAP7_75t_L g4943 ( 
.A1(n_4742),
.A2(n_175),
.B1(n_173),
.B2(n_174),
.Y(n_4943)
);

INVx4_ASAP7_75t_L g4944 ( 
.A(n_4668),
.Y(n_4944)
);

AOI21xp5_ASAP7_75t_L g4945 ( 
.A1(n_4580),
.A2(n_1867),
.B(n_1729),
.Y(n_4945)
);

INVx2_ASAP7_75t_L g4946 ( 
.A(n_4765),
.Y(n_4946)
);

INVx1_ASAP7_75t_L g4947 ( 
.A(n_4708),
.Y(n_4947)
);

INVx3_ASAP7_75t_L g4948 ( 
.A(n_4641),
.Y(n_4948)
);

OAI22xp5_ASAP7_75t_L g4949 ( 
.A1(n_4752),
.A2(n_175),
.B1(n_173),
.B2(n_174),
.Y(n_4949)
);

INVx1_ASAP7_75t_L g4950 ( 
.A(n_4734),
.Y(n_4950)
);

INVx1_ASAP7_75t_L g4951 ( 
.A(n_4596),
.Y(n_4951)
);

INVx2_ASAP7_75t_L g4952 ( 
.A(n_4763),
.Y(n_4952)
);

BUFx6f_ASAP7_75t_L g4953 ( 
.A(n_4668),
.Y(n_4953)
);

INVx1_ASAP7_75t_L g4954 ( 
.A(n_4581),
.Y(n_4954)
);

HB1xp67_ASAP7_75t_L g4955 ( 
.A(n_4725),
.Y(n_4955)
);

OAI22xp33_ASAP7_75t_L g4956 ( 
.A1(n_4742),
.A2(n_179),
.B1(n_176),
.B2(n_177),
.Y(n_4956)
);

INVx1_ASAP7_75t_SL g4957 ( 
.A(n_4618),
.Y(n_4957)
);

NAND2xp5_ASAP7_75t_L g4958 ( 
.A(n_4577),
.B(n_177),
.Y(n_4958)
);

INVx2_ASAP7_75t_L g4959 ( 
.A(n_4791),
.Y(n_4959)
);

BUFx2_ASAP7_75t_SL g4960 ( 
.A(n_4589),
.Y(n_4960)
);

CKINVDCx6p67_ASAP7_75t_R g4961 ( 
.A(n_4667),
.Y(n_4961)
);

INVx2_ASAP7_75t_L g4962 ( 
.A(n_4791),
.Y(n_4962)
);

INVx1_ASAP7_75t_L g4963 ( 
.A(n_4616),
.Y(n_4963)
);

BUFx3_ASAP7_75t_L g4964 ( 
.A(n_4675),
.Y(n_4964)
);

OAI22xp5_ASAP7_75t_L g4965 ( 
.A1(n_4735),
.A2(n_181),
.B1(n_179),
.B2(n_180),
.Y(n_4965)
);

OAI22xp5_ASAP7_75t_L g4966 ( 
.A1(n_4787),
.A2(n_185),
.B1(n_182),
.B2(n_184),
.Y(n_4966)
);

INVx5_ASAP7_75t_L g4967 ( 
.A(n_4791),
.Y(n_4967)
);

BUFx12f_ASAP7_75t_L g4968 ( 
.A(n_4652),
.Y(n_4968)
);

HB1xp67_ASAP7_75t_L g4969 ( 
.A(n_4757),
.Y(n_4969)
);

INVx6_ASAP7_75t_L g4970 ( 
.A(n_4675),
.Y(n_4970)
);

INVx2_ASAP7_75t_L g4971 ( 
.A(n_4776),
.Y(n_4971)
);

INVx1_ASAP7_75t_L g4972 ( 
.A(n_4780),
.Y(n_4972)
);

AOI22xp33_ASAP7_75t_L g4973 ( 
.A1(n_4560),
.A2(n_4629),
.B1(n_4615),
.B2(n_4793),
.Y(n_4973)
);

INVx1_ASAP7_75t_L g4974 ( 
.A(n_4800),
.Y(n_4974)
);

BUFx6f_ASAP7_75t_L g4975 ( 
.A(n_4675),
.Y(n_4975)
);

BUFx12f_ASAP7_75t_L g4976 ( 
.A(n_4760),
.Y(n_4976)
);

CKINVDCx5p33_ASAP7_75t_R g4977 ( 
.A(n_4623),
.Y(n_4977)
);

NAND2x1p5_ASAP7_75t_L g4978 ( 
.A(n_4620),
.B(n_1867),
.Y(n_4978)
);

BUFx6f_ASAP7_75t_L g4979 ( 
.A(n_4635),
.Y(n_4979)
);

INVx1_ASAP7_75t_L g4980 ( 
.A(n_4625),
.Y(n_4980)
);

AOI22xp33_ASAP7_75t_L g4981 ( 
.A1(n_4793),
.A2(n_185),
.B1(n_182),
.B2(n_184),
.Y(n_4981)
);

INVx4_ASAP7_75t_L g4982 ( 
.A(n_4620),
.Y(n_4982)
);

INVx2_ASAP7_75t_SL g4983 ( 
.A(n_4639),
.Y(n_4983)
);

INVx2_ASAP7_75t_L g4984 ( 
.A(n_4762),
.Y(n_4984)
);

AOI22xp33_ASAP7_75t_SL g4985 ( 
.A1(n_4740),
.A2(n_189),
.B1(n_186),
.B2(n_187),
.Y(n_4985)
);

INVx1_ASAP7_75t_L g4986 ( 
.A(n_4570),
.Y(n_4986)
);

INVx1_ASAP7_75t_SL g4987 ( 
.A(n_4680),
.Y(n_4987)
);

BUFx3_ASAP7_75t_L g4988 ( 
.A(n_4705),
.Y(n_4988)
);

BUFx2_ASAP7_75t_L g4989 ( 
.A(n_4705),
.Y(n_4989)
);

INVx2_ASAP7_75t_L g4990 ( 
.A(n_4726),
.Y(n_4990)
);

CKINVDCx11_ASAP7_75t_R g4991 ( 
.A(n_4674),
.Y(n_4991)
);

AOI22xp33_ASAP7_75t_L g4992 ( 
.A1(n_4789),
.A2(n_189),
.B1(n_186),
.B2(n_187),
.Y(n_4992)
);

BUFx6f_ASAP7_75t_L g4993 ( 
.A(n_4712),
.Y(n_4993)
);

INVx2_ASAP7_75t_L g4994 ( 
.A(n_4726),
.Y(n_4994)
);

INVx6_ASAP7_75t_L g4995 ( 
.A(n_4573),
.Y(n_4995)
);

OAI22xp5_ASAP7_75t_L g4996 ( 
.A1(n_4733),
.A2(n_192),
.B1(n_190),
.B2(n_191),
.Y(n_4996)
);

AOI22xp33_ASAP7_75t_L g4997 ( 
.A1(n_4779),
.A2(n_193),
.B1(n_191),
.B2(n_192),
.Y(n_4997)
);

BUFx8_ASAP7_75t_L g4998 ( 
.A(n_4695),
.Y(n_4998)
);

INVxp67_ASAP7_75t_SL g4999 ( 
.A(n_4804),
.Y(n_4999)
);

INVx3_ASAP7_75t_L g5000 ( 
.A(n_4644),
.Y(n_5000)
);

AND2x2_ASAP7_75t_L g5001 ( 
.A(n_4877),
.B(n_4563),
.Y(n_5001)
);

AOI21x1_ASAP7_75t_SL g5002 ( 
.A1(n_4832),
.A2(n_4844),
.B(n_4914),
.Y(n_5002)
);

NAND2xp5_ASAP7_75t_L g5003 ( 
.A(n_4829),
.B(n_4613),
.Y(n_5003)
);

O2A1O1Ixp33_ASAP7_75t_L g5004 ( 
.A1(n_4835),
.A2(n_4698),
.B(n_4755),
.C(n_4737),
.Y(n_5004)
);

AND2x2_ASAP7_75t_L g5005 ( 
.A(n_4825),
.B(n_4572),
.Y(n_5005)
);

AND2x2_ASAP7_75t_L g5006 ( 
.A(n_4847),
.B(n_4644),
.Y(n_5006)
);

AO21x2_ASAP7_75t_L g5007 ( 
.A1(n_4929),
.A2(n_4798),
.B(n_4715),
.Y(n_5007)
);

AND2x2_ASAP7_75t_L g5008 ( 
.A(n_4836),
.B(n_4781),
.Y(n_5008)
);

AND2x2_ASAP7_75t_L g5009 ( 
.A(n_4948),
.B(n_4775),
.Y(n_5009)
);

INVx1_ASAP7_75t_L g5010 ( 
.A(n_4811),
.Y(n_5010)
);

AND2x2_ASAP7_75t_L g5011 ( 
.A(n_4948),
.B(n_4638),
.Y(n_5011)
);

AND2x2_ASAP7_75t_L g5012 ( 
.A(n_4989),
.B(n_4638),
.Y(n_5012)
);

HB1xp67_ASAP7_75t_L g5013 ( 
.A(n_4955),
.Y(n_5013)
);

NAND2xp5_ASAP7_75t_L g5014 ( 
.A(n_4999),
.B(n_4802),
.Y(n_5014)
);

OAI22xp5_ASAP7_75t_SL g5015 ( 
.A1(n_4926),
.A2(n_4711),
.B1(n_4718),
.B2(n_4678),
.Y(n_5015)
);

AND2x2_ASAP7_75t_L g5016 ( 
.A(n_4809),
.B(n_4679),
.Y(n_5016)
);

NAND2xp5_ASAP7_75t_L g5017 ( 
.A(n_4833),
.B(n_4807),
.Y(n_5017)
);

HB1xp67_ASAP7_75t_L g5018 ( 
.A(n_4839),
.Y(n_5018)
);

AND2x2_ASAP7_75t_L g5019 ( 
.A(n_4870),
.B(n_4691),
.Y(n_5019)
);

NAND2xp5_ASAP7_75t_L g5020 ( 
.A(n_4950),
.B(n_4598),
.Y(n_5020)
);

AND2x4_ASAP7_75t_L g5021 ( 
.A(n_4870),
.B(n_4803),
.Y(n_5021)
);

HB1xp67_ASAP7_75t_L g5022 ( 
.A(n_4885),
.Y(n_5022)
);

NAND2xp5_ASAP7_75t_L g5023 ( 
.A(n_4826),
.B(n_4807),
.Y(n_5023)
);

OR2x2_ASAP7_75t_L g5024 ( 
.A(n_4827),
.B(n_4805),
.Y(n_5024)
);

AND2x2_ASAP7_75t_L g5025 ( 
.A(n_4988),
.B(n_4709),
.Y(n_5025)
);

AOI21xp5_ASAP7_75t_L g5026 ( 
.A1(n_4862),
.A2(n_4732),
.B(n_4681),
.Y(n_5026)
);

AOI21xp5_ASAP7_75t_L g5027 ( 
.A1(n_4924),
.A2(n_4575),
.B(n_4808),
.Y(n_5027)
);

INVx4_ASAP7_75t_L g5028 ( 
.A(n_4817),
.Y(n_5028)
);

AND2x4_ASAP7_75t_L g5029 ( 
.A(n_4959),
.B(n_4785),
.Y(n_5029)
);

AND2x2_ASAP7_75t_L g5030 ( 
.A(n_4837),
.B(n_4709),
.Y(n_5030)
);

AOI21xp5_ASAP7_75t_L g5031 ( 
.A1(n_4857),
.A2(n_4662),
.B(n_4806),
.Y(n_5031)
);

BUFx2_ASAP7_75t_L g5032 ( 
.A(n_4879),
.Y(n_5032)
);

AND2x2_ASAP7_75t_L g5033 ( 
.A(n_4855),
.B(n_4785),
.Y(n_5033)
);

BUFx2_ASAP7_75t_L g5034 ( 
.A(n_4979),
.Y(n_5034)
);

NAND2xp5_ASAP7_75t_L g5035 ( 
.A(n_4884),
.B(n_4807),
.Y(n_5035)
);

AND2x2_ASAP7_75t_L g5036 ( 
.A(n_4864),
.B(n_4743),
.Y(n_5036)
);

AND2x2_ASAP7_75t_L g5037 ( 
.A(n_4874),
.B(n_4743),
.Y(n_5037)
);

BUFx4f_ASAP7_75t_L g5038 ( 
.A(n_4819),
.Y(n_5038)
);

AND2x2_ASAP7_75t_L g5039 ( 
.A(n_4960),
.B(n_4617),
.Y(n_5039)
);

INVx1_ASAP7_75t_L g5040 ( 
.A(n_4811),
.Y(n_5040)
);

INVx1_ASAP7_75t_L g5041 ( 
.A(n_4863),
.Y(n_5041)
);

AND2x2_ASAP7_75t_L g5042 ( 
.A(n_4936),
.B(n_4766),
.Y(n_5042)
);

O2A1O1Ixp33_ASAP7_75t_L g5043 ( 
.A1(n_4878),
.A2(n_4659),
.B(n_4666),
.C(n_4657),
.Y(n_5043)
);

O2A1O1Ixp5_ASAP7_75t_L g5044 ( 
.A1(n_4943),
.A2(n_4587),
.B(n_4583),
.C(n_4693),
.Y(n_5044)
);

OA21x2_ASAP7_75t_L g5045 ( 
.A1(n_4990),
.A2(n_4645),
.B(n_4792),
.Y(n_5045)
);

OA21x2_ASAP7_75t_L g5046 ( 
.A1(n_4994),
.A2(n_4699),
.B(n_4720),
.Y(n_5046)
);

HB1xp67_ASAP7_75t_L g5047 ( 
.A(n_4894),
.Y(n_5047)
);

INVx1_ASAP7_75t_L g5048 ( 
.A(n_4815),
.Y(n_5048)
);

INVx2_ASAP7_75t_L g5049 ( 
.A(n_4984),
.Y(n_5049)
);

INVx2_ASAP7_75t_L g5050 ( 
.A(n_4969),
.Y(n_5050)
);

AOI21xp5_ASAP7_75t_L g5051 ( 
.A1(n_4843),
.A2(n_4759),
.B(n_4782),
.Y(n_5051)
);

AOI21x1_ASAP7_75t_SL g5052 ( 
.A1(n_4905),
.A2(n_4902),
.B(n_4891),
.Y(n_5052)
);

A2O1A1Ixp33_ASAP7_75t_L g5053 ( 
.A1(n_4883),
.A2(n_4670),
.B(n_4751),
.C(n_4590),
.Y(n_5053)
);

NAND2xp5_ASAP7_75t_L g5054 ( 
.A(n_4886),
.B(n_4892),
.Y(n_5054)
);

AOI21x1_ASAP7_75t_SL g5055 ( 
.A1(n_4840),
.A2(n_4654),
.B(n_4636),
.Y(n_5055)
);

A2O1A1Ixp33_ASAP7_75t_L g5056 ( 
.A1(n_4859),
.A2(n_4590),
.B(n_4703),
.C(n_4693),
.Y(n_5056)
);

HB1xp67_ASAP7_75t_L g5057 ( 
.A(n_4869),
.Y(n_5057)
);

CKINVDCx20_ASAP7_75t_R g5058 ( 
.A(n_4828),
.Y(n_5058)
);

INVx1_ASAP7_75t_L g5059 ( 
.A(n_4850),
.Y(n_5059)
);

BUFx3_ASAP7_75t_L g5060 ( 
.A(n_4854),
.Y(n_5060)
);

AOI21x1_ASAP7_75t_SL g5061 ( 
.A1(n_4958),
.A2(n_4663),
.B(n_4770),
.Y(n_5061)
);

AOI21xp5_ASAP7_75t_SL g5062 ( 
.A1(n_4831),
.A2(n_4605),
.B(n_4663),
.Y(n_5062)
);

AOI21xp5_ASAP7_75t_L g5063 ( 
.A1(n_4812),
.A2(n_4593),
.B(n_4568),
.Y(n_5063)
);

OAI22xp5_ASAP7_75t_L g5064 ( 
.A1(n_4882),
.A2(n_4579),
.B1(n_4703),
.B2(n_4770),
.Y(n_5064)
);

NAND2xp5_ASAP7_75t_L g5065 ( 
.A(n_4896),
.B(n_4773),
.Y(n_5065)
);

AOI21x1_ASAP7_75t_SL g5066 ( 
.A1(n_4890),
.A2(n_4579),
.B(n_4756),
.Y(n_5066)
);

INVx2_ASAP7_75t_L g5067 ( 
.A(n_4880),
.Y(n_5067)
);

OA21x2_ASAP7_75t_L g5068 ( 
.A1(n_4974),
.A2(n_4687),
.B(n_4784),
.Y(n_5068)
);

NAND2xp5_ASAP7_75t_L g5069 ( 
.A(n_4916),
.B(n_4786),
.Y(n_5069)
);

AND2x2_ASAP7_75t_SL g5070 ( 
.A(n_4831),
.B(n_4571),
.Y(n_5070)
);

O2A1O1Ixp33_ASAP7_75t_L g5071 ( 
.A1(n_4895),
.A2(n_4949),
.B(n_4956),
.C(n_4940),
.Y(n_5071)
);

INVx1_ASAP7_75t_L g5072 ( 
.A(n_4851),
.Y(n_5072)
);

NOR2xp67_ASAP7_75t_L g5073 ( 
.A(n_4867),
.B(n_4739),
.Y(n_5073)
);

OA21x2_ASAP7_75t_L g5074 ( 
.A1(n_4974),
.A2(n_4736),
.B(n_4728),
.Y(n_5074)
);

AOI21xp5_ASAP7_75t_L g5075 ( 
.A1(n_4816),
.A2(n_4756),
.B(n_4626),
.Y(n_5075)
);

AND2x2_ASAP7_75t_L g5076 ( 
.A(n_4818),
.B(n_4795),
.Y(n_5076)
);

AND2x2_ASAP7_75t_L g5077 ( 
.A(n_4856),
.B(n_4795),
.Y(n_5077)
);

O2A1O1Ixp5_ASAP7_75t_L g5078 ( 
.A1(n_4867),
.A2(n_4674),
.B(n_4684),
.C(n_4607),
.Y(n_5078)
);

INVx1_ASAP7_75t_L g5079 ( 
.A(n_4852),
.Y(n_5079)
);

INVx1_ASAP7_75t_L g5080 ( 
.A(n_4875),
.Y(n_5080)
);

CKINVDCx5p33_ASAP7_75t_R g5081 ( 
.A(n_4824),
.Y(n_5081)
);

NAND2xp5_ASAP7_75t_L g5082 ( 
.A(n_4939),
.B(n_4897),
.Y(n_5082)
);

AOI21x1_ASAP7_75t_SL g5083 ( 
.A1(n_4893),
.A2(n_4750),
.B(n_194),
.Y(n_5083)
);

AND2x2_ASAP7_75t_L g5084 ( 
.A(n_4904),
.B(n_4795),
.Y(n_5084)
);

BUFx3_ASAP7_75t_L g5085 ( 
.A(n_4860),
.Y(n_5085)
);

AND2x2_ASAP7_75t_L g5086 ( 
.A(n_4930),
.B(n_4671),
.Y(n_5086)
);

OAI22xp5_ASAP7_75t_L g5087 ( 
.A1(n_4942),
.A2(n_4771),
.B1(n_4719),
.B2(n_198),
.Y(n_5087)
);

NAND2xp5_ASAP7_75t_L g5088 ( 
.A(n_4901),
.B(n_195),
.Y(n_5088)
);

NOR2x1_ASAP7_75t_SL g5089 ( 
.A(n_4967),
.B(n_4834),
.Y(n_5089)
);

AND2x2_ASAP7_75t_L g5090 ( 
.A(n_4912),
.B(n_195),
.Y(n_5090)
);

AND2x2_ASAP7_75t_L g5091 ( 
.A(n_4954),
.B(n_197),
.Y(n_5091)
);

OAI22xp5_ASAP7_75t_L g5092 ( 
.A1(n_4913),
.A2(n_200),
.B1(n_197),
.B2(n_199),
.Y(n_5092)
);

O2A1O1Ixp33_ASAP7_75t_L g5093 ( 
.A1(n_4996),
.A2(n_202),
.B(n_199),
.C(n_200),
.Y(n_5093)
);

INVx2_ASAP7_75t_L g5094 ( 
.A(n_4909),
.Y(n_5094)
);

NOR2xp33_ASAP7_75t_R g5095 ( 
.A(n_4977),
.B(n_4991),
.Y(n_5095)
);

INVx2_ASAP7_75t_L g5096 ( 
.A(n_4917),
.Y(n_5096)
);

OAI22xp5_ASAP7_75t_L g5097 ( 
.A1(n_4920),
.A2(n_205),
.B1(n_203),
.B2(n_204),
.Y(n_5097)
);

AOI21xp5_ASAP7_75t_SL g5098 ( 
.A1(n_4841),
.A2(n_203),
.B(n_205),
.Y(n_5098)
);

AND2x2_ASAP7_75t_L g5099 ( 
.A(n_4951),
.B(n_206),
.Y(n_5099)
);

AOI21x1_ASAP7_75t_SL g5100 ( 
.A1(n_4872),
.A2(n_206),
.B(n_207),
.Y(n_5100)
);

O2A1O1Ixp33_ASAP7_75t_L g5101 ( 
.A1(n_4965),
.A2(n_211),
.B(n_209),
.C(n_210),
.Y(n_5101)
);

OAI22xp5_ASAP7_75t_L g5102 ( 
.A1(n_4922),
.A2(n_211),
.B1(n_209),
.B2(n_210),
.Y(n_5102)
);

O2A1O1Ixp33_ASAP7_75t_L g5103 ( 
.A1(n_4966),
.A2(n_215),
.B(n_212),
.C(n_214),
.Y(n_5103)
);

OA21x2_ASAP7_75t_L g5104 ( 
.A1(n_4932),
.A2(n_217),
.B(n_218),
.Y(n_5104)
);

AOI21xp5_ASAP7_75t_SL g5105 ( 
.A1(n_4982),
.A2(n_218),
.B(n_219),
.Y(n_5105)
);

INVxp33_ASAP7_75t_L g5106 ( 
.A(n_4810),
.Y(n_5106)
);

O2A1O1Ixp5_ASAP7_75t_L g5107 ( 
.A1(n_4962),
.A2(n_225),
.B(n_219),
.C(n_221),
.Y(n_5107)
);

INVx2_ASAP7_75t_L g5108 ( 
.A(n_4946),
.Y(n_5108)
);

NAND2x1_ASAP7_75t_L g5109 ( 
.A(n_5000),
.B(n_221),
.Y(n_5109)
);

AND2x2_ASAP7_75t_L g5110 ( 
.A(n_4903),
.B(n_225),
.Y(n_5110)
);

AND2x2_ASAP7_75t_L g5111 ( 
.A(n_4961),
.B(n_226),
.Y(n_5111)
);

INVx2_ASAP7_75t_L g5112 ( 
.A(n_4971),
.Y(n_5112)
);

AOI21x1_ASAP7_75t_SL g5113 ( 
.A1(n_4931),
.A2(n_226),
.B(n_230),
.Y(n_5113)
);

INVx1_ASAP7_75t_L g5114 ( 
.A(n_4881),
.Y(n_5114)
);

INVx1_ASAP7_75t_L g5115 ( 
.A(n_4868),
.Y(n_5115)
);

OAI22xp5_ASAP7_75t_L g5116 ( 
.A1(n_4985),
.A2(n_233),
.B1(n_231),
.B2(n_232),
.Y(n_5116)
);

AND2x2_ASAP7_75t_L g5117 ( 
.A(n_4937),
.B(n_234),
.Y(n_5117)
);

OA21x2_ASAP7_75t_L g5118 ( 
.A1(n_4868),
.A2(n_235),
.B(n_236),
.Y(n_5118)
);

OA21x2_ASAP7_75t_L g5119 ( 
.A1(n_4972),
.A2(n_235),
.B(n_239),
.Y(n_5119)
);

NOR3xp33_ASAP7_75t_L g5120 ( 
.A(n_4887),
.B(n_239),
.C(n_240),
.Y(n_5120)
);

CKINVDCx5p33_ASAP7_75t_R g5121 ( 
.A(n_4814),
.Y(n_5121)
);

BUFx10_ASAP7_75t_L g5122 ( 
.A(n_4819),
.Y(n_5122)
);

OR2x2_ASAP7_75t_L g5123 ( 
.A(n_4972),
.B(n_241),
.Y(n_5123)
);

AND2x2_ASAP7_75t_L g5124 ( 
.A(n_4987),
.B(n_241),
.Y(n_5124)
);

AND2x2_ASAP7_75t_L g5125 ( 
.A(n_4986),
.B(n_244),
.Y(n_5125)
);

OR2x2_ASAP7_75t_L g5126 ( 
.A(n_4925),
.B(n_244),
.Y(n_5126)
);

CKINVDCx5p33_ASAP7_75t_R g5127 ( 
.A(n_4814),
.Y(n_5127)
);

INVx1_ASAP7_75t_SL g5128 ( 
.A(n_4957),
.Y(n_5128)
);

INVx1_ASAP7_75t_L g5129 ( 
.A(n_4933),
.Y(n_5129)
);

NAND2xp5_ASAP7_75t_L g5130 ( 
.A(n_4963),
.B(n_245),
.Y(n_5130)
);

INVx1_ASAP7_75t_L g5131 ( 
.A(n_4933),
.Y(n_5131)
);

CKINVDCx5p33_ASAP7_75t_R g5132 ( 
.A(n_4853),
.Y(n_5132)
);

INVx3_ASAP7_75t_L g5133 ( 
.A(n_4982),
.Y(n_5133)
);

OA21x2_ASAP7_75t_L g5134 ( 
.A1(n_4938),
.A2(n_245),
.B(n_246),
.Y(n_5134)
);

INVx1_ASAP7_75t_L g5135 ( 
.A(n_4938),
.Y(n_5135)
);

CKINVDCx5p33_ASAP7_75t_R g5136 ( 
.A(n_4830),
.Y(n_5136)
);

AND2x2_ASAP7_75t_SL g5137 ( 
.A(n_4973),
.B(n_247),
.Y(n_5137)
);

INVx1_ASAP7_75t_L g5138 ( 
.A(n_4952),
.Y(n_5138)
);

AND2x2_ASAP7_75t_L g5139 ( 
.A(n_4993),
.B(n_247),
.Y(n_5139)
);

INVx1_ASAP7_75t_L g5140 ( 
.A(n_4947),
.Y(n_5140)
);

AOI21xp5_ASAP7_75t_SL g5141 ( 
.A1(n_4908),
.A2(n_249),
.B(n_250),
.Y(n_5141)
);

BUFx6f_ASAP7_75t_L g5142 ( 
.A(n_4823),
.Y(n_5142)
);

AND2x4_ASAP7_75t_L g5143 ( 
.A(n_5000),
.B(n_249),
.Y(n_5143)
);

AND2x2_ASAP7_75t_L g5144 ( 
.A(n_4993),
.B(n_251),
.Y(n_5144)
);

CKINVDCx20_ASAP7_75t_R g5145 ( 
.A(n_4889),
.Y(n_5145)
);

AND2x2_ASAP7_75t_L g5146 ( 
.A(n_4993),
.B(n_252),
.Y(n_5146)
);

INVx3_ASAP7_75t_L g5147 ( 
.A(n_4979),
.Y(n_5147)
);

AND2x2_ASAP7_75t_L g5148 ( 
.A(n_4838),
.B(n_253),
.Y(n_5148)
);

NOR2xp33_ASAP7_75t_R g5149 ( 
.A(n_5081),
.B(n_5145),
.Y(n_5149)
);

OR2x6_ASAP7_75t_L g5150 ( 
.A(n_5062),
.B(n_4838),
.Y(n_5150)
);

INVx1_ASAP7_75t_L g5151 ( 
.A(n_5115),
.Y(n_5151)
);

CKINVDCx14_ASAP7_75t_R g5152 ( 
.A(n_5095),
.Y(n_5152)
);

CKINVDCx16_ASAP7_75t_R g5153 ( 
.A(n_5058),
.Y(n_5153)
);

NAND2xp33_ASAP7_75t_R g5154 ( 
.A(n_5121),
.B(n_5127),
.Y(n_5154)
);

NOR2xp33_ASAP7_75t_R g5155 ( 
.A(n_5136),
.B(n_4830),
.Y(n_5155)
);

AO31x2_ASAP7_75t_L g5156 ( 
.A1(n_5089),
.A2(n_4927),
.A3(n_4944),
.B(n_4898),
.Y(n_5156)
);

HB1xp67_ASAP7_75t_L g5157 ( 
.A(n_5022),
.Y(n_5157)
);

AOI21xp33_ASAP7_75t_L g5158 ( 
.A1(n_5004),
.A2(n_4980),
.B(n_4858),
.Y(n_5158)
);

NOR2xp33_ASAP7_75t_R g5159 ( 
.A(n_5132),
.B(n_5038),
.Y(n_5159)
);

CKINVDCx5p33_ASAP7_75t_R g5160 ( 
.A(n_5060),
.Y(n_5160)
);

NOR3xp33_ASAP7_75t_SL g5161 ( 
.A(n_5031),
.B(n_4813),
.C(n_4945),
.Y(n_5161)
);

INVx1_ASAP7_75t_L g5162 ( 
.A(n_5018),
.Y(n_5162)
);

NOR3xp33_ASAP7_75t_SL g5163 ( 
.A(n_5015),
.B(n_4923),
.C(n_4899),
.Y(n_5163)
);

INVx2_ASAP7_75t_L g5164 ( 
.A(n_5108),
.Y(n_5164)
);

OR2x6_ASAP7_75t_L g5165 ( 
.A(n_5075),
.B(n_4976),
.Y(n_5165)
);

INVx1_ASAP7_75t_SL g5166 ( 
.A(n_5128),
.Y(n_5166)
);

AND3x2_ASAP7_75t_L g5167 ( 
.A(n_5098),
.B(n_4899),
.C(n_4998),
.Y(n_5167)
);

INVx2_ASAP7_75t_L g5168 ( 
.A(n_5033),
.Y(n_5168)
);

NOR2xp33_ASAP7_75t_R g5169 ( 
.A(n_5038),
.B(n_4998),
.Y(n_5169)
);

CKINVDCx16_ASAP7_75t_R g5170 ( 
.A(n_5085),
.Y(n_5170)
);

OR2x6_ASAP7_75t_L g5171 ( 
.A(n_5028),
.B(n_4935),
.Y(n_5171)
);

INVx2_ASAP7_75t_L g5172 ( 
.A(n_5024),
.Y(n_5172)
);

AND2x2_ASAP7_75t_L g5173 ( 
.A(n_5032),
.B(n_4983),
.Y(n_5173)
);

NAND2xp33_ASAP7_75t_R g5174 ( 
.A(n_5111),
.B(n_253),
.Y(n_5174)
);

INVx1_ASAP7_75t_SL g5175 ( 
.A(n_5128),
.Y(n_5175)
);

BUFx2_ASAP7_75t_L g5176 ( 
.A(n_5021),
.Y(n_5176)
);

BUFx6f_ASAP7_75t_L g5177 ( 
.A(n_5122),
.Y(n_5177)
);

AND2x4_ASAP7_75t_L g5178 ( 
.A(n_5133),
.B(n_5021),
.Y(n_5178)
);

AND2x2_ASAP7_75t_L g5179 ( 
.A(n_5006),
.B(n_4995),
.Y(n_5179)
);

NAND2x1p5_ASAP7_75t_L g5180 ( 
.A(n_5133),
.B(n_5030),
.Y(n_5180)
);

NAND3xp33_ASAP7_75t_SL g5181 ( 
.A(n_5026),
.B(n_4845),
.C(n_4907),
.Y(n_5181)
);

AND2x2_ASAP7_75t_L g5182 ( 
.A(n_5011),
.B(n_4995),
.Y(n_5182)
);

AND2x2_ASAP7_75t_L g5183 ( 
.A(n_5012),
.B(n_4979),
.Y(n_5183)
);

CKINVDCx20_ASAP7_75t_R g5184 ( 
.A(n_5028),
.Y(n_5184)
);

NOR2xp33_ASAP7_75t_R g5185 ( 
.A(n_5070),
.B(n_4968),
.Y(n_5185)
);

AND2x2_ASAP7_75t_L g5186 ( 
.A(n_5001),
.B(n_4964),
.Y(n_5186)
);

INVx2_ASAP7_75t_L g5187 ( 
.A(n_5010),
.Y(n_5187)
);

INVx2_ASAP7_75t_L g5188 ( 
.A(n_5040),
.Y(n_5188)
);

NOR3xp33_ASAP7_75t_SL g5189 ( 
.A(n_5015),
.B(n_4888),
.C(n_4820),
.Y(n_5189)
);

INVx1_ASAP7_75t_SL g5190 ( 
.A(n_5034),
.Y(n_5190)
);

INVx2_ASAP7_75t_L g5191 ( 
.A(n_5050),
.Y(n_5191)
);

INVx1_ASAP7_75t_L g5192 ( 
.A(n_5041),
.Y(n_5192)
);

INVx1_ASAP7_75t_L g5193 ( 
.A(n_5059),
.Y(n_5193)
);

CKINVDCx5p33_ASAP7_75t_R g5194 ( 
.A(n_5122),
.Y(n_5194)
);

INVx1_ASAP7_75t_L g5195 ( 
.A(n_5129),
.Y(n_5195)
);

AND2x2_ASAP7_75t_L g5196 ( 
.A(n_5019),
.B(n_4967),
.Y(n_5196)
);

NAND2xp33_ASAP7_75t_R g5197 ( 
.A(n_5117),
.B(n_254),
.Y(n_5197)
);

INVx1_ASAP7_75t_L g5198 ( 
.A(n_5072),
.Y(n_5198)
);

INVx1_ASAP7_75t_L g5199 ( 
.A(n_5079),
.Y(n_5199)
);

NOR2xp33_ASAP7_75t_L g5200 ( 
.A(n_5043),
.B(n_4927),
.Y(n_5200)
);

NAND2xp5_ASAP7_75t_L g5201 ( 
.A(n_5014),
.B(n_5020),
.Y(n_5201)
);

INVx2_ASAP7_75t_L g5202 ( 
.A(n_5112),
.Y(n_5202)
);

NOR2xp33_ASAP7_75t_R g5203 ( 
.A(n_5137),
.B(n_4906),
.Y(n_5203)
);

BUFx6f_ASAP7_75t_L g5204 ( 
.A(n_5109),
.Y(n_5204)
);

INVx1_ASAP7_75t_L g5205 ( 
.A(n_5080),
.Y(n_5205)
);

NAND2xp5_ASAP7_75t_L g5206 ( 
.A(n_5014),
.B(n_4928),
.Y(n_5206)
);

CKINVDCx5p33_ASAP7_75t_R g5207 ( 
.A(n_5142),
.Y(n_5207)
);

INVx1_ASAP7_75t_L g5208 ( 
.A(n_5114),
.Y(n_5208)
);

AND2x2_ASAP7_75t_L g5209 ( 
.A(n_5005),
.B(n_4967),
.Y(n_5209)
);

AND2x2_ASAP7_75t_L g5210 ( 
.A(n_5076),
.B(n_4934),
.Y(n_5210)
);

INVx1_ASAP7_75t_L g5211 ( 
.A(n_5131),
.Y(n_5211)
);

AOI22xp33_ASAP7_75t_L g5212 ( 
.A1(n_5120),
.A2(n_4919),
.B1(n_4871),
.B2(n_4910),
.Y(n_5212)
);

INVx2_ASAP7_75t_L g5213 ( 
.A(n_5009),
.Y(n_5213)
);

INVx2_ASAP7_75t_L g5214 ( 
.A(n_5049),
.Y(n_5214)
);

OAI22xp5_ASAP7_75t_SL g5215 ( 
.A1(n_5064),
.A2(n_4997),
.B1(n_4981),
.B2(n_4900),
.Y(n_5215)
);

INVx2_ASAP7_75t_L g5216 ( 
.A(n_5067),
.Y(n_5216)
);

NAND2xp33_ASAP7_75t_R g5217 ( 
.A(n_5143),
.B(n_254),
.Y(n_5217)
);

BUFx6f_ASAP7_75t_L g5218 ( 
.A(n_5142),
.Y(n_5218)
);

NAND2xp5_ASAP7_75t_L g5219 ( 
.A(n_5003),
.B(n_4944),
.Y(n_5219)
);

AND2x4_ASAP7_75t_L g5220 ( 
.A(n_5042),
.B(n_5077),
.Y(n_5220)
);

INVx2_ASAP7_75t_L g5221 ( 
.A(n_5094),
.Y(n_5221)
);

NOR2xp33_ASAP7_75t_R g5222 ( 
.A(n_5086),
.B(n_5139),
.Y(n_5222)
);

AND2x2_ASAP7_75t_L g5223 ( 
.A(n_5016),
.B(n_4842),
.Y(n_5223)
);

OAI21x1_ASAP7_75t_L g5224 ( 
.A1(n_5023),
.A2(n_4873),
.B(n_4846),
.Y(n_5224)
);

NAND2xp5_ASAP7_75t_L g5225 ( 
.A(n_5003),
.B(n_4823),
.Y(n_5225)
);

CKINVDCx16_ASAP7_75t_R g5226 ( 
.A(n_5039),
.Y(n_5226)
);

O2A1O1Ixp33_ASAP7_75t_L g5227 ( 
.A1(n_5071),
.A2(n_4866),
.B(n_4861),
.C(n_4992),
.Y(n_5227)
);

INVx2_ASAP7_75t_L g5228 ( 
.A(n_5096),
.Y(n_5228)
);

AOI21x1_ASAP7_75t_L g5229 ( 
.A1(n_5130),
.A2(n_4911),
.B(n_4842),
.Y(n_5229)
);

XNOR2xp5_ASAP7_75t_L g5230 ( 
.A(n_5106),
.B(n_5110),
.Y(n_5230)
);

NAND2xp5_ASAP7_75t_L g5231 ( 
.A(n_5048),
.B(n_5057),
.Y(n_5231)
);

BUFx4f_ASAP7_75t_SL g5232 ( 
.A(n_5148),
.Y(n_5232)
);

AND2x2_ASAP7_75t_L g5233 ( 
.A(n_5084),
.B(n_4911),
.Y(n_5233)
);

AO31x2_ASAP7_75t_L g5234 ( 
.A1(n_5017),
.A2(n_5023),
.A3(n_5035),
.B(n_5069),
.Y(n_5234)
);

AOI22xp33_ASAP7_75t_L g5235 ( 
.A1(n_5092),
.A2(n_4822),
.B1(n_4848),
.B2(n_4918),
.Y(n_5235)
);

AOI22xp33_ASAP7_75t_SL g5236 ( 
.A1(n_5064),
.A2(n_4921),
.B1(n_4970),
.B2(n_4915),
.Y(n_5236)
);

OR2x6_ASAP7_75t_L g5237 ( 
.A(n_5105),
.B(n_4915),
.Y(n_5237)
);

AOI21xp33_ASAP7_75t_L g5238 ( 
.A1(n_5044),
.A2(n_4876),
.B(n_4849),
.Y(n_5238)
);

INVx2_ASAP7_75t_L g5239 ( 
.A(n_5138),
.Y(n_5239)
);

OAI22xp5_ASAP7_75t_L g5240 ( 
.A1(n_5053),
.A2(n_4970),
.B1(n_4921),
.B2(n_4823),
.Y(n_5240)
);

NAND2xp5_ASAP7_75t_SL g5241 ( 
.A(n_5025),
.B(n_5142),
.Y(n_5241)
);

INVx1_ASAP7_75t_L g5242 ( 
.A(n_5135),
.Y(n_5242)
);

AOI21xp33_ASAP7_75t_L g5243 ( 
.A1(n_5093),
.A2(n_4941),
.B(n_4865),
.Y(n_5243)
);

A2O1A1Ixp33_ASAP7_75t_L g5244 ( 
.A1(n_5051),
.A2(n_5101),
.B(n_5103),
.C(n_5056),
.Y(n_5244)
);

INVx8_ASAP7_75t_L g5245 ( 
.A(n_5143),
.Y(n_5245)
);

CKINVDCx20_ASAP7_75t_R g5246 ( 
.A(n_5090),
.Y(n_5246)
);

AOI22xp33_ASAP7_75t_L g5247 ( 
.A1(n_5092),
.A2(n_4821),
.B1(n_4941),
.B2(n_4865),
.Y(n_5247)
);

NAND2xp33_ASAP7_75t_R g5248 ( 
.A(n_5144),
.B(n_256),
.Y(n_5248)
);

AOI22xp33_ASAP7_75t_L g5249 ( 
.A1(n_5097),
.A2(n_4941),
.B1(n_4953),
.B2(n_4865),
.Y(n_5249)
);

INVx1_ASAP7_75t_L g5250 ( 
.A(n_5140),
.Y(n_5250)
);

NOR2xp33_ASAP7_75t_L g5251 ( 
.A(n_5130),
.B(n_5146),
.Y(n_5251)
);

NAND2xp5_ASAP7_75t_L g5252 ( 
.A(n_5008),
.B(n_4953),
.Y(n_5252)
);

INVx2_ASAP7_75t_L g5253 ( 
.A(n_5029),
.Y(n_5253)
);

BUFx2_ASAP7_75t_L g5254 ( 
.A(n_5013),
.Y(n_5254)
);

AND2x2_ASAP7_75t_L g5255 ( 
.A(n_5036),
.B(n_4953),
.Y(n_5255)
);

AOI21xp33_ASAP7_75t_L g5256 ( 
.A1(n_5097),
.A2(n_4975),
.B(n_4978),
.Y(n_5256)
);

INVx1_ASAP7_75t_L g5257 ( 
.A(n_5082),
.Y(n_5257)
);

HB1xp67_ASAP7_75t_L g5258 ( 
.A(n_5082),
.Y(n_5258)
);

CKINVDCx5p33_ASAP7_75t_R g5259 ( 
.A(n_5147),
.Y(n_5259)
);

NAND2xp33_ASAP7_75t_SL g5260 ( 
.A(n_5124),
.B(n_4975),
.Y(n_5260)
);

AOI22xp33_ASAP7_75t_SL g5261 ( 
.A1(n_5102),
.A2(n_5116),
.B1(n_5087),
.B2(n_5027),
.Y(n_5261)
);

NOR2xp33_ASAP7_75t_R g5262 ( 
.A(n_5091),
.B(n_257),
.Y(n_5262)
);

CKINVDCx5p33_ASAP7_75t_R g5263 ( 
.A(n_5147),
.Y(n_5263)
);

INVx1_ASAP7_75t_L g5264 ( 
.A(n_5054),
.Y(n_5264)
);

INVx2_ASAP7_75t_L g5265 ( 
.A(n_5029),
.Y(n_5265)
);

OR2x6_ASAP7_75t_L g5266 ( 
.A(n_5141),
.B(n_4975),
.Y(n_5266)
);

INVx2_ASAP7_75t_L g5267 ( 
.A(n_5047),
.Y(n_5267)
);

HB1xp67_ASAP7_75t_L g5268 ( 
.A(n_5035),
.Y(n_5268)
);

INVx2_ASAP7_75t_L g5269 ( 
.A(n_5037),
.Y(n_5269)
);

NAND2xp5_ASAP7_75t_L g5270 ( 
.A(n_5088),
.B(n_257),
.Y(n_5270)
);

O2A1O1Ixp33_ASAP7_75t_SL g5271 ( 
.A1(n_5102),
.A2(n_260),
.B(n_258),
.C(n_259),
.Y(n_5271)
);

INVx2_ASAP7_75t_L g5272 ( 
.A(n_5054),
.Y(n_5272)
);

NOR3xp33_ASAP7_75t_SL g5273 ( 
.A(n_5116),
.B(n_260),
.C(n_261),
.Y(n_5273)
);

AND2x2_ASAP7_75t_L g5274 ( 
.A(n_5099),
.B(n_262),
.Y(n_5274)
);

AND2x4_ASAP7_75t_L g5275 ( 
.A(n_5126),
.B(n_263),
.Y(n_5275)
);

CKINVDCx5p33_ASAP7_75t_R g5276 ( 
.A(n_5125),
.Y(n_5276)
);

AND2x2_ASAP7_75t_L g5277 ( 
.A(n_5017),
.B(n_265),
.Y(n_5277)
);

AOI22xp5_ASAP7_75t_L g5278 ( 
.A1(n_5087),
.A2(n_268),
.B1(n_266),
.B2(n_267),
.Y(n_5278)
);

INVx1_ASAP7_75t_L g5279 ( 
.A(n_5065),
.Y(n_5279)
);

INVx1_ASAP7_75t_L g5280 ( 
.A(n_5065),
.Y(n_5280)
);

AOI22xp33_ASAP7_75t_L g5281 ( 
.A1(n_5063),
.A2(n_270),
.B1(n_266),
.B2(n_269),
.Y(n_5281)
);

NOR2xp33_ASAP7_75t_R g5282 ( 
.A(n_5123),
.B(n_269),
.Y(n_5282)
);

INVx2_ASAP7_75t_L g5283 ( 
.A(n_5069),
.Y(n_5283)
);

OR2x2_ASAP7_75t_L g5284 ( 
.A(n_5088),
.B(n_271),
.Y(n_5284)
);

NAND2x1p5_ASAP7_75t_L g5285 ( 
.A(n_5104),
.B(n_1712),
.Y(n_5285)
);

OR2x6_ASAP7_75t_SL g5286 ( 
.A(n_5052),
.B(n_272),
.Y(n_5286)
);

NOR2xp33_ASAP7_75t_R g5287 ( 
.A(n_5100),
.B(n_272),
.Y(n_5287)
);

OR2x2_ASAP7_75t_L g5288 ( 
.A(n_5007),
.B(n_5134),
.Y(n_5288)
);

INVx2_ASAP7_75t_L g5289 ( 
.A(n_5104),
.Y(n_5289)
);

HB1xp67_ASAP7_75t_L g5290 ( 
.A(n_5134),
.Y(n_5290)
);

BUFx6f_ASAP7_75t_L g5291 ( 
.A(n_5119),
.Y(n_5291)
);

INVx2_ASAP7_75t_L g5292 ( 
.A(n_5119),
.Y(n_5292)
);

AND2x2_ASAP7_75t_L g5293 ( 
.A(n_5220),
.B(n_5118),
.Y(n_5293)
);

AND2x2_ASAP7_75t_L g5294 ( 
.A(n_5220),
.B(n_5180),
.Y(n_5294)
);

OR2x2_ASAP7_75t_L g5295 ( 
.A(n_5201),
.B(n_5118),
.Y(n_5295)
);

AOI22xp33_ASAP7_75t_SL g5296 ( 
.A1(n_5215),
.A2(n_5113),
.B1(n_5007),
.B2(n_5074),
.Y(n_5296)
);

INVx1_ASAP7_75t_L g5297 ( 
.A(n_5151),
.Y(n_5297)
);

NOR2x1_ASAP7_75t_L g5298 ( 
.A(n_5150),
.B(n_5073),
.Y(n_5298)
);

INVx2_ASAP7_75t_L g5299 ( 
.A(n_5218),
.Y(n_5299)
);

AOI22xp33_ASAP7_75t_L g5300 ( 
.A1(n_5261),
.A2(n_5074),
.B1(n_5046),
.B2(n_5045),
.Y(n_5300)
);

AND2x4_ASAP7_75t_L g5301 ( 
.A(n_5150),
.B(n_5061),
.Y(n_5301)
);

OR2x2_ASAP7_75t_L g5302 ( 
.A(n_5258),
.B(n_5257),
.Y(n_5302)
);

OA21x2_ASAP7_75t_L g5303 ( 
.A1(n_5224),
.A2(n_5078),
.B(n_5107),
.Y(n_5303)
);

AND2x2_ASAP7_75t_L g5304 ( 
.A(n_5226),
.B(n_5068),
.Y(n_5304)
);

INVx1_ASAP7_75t_L g5305 ( 
.A(n_5250),
.Y(n_5305)
);

AND2x2_ASAP7_75t_L g5306 ( 
.A(n_5176),
.B(n_5068),
.Y(n_5306)
);

INVx1_ASAP7_75t_L g5307 ( 
.A(n_5192),
.Y(n_5307)
);

NOR2xp33_ASAP7_75t_L g5308 ( 
.A(n_5152),
.B(n_273),
.Y(n_5308)
);

AND2x2_ASAP7_75t_L g5309 ( 
.A(n_5178),
.B(n_5045),
.Y(n_5309)
);

OR2x2_ASAP7_75t_L g5310 ( 
.A(n_5267),
.B(n_5046),
.Y(n_5310)
);

OAI221xp5_ASAP7_75t_L g5311 ( 
.A1(n_5244),
.A2(n_5083),
.B1(n_5002),
.B2(n_5055),
.C(n_5066),
.Y(n_5311)
);

OA21x2_ASAP7_75t_L g5312 ( 
.A1(n_5292),
.A2(n_273),
.B(n_274),
.Y(n_5312)
);

AO21x1_ASAP7_75t_L g5313 ( 
.A1(n_5174),
.A2(n_275),
.B(n_276),
.Y(n_5313)
);

BUFx2_ASAP7_75t_L g5314 ( 
.A(n_5185),
.Y(n_5314)
);

OR2x2_ASAP7_75t_L g5315 ( 
.A(n_5166),
.B(n_275),
.Y(n_5315)
);

OAI21xp5_ASAP7_75t_L g5316 ( 
.A1(n_5189),
.A2(n_276),
.B(n_277),
.Y(n_5316)
);

AO21x2_ASAP7_75t_L g5317 ( 
.A1(n_5290),
.A2(n_279),
.B(n_280),
.Y(n_5317)
);

INVx1_ASAP7_75t_L g5318 ( 
.A(n_5193),
.Y(n_5318)
);

INVx2_ASAP7_75t_L g5319 ( 
.A(n_5218),
.Y(n_5319)
);

AND2x2_ASAP7_75t_L g5320 ( 
.A(n_5178),
.B(n_279),
.Y(n_5320)
);

AND2x2_ASAP7_75t_L g5321 ( 
.A(n_5196),
.B(n_280),
.Y(n_5321)
);

INVx2_ASAP7_75t_L g5322 ( 
.A(n_5218),
.Y(n_5322)
);

NAND3xp33_ASAP7_75t_L g5323 ( 
.A(n_5273),
.B(n_5278),
.C(n_5158),
.Y(n_5323)
);

INVx1_ASAP7_75t_L g5324 ( 
.A(n_5198),
.Y(n_5324)
);

OA21x2_ASAP7_75t_L g5325 ( 
.A1(n_5289),
.A2(n_281),
.B(n_282),
.Y(n_5325)
);

AOI21xp5_ASAP7_75t_L g5326 ( 
.A1(n_5238),
.A2(n_281),
.B(n_282),
.Y(n_5326)
);

AND2x2_ASAP7_75t_L g5327 ( 
.A(n_5165),
.B(n_283),
.Y(n_5327)
);

INVx2_ASAP7_75t_L g5328 ( 
.A(n_5253),
.Y(n_5328)
);

INVx4_ASAP7_75t_L g5329 ( 
.A(n_5177),
.Y(n_5329)
);

HB1xp67_ASAP7_75t_L g5330 ( 
.A(n_5291),
.Y(n_5330)
);

INVx2_ASAP7_75t_L g5331 ( 
.A(n_5265),
.Y(n_5331)
);

INVx1_ASAP7_75t_L g5332 ( 
.A(n_5199),
.Y(n_5332)
);

INVx3_ASAP7_75t_L g5333 ( 
.A(n_5177),
.Y(n_5333)
);

OAI221xp5_ASAP7_75t_L g5334 ( 
.A1(n_5197),
.A2(n_285),
.B1(n_283),
.B2(n_284),
.C(n_286),
.Y(n_5334)
);

AND2x2_ASAP7_75t_L g5335 ( 
.A(n_5165),
.B(n_284),
.Y(n_5335)
);

INVx2_ASAP7_75t_L g5336 ( 
.A(n_5204),
.Y(n_5336)
);

INVx4_ASAP7_75t_L g5337 ( 
.A(n_5177),
.Y(n_5337)
);

BUFx3_ASAP7_75t_L g5338 ( 
.A(n_5184),
.Y(n_5338)
);

AO21x2_ASAP7_75t_L g5339 ( 
.A1(n_5288),
.A2(n_5277),
.B(n_5282),
.Y(n_5339)
);

INVx1_ASAP7_75t_L g5340 ( 
.A(n_5205),
.Y(n_5340)
);

OAI322xp33_ASAP7_75t_L g5341 ( 
.A1(n_5248),
.A2(n_285),
.A3(n_287),
.B1(n_288),
.B2(n_289),
.C1(n_290),
.C2(n_291),
.Y(n_5341)
);

INVx3_ASAP7_75t_L g5342 ( 
.A(n_5156),
.Y(n_5342)
);

AND2x2_ASAP7_75t_L g5343 ( 
.A(n_5209),
.B(n_287),
.Y(n_5343)
);

INVx2_ASAP7_75t_L g5344 ( 
.A(n_5204),
.Y(n_5344)
);

AOI33xp33_ASAP7_75t_L g5345 ( 
.A1(n_5167),
.A2(n_288),
.A3(n_289),
.B1(n_291),
.B2(n_292),
.B3(n_293),
.Y(n_5345)
);

OAI22xp5_ASAP7_75t_L g5346 ( 
.A1(n_5286),
.A2(n_295),
.B1(n_293),
.B2(n_294),
.Y(n_5346)
);

INVx1_ASAP7_75t_L g5347 ( 
.A(n_5208),
.Y(n_5347)
);

OR2x6_ASAP7_75t_L g5348 ( 
.A(n_5171),
.B(n_295),
.Y(n_5348)
);

AND2x4_ASAP7_75t_L g5349 ( 
.A(n_5156),
.B(n_296),
.Y(n_5349)
);

INVx1_ASAP7_75t_L g5350 ( 
.A(n_5195),
.Y(n_5350)
);

AND2x2_ASAP7_75t_L g5351 ( 
.A(n_5190),
.B(n_297),
.Y(n_5351)
);

AND2x2_ASAP7_75t_L g5352 ( 
.A(n_5213),
.B(n_297),
.Y(n_5352)
);

INVx2_ASAP7_75t_L g5353 ( 
.A(n_5204),
.Y(n_5353)
);

NAND2xp5_ASAP7_75t_SL g5354 ( 
.A(n_5236),
.B(n_1867),
.Y(n_5354)
);

INVxp67_ASAP7_75t_SL g5355 ( 
.A(n_5291),
.Y(n_5355)
);

INVx2_ASAP7_75t_L g5356 ( 
.A(n_5229),
.Y(n_5356)
);

INVx2_ASAP7_75t_L g5357 ( 
.A(n_5164),
.Y(n_5357)
);

OA21x2_ASAP7_75t_L g5358 ( 
.A1(n_5163),
.A2(n_298),
.B(n_299),
.Y(n_5358)
);

INVx1_ASAP7_75t_L g5359 ( 
.A(n_5195),
.Y(n_5359)
);

AND2x2_ASAP7_75t_L g5360 ( 
.A(n_5269),
.B(n_5168),
.Y(n_5360)
);

INVx1_ASAP7_75t_L g5361 ( 
.A(n_5211),
.Y(n_5361)
);

OR2x2_ASAP7_75t_L g5362 ( 
.A(n_5175),
.B(n_298),
.Y(n_5362)
);

INVx2_ASAP7_75t_L g5363 ( 
.A(n_5216),
.Y(n_5363)
);

INVx1_ASAP7_75t_L g5364 ( 
.A(n_5242),
.Y(n_5364)
);

BUFx2_ASAP7_75t_L g5365 ( 
.A(n_5171),
.Y(n_5365)
);

INVx1_ASAP7_75t_SL g5366 ( 
.A(n_5260),
.Y(n_5366)
);

AND2x2_ASAP7_75t_L g5367 ( 
.A(n_5233),
.B(n_299),
.Y(n_5367)
);

AO21x2_ASAP7_75t_L g5368 ( 
.A1(n_5268),
.A2(n_5270),
.B(n_5181),
.Y(n_5368)
);

HB1xp67_ASAP7_75t_L g5369 ( 
.A(n_5291),
.Y(n_5369)
);

OA21x2_ASAP7_75t_L g5370 ( 
.A1(n_5219),
.A2(n_301),
.B(n_302),
.Y(n_5370)
);

NOR2xp33_ASAP7_75t_L g5371 ( 
.A(n_5170),
.B(n_301),
.Y(n_5371)
);

INVx1_ASAP7_75t_L g5372 ( 
.A(n_5231),
.Y(n_5372)
);

OR2x6_ASAP7_75t_L g5373 ( 
.A(n_5237),
.B(n_302),
.Y(n_5373)
);

INVx1_ASAP7_75t_L g5374 ( 
.A(n_5187),
.Y(n_5374)
);

AO21x2_ASAP7_75t_L g5375 ( 
.A1(n_5262),
.A2(n_303),
.B(n_304),
.Y(n_5375)
);

HB1xp67_ASAP7_75t_L g5376 ( 
.A(n_5157),
.Y(n_5376)
);

INVx2_ASAP7_75t_L g5377 ( 
.A(n_5221),
.Y(n_5377)
);

INVx5_ASAP7_75t_L g5378 ( 
.A(n_5237),
.Y(n_5378)
);

NAND2xp5_ASAP7_75t_L g5379 ( 
.A(n_5264),
.B(n_305),
.Y(n_5379)
);

AO21x2_ASAP7_75t_L g5380 ( 
.A1(n_5241),
.A2(n_306),
.B(n_307),
.Y(n_5380)
);

AND2x2_ASAP7_75t_L g5381 ( 
.A(n_5254),
.B(n_308),
.Y(n_5381)
);

OR2x6_ASAP7_75t_L g5382 ( 
.A(n_5266),
.B(n_309),
.Y(n_5382)
);

INVx2_ASAP7_75t_SL g5383 ( 
.A(n_5155),
.Y(n_5383)
);

INVx1_ASAP7_75t_L g5384 ( 
.A(n_5188),
.Y(n_5384)
);

OR2x2_ASAP7_75t_L g5385 ( 
.A(n_5172),
.B(n_309),
.Y(n_5385)
);

AOI322xp5_ASAP7_75t_L g5386 ( 
.A1(n_5212),
.A2(n_311),
.A3(n_312),
.B1(n_313),
.B2(n_314),
.C1(n_315),
.C2(n_316),
.Y(n_5386)
);

INVx1_ASAP7_75t_L g5387 ( 
.A(n_5162),
.Y(n_5387)
);

AOI21xp5_ASAP7_75t_SL g5388 ( 
.A1(n_5266),
.A2(n_5200),
.B(n_5240),
.Y(n_5388)
);

INVxp67_ASAP7_75t_L g5389 ( 
.A(n_5217),
.Y(n_5389)
);

HB1xp67_ASAP7_75t_L g5390 ( 
.A(n_5234),
.Y(n_5390)
);

AOI22xp33_ASAP7_75t_L g5391 ( 
.A1(n_5203),
.A2(n_314),
.B1(n_311),
.B2(n_313),
.Y(n_5391)
);

INVx2_ASAP7_75t_L g5392 ( 
.A(n_5228),
.Y(n_5392)
);

OR2x6_ASAP7_75t_L g5393 ( 
.A(n_5245),
.B(n_316),
.Y(n_5393)
);

NOR2xp33_ASAP7_75t_L g5394 ( 
.A(n_5153),
.B(n_317),
.Y(n_5394)
);

INVx2_ASAP7_75t_L g5395 ( 
.A(n_5202),
.Y(n_5395)
);

INVx3_ASAP7_75t_L g5396 ( 
.A(n_5156),
.Y(n_5396)
);

OA21x2_ASAP7_75t_L g5397 ( 
.A1(n_5279),
.A2(n_5280),
.B(n_5225),
.Y(n_5397)
);

INVx1_ASAP7_75t_L g5398 ( 
.A(n_5239),
.Y(n_5398)
);

AO21x2_ASAP7_75t_L g5399 ( 
.A1(n_5287),
.A2(n_318),
.B(n_320),
.Y(n_5399)
);

INVx2_ASAP7_75t_SL g5400 ( 
.A(n_5245),
.Y(n_5400)
);

OAI21xp5_ASAP7_75t_L g5401 ( 
.A1(n_5227),
.A2(n_5247),
.B(n_5281),
.Y(n_5401)
);

INVx1_ASAP7_75t_L g5402 ( 
.A(n_5272),
.Y(n_5402)
);

AOI22xp33_ASAP7_75t_L g5403 ( 
.A1(n_5235),
.A2(n_324),
.B1(n_320),
.B2(n_323),
.Y(n_5403)
);

INVx1_ASAP7_75t_L g5404 ( 
.A(n_5214),
.Y(n_5404)
);

OR2x2_ASAP7_75t_L g5405 ( 
.A(n_5372),
.B(n_5206),
.Y(n_5405)
);

INVx1_ASAP7_75t_L g5406 ( 
.A(n_5350),
.Y(n_5406)
);

AOI22xp33_ASAP7_75t_L g5407 ( 
.A1(n_5323),
.A2(n_5251),
.B1(n_5249),
.B2(n_5284),
.Y(n_5407)
);

OR2x2_ASAP7_75t_L g5408 ( 
.A(n_5339),
.B(n_5191),
.Y(n_5408)
);

AOI22xp33_ASAP7_75t_L g5409 ( 
.A1(n_5323),
.A2(n_5401),
.B1(n_5339),
.B2(n_5316),
.Y(n_5409)
);

INVx2_ASAP7_75t_L g5410 ( 
.A(n_5349),
.Y(n_5410)
);

OR2x2_ASAP7_75t_L g5411 ( 
.A(n_5328),
.B(n_5283),
.Y(n_5411)
);

AOI22xp33_ASAP7_75t_L g5412 ( 
.A1(n_5401),
.A2(n_5243),
.B1(n_5275),
.B2(n_5246),
.Y(n_5412)
);

AND2x2_ASAP7_75t_L g5413 ( 
.A(n_5365),
.B(n_5255),
.Y(n_5413)
);

NAND2xp5_ASAP7_75t_L g5414 ( 
.A(n_5326),
.B(n_5275),
.Y(n_5414)
);

INVx1_ASAP7_75t_L g5415 ( 
.A(n_5359),
.Y(n_5415)
);

INVx1_ASAP7_75t_L g5416 ( 
.A(n_5376),
.Y(n_5416)
);

AND2x4_ASAP7_75t_L g5417 ( 
.A(n_5378),
.B(n_5179),
.Y(n_5417)
);

INVx1_ASAP7_75t_L g5418 ( 
.A(n_5376),
.Y(n_5418)
);

INVx2_ASAP7_75t_L g5419 ( 
.A(n_5349),
.Y(n_5419)
);

BUFx2_ASAP7_75t_L g5420 ( 
.A(n_5314),
.Y(n_5420)
);

INVxp67_ASAP7_75t_SL g5421 ( 
.A(n_5313),
.Y(n_5421)
);

INVx2_ASAP7_75t_SL g5422 ( 
.A(n_5383),
.Y(n_5422)
);

INVx2_ASAP7_75t_L g5423 ( 
.A(n_5330),
.Y(n_5423)
);

AND2x2_ASAP7_75t_L g5424 ( 
.A(n_5294),
.B(n_5183),
.Y(n_5424)
);

OR2x2_ASAP7_75t_L g5425 ( 
.A(n_5331),
.B(n_5234),
.Y(n_5425)
);

NOR2xp33_ASAP7_75t_L g5426 ( 
.A(n_5389),
.B(n_5194),
.Y(n_5426)
);

INVx2_ASAP7_75t_L g5427 ( 
.A(n_5330),
.Y(n_5427)
);

INVx2_ASAP7_75t_L g5428 ( 
.A(n_5369),
.Y(n_5428)
);

HB1xp67_ASAP7_75t_L g5429 ( 
.A(n_5390),
.Y(n_5429)
);

INVx2_ASAP7_75t_SL g5430 ( 
.A(n_5378),
.Y(n_5430)
);

CKINVDCx20_ASAP7_75t_R g5431 ( 
.A(n_5338),
.Y(n_5431)
);

INVx2_ASAP7_75t_L g5432 ( 
.A(n_5369),
.Y(n_5432)
);

INVx2_ASAP7_75t_L g5433 ( 
.A(n_5342),
.Y(n_5433)
);

AOI22xp33_ASAP7_75t_L g5434 ( 
.A1(n_5316),
.A2(n_5232),
.B1(n_5256),
.B2(n_5285),
.Y(n_5434)
);

INVx1_ASAP7_75t_L g5435 ( 
.A(n_5297),
.Y(n_5435)
);

INVx1_ASAP7_75t_L g5436 ( 
.A(n_5361),
.Y(n_5436)
);

INVx2_ASAP7_75t_SL g5437 ( 
.A(n_5378),
.Y(n_5437)
);

INVx2_ASAP7_75t_L g5438 ( 
.A(n_5342),
.Y(n_5438)
);

INVx1_ASAP7_75t_L g5439 ( 
.A(n_5364),
.Y(n_5439)
);

INVx1_ASAP7_75t_L g5440 ( 
.A(n_5305),
.Y(n_5440)
);

INVx1_ASAP7_75t_L g5441 ( 
.A(n_5307),
.Y(n_5441)
);

INVx2_ASAP7_75t_SL g5442 ( 
.A(n_5378),
.Y(n_5442)
);

AND2x4_ASAP7_75t_L g5443 ( 
.A(n_5355),
.B(n_5182),
.Y(n_5443)
);

NAND2xp5_ASAP7_75t_L g5444 ( 
.A(n_5326),
.B(n_5274),
.Y(n_5444)
);

AND2x2_ASAP7_75t_L g5445 ( 
.A(n_5366),
.B(n_5210),
.Y(n_5445)
);

BUFx2_ASAP7_75t_L g5446 ( 
.A(n_5329),
.Y(n_5446)
);

AND2x4_ASAP7_75t_L g5447 ( 
.A(n_5336),
.B(n_5173),
.Y(n_5447)
);

INVx1_ASAP7_75t_L g5448 ( 
.A(n_5318),
.Y(n_5448)
);

INVx1_ASAP7_75t_L g5449 ( 
.A(n_5324),
.Y(n_5449)
);

NAND4xp25_ASAP7_75t_L g5450 ( 
.A(n_5386),
.B(n_5271),
.C(n_5154),
.D(n_5252),
.Y(n_5450)
);

INVx1_ASAP7_75t_L g5451 ( 
.A(n_5332),
.Y(n_5451)
);

NOR2xp67_ASAP7_75t_L g5452 ( 
.A(n_5389),
.B(n_5230),
.Y(n_5452)
);

INVx1_ASAP7_75t_SL g5453 ( 
.A(n_5366),
.Y(n_5453)
);

OR2x2_ASAP7_75t_L g5454 ( 
.A(n_5302),
.B(n_5234),
.Y(n_5454)
);

AND2x2_ASAP7_75t_L g5455 ( 
.A(n_5344),
.B(n_5223),
.Y(n_5455)
);

INVx2_ASAP7_75t_L g5456 ( 
.A(n_5396),
.Y(n_5456)
);

INVx2_ASAP7_75t_L g5457 ( 
.A(n_5396),
.Y(n_5457)
);

NAND2xp5_ASAP7_75t_L g5458 ( 
.A(n_5370),
.B(n_5276),
.Y(n_5458)
);

AND2x2_ASAP7_75t_L g5459 ( 
.A(n_5353),
.B(n_5186),
.Y(n_5459)
);

BUFx2_ASAP7_75t_L g5460 ( 
.A(n_5329),
.Y(n_5460)
);

AOI22xp33_ASAP7_75t_L g5461 ( 
.A1(n_5399),
.A2(n_5169),
.B1(n_5222),
.B2(n_5159),
.Y(n_5461)
);

AND2x4_ASAP7_75t_L g5462 ( 
.A(n_5333),
.B(n_5161),
.Y(n_5462)
);

INVxp67_ASAP7_75t_SL g5463 ( 
.A(n_5390),
.Y(n_5463)
);

INVx1_ASAP7_75t_L g5464 ( 
.A(n_5340),
.Y(n_5464)
);

AND2x2_ASAP7_75t_L g5465 ( 
.A(n_5301),
.B(n_5207),
.Y(n_5465)
);

NAND2xp5_ASAP7_75t_L g5466 ( 
.A(n_5370),
.B(n_5259),
.Y(n_5466)
);

AND2x2_ASAP7_75t_L g5467 ( 
.A(n_5301),
.B(n_5263),
.Y(n_5467)
);

AND2x2_ASAP7_75t_L g5468 ( 
.A(n_5400),
.B(n_5160),
.Y(n_5468)
);

AND2x2_ASAP7_75t_L g5469 ( 
.A(n_5293),
.B(n_5149),
.Y(n_5469)
);

INVx1_ASAP7_75t_L g5470 ( 
.A(n_5347),
.Y(n_5470)
);

INVx2_ASAP7_75t_L g5471 ( 
.A(n_5299),
.Y(n_5471)
);

AND2x4_ASAP7_75t_L g5472 ( 
.A(n_5333),
.B(n_325),
.Y(n_5472)
);

NOR2xp33_ASAP7_75t_L g5473 ( 
.A(n_5337),
.B(n_327),
.Y(n_5473)
);

INVx2_ASAP7_75t_L g5474 ( 
.A(n_5319),
.Y(n_5474)
);

INVx2_ASAP7_75t_L g5475 ( 
.A(n_5322),
.Y(n_5475)
);

OAI22xp5_ASAP7_75t_L g5476 ( 
.A1(n_5296),
.A2(n_330),
.B1(n_328),
.B2(n_329),
.Y(n_5476)
);

INVx2_ASAP7_75t_L g5477 ( 
.A(n_5325),
.Y(n_5477)
);

OR2x2_ASAP7_75t_L g5478 ( 
.A(n_5295),
.B(n_331),
.Y(n_5478)
);

AOI22xp33_ASAP7_75t_L g5479 ( 
.A1(n_5399),
.A2(n_333),
.B1(n_331),
.B2(n_332),
.Y(n_5479)
);

HB1xp67_ASAP7_75t_L g5480 ( 
.A(n_5420),
.Y(n_5480)
);

OR2x2_ASAP7_75t_L g5481 ( 
.A(n_5453),
.B(n_5368),
.Y(n_5481)
);

HB1xp67_ASAP7_75t_L g5482 ( 
.A(n_5452),
.Y(n_5482)
);

OAI33xp33_ASAP7_75t_L g5483 ( 
.A1(n_5476),
.A2(n_5346),
.A3(n_5379),
.B1(n_5387),
.B2(n_5354),
.B3(n_5356),
.Y(n_5483)
);

AOI21xp5_ASAP7_75t_L g5484 ( 
.A1(n_5421),
.A2(n_5388),
.B(n_5368),
.Y(n_5484)
);

AND2x2_ASAP7_75t_L g5485 ( 
.A(n_5469),
.B(n_5337),
.Y(n_5485)
);

AOI31xp33_ASAP7_75t_L g5486 ( 
.A1(n_5409),
.A2(n_5346),
.A3(n_5391),
.B(n_5334),
.Y(n_5486)
);

AOI21xp33_ASAP7_75t_SL g5487 ( 
.A1(n_5409),
.A2(n_5334),
.B(n_5375),
.Y(n_5487)
);

OAI22xp33_ASAP7_75t_L g5488 ( 
.A1(n_5421),
.A2(n_5311),
.B1(n_5373),
.B2(n_5382),
.Y(n_5488)
);

OR2x2_ASAP7_75t_L g5489 ( 
.A(n_5478),
.B(n_5355),
.Y(n_5489)
);

INVx2_ASAP7_75t_L g5490 ( 
.A(n_5422),
.Y(n_5490)
);

AOI33xp33_ASAP7_75t_L g5491 ( 
.A1(n_5412),
.A2(n_5391),
.A3(n_5296),
.B1(n_5403),
.B2(n_5300),
.B3(n_5381),
.Y(n_5491)
);

BUFx3_ASAP7_75t_L g5492 ( 
.A(n_5431),
.Y(n_5492)
);

CKINVDCx20_ASAP7_75t_R g5493 ( 
.A(n_5431),
.Y(n_5493)
);

AOI22xp5_ASAP7_75t_L g5494 ( 
.A1(n_5426),
.A2(n_5358),
.B1(n_5311),
.B2(n_5373),
.Y(n_5494)
);

AND2x2_ASAP7_75t_L g5495 ( 
.A(n_5465),
.B(n_5373),
.Y(n_5495)
);

INVxp67_ASAP7_75t_SL g5496 ( 
.A(n_5426),
.Y(n_5496)
);

OAI221xp5_ASAP7_75t_L g5497 ( 
.A1(n_5461),
.A2(n_5412),
.B1(n_5407),
.B2(n_5434),
.C(n_5479),
.Y(n_5497)
);

AND2x2_ASAP7_75t_L g5498 ( 
.A(n_5467),
.B(n_5382),
.Y(n_5498)
);

OAI221xp5_ASAP7_75t_L g5499 ( 
.A1(n_5461),
.A2(n_5348),
.B1(n_5382),
.B2(n_5386),
.C(n_5371),
.Y(n_5499)
);

AND2x2_ASAP7_75t_L g5500 ( 
.A(n_5413),
.B(n_5327),
.Y(n_5500)
);

AOI221x1_ASAP7_75t_SL g5501 ( 
.A1(n_5450),
.A2(n_5308),
.B1(n_5379),
.B2(n_5394),
.C(n_5341),
.Y(n_5501)
);

INVx3_ASAP7_75t_L g5502 ( 
.A(n_5417),
.Y(n_5502)
);

INVx1_ASAP7_75t_L g5503 ( 
.A(n_5429),
.Y(n_5503)
);

INVx1_ASAP7_75t_L g5504 ( 
.A(n_5429),
.Y(n_5504)
);

AOI222xp33_ASAP7_75t_L g5505 ( 
.A1(n_5407),
.A2(n_5335),
.B1(n_5351),
.B2(n_5300),
.C1(n_5341),
.C2(n_5345),
.Y(n_5505)
);

AND2x2_ASAP7_75t_L g5506 ( 
.A(n_5445),
.B(n_5360),
.Y(n_5506)
);

INVx1_ASAP7_75t_L g5507 ( 
.A(n_5463),
.Y(n_5507)
);

OAI22xp5_ASAP7_75t_L g5508 ( 
.A1(n_5434),
.A2(n_5358),
.B1(n_5393),
.B2(n_5348),
.Y(n_5508)
);

INVx1_ASAP7_75t_L g5509 ( 
.A(n_5463),
.Y(n_5509)
);

INVx1_ASAP7_75t_L g5510 ( 
.A(n_5416),
.Y(n_5510)
);

AND2x2_ASAP7_75t_L g5511 ( 
.A(n_5424),
.B(n_5320),
.Y(n_5511)
);

OAI221xp5_ASAP7_75t_L g5512 ( 
.A1(n_5479),
.A2(n_5348),
.B1(n_5298),
.B2(n_5303),
.C(n_5393),
.Y(n_5512)
);

INVx1_ASAP7_75t_L g5513 ( 
.A(n_5418),
.Y(n_5513)
);

INVx1_ASAP7_75t_L g5514 ( 
.A(n_5406),
.Y(n_5514)
);

INVx1_ASAP7_75t_L g5515 ( 
.A(n_5415),
.Y(n_5515)
);

NAND2xp33_ASAP7_75t_SL g5516 ( 
.A(n_5414),
.B(n_5375),
.Y(n_5516)
);

INVx1_ASAP7_75t_L g5517 ( 
.A(n_5423),
.Y(n_5517)
);

BUFx2_ASAP7_75t_L g5518 ( 
.A(n_5446),
.Y(n_5518)
);

NOR4xp25_ASAP7_75t_L g5519 ( 
.A(n_5477),
.B(n_5315),
.C(n_5362),
.D(n_5385),
.Y(n_5519)
);

INVx1_ASAP7_75t_L g5520 ( 
.A(n_5423),
.Y(n_5520)
);

AOI21xp5_ASAP7_75t_L g5521 ( 
.A1(n_5444),
.A2(n_5317),
.B(n_5393),
.Y(n_5521)
);

INVx1_ASAP7_75t_L g5522 ( 
.A(n_5427),
.Y(n_5522)
);

AO21x2_ASAP7_75t_L g5523 ( 
.A1(n_5477),
.A2(n_5317),
.B(n_5380),
.Y(n_5523)
);

BUFx2_ASAP7_75t_SL g5524 ( 
.A(n_5430),
.Y(n_5524)
);

BUFx3_ASAP7_75t_L g5525 ( 
.A(n_5460),
.Y(n_5525)
);

OAI22xp5_ASAP7_75t_L g5526 ( 
.A1(n_5458),
.A2(n_5303),
.B1(n_5312),
.B2(n_5325),
.Y(n_5526)
);

NAND2xp5_ASAP7_75t_L g5527 ( 
.A(n_5501),
.B(n_5410),
.Y(n_5527)
);

INVx1_ASAP7_75t_L g5528 ( 
.A(n_5480),
.Y(n_5528)
);

NAND2xp5_ASAP7_75t_L g5529 ( 
.A(n_5501),
.B(n_5410),
.Y(n_5529)
);

AND2x2_ASAP7_75t_L g5530 ( 
.A(n_5524),
.B(n_5417),
.Y(n_5530)
);

INVx1_ASAP7_75t_L g5531 ( 
.A(n_5507),
.Y(n_5531)
);

INVx1_ASAP7_75t_L g5532 ( 
.A(n_5509),
.Y(n_5532)
);

INVxp67_ASAP7_75t_L g5533 ( 
.A(n_5482),
.Y(n_5533)
);

INVx2_ASAP7_75t_L g5534 ( 
.A(n_5492),
.Y(n_5534)
);

AND2x4_ASAP7_75t_L g5535 ( 
.A(n_5502),
.B(n_5419),
.Y(n_5535)
);

INVx2_ASAP7_75t_L g5536 ( 
.A(n_5502),
.Y(n_5536)
);

AND2x2_ASAP7_75t_L g5537 ( 
.A(n_5495),
.B(n_5417),
.Y(n_5537)
);

INVx2_ASAP7_75t_L g5538 ( 
.A(n_5493),
.Y(n_5538)
);

AND2x2_ASAP7_75t_L g5539 ( 
.A(n_5498),
.B(n_5518),
.Y(n_5539)
);

INVx1_ASAP7_75t_L g5540 ( 
.A(n_5503),
.Y(n_5540)
);

INVx1_ASAP7_75t_SL g5541 ( 
.A(n_5525),
.Y(n_5541)
);

NAND3xp33_ASAP7_75t_L g5542 ( 
.A(n_5487),
.B(n_5442),
.C(n_5437),
.Y(n_5542)
);

INVxp67_ASAP7_75t_SL g5543 ( 
.A(n_5484),
.Y(n_5543)
);

OR2x2_ASAP7_75t_L g5544 ( 
.A(n_5519),
.B(n_5427),
.Y(n_5544)
);

BUFx2_ASAP7_75t_L g5545 ( 
.A(n_5516),
.Y(n_5545)
);

AND2x2_ASAP7_75t_L g5546 ( 
.A(n_5485),
.B(n_5443),
.Y(n_5546)
);

INVx1_ASAP7_75t_L g5547 ( 
.A(n_5504),
.Y(n_5547)
);

NAND2xp5_ASAP7_75t_L g5548 ( 
.A(n_5505),
.B(n_5419),
.Y(n_5548)
);

NAND2xp5_ASAP7_75t_L g5549 ( 
.A(n_5505),
.B(n_5473),
.Y(n_5549)
);

INVx3_ASAP7_75t_L g5550 ( 
.A(n_5523),
.Y(n_5550)
);

HB1xp67_ASAP7_75t_L g5551 ( 
.A(n_5523),
.Y(n_5551)
);

INVx1_ASAP7_75t_L g5552 ( 
.A(n_5517),
.Y(n_5552)
);

AND2x2_ASAP7_75t_L g5553 ( 
.A(n_5500),
.B(n_5443),
.Y(n_5553)
);

HB1xp67_ASAP7_75t_L g5554 ( 
.A(n_5490),
.Y(n_5554)
);

CKINVDCx20_ASAP7_75t_R g5555 ( 
.A(n_5494),
.Y(n_5555)
);

AND2x4_ASAP7_75t_SL g5556 ( 
.A(n_5511),
.B(n_5468),
.Y(n_5556)
);

INVx1_ASAP7_75t_L g5557 ( 
.A(n_5520),
.Y(n_5557)
);

INVx1_ASAP7_75t_L g5558 ( 
.A(n_5522),
.Y(n_5558)
);

AND2x2_ASAP7_75t_L g5559 ( 
.A(n_5538),
.B(n_5506),
.Y(n_5559)
);

INVx1_ASAP7_75t_L g5560 ( 
.A(n_5550),
.Y(n_5560)
);

AOI22xp5_ASAP7_75t_L g5561 ( 
.A1(n_5555),
.A2(n_5488),
.B1(n_5508),
.B2(n_5497),
.Y(n_5561)
);

AND2x2_ASAP7_75t_L g5562 ( 
.A(n_5530),
.B(n_5496),
.Y(n_5562)
);

AND2x2_ASAP7_75t_L g5563 ( 
.A(n_5530),
.B(n_5443),
.Y(n_5563)
);

INVx1_ASAP7_75t_L g5564 ( 
.A(n_5550),
.Y(n_5564)
);

AND2x2_ASAP7_75t_L g5565 ( 
.A(n_5539),
.B(n_5471),
.Y(n_5565)
);

INVx2_ASAP7_75t_L g5566 ( 
.A(n_5550),
.Y(n_5566)
);

AND2x2_ASAP7_75t_L g5567 ( 
.A(n_5539),
.B(n_5471),
.Y(n_5567)
);

OR2x2_ASAP7_75t_L g5568 ( 
.A(n_5534),
.B(n_5489),
.Y(n_5568)
);

AND2x2_ASAP7_75t_L g5569 ( 
.A(n_5538),
.B(n_5455),
.Y(n_5569)
);

INVx1_ASAP7_75t_L g5570 ( 
.A(n_5551),
.Y(n_5570)
);

NAND2xp5_ASAP7_75t_L g5571 ( 
.A(n_5535),
.B(n_5486),
.Y(n_5571)
);

AND2x2_ASAP7_75t_L g5572 ( 
.A(n_5546),
.B(n_5474),
.Y(n_5572)
);

AND2x2_ASAP7_75t_L g5573 ( 
.A(n_5546),
.B(n_5474),
.Y(n_5573)
);

INVx1_ASAP7_75t_L g5574 ( 
.A(n_5528),
.Y(n_5574)
);

INVx2_ASAP7_75t_SL g5575 ( 
.A(n_5535),
.Y(n_5575)
);

NAND2xp5_ASAP7_75t_L g5576 ( 
.A(n_5535),
.B(n_5486),
.Y(n_5576)
);

NAND2xp5_ASAP7_75t_L g5577 ( 
.A(n_5534),
.B(n_5541),
.Y(n_5577)
);

INVx1_ASAP7_75t_L g5578 ( 
.A(n_5536),
.Y(n_5578)
);

INVx2_ASAP7_75t_L g5579 ( 
.A(n_5536),
.Y(n_5579)
);

AND2x4_ASAP7_75t_SL g5580 ( 
.A(n_5537),
.B(n_5472),
.Y(n_5580)
);

AND2x2_ASAP7_75t_L g5581 ( 
.A(n_5553),
.B(n_5447),
.Y(n_5581)
);

AND2x2_ASAP7_75t_L g5582 ( 
.A(n_5563),
.B(n_5553),
.Y(n_5582)
);

NAND2xp5_ASAP7_75t_L g5583 ( 
.A(n_5562),
.B(n_5533),
.Y(n_5583)
);

AND2x2_ASAP7_75t_L g5584 ( 
.A(n_5563),
.B(n_5562),
.Y(n_5584)
);

BUFx2_ASAP7_75t_L g5585 ( 
.A(n_5575),
.Y(n_5585)
);

NAND2xp5_ASAP7_75t_L g5586 ( 
.A(n_5565),
.B(n_5554),
.Y(n_5586)
);

OR2x2_ASAP7_75t_L g5587 ( 
.A(n_5571),
.B(n_5544),
.Y(n_5587)
);

NOR3x1_ASAP7_75t_L g5588 ( 
.A(n_5576),
.B(n_5497),
.C(n_5542),
.Y(n_5588)
);

NAND4xp25_ASAP7_75t_L g5589 ( 
.A(n_5561),
.B(n_5549),
.C(n_5548),
.D(n_5527),
.Y(n_5589)
);

INVx1_ASAP7_75t_L g5590 ( 
.A(n_5575),
.Y(n_5590)
);

INVx1_ASAP7_75t_L g5591 ( 
.A(n_5566),
.Y(n_5591)
);

OR2x2_ASAP7_75t_L g5592 ( 
.A(n_5568),
.B(n_5544),
.Y(n_5592)
);

NAND2xp5_ASAP7_75t_L g5593 ( 
.A(n_5579),
.B(n_5529),
.Y(n_5593)
);

NAND2xp5_ASAP7_75t_L g5594 ( 
.A(n_5579),
.B(n_5543),
.Y(n_5594)
);

INVx1_ASAP7_75t_L g5595 ( 
.A(n_5566),
.Y(n_5595)
);

INVx2_ASAP7_75t_L g5596 ( 
.A(n_5580),
.Y(n_5596)
);

AND2x2_ASAP7_75t_L g5597 ( 
.A(n_5580),
.B(n_5537),
.Y(n_5597)
);

AND2x4_ASAP7_75t_L g5598 ( 
.A(n_5565),
.B(n_5556),
.Y(n_5598)
);

INVx1_ASAP7_75t_L g5599 ( 
.A(n_5560),
.Y(n_5599)
);

AND2x2_ASAP7_75t_L g5600 ( 
.A(n_5581),
.B(n_5556),
.Y(n_5600)
);

INVx1_ASAP7_75t_L g5601 ( 
.A(n_5564),
.Y(n_5601)
);

INVx2_ASAP7_75t_L g5602 ( 
.A(n_5567),
.Y(n_5602)
);

INVx2_ASAP7_75t_L g5603 ( 
.A(n_5567),
.Y(n_5603)
);

AOI22xp5_ASAP7_75t_L g5604 ( 
.A1(n_5569),
.A2(n_5555),
.B1(n_5508),
.B2(n_5499),
.Y(n_5604)
);

INVx1_ASAP7_75t_L g5605 ( 
.A(n_5585),
.Y(n_5605)
);

AOI21xp5_ASAP7_75t_L g5606 ( 
.A1(n_5604),
.A2(n_5545),
.B(n_5521),
.Y(n_5606)
);

INVxp67_ASAP7_75t_L g5607 ( 
.A(n_5584),
.Y(n_5607)
);

NAND2xp5_ASAP7_75t_L g5608 ( 
.A(n_5582),
.B(n_5572),
.Y(n_5608)
);

AOI32xp33_ASAP7_75t_L g5609 ( 
.A1(n_5587),
.A2(n_5545),
.A3(n_5499),
.B1(n_5512),
.B2(n_5526),
.Y(n_5609)
);

INVx2_ASAP7_75t_SL g5610 ( 
.A(n_5598),
.Y(n_5610)
);

INVx3_ASAP7_75t_L g5611 ( 
.A(n_5598),
.Y(n_5611)
);

AND2x4_ASAP7_75t_L g5612 ( 
.A(n_5597),
.B(n_5559),
.Y(n_5612)
);

NOR2xp33_ASAP7_75t_L g5613 ( 
.A(n_5583),
.B(n_5577),
.Y(n_5613)
);

INVx1_ASAP7_75t_L g5614 ( 
.A(n_5590),
.Y(n_5614)
);

NOR2xp33_ASAP7_75t_SL g5615 ( 
.A(n_5600),
.B(n_5473),
.Y(n_5615)
);

OAI32xp33_ASAP7_75t_L g5616 ( 
.A1(n_5592),
.A2(n_5481),
.A3(n_5526),
.B1(n_5408),
.B2(n_5574),
.Y(n_5616)
);

NOR2xp33_ASAP7_75t_L g5617 ( 
.A(n_5589),
.B(n_5483),
.Y(n_5617)
);

NAND2xp5_ASAP7_75t_L g5618 ( 
.A(n_5596),
.B(n_5572),
.Y(n_5618)
);

INVxp67_ASAP7_75t_SL g5619 ( 
.A(n_5586),
.Y(n_5619)
);

HB1xp67_ASAP7_75t_L g5620 ( 
.A(n_5610),
.Y(n_5620)
);

NAND2xp5_ASAP7_75t_L g5621 ( 
.A(n_5612),
.B(n_5604),
.Y(n_5621)
);

INVx1_ASAP7_75t_SL g5622 ( 
.A(n_5612),
.Y(n_5622)
);

NOR2xp33_ASAP7_75t_L g5623 ( 
.A(n_5615),
.B(n_5589),
.Y(n_5623)
);

INVx1_ASAP7_75t_L g5624 ( 
.A(n_5618),
.Y(n_5624)
);

OR2x2_ASAP7_75t_L g5625 ( 
.A(n_5608),
.B(n_5602),
.Y(n_5625)
);

INVx2_ASAP7_75t_L g5626 ( 
.A(n_5611),
.Y(n_5626)
);

NAND2x1p5_ASAP7_75t_L g5627 ( 
.A(n_5605),
.B(n_5472),
.Y(n_5627)
);

AOI22xp33_ASAP7_75t_L g5628 ( 
.A1(n_5617),
.A2(n_5573),
.B1(n_5603),
.B2(n_5593),
.Y(n_5628)
);

AND2x2_ASAP7_75t_L g5629 ( 
.A(n_5607),
.B(n_5573),
.Y(n_5629)
);

NOR2xp33_ASAP7_75t_L g5630 ( 
.A(n_5613),
.B(n_5594),
.Y(n_5630)
);

INVx1_ASAP7_75t_L g5631 ( 
.A(n_5620),
.Y(n_5631)
);

AOI22xp5_ASAP7_75t_L g5632 ( 
.A1(n_5623),
.A2(n_5626),
.B1(n_5622),
.B2(n_5621),
.Y(n_5632)
);

OAI332xp33_ASAP7_75t_L g5633 ( 
.A1(n_5622),
.A2(n_5593),
.A3(n_5594),
.B1(n_5614),
.B2(n_5619),
.B3(n_5588),
.C1(n_5578),
.C2(n_5609),
.Y(n_5633)
);

INVx2_ASAP7_75t_SL g5634 ( 
.A(n_5627),
.Y(n_5634)
);

XOR2x2_ASAP7_75t_L g5635 ( 
.A(n_5630),
.B(n_5606),
.Y(n_5635)
);

INVxp67_ASAP7_75t_L g5636 ( 
.A(n_5629),
.Y(n_5636)
);

INVx1_ASAP7_75t_L g5637 ( 
.A(n_5625),
.Y(n_5637)
);

AOI21xp5_ASAP7_75t_L g5638 ( 
.A1(n_5624),
.A2(n_5616),
.B(n_5570),
.Y(n_5638)
);

NAND2xp33_ASAP7_75t_L g5639 ( 
.A(n_5628),
.B(n_5540),
.Y(n_5639)
);

INVx2_ASAP7_75t_SL g5640 ( 
.A(n_5627),
.Y(n_5640)
);

AOI22xp5_ASAP7_75t_L g5641 ( 
.A1(n_5623),
.A2(n_5462),
.B1(n_5547),
.B2(n_5513),
.Y(n_5641)
);

AOI221xp5_ASAP7_75t_L g5642 ( 
.A1(n_5623),
.A2(n_5532),
.B1(n_5531),
.B2(n_5557),
.C(n_5552),
.Y(n_5642)
);

AOI22xp5_ASAP7_75t_L g5643 ( 
.A1(n_5623),
.A2(n_5462),
.B1(n_5510),
.B2(n_5475),
.Y(n_5643)
);

INVx1_ASAP7_75t_L g5644 ( 
.A(n_5620),
.Y(n_5644)
);

INVx2_ASAP7_75t_L g5645 ( 
.A(n_5634),
.Y(n_5645)
);

AND2x4_ASAP7_75t_L g5646 ( 
.A(n_5640),
.B(n_5591),
.Y(n_5646)
);

NOR2xp33_ASAP7_75t_SL g5647 ( 
.A(n_5631),
.B(n_5595),
.Y(n_5647)
);

OAI22xp5_ASAP7_75t_L g5648 ( 
.A1(n_5632),
.A2(n_5466),
.B1(n_5475),
.B2(n_5428),
.Y(n_5648)
);

OAI221xp5_ASAP7_75t_L g5649 ( 
.A1(n_5641),
.A2(n_5558),
.B1(n_5601),
.B2(n_5599),
.C(n_5432),
.Y(n_5649)
);

OAI21xp33_ASAP7_75t_L g5650 ( 
.A1(n_5644),
.A2(n_5491),
.B(n_5432),
.Y(n_5650)
);

INVx1_ASAP7_75t_L g5651 ( 
.A(n_5637),
.Y(n_5651)
);

INVx2_ASAP7_75t_L g5652 ( 
.A(n_5636),
.Y(n_5652)
);

OAI32xp33_ASAP7_75t_L g5653 ( 
.A1(n_5633),
.A2(n_5428),
.A3(n_5515),
.B1(n_5514),
.B2(n_5438),
.Y(n_5653)
);

AOI21xp33_ASAP7_75t_SL g5654 ( 
.A1(n_5643),
.A2(n_5454),
.B(n_5312),
.Y(n_5654)
);

OAI32xp33_ASAP7_75t_L g5655 ( 
.A1(n_5635),
.A2(n_5456),
.A3(n_5457),
.B1(n_5438),
.B2(n_5433),
.Y(n_5655)
);

INVx1_ASAP7_75t_L g5656 ( 
.A(n_5646),
.Y(n_5656)
);

NAND3x1_ASAP7_75t_L g5657 ( 
.A(n_5651),
.B(n_5638),
.C(n_5642),
.Y(n_5657)
);

NAND2xp5_ASAP7_75t_L g5658 ( 
.A(n_5645),
.B(n_5639),
.Y(n_5658)
);

INVxp67_ASAP7_75t_SL g5659 ( 
.A(n_5647),
.Y(n_5659)
);

NOR2x1_ASAP7_75t_L g5660 ( 
.A(n_5652),
.B(n_5649),
.Y(n_5660)
);

OR2x2_ASAP7_75t_L g5661 ( 
.A(n_5648),
.B(n_5435),
.Y(n_5661)
);

AND2x2_ASAP7_75t_L g5662 ( 
.A(n_5650),
.B(n_5447),
.Y(n_5662)
);

NOR2xp33_ASAP7_75t_L g5663 ( 
.A(n_5653),
.B(n_5436),
.Y(n_5663)
);

HB1xp67_ASAP7_75t_L g5664 ( 
.A(n_5655),
.Y(n_5664)
);

INVx1_ASAP7_75t_L g5665 ( 
.A(n_5654),
.Y(n_5665)
);

AOI21xp5_ASAP7_75t_L g5666 ( 
.A1(n_5659),
.A2(n_5658),
.B(n_5665),
.Y(n_5666)
);

NAND2x1_ASAP7_75t_L g5667 ( 
.A(n_5656),
.B(n_5433),
.Y(n_5667)
);

OAI21xp5_ASAP7_75t_L g5668 ( 
.A1(n_5657),
.A2(n_5321),
.B(n_5343),
.Y(n_5668)
);

A2O1A1Ixp33_ASAP7_75t_L g5669 ( 
.A1(n_5663),
.A2(n_5457),
.B(n_5456),
.C(n_5440),
.Y(n_5669)
);

NAND4xp25_ASAP7_75t_L g5670 ( 
.A(n_5660),
.B(n_5367),
.C(n_5352),
.D(n_5439),
.Y(n_5670)
);

O2A1O1Ixp33_ASAP7_75t_L g5671 ( 
.A1(n_5664),
.A2(n_5441),
.B(n_5449),
.C(n_5448),
.Y(n_5671)
);

AOI21xp5_ASAP7_75t_L g5672 ( 
.A1(n_5661),
.A2(n_5464),
.B(n_5451),
.Y(n_5672)
);

NOR3xp33_ASAP7_75t_L g5673 ( 
.A(n_5662),
.B(n_5470),
.C(n_5405),
.Y(n_5673)
);

OAI211xp5_ASAP7_75t_L g5674 ( 
.A1(n_5659),
.A2(n_5425),
.B(n_5397),
.C(n_5304),
.Y(n_5674)
);

NAND4xp75_ASAP7_75t_L g5675 ( 
.A(n_5660),
.B(n_5397),
.C(n_5459),
.D(n_5306),
.Y(n_5675)
);

NAND2xp5_ASAP7_75t_L g5676 ( 
.A(n_5656),
.B(n_5380),
.Y(n_5676)
);

INVxp67_ASAP7_75t_L g5677 ( 
.A(n_5663),
.Y(n_5677)
);

NAND4xp75_ASAP7_75t_L g5678 ( 
.A(n_5660),
.B(n_5309),
.C(n_5398),
.D(n_5402),
.Y(n_5678)
);

NOR4xp25_ASAP7_75t_L g5679 ( 
.A(n_5657),
.B(n_5411),
.C(n_5310),
.D(n_5404),
.Y(n_5679)
);

NAND3xp33_ASAP7_75t_L g5680 ( 
.A(n_5665),
.B(n_5384),
.C(n_5374),
.Y(n_5680)
);

INVx1_ASAP7_75t_L g5681 ( 
.A(n_5662),
.Y(n_5681)
);

NOR3xp33_ASAP7_75t_L g5682 ( 
.A(n_5659),
.B(n_5363),
.C(n_5357),
.Y(n_5682)
);

NAND2xp5_ASAP7_75t_L g5683 ( 
.A(n_5656),
.B(n_5377),
.Y(n_5683)
);

AND2x2_ASAP7_75t_L g5684 ( 
.A(n_5668),
.B(n_5395),
.Y(n_5684)
);

NOR2xp33_ASAP7_75t_L g5685 ( 
.A(n_5670),
.B(n_5392),
.Y(n_5685)
);

NOR4xp25_ASAP7_75t_SL g5686 ( 
.A(n_5681),
.B(n_337),
.C(n_334),
.D(n_336),
.Y(n_5686)
);

NOR2xp33_ASAP7_75t_L g5687 ( 
.A(n_5677),
.B(n_336),
.Y(n_5687)
);

NAND4xp25_ASAP7_75t_L g5688 ( 
.A(n_5666),
.B(n_339),
.C(n_337),
.D(n_338),
.Y(n_5688)
);

NAND2xp5_ASAP7_75t_L g5689 ( 
.A(n_5679),
.B(n_339),
.Y(n_5689)
);

INVx1_ASAP7_75t_L g5690 ( 
.A(n_5667),
.Y(n_5690)
);

INVx1_ASAP7_75t_L g5691 ( 
.A(n_5676),
.Y(n_5691)
);

INVx1_ASAP7_75t_L g5692 ( 
.A(n_5678),
.Y(n_5692)
);

INVx1_ASAP7_75t_L g5693 ( 
.A(n_5683),
.Y(n_5693)
);

INVx1_ASAP7_75t_L g5694 ( 
.A(n_5671),
.Y(n_5694)
);

INVx1_ASAP7_75t_L g5695 ( 
.A(n_5673),
.Y(n_5695)
);

CKINVDCx16_ASAP7_75t_R g5696 ( 
.A(n_5682),
.Y(n_5696)
);

AOI21xp5_ASAP7_75t_L g5697 ( 
.A1(n_5672),
.A2(n_340),
.B(n_341),
.Y(n_5697)
);

AOI221xp5_ASAP7_75t_L g5698 ( 
.A1(n_5669),
.A2(n_340),
.B1(n_341),
.B2(n_342),
.C(n_343),
.Y(n_5698)
);

NOR3xp33_ASAP7_75t_SL g5699 ( 
.A(n_5680),
.B(n_5675),
.C(n_5674),
.Y(n_5699)
);

XNOR2xp5_ASAP7_75t_L g5700 ( 
.A(n_5681),
.B(n_343),
.Y(n_5700)
);

AOI21xp5_ASAP7_75t_L g5701 ( 
.A1(n_5666),
.A2(n_344),
.B(n_345),
.Y(n_5701)
);

NAND2xp5_ASAP7_75t_L g5702 ( 
.A(n_5668),
.B(n_345),
.Y(n_5702)
);

NAND2xp5_ASAP7_75t_L g5703 ( 
.A(n_5668),
.B(n_346),
.Y(n_5703)
);

AND2x2_ASAP7_75t_L g5704 ( 
.A(n_5668),
.B(n_347),
.Y(n_5704)
);

OAI21xp5_ASAP7_75t_SL g5705 ( 
.A1(n_5668),
.A2(n_347),
.B(n_348),
.Y(n_5705)
);

INVx1_ASAP7_75t_L g5706 ( 
.A(n_5667),
.Y(n_5706)
);

NOR3xp33_ASAP7_75t_L g5707 ( 
.A(n_5681),
.B(n_349),
.C(n_352),
.Y(n_5707)
);

OAI211xp5_ASAP7_75t_SL g5708 ( 
.A1(n_5677),
.A2(n_356),
.B(n_353),
.C(n_355),
.Y(n_5708)
);

NOR3xp33_ASAP7_75t_L g5709 ( 
.A(n_5696),
.B(n_353),
.C(n_358),
.Y(n_5709)
);

NAND4xp25_ASAP7_75t_SL g5710 ( 
.A(n_5692),
.B(n_5701),
.C(n_5703),
.D(n_5702),
.Y(n_5710)
);

NAND4xp75_ASAP7_75t_L g5711 ( 
.A(n_5704),
.B(n_362),
.C(n_359),
.D(n_361),
.Y(n_5711)
);

AOI221xp5_ASAP7_75t_SL g5712 ( 
.A1(n_5689),
.A2(n_359),
.B1(n_361),
.B2(n_362),
.C(n_363),
.Y(n_5712)
);

NAND2xp5_ASAP7_75t_L g5713 ( 
.A(n_5700),
.B(n_363),
.Y(n_5713)
);

AOI21xp5_ASAP7_75t_L g5714 ( 
.A1(n_5690),
.A2(n_364),
.B(n_365),
.Y(n_5714)
);

OAI21xp33_ASAP7_75t_SL g5715 ( 
.A1(n_5706),
.A2(n_364),
.B(n_365),
.Y(n_5715)
);

OA211x2_ASAP7_75t_L g5716 ( 
.A1(n_5698),
.A2(n_368),
.B(n_366),
.C(n_367),
.Y(n_5716)
);

INVx1_ASAP7_75t_SL g5717 ( 
.A(n_5684),
.Y(n_5717)
);

NOR3x1_ASAP7_75t_SL g5718 ( 
.A(n_5688),
.B(n_366),
.C(n_367),
.Y(n_5718)
);

AND2x2_ASAP7_75t_L g5719 ( 
.A(n_5686),
.B(n_370),
.Y(n_5719)
);

NOR2xp33_ASAP7_75t_L g5720 ( 
.A(n_5708),
.B(n_370),
.Y(n_5720)
);

NOR2xp33_ASAP7_75t_SL g5721 ( 
.A(n_5705),
.B(n_371),
.Y(n_5721)
);

NOR4xp25_ASAP7_75t_L g5722 ( 
.A(n_5694),
.B(n_374),
.C(n_371),
.D(n_372),
.Y(n_5722)
);

OAI211xp5_ASAP7_75t_SL g5723 ( 
.A1(n_5699),
.A2(n_376),
.B(n_374),
.C(n_375),
.Y(n_5723)
);

NAND4xp25_ASAP7_75t_L g5724 ( 
.A(n_5687),
.B(n_378),
.C(n_375),
.D(n_376),
.Y(n_5724)
);

INVxp67_ASAP7_75t_SL g5725 ( 
.A(n_5707),
.Y(n_5725)
);

NAND3xp33_ASAP7_75t_L g5726 ( 
.A(n_5697),
.B(n_379),
.C(n_380),
.Y(n_5726)
);

AND4x1_ASAP7_75t_L g5727 ( 
.A(n_5695),
.B(n_384),
.C(n_381),
.D(n_383),
.Y(n_5727)
);

NOR3xp33_ASAP7_75t_L g5728 ( 
.A(n_5693),
.B(n_381),
.C(n_383),
.Y(n_5728)
);

OAI211xp5_ASAP7_75t_L g5729 ( 
.A1(n_5691),
.A2(n_388),
.B(n_385),
.C(n_386),
.Y(n_5729)
);

INVx1_ASAP7_75t_L g5730 ( 
.A(n_5685),
.Y(n_5730)
);

NOR4xp25_ASAP7_75t_SL g5731 ( 
.A(n_5705),
.B(n_390),
.C(n_386),
.D(n_388),
.Y(n_5731)
);

NAND2xp5_ASAP7_75t_L g5732 ( 
.A(n_5700),
.B(n_390),
.Y(n_5732)
);

NOR3x1_ASAP7_75t_L g5733 ( 
.A(n_5705),
.B(n_391),
.C(n_392),
.Y(n_5733)
);

INVx1_ASAP7_75t_L g5734 ( 
.A(n_5700),
.Y(n_5734)
);

NOR2x1_ASAP7_75t_L g5735 ( 
.A(n_5688),
.B(n_391),
.Y(n_5735)
);

NAND3xp33_ASAP7_75t_L g5736 ( 
.A(n_5699),
.B(n_392),
.C(n_393),
.Y(n_5736)
);

OAI21xp5_ASAP7_75t_L g5737 ( 
.A1(n_5736),
.A2(n_394),
.B(n_395),
.Y(n_5737)
);

NAND4xp25_ASAP7_75t_SL g5738 ( 
.A(n_5712),
.B(n_396),
.C(n_397),
.D(n_398),
.Y(n_5738)
);

NAND4xp25_ASAP7_75t_SL g5739 ( 
.A(n_5715),
.B(n_398),
.C(n_400),
.D(n_401),
.Y(n_5739)
);

INVx2_ASAP7_75t_SL g5740 ( 
.A(n_5719),
.Y(n_5740)
);

NAND4xp25_ASAP7_75t_L g5741 ( 
.A(n_5733),
.B(n_400),
.C(n_401),
.D(n_402),
.Y(n_5741)
);

OAI321xp33_ASAP7_75t_L g5742 ( 
.A1(n_5723),
.A2(n_5730),
.A3(n_5734),
.B1(n_5725),
.B2(n_5726),
.C(n_5720),
.Y(n_5742)
);

NAND2xp5_ASAP7_75t_SL g5743 ( 
.A(n_5722),
.B(n_403),
.Y(n_5743)
);

NAND2xp5_ASAP7_75t_L g5744 ( 
.A(n_5727),
.B(n_403),
.Y(n_5744)
);

NOR3xp33_ASAP7_75t_L g5745 ( 
.A(n_5710),
.B(n_404),
.C(n_405),
.Y(n_5745)
);

AND2x2_ASAP7_75t_L g5746 ( 
.A(n_5731),
.B(n_404),
.Y(n_5746)
);

NOR3x1_ASAP7_75t_L g5747 ( 
.A(n_5711),
.B(n_405),
.C(n_406),
.Y(n_5747)
);

NOR2xp33_ASAP7_75t_L g5748 ( 
.A(n_5724),
.B(n_5721),
.Y(n_5748)
);

NOR3xp33_ASAP7_75t_L g5749 ( 
.A(n_5713),
.B(n_407),
.C(n_409),
.Y(n_5749)
);

NAND4xp25_ASAP7_75t_L g5750 ( 
.A(n_5716),
.B(n_407),
.C(n_409),
.D(n_410),
.Y(n_5750)
);

OAI221xp5_ASAP7_75t_L g5751 ( 
.A1(n_5717),
.A2(n_411),
.B1(n_412),
.B2(n_413),
.C(n_414),
.Y(n_5751)
);

INVx1_ASAP7_75t_L g5752 ( 
.A(n_5718),
.Y(n_5752)
);

AOI211xp5_ASAP7_75t_L g5753 ( 
.A1(n_5729),
.A2(n_411),
.B(n_414),
.C(n_415),
.Y(n_5753)
);

AOI221x1_ASAP7_75t_L g5754 ( 
.A1(n_5709),
.A2(n_416),
.B1(n_417),
.B2(n_418),
.C(n_419),
.Y(n_5754)
);

AOI211xp5_ASAP7_75t_L g5755 ( 
.A1(n_5732),
.A2(n_417),
.B(n_418),
.C(n_420),
.Y(n_5755)
);

AND3x2_ASAP7_75t_L g5756 ( 
.A(n_5728),
.B(n_422),
.C(n_423),
.Y(n_5756)
);

OAI211xp5_ASAP7_75t_SL g5757 ( 
.A1(n_5735),
.A2(n_424),
.B(n_425),
.C(n_426),
.Y(n_5757)
);

AOI221xp5_ASAP7_75t_L g5758 ( 
.A1(n_5714),
.A2(n_424),
.B1(n_426),
.B2(n_427),
.C(n_428),
.Y(n_5758)
);

NOR2x1_ASAP7_75t_L g5759 ( 
.A(n_5711),
.B(n_427),
.Y(n_5759)
);

OAI211xp5_ASAP7_75t_SL g5760 ( 
.A1(n_5717),
.A2(n_429),
.B(n_430),
.C(n_432),
.Y(n_5760)
);

AOI321xp33_ASAP7_75t_L g5761 ( 
.A1(n_5725),
.A2(n_430),
.A3(n_433),
.B1(n_434),
.B2(n_435),
.C(n_436),
.Y(n_5761)
);

NAND4xp75_ASAP7_75t_L g5762 ( 
.A(n_5747),
.B(n_434),
.C(n_436),
.D(n_438),
.Y(n_5762)
);

HB1xp67_ASAP7_75t_L g5763 ( 
.A(n_5746),
.Y(n_5763)
);

INVx1_ASAP7_75t_L g5764 ( 
.A(n_5744),
.Y(n_5764)
);

INVx1_ASAP7_75t_L g5765 ( 
.A(n_5740),
.Y(n_5765)
);

INVx1_ASAP7_75t_L g5766 ( 
.A(n_5752),
.Y(n_5766)
);

AND2x2_ASAP7_75t_SL g5767 ( 
.A(n_5745),
.B(n_439),
.Y(n_5767)
);

OAI221xp5_ASAP7_75t_L g5768 ( 
.A1(n_5737),
.A2(n_439),
.B1(n_442),
.B2(n_443),
.C(n_444),
.Y(n_5768)
);

NAND3xp33_ASAP7_75t_L g5769 ( 
.A(n_5753),
.B(n_442),
.C(n_446),
.Y(n_5769)
);

AOI221xp5_ASAP7_75t_L g5770 ( 
.A1(n_5739),
.A2(n_447),
.B1(n_450),
.B2(n_451),
.C(n_452),
.Y(n_5770)
);

NAND2xp33_ASAP7_75t_R g5771 ( 
.A(n_5756),
.B(n_447),
.Y(n_5771)
);

OAI22xp5_ASAP7_75t_L g5772 ( 
.A1(n_5751),
.A2(n_5755),
.B1(n_5759),
.B2(n_5748),
.Y(n_5772)
);

NAND2xp5_ASAP7_75t_L g5773 ( 
.A(n_5754),
.B(n_5749),
.Y(n_5773)
);

NAND2xp5_ASAP7_75t_SL g5774 ( 
.A(n_5761),
.B(n_450),
.Y(n_5774)
);

AOI21xp33_ASAP7_75t_L g5775 ( 
.A1(n_5757),
.A2(n_451),
.B(n_452),
.Y(n_5775)
);

AO22x2_ASAP7_75t_L g5776 ( 
.A1(n_5743),
.A2(n_454),
.B1(n_455),
.B2(n_456),
.Y(n_5776)
);

INVx1_ASAP7_75t_L g5777 ( 
.A(n_5750),
.Y(n_5777)
);

HB1xp67_ASAP7_75t_L g5778 ( 
.A(n_5738),
.Y(n_5778)
);

AOI22xp5_ASAP7_75t_L g5779 ( 
.A1(n_5741),
.A2(n_455),
.B1(n_457),
.B2(n_458),
.Y(n_5779)
);

OAI221xp5_ASAP7_75t_SL g5780 ( 
.A1(n_5758),
.A2(n_457),
.B1(n_462),
.B2(n_464),
.C(n_465),
.Y(n_5780)
);

XNOR2xp5_ASAP7_75t_L g5781 ( 
.A(n_5762),
.B(n_5742),
.Y(n_5781)
);

INVx1_ASAP7_75t_L g5782 ( 
.A(n_5776),
.Y(n_5782)
);

NAND4xp75_ASAP7_75t_L g5783 ( 
.A(n_5766),
.B(n_5760),
.C(n_464),
.D(n_466),
.Y(n_5783)
);

INVx1_ASAP7_75t_L g5784 ( 
.A(n_5776),
.Y(n_5784)
);

INVx1_ASAP7_75t_L g5785 ( 
.A(n_5763),
.Y(n_5785)
);

NOR2x1_ASAP7_75t_L g5786 ( 
.A(n_5777),
.B(n_462),
.Y(n_5786)
);

AND2x4_ASAP7_75t_L g5787 ( 
.A(n_5765),
.B(n_466),
.Y(n_5787)
);

NOR2x1_ASAP7_75t_L g5788 ( 
.A(n_5769),
.B(n_467),
.Y(n_5788)
);

INVx1_ASAP7_75t_L g5789 ( 
.A(n_5767),
.Y(n_5789)
);

OR2x2_ASAP7_75t_L g5790 ( 
.A(n_5774),
.B(n_467),
.Y(n_5790)
);

INVx1_ASAP7_75t_L g5791 ( 
.A(n_5779),
.Y(n_5791)
);

INVx1_ASAP7_75t_L g5792 ( 
.A(n_5778),
.Y(n_5792)
);

NOR3xp33_ASAP7_75t_L g5793 ( 
.A(n_5772),
.B(n_468),
.C(n_469),
.Y(n_5793)
);

XNOR2xp5_ASAP7_75t_L g5794 ( 
.A(n_5770),
.B(n_5768),
.Y(n_5794)
);

AOI22xp5_ASAP7_75t_L g5795 ( 
.A1(n_5771),
.A2(n_468),
.B1(n_470),
.B2(n_471),
.Y(n_5795)
);

AND2x4_ASAP7_75t_L g5796 ( 
.A(n_5764),
.B(n_472),
.Y(n_5796)
);

NOR3xp33_ASAP7_75t_L g5797 ( 
.A(n_5792),
.B(n_5773),
.C(n_5780),
.Y(n_5797)
);

AND2x4_ASAP7_75t_L g5798 ( 
.A(n_5785),
.B(n_5775),
.Y(n_5798)
);

NOR4xp25_ASAP7_75t_L g5799 ( 
.A(n_5782),
.B(n_472),
.C(n_474),
.D(n_475),
.Y(n_5799)
);

INVx2_ASAP7_75t_L g5800 ( 
.A(n_5787),
.Y(n_5800)
);

NAND2xp5_ASAP7_75t_SL g5801 ( 
.A(n_5795),
.B(n_476),
.Y(n_5801)
);

NAND3xp33_ASAP7_75t_SL g5802 ( 
.A(n_5793),
.B(n_476),
.C(n_477),
.Y(n_5802)
);

OR2x2_ASAP7_75t_L g5803 ( 
.A(n_5790),
.B(n_477),
.Y(n_5803)
);

NAND2xp5_ASAP7_75t_L g5804 ( 
.A(n_5786),
.B(n_5784),
.Y(n_5804)
);

NAND4xp25_ASAP7_75t_SL g5805 ( 
.A(n_5788),
.B(n_478),
.C(n_479),
.D(n_480),
.Y(n_5805)
);

NOR2xp33_ASAP7_75t_L g5806 ( 
.A(n_5783),
.B(n_478),
.Y(n_5806)
);

NAND2xp5_ASAP7_75t_L g5807 ( 
.A(n_5796),
.B(n_480),
.Y(n_5807)
);

OAI21xp33_ASAP7_75t_L g5808 ( 
.A1(n_5781),
.A2(n_5791),
.B(n_5794),
.Y(n_5808)
);

NOR3xp33_ASAP7_75t_L g5809 ( 
.A(n_5789),
.B(n_481),
.C(n_482),
.Y(n_5809)
);

OR2x6_ASAP7_75t_L g5810 ( 
.A(n_5789),
.B(n_481),
.Y(n_5810)
);

INVx1_ASAP7_75t_L g5811 ( 
.A(n_5786),
.Y(n_5811)
);

OR5x1_ASAP7_75t_L g5812 ( 
.A(n_5781),
.B(n_483),
.C(n_484),
.D(n_487),
.E(n_489),
.Y(n_5812)
);

XNOR2xp5_ASAP7_75t_L g5813 ( 
.A(n_5781),
.B(n_483),
.Y(n_5813)
);

NOR3xp33_ASAP7_75t_L g5814 ( 
.A(n_5792),
.B(n_487),
.C(n_489),
.Y(n_5814)
);

HB1xp67_ASAP7_75t_L g5815 ( 
.A(n_5812),
.Y(n_5815)
);

HB1xp67_ASAP7_75t_L g5816 ( 
.A(n_5813),
.Y(n_5816)
);

OR2x2_ASAP7_75t_L g5817 ( 
.A(n_5799),
.B(n_490),
.Y(n_5817)
);

CKINVDCx5p33_ASAP7_75t_R g5818 ( 
.A(n_5800),
.Y(n_5818)
);

CKINVDCx5p33_ASAP7_75t_R g5819 ( 
.A(n_5798),
.Y(n_5819)
);

INVxp33_ASAP7_75t_L g5820 ( 
.A(n_5806),
.Y(n_5820)
);

INVx1_ASAP7_75t_L g5821 ( 
.A(n_5807),
.Y(n_5821)
);

NOR2xp33_ASAP7_75t_R g5822 ( 
.A(n_5805),
.B(n_491),
.Y(n_5822)
);

CKINVDCx5p33_ASAP7_75t_R g5823 ( 
.A(n_5808),
.Y(n_5823)
);

BUFx2_ASAP7_75t_L g5824 ( 
.A(n_5811),
.Y(n_5824)
);

INVxp67_ASAP7_75t_SL g5825 ( 
.A(n_5814),
.Y(n_5825)
);

INVx1_ASAP7_75t_SL g5826 ( 
.A(n_5803),
.Y(n_5826)
);

INVx1_ASAP7_75t_SL g5827 ( 
.A(n_5810),
.Y(n_5827)
);

AOI21xp5_ASAP7_75t_L g5828 ( 
.A1(n_5804),
.A2(n_491),
.B(n_492),
.Y(n_5828)
);

NAND2xp5_ASAP7_75t_L g5829 ( 
.A(n_5828),
.B(n_5809),
.Y(n_5829)
);

OAI31xp33_ASAP7_75t_L g5830 ( 
.A1(n_5817),
.A2(n_5801),
.A3(n_5797),
.B(n_5802),
.Y(n_5830)
);

NOR3xp33_ASAP7_75t_L g5831 ( 
.A(n_5824),
.B(n_5810),
.C(n_493),
.Y(n_5831)
);

OAI32xp33_ASAP7_75t_L g5832 ( 
.A1(n_5820),
.A2(n_492),
.A3(n_493),
.B1(n_494),
.B2(n_495),
.Y(n_5832)
);

AOI221xp5_ASAP7_75t_L g5833 ( 
.A1(n_5823),
.A2(n_494),
.B1(n_496),
.B2(n_497),
.C(n_498),
.Y(n_5833)
);

AOI322xp5_ASAP7_75t_L g5834 ( 
.A1(n_5827),
.A2(n_5815),
.A3(n_5825),
.B1(n_5826),
.B2(n_5816),
.C1(n_5818),
.C2(n_5821),
.Y(n_5834)
);

AOI322xp5_ASAP7_75t_L g5835 ( 
.A1(n_5819),
.A2(n_496),
.A3(n_498),
.B1(n_499),
.B2(n_500),
.C1(n_501),
.C2(n_502),
.Y(n_5835)
);

AO22x2_ASAP7_75t_L g5836 ( 
.A1(n_5831),
.A2(n_5822),
.B1(n_500),
.B2(n_503),
.Y(n_5836)
);

INVx1_ASAP7_75t_L g5837 ( 
.A(n_5829),
.Y(n_5837)
);

OAI22xp5_ASAP7_75t_L g5838 ( 
.A1(n_5833),
.A2(n_499),
.B1(n_503),
.B2(n_505),
.Y(n_5838)
);

HB1xp67_ASAP7_75t_L g5839 ( 
.A(n_5832),
.Y(n_5839)
);

AOI22xp5_ASAP7_75t_L g5840 ( 
.A1(n_5834),
.A2(n_505),
.B1(n_506),
.B2(n_507),
.Y(n_5840)
);

INVx1_ASAP7_75t_L g5841 ( 
.A(n_5830),
.Y(n_5841)
);

AO22x2_ASAP7_75t_L g5842 ( 
.A1(n_5835),
.A2(n_507),
.B1(n_508),
.B2(n_509),
.Y(n_5842)
);

INVx3_ASAP7_75t_L g5843 ( 
.A(n_5836),
.Y(n_5843)
);

OAI222xp33_ASAP7_75t_L g5844 ( 
.A1(n_5841),
.A2(n_508),
.B1(n_510),
.B2(n_511),
.C1(n_512),
.C2(n_513),
.Y(n_5844)
);

NAND4xp25_ASAP7_75t_SL g5845 ( 
.A(n_5840),
.B(n_511),
.C(n_513),
.D(n_515),
.Y(n_5845)
);

AND2x2_ASAP7_75t_L g5846 ( 
.A(n_5842),
.B(n_515),
.Y(n_5846)
);

O2A1O1Ixp33_ASAP7_75t_L g5847 ( 
.A1(n_5839),
.A2(n_516),
.B(n_517),
.C(n_519),
.Y(n_5847)
);

NOR2xp67_ASAP7_75t_L g5848 ( 
.A(n_5838),
.B(n_516),
.Y(n_5848)
);

OAI22xp33_ASAP7_75t_L g5849 ( 
.A1(n_5848),
.A2(n_5837),
.B1(n_520),
.B2(n_521),
.Y(n_5849)
);

AOI22xp5_ASAP7_75t_L g5850 ( 
.A1(n_5845),
.A2(n_519),
.B1(n_520),
.B2(n_524),
.Y(n_5850)
);

OAI21xp5_ASAP7_75t_L g5851 ( 
.A1(n_5846),
.A2(n_525),
.B(n_527),
.Y(n_5851)
);

NAND2xp5_ASAP7_75t_L g5852 ( 
.A(n_5847),
.B(n_5843),
.Y(n_5852)
);

OAI22xp5_ASAP7_75t_L g5853 ( 
.A1(n_5844),
.A2(n_525),
.B1(n_527),
.B2(n_528),
.Y(n_5853)
);

INVx2_ASAP7_75t_L g5854 ( 
.A(n_5850),
.Y(n_5854)
);

AO21x2_ASAP7_75t_L g5855 ( 
.A1(n_5852),
.A2(n_528),
.B(n_529),
.Y(n_5855)
);

AOI21xp5_ASAP7_75t_L g5856 ( 
.A1(n_5849),
.A2(n_530),
.B(n_532),
.Y(n_5856)
);

NAND2xp5_ASAP7_75t_L g5857 ( 
.A(n_5851),
.B(n_5853),
.Y(n_5857)
);

AOI21xp5_ASAP7_75t_L g5858 ( 
.A1(n_5857),
.A2(n_533),
.B(n_535),
.Y(n_5858)
);

INVx2_ASAP7_75t_L g5859 ( 
.A(n_5855),
.Y(n_5859)
);

INVx1_ASAP7_75t_L g5860 ( 
.A(n_5856),
.Y(n_5860)
);

OAI21xp5_ASAP7_75t_L g5861 ( 
.A1(n_5854),
.A2(n_536),
.B(n_538),
.Y(n_5861)
);

OAI22xp5_ASAP7_75t_L g5862 ( 
.A1(n_5854),
.A2(n_540),
.B1(n_541),
.B2(n_543),
.Y(n_5862)
);

AOI21xp5_ASAP7_75t_L g5863 ( 
.A1(n_5859),
.A2(n_540),
.B(n_541),
.Y(n_5863)
);

NAND2xp5_ASAP7_75t_L g5864 ( 
.A(n_5858),
.B(n_544),
.Y(n_5864)
);

AOI22xp33_ASAP7_75t_L g5865 ( 
.A1(n_5860),
.A2(n_545),
.B1(n_546),
.B2(n_547),
.Y(n_5865)
);

OR2x2_ASAP7_75t_L g5866 ( 
.A(n_5861),
.B(n_546),
.Y(n_5866)
);

AOI21xp5_ASAP7_75t_L g5867 ( 
.A1(n_5862),
.A2(n_547),
.B(n_549),
.Y(n_5867)
);

AOI22xp33_ASAP7_75t_L g5868 ( 
.A1(n_5860),
.A2(n_549),
.B1(n_552),
.B2(n_553),
.Y(n_5868)
);

NAND2xp5_ASAP7_75t_L g5869 ( 
.A(n_5859),
.B(n_552),
.Y(n_5869)
);

INVx1_ASAP7_75t_L g5870 ( 
.A(n_5859),
.Y(n_5870)
);

OAI221xp5_ASAP7_75t_L g5871 ( 
.A1(n_5859),
.A2(n_553),
.B1(n_554),
.B2(n_555),
.C(n_556),
.Y(n_5871)
);

INVxp67_ASAP7_75t_SL g5872 ( 
.A(n_5859),
.Y(n_5872)
);

OAI22xp33_ASAP7_75t_L g5873 ( 
.A1(n_5866),
.A2(n_554),
.B1(n_555),
.B2(n_556),
.Y(n_5873)
);

OAI22xp33_ASAP7_75t_L g5874 ( 
.A1(n_5864),
.A2(n_557),
.B1(n_559),
.B2(n_560),
.Y(n_5874)
);

OA22x2_ASAP7_75t_L g5875 ( 
.A1(n_5870),
.A2(n_557),
.B1(n_559),
.B2(n_561),
.Y(n_5875)
);

OAI22xp5_ASAP7_75t_L g5876 ( 
.A1(n_5872),
.A2(n_561),
.B1(n_562),
.B2(n_564),
.Y(n_5876)
);

OAI22xp5_ASAP7_75t_L g5877 ( 
.A1(n_5867),
.A2(n_565),
.B1(n_567),
.B2(n_568),
.Y(n_5877)
);

AO22x2_ASAP7_75t_L g5878 ( 
.A1(n_5863),
.A2(n_565),
.B1(n_567),
.B2(n_569),
.Y(n_5878)
);

AOI22xp33_ASAP7_75t_L g5879 ( 
.A1(n_5871),
.A2(n_569),
.B1(n_570),
.B2(n_571),
.Y(n_5879)
);

AOI22xp5_ASAP7_75t_L g5880 ( 
.A1(n_5865),
.A2(n_571),
.B1(n_572),
.B2(n_573),
.Y(n_5880)
);

AOI22xp33_ASAP7_75t_L g5881 ( 
.A1(n_5868),
.A2(n_573),
.B1(n_574),
.B2(n_576),
.Y(n_5881)
);

OA22x2_ASAP7_75t_L g5882 ( 
.A1(n_5869),
.A2(n_574),
.B1(n_578),
.B2(n_580),
.Y(n_5882)
);

AND2x2_ASAP7_75t_L g5883 ( 
.A(n_5879),
.B(n_578),
.Y(n_5883)
);

OAI21xp5_ASAP7_75t_L g5884 ( 
.A1(n_5877),
.A2(n_581),
.B(n_582),
.Y(n_5884)
);

OAI221xp5_ASAP7_75t_L g5885 ( 
.A1(n_5881),
.A2(n_582),
.B1(n_583),
.B2(n_584),
.C(n_586),
.Y(n_5885)
);

NAND2xp5_ASAP7_75t_L g5886 ( 
.A(n_5878),
.B(n_584),
.Y(n_5886)
);

OR2x6_ASAP7_75t_L g5887 ( 
.A(n_5882),
.B(n_586),
.Y(n_5887)
);

AND2x2_ASAP7_75t_L g5888 ( 
.A(n_5880),
.B(n_587),
.Y(n_5888)
);

XNOR2xp5_ASAP7_75t_L g5889 ( 
.A(n_5886),
.B(n_5873),
.Y(n_5889)
);

XNOR2xp5_ASAP7_75t_L g5890 ( 
.A(n_5883),
.B(n_5874),
.Y(n_5890)
);

AOI22xp5_ASAP7_75t_L g5891 ( 
.A1(n_5887),
.A2(n_5876),
.B1(n_5875),
.B2(n_589),
.Y(n_5891)
);

AOI21xp33_ASAP7_75t_L g5892 ( 
.A1(n_5888),
.A2(n_587),
.B(n_588),
.Y(n_5892)
);

AOI221xp5_ASAP7_75t_L g5893 ( 
.A1(n_5891),
.A2(n_5884),
.B1(n_5885),
.B2(n_593),
.C(n_594),
.Y(n_5893)
);

AOI221xp5_ASAP7_75t_L g5894 ( 
.A1(n_5893),
.A2(n_5889),
.B1(n_5890),
.B2(n_5892),
.C(n_595),
.Y(n_5894)
);

AOI211xp5_ASAP7_75t_L g5895 ( 
.A1(n_5894),
.A2(n_588),
.B(n_592),
.C(n_593),
.Y(n_5895)
);


endmodule