module fake_jpeg_3166_n_142 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_142);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_142;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx10_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx2_ASAP7_75t_SL g42 ( 
.A(n_30),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_6),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_31),
.B(n_32),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_16),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_15),
.B(n_6),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_37),
.B(n_39),
.Y(n_40)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_19),
.B(n_4),
.Y(n_39)
);

OAI22xp33_ASAP7_75t_L g43 ( 
.A1(n_33),
.A2(n_35),
.B1(n_38),
.B2(n_32),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_43),
.A2(n_35),
.B1(n_34),
.B2(n_30),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_29),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_49),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_29),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_31),
.B(n_26),
.Y(n_50)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_18),
.Y(n_59)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

BUFx2_ASAP7_75t_SL g56 ( 
.A(n_51),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

OA22x2_ASAP7_75t_L g57 ( 
.A1(n_48),
.A2(n_33),
.B1(n_38),
.B2(n_30),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_58),
.A2(n_34),
.B1(n_36),
.B2(n_25),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_60),
.Y(n_73)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_62),
.Y(n_76)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_63),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_18),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_64),
.B(n_67),
.Y(n_75)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_65),
.B(n_66),
.Y(n_71)
);

CKINVDCx14_ASAP7_75t_R g66 ( 
.A(n_47),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_45),
.Y(n_67)
);

OA22x2_ASAP7_75t_L g68 ( 
.A1(n_43),
.A2(n_30),
.B1(n_36),
.B2(n_26),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_57),
.Y(n_83)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_69),
.B(n_70),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_45),
.Y(n_70)
);

A2O1A1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_66),
.A2(n_47),
.B(n_50),
.C(n_22),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_74),
.B(n_17),
.Y(n_94)
);

NOR2xp67_ASAP7_75t_L g79 ( 
.A(n_54),
.B(n_59),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_79),
.B(n_21),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_80),
.A2(n_83),
.B1(n_55),
.B2(n_65),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_68),
.A2(n_34),
.B1(n_17),
.B2(n_23),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_86),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_62),
.B(n_23),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_71),
.A2(n_68),
.B(n_61),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_89),
.A2(n_90),
.B(n_95),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_83),
.A2(n_57),
.B(n_24),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_87),
.A2(n_24),
.B1(n_20),
.B2(n_17),
.Y(n_91)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_91),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_71),
.B(n_20),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_84),
.C(n_72),
.Y(n_107)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_93),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_94),
.B(n_98),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_87),
.A2(n_16),
.B(n_17),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_73),
.A2(n_21),
.B1(n_16),
.B2(n_2),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_96),
.B(n_99),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_80),
.A2(n_21),
.B1(n_16),
.B2(n_2),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_72),
.B(n_0),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_100),
.B(n_86),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_75),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_101),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_103),
.B(n_112),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_74),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_105),
.B(n_90),
.C(n_97),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_107),
.B(n_85),
.C(n_78),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_100),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_109),
.B(n_93),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_114),
.B(n_115),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_102),
.A2(n_110),
.B1(n_108),
.B2(n_104),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_116),
.B(n_117),
.C(n_118),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_105),
.B(n_97),
.C(n_76),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_102),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_119),
.Y(n_126)
);

AOI322xp5_ASAP7_75t_SL g120 ( 
.A1(n_106),
.A2(n_95),
.A3(n_89),
.B1(n_81),
.B2(n_99),
.C1(n_84),
.C2(n_85),
.Y(n_120)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_120),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_113),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_124),
.A2(n_107),
.B(n_111),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_117),
.A2(n_111),
.B1(n_104),
.B2(n_103),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_125),
.A2(n_78),
.B1(n_82),
.B2(n_7),
.Y(n_129)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_127),
.Y(n_134)
);

NOR3xp33_ASAP7_75t_SL g128 ( 
.A(n_123),
.B(n_120),
.C(n_82),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_128),
.B(n_123),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_129),
.B(n_130),
.C(n_122),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_121),
.B(n_8),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_131),
.A2(n_125),
.B1(n_124),
.B2(n_126),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_132),
.B(n_133),
.C(n_12),
.Y(n_137)
);

BUFx24_ASAP7_75t_SL g133 ( 
.A(n_127),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_135),
.B(n_136),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_134),
.A2(n_121),
.B(n_8),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_137),
.B(n_12),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_139),
.A2(n_13),
.B(n_1),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_138),
.C(n_1),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_3),
.Y(n_142)
);


endmodule