module fake_jpeg_6159_n_271 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_271);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_271;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx5_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_13),
.B(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

CKINVDCx14_ASAP7_75t_R g63 ( 
.A(n_34),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_30),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_38),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_37),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_30),
.Y(n_38)
);

INVx8_ASAP7_75t_SL g39 ( 
.A(n_18),
.Y(n_39)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_39),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_42),
.Y(n_57)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_44),
.B(n_16),
.Y(n_86)
);

BUFx16f_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_45),
.B(n_48),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_24),
.B(n_7),
.Y(n_47)
);

A2O1A1Ixp33_ASAP7_75t_L g55 ( 
.A1(n_47),
.A2(n_24),
.B(n_17),
.C(n_20),
.Y(n_55)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_50),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_52),
.B(n_54),
.Y(n_101)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_55),
.B(n_60),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_41),
.A2(n_28),
.B1(n_20),
.B2(n_29),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_56),
.A2(n_67),
.B(n_69),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_36),
.A2(n_20),
.B1(n_33),
.B2(n_28),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_58),
.A2(n_59),
.B1(n_66),
.B2(n_21),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_38),
.A2(n_33),
.B1(n_28),
.B2(n_17),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_62),
.B(n_65),
.Y(n_113)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_64),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_41),
.A2(n_32),
.B1(n_19),
.B2(n_15),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_42),
.A2(n_32),
.B1(n_19),
.B2(n_15),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_68),
.B(n_71),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_44),
.A2(n_25),
.B1(n_26),
.B2(n_22),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_70),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g73 ( 
.A(n_37),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_73),
.B(n_74),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_43),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_78),
.B(n_80),
.Y(n_120)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_47),
.B(n_16),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_79),
.B(n_81),
.Y(n_108)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_43),
.B(n_26),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_37),
.Y(n_82)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_40),
.Y(n_83)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_83),
.Y(n_114)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_84),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_40),
.B(n_22),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_86),
.Y(n_97)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_34),
.Y(n_87)
);

BUFx5_ASAP7_75t_L g119 ( 
.A(n_87),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_43),
.A2(n_25),
.B1(n_21),
.B2(n_27),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_88),
.A2(n_93),
.B1(n_2),
.B2(n_3),
.Y(n_105)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_35),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_89),
.A2(n_96),
.B1(n_4),
.B2(n_5),
.Y(n_118)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_34),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_91),
.Y(n_103)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_34),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_43),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_94),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_35),
.A2(n_27),
.B1(n_21),
.B2(n_3),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_34),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_35),
.B(n_27),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_95),
.B(n_49),
.Y(n_107)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_35),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_99),
.A2(n_100),
.B1(n_111),
.B2(n_121),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_56),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_0),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_107),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_105),
.A2(n_76),
.B1(n_61),
.B2(n_121),
.Y(n_128)
);

OAI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_61),
.A2(n_9),
.B1(n_4),
.B2(n_5),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_51),
.B(n_2),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_116),
.B(n_123),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_118),
.B(n_10),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_88),
.A2(n_6),
.B1(n_8),
.B2(n_10),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_69),
.B(n_67),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_79),
.B(n_8),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_125),
.B(n_10),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_123),
.A2(n_57),
.B(n_77),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_126),
.A2(n_128),
.B(n_100),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_104),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_127),
.Y(n_178)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_119),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_130),
.B(n_131),
.Y(n_164)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_119),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_SL g132 ( 
.A(n_108),
.B(n_72),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_132),
.B(n_151),
.C(n_152),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_97),
.B(n_96),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_133),
.B(n_138),
.Y(n_179)
);

O2A1O1Ixp33_ASAP7_75t_L g135 ( 
.A1(n_105),
.A2(n_93),
.B(n_80),
.C(n_76),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_135),
.A2(n_101),
.B(n_109),
.Y(n_173)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_117),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_136),
.B(n_137),
.Y(n_165)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_117),
.Y(n_137)
);

AOI21xp33_ASAP7_75t_L g139 ( 
.A1(n_116),
.A2(n_52),
.B(n_65),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_SL g158 ( 
.A(n_139),
.B(n_145),
.C(n_97),
.Y(n_158)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_104),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_140),
.B(n_141),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_103),
.B(n_82),
.Y(n_142)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_142),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_103),
.B(n_73),
.Y(n_143)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_143),
.Y(n_168)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_115),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_144),
.B(n_148),
.Y(n_162)
);

OAI21xp33_ASAP7_75t_L g145 ( 
.A1(n_106),
.A2(n_89),
.B(n_53),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_113),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_147),
.Y(n_175)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_115),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_108),
.B(n_63),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_149),
.B(n_156),
.Y(n_171)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_114),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_150),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_112),
.B(n_53),
.C(n_68),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_112),
.B(n_62),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g153 ( 
.A(n_113),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_153),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_122),
.B(n_71),
.Y(n_154)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_154),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_106),
.A2(n_78),
.B(n_75),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_155),
.A2(n_98),
.B(n_122),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_108),
.B(n_11),
.Y(n_156)
);

INVx2_ASAP7_75t_SL g157 ( 
.A(n_114),
.Y(n_157)
);

AO22x1_ASAP7_75t_L g169 ( 
.A1(n_157),
.A2(n_98),
.B1(n_120),
.B2(n_110),
.Y(n_169)
);

CKINVDCx14_ASAP7_75t_R g192 ( 
.A(n_158),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_159),
.A2(n_173),
.B(n_182),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_135),
.A2(n_99),
.B1(n_75),
.B2(n_107),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_161),
.A2(n_163),
.B1(n_184),
.B2(n_144),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_146),
.A2(n_120),
.B1(n_110),
.B2(n_102),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_152),
.B(n_102),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_166),
.B(n_185),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_149),
.B(n_125),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_167),
.B(n_129),
.Y(n_197)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_169),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_134),
.B(n_124),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_176),
.B(n_147),
.Y(n_188)
);

A2O1A1O1Ixp25_ASAP7_75t_L g180 ( 
.A1(n_126),
.A2(n_125),
.B(n_101),
.C(n_124),
.D(n_109),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_180),
.B(n_183),
.Y(n_194)
);

NAND2xp33_ASAP7_75t_L g183 ( 
.A(n_155),
.B(n_11),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_134),
.A2(n_12),
.B1(n_13),
.B2(n_151),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_127),
.B(n_13),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_140),
.A2(n_132),
.B1(n_136),
.B2(n_137),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_186),
.A2(n_157),
.B1(n_150),
.B2(n_131),
.Y(n_205)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_188),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_164),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_191),
.B(n_202),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_176),
.A2(n_156),
.B(n_129),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_193),
.B(n_197),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_174),
.B(n_186),
.C(n_166),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_195),
.B(n_201),
.C(n_184),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_166),
.B(n_129),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_196),
.B(n_167),
.C(n_171),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_198),
.B(n_203),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_178),
.B(n_148),
.Y(n_199)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_199),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_182),
.A2(n_138),
.B(n_157),
.Y(n_200)
);

OAI21xp33_ASAP7_75t_L g209 ( 
.A1(n_200),
.A2(n_175),
.B(n_179),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_174),
.B(n_159),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_165),
.B(n_138),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_169),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_169),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_204),
.B(n_207),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_205),
.B(n_206),
.Y(n_225)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_162),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_162),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_208),
.B(n_212),
.C(n_214),
.Y(n_231)
);

O2A1O1Ixp33_ASAP7_75t_L g226 ( 
.A1(n_209),
.A2(n_188),
.B(n_187),
.C(n_197),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_201),
.B(n_173),
.C(n_171),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_195),
.B(n_161),
.C(n_160),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_215),
.B(n_222),
.C(n_224),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_199),
.B(n_160),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_216),
.B(n_219),
.Y(n_228)
);

AO32x1_ASAP7_75t_L g217 ( 
.A1(n_200),
.A2(n_180),
.A3(n_158),
.B1(n_185),
.B2(n_175),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_217),
.A2(n_194),
.B(n_172),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_191),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_193),
.B(n_168),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_221),
.B(n_205),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_196),
.B(n_163),
.C(n_168),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_192),
.B(n_181),
.C(n_177),
.Y(n_224)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_226),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_211),
.B(n_187),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_227),
.B(n_233),
.Y(n_239)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_229),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_223),
.A2(n_198),
.B1(n_190),
.B2(n_204),
.Y(n_230)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_230),
.Y(n_246)
);

OA22x2_ASAP7_75t_L g232 ( 
.A1(n_217),
.A2(n_190),
.B1(n_194),
.B2(n_189),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_232),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_208),
.B(n_189),
.Y(n_233)
);

XOR2x2_ASAP7_75t_L g235 ( 
.A(n_209),
.B(n_189),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_235),
.B(n_236),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_225),
.A2(n_170),
.B1(n_185),
.B2(n_130),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_237),
.B(n_224),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_233),
.B(n_214),
.C(n_222),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_238),
.B(n_231),
.C(n_234),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_240),
.B(n_244),
.Y(n_249)
);

NOR3xp33_ASAP7_75t_SL g244 ( 
.A(n_232),
.B(n_218),
.C(n_220),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_247),
.B(n_248),
.Y(n_260)
);

BUFx24_ASAP7_75t_SL g248 ( 
.A(n_245),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_238),
.B(n_231),
.C(n_234),
.Y(n_250)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_250),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_241),
.A2(n_246),
.B(n_243),
.Y(n_251)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_251),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_227),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_252),
.B(n_254),
.Y(n_256)
);

INVx11_ASAP7_75t_L g253 ( 
.A(n_244),
.Y(n_253)
);

AOI322xp5_ASAP7_75t_L g259 ( 
.A1(n_253),
.A2(n_232),
.A3(n_210),
.B1(n_230),
.B2(n_219),
.C1(n_226),
.C2(n_242),
.Y(n_259)
);

OR2x2_ASAP7_75t_L g254 ( 
.A(n_241),
.B(n_235),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_249),
.B(n_213),
.Y(n_257)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_257),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_259),
.A2(n_228),
.B(n_232),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_255),
.B(n_170),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_261),
.B(n_256),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_262),
.A2(n_257),
.B(n_258),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_256),
.A2(n_254),
.B(n_252),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_264),
.A2(n_253),
.B(n_239),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_265),
.B(n_263),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_266),
.B(n_267),
.C(n_260),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_268),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_270),
.B(n_269),
.Y(n_271)
);


endmodule