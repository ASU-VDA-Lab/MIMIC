module fake_jpeg_29025_n_72 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_72);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_72;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_71;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;
wire n_70;
wire n_66;

INVx13_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_12),
.B(n_21),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

HAxp5_ASAP7_75t_SL g32 ( 
.A(n_11),
.B(n_0),
.CON(n_32),
.SN(n_32)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_13),
.C(n_24),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_32),
.C(n_29),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_30),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_30),
.Y(n_35)
);

CKINVDCx14_ASAP7_75t_R g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_29),
.A2(n_10),
.B1(n_23),
.B2(n_22),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_37),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_40)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_29),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_39),
.A2(n_4),
.B(n_5),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_40),
.A2(n_42),
.B(n_15),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_44),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_35),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_43),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_26),
.Y(n_45)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_46),
.A2(n_37),
.B1(n_28),
.B2(n_38),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_53),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_48),
.A2(n_36),
.B1(n_26),
.B2(n_31),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_SL g53 ( 
.A1(n_44),
.A2(n_31),
.B(n_7),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g54 ( 
.A1(n_47),
.A2(n_6),
.B(n_9),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_17),
.C(n_19),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_55),
.Y(n_58)
);

XNOR2x1_ASAP7_75t_L g61 ( 
.A(n_57),
.B(n_16),
.Y(n_61)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_64),
.C(n_56),
.Y(n_65)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_63),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_65),
.B(n_49),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_68),
.B(n_69),
.C(n_67),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_66),
.A2(n_62),
.B1(n_59),
.B2(n_51),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_70),
.B(n_58),
.C(n_62),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_71),
.B(n_20),
.C(n_25),
.Y(n_72)
);


endmodule