module fake_jpeg_23459_n_177 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_177);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_177;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_SL g14 ( 
.A(n_5),
.B(n_10),
.Y(n_14)
);

BUFx12_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_4),
.B(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx11_ASAP7_75t_SL g23 ( 
.A(n_9),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_29),
.B(n_34),
.Y(n_42)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_37),
.Y(n_38)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_40),
.B(n_43),
.Y(n_55)
);

CKINVDCx12_ASAP7_75t_R g41 ( 
.A(n_36),
.Y(n_41)
);

INVx4_ASAP7_75t_SL g56 ( 
.A(n_41),
.Y(n_56)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_34),
.B(n_14),
.Y(n_45)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_35),
.A2(n_22),
.B1(n_26),
.B2(n_25),
.Y(n_46)
);

OAI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_46),
.A2(n_25),
.B1(n_22),
.B2(n_24),
.Y(n_65)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_50),
.Y(n_59)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_53),
.Y(n_64)
);

OA22x2_ASAP7_75t_L g54 ( 
.A1(n_46),
.A2(n_30),
.B1(n_16),
.B2(n_18),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_54),
.A2(n_57),
.B1(n_65),
.B2(n_35),
.Y(n_73)
);

OA22x2_ASAP7_75t_L g57 ( 
.A1(n_47),
.A2(n_30),
.B1(n_16),
.B2(n_18),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_18),
.Y(n_58)
);

OAI21xp33_ASAP7_75t_L g78 ( 
.A1(n_58),
.A2(n_13),
.B(n_27),
.Y(n_78)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_61),
.Y(n_71)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_32),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_68),
.B(n_38),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_51),
.A2(n_24),
.B1(n_26),
.B2(n_23),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_69),
.A2(n_61),
.B1(n_60),
.B2(n_29),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_62),
.B(n_14),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_70),
.Y(n_95)
);

AO21x1_ASAP7_75t_SL g91 ( 
.A1(n_73),
.A2(n_54),
.B(n_57),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_62),
.A2(n_39),
.B1(n_33),
.B2(n_49),
.Y(n_74)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_78),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_54),
.A2(n_39),
.B1(n_33),
.B2(n_49),
.Y(n_76)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_68),
.A2(n_52),
.B(n_13),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_79),
.B(n_83),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_80),
.A2(n_37),
.B1(n_67),
.B2(n_66),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_58),
.B(n_32),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_82),
.B(n_86),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_58),
.B(n_52),
.C(n_37),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_64),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_84),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_64),
.B(n_20),
.Y(n_85)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_59),
.B(n_27),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_71),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_71),
.Y(n_105)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_81),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_91),
.A2(n_98),
.B1(n_77),
.B2(n_56),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_55),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_94),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_70),
.B(n_17),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_82),
.A2(n_54),
.B1(n_57),
.B2(n_56),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_96),
.A2(n_77),
.B1(n_17),
.B2(n_20),
.Y(n_118)
);

AND2x2_ASAP7_75t_SL g101 ( 
.A(n_86),
.B(n_67),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_101),
.A2(n_72),
.B(n_66),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_87),
.A2(n_79),
.B(n_83),
.Y(n_103)
);

OAI21xp33_ASAP7_75t_L g121 ( 
.A1(n_103),
.A2(n_106),
.B(n_112),
.Y(n_121)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_105),
.Y(n_125)
);

A2O1A1Ixp33_ASAP7_75t_SL g106 ( 
.A1(n_91),
.A2(n_76),
.B(n_80),
.C(n_57),
.Y(n_106)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_107),
.Y(n_132)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_108),
.B(n_109),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_102),
.Y(n_109)
);

AOI322xp5_ASAP7_75t_L g110 ( 
.A1(n_93),
.A2(n_83),
.A3(n_73),
.B1(n_84),
.B2(n_85),
.C1(n_74),
.C2(n_63),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_110),
.B(n_116),
.C(n_101),
.Y(n_119)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_111),
.B(n_114),
.Y(n_120)
);

OAI21xp33_ASAP7_75t_L g112 ( 
.A1(n_88),
.A2(n_1),
.B(n_2),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_101),
.B(n_72),
.Y(n_113)
);

OAI21xp33_ASAP7_75t_L g128 ( 
.A1(n_113),
.A2(n_115),
.B(n_89),
.Y(n_128)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_102),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_90),
.B(n_81),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_117),
.A2(n_118),
.B1(n_99),
.B2(n_90),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_126),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_111),
.B(n_97),
.C(n_93),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_122),
.B(n_123),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_97),
.C(n_93),
.Y(n_123)
);

MAJx2_ASAP7_75t_L g126 ( 
.A(n_108),
.B(n_96),
.C(n_95),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_99),
.C(n_89),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_127),
.B(n_105),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_128),
.B(n_131),
.Y(n_140)
);

NOR2x1_ASAP7_75t_L g129 ( 
.A(n_118),
.B(n_100),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_129),
.B(n_100),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_130),
.A2(n_106),
.B1(n_109),
.B2(n_104),
.Y(n_136)
);

MAJx2_ASAP7_75t_L g131 ( 
.A(n_104),
.B(n_115),
.C(n_106),
.Y(n_131)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_133),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_124),
.B(n_114),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_134),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_135),
.B(n_136),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_129),
.B(n_94),
.Y(n_138)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_138),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_125),
.A2(n_77),
.B1(n_106),
.B2(n_3),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_139),
.A2(n_142),
.B1(n_121),
.B2(n_15),
.Y(n_152)
);

INVxp33_ASAP7_75t_L g141 ( 
.A(n_120),
.Y(n_141)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_141),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_131),
.A2(n_106),
.B1(n_123),
.B2(n_128),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_132),
.B(n_19),
.Y(n_143)
);

OAI322xp33_ASAP7_75t_L g149 ( 
.A1(n_143),
.A2(n_126),
.A3(n_19),
.B1(n_121),
.B2(n_11),
.C1(n_6),
.C2(n_7),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_144),
.B(n_122),
.Y(n_146)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_146),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_149),
.B(n_1),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_152),
.B(n_137),
.Y(n_157)
);

AO21x1_ASAP7_75t_L g153 ( 
.A1(n_140),
.A2(n_139),
.B(n_141),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_153),
.B(n_140),
.Y(n_154)
);

AOI322xp5_ASAP7_75t_L g162 ( 
.A1(n_154),
.A2(n_151),
.A3(n_152),
.B1(n_147),
.B2(n_146),
.C1(n_7),
.C2(n_8),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_155),
.B(n_159),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_145),
.B(n_137),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_156),
.B(n_1),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_157),
.A2(n_160),
.B1(n_147),
.B2(n_3),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_150),
.B(n_15),
.Y(n_159)
);

OAI31xp33_ASAP7_75t_L g160 ( 
.A1(n_153),
.A2(n_144),
.A3(n_2),
.B(n_3),
.Y(n_160)
);

NOR3xp33_ASAP7_75t_SL g161 ( 
.A(n_160),
.B(n_145),
.C(n_148),
.Y(n_161)
);

OR2x2_ASAP7_75t_L g170 ( 
.A(n_161),
.B(n_162),
.Y(n_170)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_164),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_165),
.B(n_166),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_158),
.B(n_4),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_162),
.A2(n_6),
.B(n_8),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_168),
.Y(n_171)
);

OR2x2_ASAP7_75t_L g172 ( 
.A(n_170),
.B(n_163),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_172),
.A2(n_9),
.B1(n_10),
.B2(n_171),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_167),
.B(n_169),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_173),
.A2(n_9),
.B(n_10),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_174),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_175),
.Y(n_177)
);


endmodule