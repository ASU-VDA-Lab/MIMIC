module fake_jpeg_1931_n_153 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_153);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_153;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_32),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_9),
.B(n_14),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_15),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_6),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_24),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_34),
.Y(n_50)
);

BUFx4f_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_6),
.Y(n_52)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_38),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_55),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

INVx2_ASAP7_75t_R g57 ( 
.A(n_53),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_46),
.Y(n_68)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_39),
.Y(n_59)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_59),
.Y(n_64)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_58),
.A2(n_42),
.B1(n_41),
.B2(n_51),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_L g82 ( 
.A1(n_61),
.A2(n_43),
.B1(n_44),
.B2(n_48),
.Y(n_82)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_60),
.Y(n_62)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

OR2x4_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_53),
.Y(n_66)
);

NAND3xp33_ASAP7_75t_L g73 ( 
.A(n_66),
.B(n_68),
.C(n_42),
.Y(n_73)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_54),
.A2(n_48),
.B1(n_44),
.B2(n_43),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_71),
.B(n_51),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_63),
.B(n_68),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_72),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_73),
.A2(n_76),
.B(n_77),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_70),
.Y(n_75)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_75),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_68),
.B(n_55),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_49),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_49),
.Y(n_79)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_81),
.A2(n_82),
.B1(n_3),
.B2(n_4),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_45),
.Y(n_83)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_65),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_19),
.C(n_35),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_82),
.A2(n_51),
.B1(n_56),
.B2(n_69),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_89),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_84),
.A2(n_50),
.B1(n_47),
.B2(n_2),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_88),
.A2(n_91),
.B1(n_92),
.B2(n_93),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_80),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_SL g90 ( 
.A(n_74),
.B(n_17),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_90),
.B(n_99),
.C(n_9),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_74),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_75),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_93)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_100),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_96),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_104),
.A2(n_12),
.B1(n_13),
.B2(n_37),
.Y(n_123)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_105),
.B(n_106),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_99),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_109),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_98),
.B(n_10),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_96),
.A2(n_10),
.B(n_11),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_110),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_101),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_111),
.B(n_112),
.Y(n_127)
);

AOI322xp5_ASAP7_75t_L g112 ( 
.A1(n_97),
.A2(n_25),
.A3(n_33),
.B1(n_28),
.B2(n_18),
.C1(n_20),
.C2(n_23),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_26),
.C(n_27),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_113),
.B(n_108),
.C(n_106),
.Y(n_119)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_101),
.Y(n_114)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_114),
.Y(n_121)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_115),
.Y(n_124)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_116),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_87),
.Y(n_117)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_117),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_11),
.Y(n_118)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_118),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_128),
.C(n_129),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_111),
.A2(n_103),
.B(n_102),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_122),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_123),
.B(n_126),
.Y(n_133)
);

INVx1_ASAP7_75t_SL g126 ( 
.A(n_103),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_110),
.A2(n_12),
.B(n_13),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_132),
.A2(n_104),
.B(n_113),
.Y(n_135)
);

XNOR2x1_ASAP7_75t_L g134 ( 
.A(n_120),
.B(n_107),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_134),
.B(n_136),
.C(n_138),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_135),
.Y(n_142)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_121),
.Y(n_137)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_137),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_131),
.B(n_119),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_134),
.B(n_127),
.C(n_130),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_143),
.B(n_130),
.Y(n_145)
);

OR2x2_ASAP7_75t_L g144 ( 
.A(n_142),
.B(n_133),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_144),
.A2(n_145),
.B(n_146),
.Y(n_147)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_140),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_147),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_141),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_149),
.A2(n_139),
.B(n_125),
.Y(n_150)
);

BUFx24_ASAP7_75t_SL g151 ( 
.A(n_150),
.Y(n_151)
);

XNOR2x2_ASAP7_75t_SL g152 ( 
.A(n_151),
.B(n_139),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_124),
.Y(n_153)
);


endmodule