module real_aes_7143_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_666;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_504;
wire n_310;
wire n_455;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_417;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_617;
wire n_602;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
AOI222xp33_ASAP7_75t_SL g128 ( .A1(n_0), .A2(n_129), .B1(n_135), .B2(n_724), .C1(n_725), .C2(n_728), .Y(n_128) );
INVx1_ASAP7_75t_L g109 ( .A(n_1), .Y(n_109) );
INVx1_ASAP7_75t_L g465 ( .A(n_2), .Y(n_465) );
INVx1_ASAP7_75t_L g268 ( .A(n_3), .Y(n_268) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_4), .A2(n_38), .B1(n_218), .B2(n_504), .Y(n_540) );
AOI21xp33_ASAP7_75t_L g229 ( .A1(n_5), .A2(n_151), .B(n_230), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_6), .B(n_173), .Y(n_490) );
AND2x6_ASAP7_75t_L g156 ( .A(n_7), .B(n_157), .Y(n_156) );
AOI21xp5_ASAP7_75t_L g149 ( .A1(n_8), .A2(n_150), .B(n_158), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_9), .B(n_115), .Y(n_114) );
NOR2xp33_ASAP7_75t_L g126 ( .A(n_9), .B(n_39), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_10), .B(n_216), .Y(n_215) );
INVx1_ASAP7_75t_L g235 ( .A(n_11), .Y(n_235) );
INVx1_ASAP7_75t_L g148 ( .A(n_12), .Y(n_148) );
INVx1_ASAP7_75t_L g459 ( .A(n_13), .Y(n_459) );
INVx1_ASAP7_75t_L g168 ( .A(n_14), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_15), .B(n_242), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_16), .B(n_174), .Y(n_492) );
AO32x2_ASAP7_75t_L g538 ( .A1(n_17), .A2(n_173), .A3(n_189), .B1(n_478), .B2(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_18), .B(n_218), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_19), .B(n_185), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_20), .B(n_174), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_21), .A2(n_49), .B1(n_218), .B2(n_504), .Y(n_541) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_22), .B(n_151), .Y(n_178) );
AOI22xp33_ASAP7_75t_SL g505 ( .A1(n_23), .A2(n_77), .B1(n_218), .B2(n_242), .Y(n_505) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_24), .B(n_218), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_25), .B(n_228), .Y(n_258) );
A2O1A1Ixp33_ASAP7_75t_L g164 ( .A1(n_26), .A2(n_165), .B(n_167), .C(n_169), .Y(n_164) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_27), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_28), .B(n_144), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_29), .B(n_200), .Y(n_269) );
OAI22xp5_ASAP7_75t_L g130 ( .A1(n_30), .A2(n_101), .B1(n_131), .B2(n_132), .Y(n_130) );
INVx1_ASAP7_75t_L g132 ( .A(n_30), .Y(n_132) );
INVx1_ASAP7_75t_L g247 ( .A(n_31), .Y(n_247) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_32), .A2(n_104), .B1(n_116), .B2(n_744), .Y(n_103) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_33), .B(n_144), .Y(n_516) );
INVx2_ASAP7_75t_L g154 ( .A(n_34), .Y(n_154) );
NAND2xp5_ASAP7_75t_SL g473 ( .A(n_35), .B(n_218), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_36), .B(n_144), .Y(n_526) );
A2O1A1Ixp33_ASAP7_75t_L g179 ( .A1(n_37), .A2(n_156), .B(n_161), .C(n_180), .Y(n_179) );
INVx1_ASAP7_75t_L g115 ( .A(n_39), .Y(n_115) );
INVx1_ASAP7_75t_L g245 ( .A(n_40), .Y(n_245) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_41), .B(n_200), .Y(n_199) );
NAND2xp5_ASAP7_75t_SL g485 ( .A(n_42), .B(n_218), .Y(n_485) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_43), .A2(n_87), .B1(n_170), .B2(n_504), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g488 ( .A(n_44), .B(n_218), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_45), .B(n_218), .Y(n_460) );
CKINVDCx16_ASAP7_75t_R g248 ( .A(n_46), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_47), .B(n_464), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_48), .B(n_151), .Y(n_219) );
AOI22xp33_ASAP7_75t_SL g496 ( .A1(n_50), .A2(n_60), .B1(n_218), .B2(n_242), .Y(n_496) );
OAI22xp5_ASAP7_75t_SL g736 ( .A1(n_51), .A2(n_737), .B1(n_740), .B2(n_741), .Y(n_736) );
CKINVDCx20_ASAP7_75t_R g740 ( .A(n_51), .Y(n_740) );
AOI22xp5_ASAP7_75t_L g241 ( .A1(n_52), .A2(n_161), .B1(n_242), .B2(n_244), .Y(n_241) );
CKINVDCx20_ASAP7_75t_R g191 ( .A(n_53), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g477 ( .A(n_54), .B(n_218), .Y(n_477) );
CKINVDCx16_ASAP7_75t_R g265 ( .A(n_55), .Y(n_265) );
NAND2xp5_ASAP7_75t_SL g520 ( .A(n_56), .B(n_218), .Y(n_520) );
A2O1A1Ixp33_ASAP7_75t_L g232 ( .A1(n_57), .A2(n_233), .B(n_234), .C(n_236), .Y(n_232) );
CKINVDCx20_ASAP7_75t_R g204 ( .A(n_58), .Y(n_204) );
INVx1_ASAP7_75t_L g231 ( .A(n_59), .Y(n_231) );
INVx1_ASAP7_75t_L g157 ( .A(n_61), .Y(n_157) );
OAI22xp5_ASAP7_75t_SL g129 ( .A1(n_62), .A2(n_130), .B1(n_133), .B2(n_134), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g134 ( .A(n_62), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_63), .B(n_218), .Y(n_466) );
INVx1_ASAP7_75t_L g147 ( .A(n_64), .Y(n_147) );
OAI22xp5_ASAP7_75t_SL g737 ( .A1(n_65), .A2(n_76), .B1(n_738), .B2(n_739), .Y(n_737) );
CKINVDCx20_ASAP7_75t_R g738 ( .A(n_65), .Y(n_738) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_66), .Y(n_120) );
AO32x2_ASAP7_75t_L g501 ( .A1(n_67), .A2(n_173), .A3(n_210), .B1(n_478), .B2(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g476 ( .A(n_68), .Y(n_476) );
INVx1_ASAP7_75t_L g511 ( .A(n_69), .Y(n_511) );
A2O1A1Ixp33_ASAP7_75t_SL g255 ( .A1(n_70), .A2(n_185), .B(n_236), .C(n_256), .Y(n_255) );
INVxp67_ASAP7_75t_L g257 ( .A(n_71), .Y(n_257) );
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_72), .B(n_242), .Y(n_512) );
INVx1_ASAP7_75t_L g112 ( .A(n_73), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g250 ( .A(n_74), .Y(n_250) );
INVx1_ASAP7_75t_L g195 ( .A(n_75), .Y(n_195) );
CKINVDCx20_ASAP7_75t_R g739 ( .A(n_76), .Y(n_739) );
A2O1A1Ixp33_ASAP7_75t_L g197 ( .A1(n_78), .A2(n_156), .B(n_161), .C(n_198), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_79), .B(n_504), .Y(n_525) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_80), .B(n_242), .Y(n_515) );
NAND2xp5_ASAP7_75t_SL g181 ( .A(n_81), .B(n_182), .Y(n_181) );
INVx2_ASAP7_75t_L g145 ( .A(n_82), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_83), .B(n_185), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_84), .B(n_242), .Y(n_486) );
A2O1A1Ixp33_ASAP7_75t_L g266 ( .A1(n_85), .A2(n_156), .B(n_161), .C(n_267), .Y(n_266) );
NAND3xp33_ASAP7_75t_SL g108 ( .A(n_86), .B(n_109), .C(n_110), .Y(n_108) );
OR2x2_ASAP7_75t_L g123 ( .A(n_86), .B(n_124), .Y(n_123) );
OR2x2_ASAP7_75t_L g136 ( .A(n_86), .B(n_125), .Y(n_136) );
INVx2_ASAP7_75t_L g448 ( .A(n_86), .Y(n_448) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_88), .A2(n_102), .B1(n_242), .B2(n_243), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_89), .B(n_144), .Y(n_237) );
CKINVDCx20_ASAP7_75t_R g272 ( .A(n_90), .Y(n_272) );
A2O1A1Ixp33_ASAP7_75t_L g212 ( .A1(n_91), .A2(n_156), .B(n_161), .C(n_213), .Y(n_212) );
CKINVDCx20_ASAP7_75t_R g221 ( .A(n_92), .Y(n_221) );
INVx1_ASAP7_75t_L g254 ( .A(n_93), .Y(n_254) );
CKINVDCx16_ASAP7_75t_R g159 ( .A(n_94), .Y(n_159) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_95), .Y(n_127) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_96), .B(n_182), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_97), .B(n_242), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_98), .B(n_173), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_99), .B(n_112), .Y(n_111) );
AOI21xp5_ASAP7_75t_L g252 ( .A1(n_100), .A2(n_151), .B(n_253), .Y(n_252) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_101), .Y(n_131) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx2_ASAP7_75t_SL g746 ( .A(n_106), .Y(n_746) );
AND2x2_ASAP7_75t_SL g106 ( .A(n_107), .B(n_113), .Y(n_106) );
CKINVDCx16_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
AND2x2_ASAP7_75t_L g125 ( .A(n_109), .B(n_126), .Y(n_125) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
INVxp67_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
AOI22x1_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_128), .B1(n_731), .B2(n_733), .Y(n_116) );
NOR2xp33_ASAP7_75t_L g117 ( .A(n_118), .B(n_121), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx2_ASAP7_75t_L g732 ( .A(n_120), .Y(n_732) );
AOI21xp5_ASAP7_75t_L g733 ( .A1(n_121), .A2(n_734), .B(n_742), .Y(n_733) );
NOR2xp33_ASAP7_75t_SL g121 ( .A(n_122), .B(n_127), .Y(n_121) );
HB1xp67_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx1_ASAP7_75t_SL g743 ( .A(n_123), .Y(n_743) );
NOR2x2_ASAP7_75t_L g730 ( .A(n_124), .B(n_448), .Y(n_730) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
OR2x2_ASAP7_75t_L g447 ( .A(n_125), .B(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g724 ( .A(n_129), .Y(n_724) );
INVx1_ASAP7_75t_L g133 ( .A(n_130), .Y(n_133) );
OAI22xp5_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_137), .B1(n_445), .B2(n_449), .Y(n_135) );
OAI22xp5_ASAP7_75t_SL g725 ( .A1(n_136), .A2(n_447), .B1(n_726), .B2(n_727), .Y(n_725) );
INVx2_ASAP7_75t_SL g726 ( .A(n_137), .Y(n_726) );
OAI22xp5_ASAP7_75t_SL g734 ( .A1(n_137), .A2(n_726), .B1(n_735), .B2(n_736), .Y(n_734) );
OR4x2_ASAP7_75t_L g137 ( .A(n_138), .B(n_341), .C(n_400), .D(n_427), .Y(n_137) );
NAND3xp33_ASAP7_75t_SL g138 ( .A(n_139), .B(n_283), .C(n_308), .Y(n_138) );
O2A1O1Ixp33_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_206), .B(n_226), .C(n_259), .Y(n_139) );
AOI211xp5_ASAP7_75t_SL g431 ( .A1(n_140), .A2(n_432), .B(n_434), .C(n_437), .Y(n_431) );
AND2x2_ASAP7_75t_L g140 ( .A(n_141), .B(n_175), .Y(n_140) );
INVx1_ASAP7_75t_L g306 ( .A(n_141), .Y(n_306) );
INVx1_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
OR2x2_ASAP7_75t_L g281 ( .A(n_142), .B(n_282), .Y(n_281) );
INVx2_ASAP7_75t_L g313 ( .A(n_142), .Y(n_313) );
AND2x2_ASAP7_75t_L g368 ( .A(n_142), .B(n_337), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_142), .B(n_224), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_142), .B(n_225), .Y(n_426) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx1_ASAP7_75t_L g287 ( .A(n_143), .Y(n_287) );
AND2x2_ASAP7_75t_L g330 ( .A(n_143), .B(n_193), .Y(n_330) );
AND2x2_ASAP7_75t_L g348 ( .A(n_143), .B(n_225), .Y(n_348) );
OA21x2_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_149), .B(n_172), .Y(n_143) );
INVx1_ASAP7_75t_L g205 ( .A(n_144), .Y(n_205) );
INVx2_ASAP7_75t_L g210 ( .A(n_144), .Y(n_210) );
OA21x2_ASAP7_75t_L g508 ( .A1(n_144), .A2(n_509), .B(n_516), .Y(n_508) );
OA21x2_ASAP7_75t_L g517 ( .A1(n_144), .A2(n_518), .B(n_526), .Y(n_517) );
AND2x2_ASAP7_75t_SL g144 ( .A(n_145), .B(n_146), .Y(n_144) );
AND2x2_ASAP7_75t_L g174 ( .A(n_145), .B(n_146), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_147), .B(n_148), .Y(n_146) );
BUFx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
AND2x4_ASAP7_75t_L g151 ( .A(n_152), .B(n_156), .Y(n_151) );
NAND2x1p5_ASAP7_75t_L g196 ( .A(n_152), .B(n_156), .Y(n_196) );
AND2x2_ASAP7_75t_L g152 ( .A(n_153), .B(n_155), .Y(n_152) );
INVx1_ASAP7_75t_L g464 ( .A(n_153), .Y(n_464) );
INVx1_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g162 ( .A(n_154), .Y(n_162) );
INVx1_ASAP7_75t_L g243 ( .A(n_154), .Y(n_243) );
INVx1_ASAP7_75t_L g163 ( .A(n_155), .Y(n_163) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_155), .Y(n_166) );
INVx3_ASAP7_75t_L g183 ( .A(n_155), .Y(n_183) );
INVx1_ASAP7_75t_L g185 ( .A(n_155), .Y(n_185) );
BUFx6f_ASAP7_75t_L g200 ( .A(n_155), .Y(n_200) );
INVx4_ASAP7_75t_SL g171 ( .A(n_156), .Y(n_171) );
OAI21xp5_ASAP7_75t_L g457 ( .A1(n_156), .A2(n_458), .B(n_462), .Y(n_457) );
BUFx3_ASAP7_75t_L g478 ( .A(n_156), .Y(n_478) );
OAI21xp5_ASAP7_75t_L g483 ( .A1(n_156), .A2(n_484), .B(n_487), .Y(n_483) );
OAI21xp5_ASAP7_75t_L g509 ( .A1(n_156), .A2(n_510), .B(n_513), .Y(n_509) );
OAI21xp5_ASAP7_75t_L g518 ( .A1(n_156), .A2(n_519), .B(n_523), .Y(n_518) );
O2A1O1Ixp33_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_160), .B(n_164), .C(n_171), .Y(n_158) );
O2A1O1Ixp33_ASAP7_75t_L g230 ( .A1(n_160), .A2(n_171), .B(n_231), .C(n_232), .Y(n_230) );
O2A1O1Ixp33_ASAP7_75t_L g253 ( .A1(n_160), .A2(n_171), .B(n_254), .C(n_255), .Y(n_253) );
INVx5_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
AND2x6_ASAP7_75t_L g161 ( .A(n_162), .B(n_163), .Y(n_161) );
BUFx3_ASAP7_75t_L g170 ( .A(n_162), .Y(n_170) );
BUFx6f_ASAP7_75t_L g218 ( .A(n_162), .Y(n_218) );
INVx1_ASAP7_75t_L g504 ( .A(n_162), .Y(n_504) );
NOR2xp33_ASAP7_75t_L g167 ( .A(n_165), .B(n_168), .Y(n_167) );
INVx1_ASAP7_75t_L g461 ( .A(n_165), .Y(n_461) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_165), .A2(n_514), .B(n_515), .Y(n_513) );
INVx4_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
OAI22xp5_ASAP7_75t_SL g244 ( .A1(n_166), .A2(n_245), .B1(n_246), .B2(n_247), .Y(n_244) );
INVx2_ASAP7_75t_L g246 ( .A(n_166), .Y(n_246) );
INVx1_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx2_ASAP7_75t_L g187 ( .A(n_170), .Y(n_187) );
OAI22xp33_ASAP7_75t_L g240 ( .A1(n_171), .A2(n_196), .B1(n_241), .B2(n_248), .Y(n_240) );
INVx4_ASAP7_75t_L g192 ( .A(n_173), .Y(n_192) );
OA21x2_ASAP7_75t_L g251 ( .A1(n_173), .A2(n_252), .B(n_258), .Y(n_251) );
OA21x2_ASAP7_75t_L g482 ( .A1(n_173), .A2(n_483), .B(n_490), .Y(n_482) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx1_ASAP7_75t_L g189 ( .A(n_174), .Y(n_189) );
INVx4_ASAP7_75t_L g280 ( .A(n_175), .Y(n_280) );
OAI21xp5_ASAP7_75t_L g335 ( .A1(n_175), .A2(n_336), .B(n_338), .Y(n_335) );
AND2x2_ASAP7_75t_L g416 ( .A(n_175), .B(n_417), .Y(n_416) );
AND2x2_ASAP7_75t_L g175 ( .A(n_176), .B(n_193), .Y(n_175) );
INVx1_ASAP7_75t_L g223 ( .A(n_176), .Y(n_223) );
AND2x2_ASAP7_75t_L g285 ( .A(n_176), .B(n_225), .Y(n_285) );
OR2x2_ASAP7_75t_L g314 ( .A(n_176), .B(n_315), .Y(n_314) );
INVx2_ASAP7_75t_L g328 ( .A(n_176), .Y(n_328) );
INVx3_ASAP7_75t_L g337 ( .A(n_176), .Y(n_337) );
AND2x2_ASAP7_75t_L g347 ( .A(n_176), .B(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g380 ( .A(n_176), .B(n_286), .Y(n_380) );
AND2x2_ASAP7_75t_L g404 ( .A(n_176), .B(n_360), .Y(n_404) );
OR2x6_ASAP7_75t_L g176 ( .A(n_177), .B(n_190), .Y(n_176) );
AOI21xp5_ASAP7_75t_SL g177 ( .A1(n_178), .A2(n_179), .B(n_188), .Y(n_177) );
AOI21xp5_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_184), .B(n_186), .Y(n_180) );
O2A1O1Ixp33_ASAP7_75t_L g267 ( .A1(n_182), .A2(n_268), .B(n_269), .C(n_270), .Y(n_267) );
INVx2_ASAP7_75t_L g467 ( .A(n_182), .Y(n_467) );
AOI21xp5_ASAP7_75t_L g472 ( .A1(n_182), .A2(n_473), .B(n_474), .Y(n_472) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_182), .A2(n_485), .B(n_486), .Y(n_484) );
O2A1O1Ixp5_ASAP7_75t_SL g510 ( .A1(n_182), .A2(n_236), .B(n_511), .C(n_512), .Y(n_510) );
INVx5_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g234 ( .A(n_183), .B(n_235), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_183), .B(n_257), .Y(n_256) );
OAI22xp5_ASAP7_75t_SL g502 ( .A1(n_183), .A2(n_200), .B1(n_503), .B2(n_505), .Y(n_502) );
INVx1_ASAP7_75t_L g522 ( .A(n_185), .Y(n_522) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_186), .A2(n_199), .B(n_201), .Y(n_198) );
INVx2_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
INVx1_ASAP7_75t_L g202 ( .A(n_188), .Y(n_202) );
OA21x2_ASAP7_75t_L g456 ( .A1(n_188), .A2(n_457), .B(n_468), .Y(n_456) );
OA21x2_ASAP7_75t_L g470 ( .A1(n_188), .A2(n_471), .B(n_479), .Y(n_470) );
INVx2_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
AO21x2_ASAP7_75t_L g239 ( .A1(n_189), .A2(n_240), .B(n_249), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_189), .B(n_250), .Y(n_249) );
AO21x2_ASAP7_75t_L g263 ( .A1(n_189), .A2(n_264), .B(n_271), .Y(n_263) );
NOR2xp33_ASAP7_75t_SL g190 ( .A(n_191), .B(n_192), .Y(n_190) );
INVx3_ASAP7_75t_L g228 ( .A(n_192), .Y(n_228) );
NAND3xp33_ASAP7_75t_L g493 ( .A(n_192), .B(n_478), .C(n_494), .Y(n_493) );
AO21x1_ASAP7_75t_L g572 ( .A1(n_192), .A2(n_494), .B(n_573), .Y(n_572) );
INVx2_ASAP7_75t_L g225 ( .A(n_193), .Y(n_225) );
AND2x2_ASAP7_75t_L g440 ( .A(n_193), .B(n_282), .Y(n_440) );
AO21x2_ASAP7_75t_L g193 ( .A1(n_194), .A2(n_202), .B(n_203), .Y(n_193) );
OAI21xp5_ASAP7_75t_L g194 ( .A1(n_195), .A2(n_196), .B(n_197), .Y(n_194) );
OAI21xp5_ASAP7_75t_L g264 ( .A1(n_196), .A2(n_265), .B(n_266), .Y(n_264) );
INVx4_ASAP7_75t_L g216 ( .A(n_200), .Y(n_216) );
INVx2_ASAP7_75t_L g233 ( .A(n_200), .Y(n_233) );
OAI22xp5_ASAP7_75t_L g494 ( .A1(n_200), .A2(n_467), .B1(n_495), .B2(n_496), .Y(n_494) );
OAI22xp5_ASAP7_75t_L g539 ( .A1(n_200), .A2(n_467), .B1(n_540), .B2(n_541), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_204), .B(n_205), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g220 ( .A(n_205), .B(n_221), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g271 ( .A(n_205), .B(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_222), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g336 ( .A(n_208), .B(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g360 ( .A(n_208), .B(n_348), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_208), .B(n_337), .Y(n_422) );
INVx1_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx2_ASAP7_75t_L g282 ( .A(n_209), .Y(n_282) );
AND2x2_ASAP7_75t_L g286 ( .A(n_209), .B(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g327 ( .A(n_209), .B(n_328), .Y(n_327) );
AO21x2_ASAP7_75t_L g209 ( .A1(n_210), .A2(n_211), .B(n_220), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_212), .B(n_219), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_214), .A2(n_215), .B(n_217), .Y(n_213) );
HB1xp67_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVx3_ASAP7_75t_L g236 ( .A(n_218), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_222), .B(n_323), .Y(n_345) );
INVx1_ASAP7_75t_L g384 ( .A(n_222), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_222), .B(n_311), .Y(n_428) );
AND2x2_ASAP7_75t_L g222 ( .A(n_223), .B(n_224), .Y(n_222) );
AND2x2_ASAP7_75t_L g291 ( .A(n_223), .B(n_286), .Y(n_291) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_225), .B(n_282), .Y(n_315) );
INVx1_ASAP7_75t_L g394 ( .A(n_225), .Y(n_394) );
AOI322xp5_ASAP7_75t_L g418 ( .A1(n_226), .A2(n_333), .A3(n_393), .B1(n_419), .B2(n_421), .C1(n_423), .C2(n_425), .Y(n_418) );
AND2x2_ASAP7_75t_SL g226 ( .A(n_227), .B(n_238), .Y(n_226) );
AND2x2_ASAP7_75t_L g273 ( .A(n_227), .B(n_251), .Y(n_273) );
INVx1_ASAP7_75t_SL g276 ( .A(n_227), .Y(n_276) );
AND2x2_ASAP7_75t_L g278 ( .A(n_227), .B(n_239), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_227), .B(n_295), .Y(n_301) );
INVx2_ASAP7_75t_L g320 ( .A(n_227), .Y(n_320) );
AND2x2_ASAP7_75t_L g333 ( .A(n_227), .B(n_334), .Y(n_333) );
OR2x2_ASAP7_75t_L g371 ( .A(n_227), .B(n_295), .Y(n_371) );
BUFx2_ASAP7_75t_L g388 ( .A(n_227), .Y(n_388) );
AND2x2_ASAP7_75t_L g402 ( .A(n_227), .B(n_262), .Y(n_402) );
OA21x2_ASAP7_75t_L g227 ( .A1(n_228), .A2(n_229), .B(n_237), .Y(n_227) );
O2A1O1Ixp5_ASAP7_75t_L g475 ( .A1(n_233), .A2(n_463), .B(n_476), .C(n_477), .Y(n_475) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_233), .A2(n_524), .B(n_525), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_238), .B(n_290), .Y(n_317) );
AND2x2_ASAP7_75t_L g444 ( .A(n_238), .B(n_320), .Y(n_444) );
AND2x2_ASAP7_75t_L g238 ( .A(n_239), .B(n_251), .Y(n_238) );
OR2x2_ASAP7_75t_L g289 ( .A(n_239), .B(n_290), .Y(n_289) );
INVx3_ASAP7_75t_L g295 ( .A(n_239), .Y(n_295) );
AND2x2_ASAP7_75t_L g340 ( .A(n_239), .B(n_263), .Y(n_340) );
NOR2xp33_ASAP7_75t_L g387 ( .A(n_239), .B(n_388), .Y(n_387) );
HB1xp67_ASAP7_75t_L g424 ( .A(n_239), .Y(n_424) );
INVx2_ASAP7_75t_L g270 ( .A(n_242), .Y(n_270) );
INVx3_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_L g275 ( .A(n_251), .B(n_276), .Y(n_275) );
INVx1_ASAP7_75t_L g297 ( .A(n_251), .Y(n_297) );
BUFx2_ASAP7_75t_L g303 ( .A(n_251), .Y(n_303) );
AND2x2_ASAP7_75t_L g322 ( .A(n_251), .B(n_295), .Y(n_322) );
INVx3_ASAP7_75t_L g334 ( .A(n_251), .Y(n_334) );
OR2x2_ASAP7_75t_L g344 ( .A(n_251), .B(n_295), .Y(n_344) );
AOI31xp33_ASAP7_75t_SL g259 ( .A1(n_260), .A2(n_274), .A3(n_277), .B(n_279), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_261), .B(n_273), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_261), .B(n_296), .Y(n_307) );
OR2x2_ASAP7_75t_L g331 ( .A(n_261), .B(n_301), .Y(n_331) );
INVx1_ASAP7_75t_SL g261 ( .A(n_262), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_262), .B(n_275), .Y(n_274) );
OR2x2_ASAP7_75t_L g352 ( .A(n_262), .B(n_344), .Y(n_352) );
NOR2xp33_ASAP7_75t_L g362 ( .A(n_262), .B(n_334), .Y(n_362) );
AND2x2_ASAP7_75t_L g369 ( .A(n_262), .B(n_370), .Y(n_369) );
NAND2x1_ASAP7_75t_L g397 ( .A(n_262), .B(n_333), .Y(n_397) );
NOR2xp33_ASAP7_75t_L g398 ( .A(n_262), .B(n_388), .Y(n_398) );
AND2x2_ASAP7_75t_L g410 ( .A(n_262), .B(n_295), .Y(n_410) );
INVx3_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
INVx3_ASAP7_75t_L g290 ( .A(n_263), .Y(n_290) );
O2A1O1Ixp33_ASAP7_75t_L g458 ( .A1(n_270), .A2(n_459), .B(n_460), .C(n_461), .Y(n_458) );
INVx1_ASAP7_75t_L g356 ( .A(n_273), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_273), .B(n_410), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_275), .B(n_351), .Y(n_385) );
AND2x4_ASAP7_75t_L g296 ( .A(n_276), .B(n_297), .Y(n_296) );
CKINVDCx16_ASAP7_75t_R g277 ( .A(n_278), .Y(n_277) );
OR2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
INVx2_ASAP7_75t_L g375 ( .A(n_281), .Y(n_375) );
NOR2xp33_ASAP7_75t_L g392 ( .A(n_281), .B(n_393), .Y(n_392) );
AND2x2_ASAP7_75t_L g323 ( .A(n_282), .B(n_313), .Y(n_323) );
AND2x2_ASAP7_75t_L g417 ( .A(n_282), .B(n_287), .Y(n_417) );
INVx1_ASAP7_75t_L g442 ( .A(n_282), .Y(n_442) );
AOI221xp5_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_288), .B1(n_291), .B2(n_292), .C(n_298), .Y(n_283) );
CKINVDCx14_ASAP7_75t_R g304 ( .A(n_284), .Y(n_304) );
AND2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_285), .B(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_288), .B(n_339), .Y(n_358) );
INVx3_ASAP7_75t_SL g288 ( .A(n_289), .Y(n_288) );
OR2x2_ASAP7_75t_L g407 ( .A(n_289), .B(n_303), .Y(n_407) );
AND2x2_ASAP7_75t_L g321 ( .A(n_290), .B(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g351 ( .A(n_290), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_290), .B(n_334), .Y(n_379) );
NOR3xp33_ASAP7_75t_L g421 ( .A(n_290), .B(n_391), .C(n_422), .Y(n_421) );
AOI211xp5_ASAP7_75t_SL g354 ( .A1(n_291), .A2(n_355), .B(n_357), .C(n_365), .Y(n_354) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
OAI22xp33_ASAP7_75t_L g343 ( .A1(n_293), .A2(n_344), .B1(n_345), .B2(n_346), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_294), .B(n_296), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_294), .B(n_333), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_294), .B(n_378), .Y(n_377) );
BUFx2_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g436 ( .A(n_296), .B(n_410), .Y(n_436) );
OAI22xp5_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_304), .B1(n_305), .B2(n_307), .Y(n_298) );
NOR2xp33_ASAP7_75t_SL g299 ( .A(n_300), .B(n_302), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_302), .B(n_351), .Y(n_382) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
OAI22xp5_ASAP7_75t_L g434 ( .A1(n_305), .A2(n_397), .B1(n_428), .B2(n_435), .Y(n_434) );
AOI221xp5_ASAP7_75t_L g308 ( .A1(n_309), .A2(n_316), .B1(n_318), .B2(n_323), .C(n_324), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
OR2x2_ASAP7_75t_L g310 ( .A(n_311), .B(n_314), .Y(n_310) );
HB1xp67_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVxp67_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
OAI221xp5_ASAP7_75t_L g324 ( .A1(n_314), .A2(n_325), .B1(n_331), .B2(n_332), .C(n_335), .Y(n_324) );
INVx1_ASAP7_75t_L g367 ( .A(n_315), .Y(n_367) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
INVx1_ASAP7_75t_SL g339 ( .A(n_320), .Y(n_339) );
OR2x2_ASAP7_75t_L g412 ( .A(n_320), .B(n_344), .Y(n_412) );
AND2x2_ASAP7_75t_L g414 ( .A(n_320), .B(n_322), .Y(n_414) );
INVx1_ASAP7_75t_L g353 ( .A(n_323), .Y(n_353) );
OR2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_329), .Y(n_325) );
AOI21xp33_ASAP7_75t_SL g383 ( .A1(n_326), .A2(n_384), .B(n_385), .Y(n_383) );
OR2x2_ASAP7_75t_L g390 ( .A(n_326), .B(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g364 ( .A(n_327), .B(n_348), .Y(n_364) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
NAND2xp33_ASAP7_75t_SL g381 ( .A(n_332), .B(n_382), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_333), .B(n_351), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_334), .B(n_370), .Y(n_433) );
O2A1O1Ixp33_ASAP7_75t_L g349 ( .A1(n_337), .A2(n_350), .B(n_352), .C(n_353), .Y(n_349) );
NAND2x1_ASAP7_75t_SL g374 ( .A(n_337), .B(n_375), .Y(n_374) );
AOI22xp5_ASAP7_75t_L g386 ( .A1(n_338), .A2(n_387), .B1(n_389), .B2(n_392), .Y(n_386) );
AND2x2_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_340), .B(n_430), .Y(n_429) );
NAND5xp2_ASAP7_75t_L g341 ( .A(n_342), .B(n_354), .C(n_372), .D(n_386), .E(n_395), .Y(n_341) );
NOR2xp33_ASAP7_75t_L g342 ( .A(n_343), .B(n_349), .Y(n_342) );
INVx1_ASAP7_75t_L g399 ( .A(n_345), .Y(n_399) );
INVx1_ASAP7_75t_SL g346 ( .A(n_347), .Y(n_346) );
AOI221xp5_ASAP7_75t_L g405 ( .A1(n_347), .A2(n_366), .B1(n_406), .B2(n_408), .C(n_411), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_348), .B(n_442), .Y(n_441) );
NOR2xp33_ASAP7_75t_L g355 ( .A(n_351), .B(n_356), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_351), .B(n_417), .Y(n_420) );
OAI22xp5_ASAP7_75t_L g357 ( .A1(n_358), .A2(n_359), .B1(n_361), .B2(n_363), .Y(n_357) );
INVx1_ASAP7_75t_SL g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g365 ( .A(n_366), .B(n_369), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_367), .B(n_368), .Y(n_366) );
AND2x2_ASAP7_75t_L g439 ( .A(n_368), .B(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
AOI221xp5_ASAP7_75t_L g372 ( .A1(n_373), .A2(n_376), .B1(n_380), .B2(n_381), .C(n_383), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_L g423 ( .A(n_378), .B(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_SL g430 ( .A(n_388), .Y(n_430) );
INVx1_ASAP7_75t_SL g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
OAI21xp5_ASAP7_75t_SL g395 ( .A1(n_396), .A2(n_398), .B(n_399), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
OAI211xp5_ASAP7_75t_SL g400 ( .A1(n_401), .A2(n_403), .B(n_405), .C(n_418), .Y(n_400) );
INVx1_ASAP7_75t_SL g401 ( .A(n_402), .Y(n_401) );
A2O1A1Ixp33_ASAP7_75t_L g427 ( .A1(n_403), .A2(n_428), .B(n_429), .C(n_431), .Y(n_427) );
INVx1_ASAP7_75t_SL g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
NAND2xp5_ASAP7_75t_SL g408 ( .A(n_407), .B(n_409), .Y(n_408) );
AOI21xp33_ASAP7_75t_L g411 ( .A1(n_412), .A2(n_413), .B(n_415), .Y(n_411) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
AOI21xp33_ASAP7_75t_L g437 ( .A1(n_438), .A2(n_441), .B(n_443), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g727 ( .A(n_449), .Y(n_727) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
OR5x1_ASAP7_75t_L g451 ( .A(n_452), .B(n_615), .C(n_673), .D(n_709), .E(n_716), .Y(n_451) );
NAND3xp33_ASAP7_75t_SL g452 ( .A(n_453), .B(n_561), .C(n_585), .Y(n_452) );
AOI221xp5_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_497), .B1(n_527), .B2(n_532), .C(n_542), .Y(n_453) );
OAI21xp5_ASAP7_75t_SL g695 ( .A1(n_454), .A2(n_696), .B(n_698), .Y(n_695) );
AND2x2_ASAP7_75t_L g454 ( .A(n_455), .B(n_480), .Y(n_454) );
NAND2x1p5_ASAP7_75t_L g685 ( .A(n_455), .B(n_686), .Y(n_685) );
AND2x2_ASAP7_75t_L g455 ( .A(n_456), .B(n_469), .Y(n_455) );
INVx2_ASAP7_75t_L g531 ( .A(n_456), .Y(n_531) );
AND2x2_ASAP7_75t_L g544 ( .A(n_456), .B(n_482), .Y(n_544) );
AND2x2_ASAP7_75t_L g598 ( .A(n_456), .B(n_481), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_456), .B(n_470), .Y(n_613) );
O2A1O1Ixp33_ASAP7_75t_L g462 ( .A1(n_463), .A2(n_465), .B(n_466), .C(n_467), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_467), .A2(n_488), .B(n_489), .Y(n_487) );
AND2x2_ASAP7_75t_L g631 ( .A(n_469), .B(n_572), .Y(n_631) );
AND2x2_ASAP7_75t_L g664 ( .A(n_469), .B(n_482), .Y(n_664) );
INVx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
OR2x2_ASAP7_75t_L g571 ( .A(n_470), .B(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g584 ( .A(n_470), .B(n_482), .Y(n_584) );
AND2x2_ASAP7_75t_L g591 ( .A(n_470), .B(n_572), .Y(n_591) );
HB1xp67_ASAP7_75t_L g600 ( .A(n_470), .Y(n_600) );
AND2x2_ASAP7_75t_L g607 ( .A(n_470), .B(n_481), .Y(n_607) );
INVx1_ASAP7_75t_L g638 ( .A(n_470), .Y(n_638) );
OAI21xp5_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_475), .B(n_478), .Y(n_471) );
INVx1_ASAP7_75t_L g614 ( .A(n_480), .Y(n_614) );
AND2x2_ASAP7_75t_L g480 ( .A(n_481), .B(n_491), .Y(n_480) );
INVx2_ASAP7_75t_L g570 ( .A(n_481), .Y(n_570) );
AND2x2_ASAP7_75t_L g592 ( .A(n_481), .B(n_531), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_481), .B(n_638), .Y(n_643) );
INVx3_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_482), .B(n_531), .Y(n_530) );
AND2x2_ASAP7_75t_L g715 ( .A(n_482), .B(n_679), .Y(n_715) );
INVx2_ASAP7_75t_L g529 ( .A(n_491), .Y(n_529) );
INVx3_ASAP7_75t_L g630 ( .A(n_491), .Y(n_630) );
OR2x2_ASAP7_75t_L g660 ( .A(n_491), .B(n_661), .Y(n_660) );
NOR2x1_ASAP7_75t_L g686 ( .A(n_491), .B(n_570), .Y(n_686) );
AND2x4_ASAP7_75t_L g491 ( .A(n_492), .B(n_493), .Y(n_491) );
INVx1_ASAP7_75t_L g573 ( .A(n_492), .Y(n_573) );
AOI33xp33_ASAP7_75t_L g706 ( .A1(n_497), .A2(n_544), .A3(n_558), .B1(n_630), .B2(n_707), .B3(n_708), .Y(n_706) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
OR2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_506), .Y(n_498) );
OR2x2_ASAP7_75t_L g559 ( .A(n_499), .B(n_560), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g618 ( .A(n_499), .B(n_556), .Y(n_618) );
OR2x2_ASAP7_75t_L g671 ( .A(n_499), .B(n_672), .Y(n_671) );
INVx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
AND2x2_ASAP7_75t_L g597 ( .A(n_500), .B(n_598), .Y(n_597) );
OR2x2_ASAP7_75t_L g622 ( .A(n_500), .B(n_506), .Y(n_622) );
AND2x2_ASAP7_75t_L g689 ( .A(n_500), .B(n_534), .Y(n_689) );
AOI21xp5_ASAP7_75t_L g714 ( .A1(n_500), .A2(n_589), .B(n_715), .Y(n_714) );
BUFx6f_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g536 ( .A(n_501), .Y(n_536) );
INVx1_ASAP7_75t_L g549 ( .A(n_501), .Y(n_549) );
AND2x2_ASAP7_75t_L g568 ( .A(n_501), .B(n_538), .Y(n_568) );
AND2x2_ASAP7_75t_L g617 ( .A(n_501), .B(n_537), .Y(n_617) );
INVx2_ASAP7_75t_SL g659 ( .A(n_506), .Y(n_659) );
OR2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_517), .Y(n_506) );
INVx2_ASAP7_75t_L g579 ( .A(n_507), .Y(n_579) );
INVx1_ASAP7_75t_L g710 ( .A(n_507), .Y(n_710) );
AND2x2_ASAP7_75t_L g723 ( .A(n_507), .B(n_604), .Y(n_723) );
INVx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx2_ASAP7_75t_L g550 ( .A(n_508), .Y(n_550) );
OR2x2_ASAP7_75t_L g556 ( .A(n_508), .B(n_557), .Y(n_556) );
HB1xp67_ASAP7_75t_L g567 ( .A(n_508), .Y(n_567) );
HB1xp67_ASAP7_75t_L g534 ( .A(n_517), .Y(n_534) );
AND2x2_ASAP7_75t_L g551 ( .A(n_517), .B(n_537), .Y(n_551) );
INVx1_ASAP7_75t_L g557 ( .A(n_517), .Y(n_557) );
INVx1_ASAP7_75t_L g564 ( .A(n_517), .Y(n_564) );
AND2x2_ASAP7_75t_L g589 ( .A(n_517), .B(n_538), .Y(n_589) );
INVx2_ASAP7_75t_L g605 ( .A(n_517), .Y(n_605) );
AND2x2_ASAP7_75t_L g698 ( .A(n_517), .B(n_699), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_517), .B(n_579), .Y(n_719) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_520), .A2(n_521), .B(n_522), .Y(n_519) );
INVx1_ASAP7_75t_SL g527 ( .A(n_528), .Y(n_527) );
OR2x2_ASAP7_75t_L g528 ( .A(n_529), .B(n_530), .Y(n_528) );
INVx2_ASAP7_75t_L g553 ( .A(n_529), .Y(n_553) );
INVx1_ASAP7_75t_L g582 ( .A(n_529), .Y(n_582) );
NOR2xp33_ASAP7_75t_L g679 ( .A(n_529), .B(n_613), .Y(n_679) );
INVx1_ASAP7_75t_SL g639 ( .A(n_530), .Y(n_639) );
INVx2_ASAP7_75t_L g560 ( .A(n_531), .Y(n_560) );
AND2x2_ASAP7_75t_L g629 ( .A(n_531), .B(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g645 ( .A(n_531), .B(n_646), .Y(n_645) );
AND2x2_ASAP7_75t_L g532 ( .A(n_533), .B(n_535), .Y(n_532) );
INVx1_ASAP7_75t_L g707 ( .A(n_533), .Y(n_707) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
AND2x2_ASAP7_75t_L g562 ( .A(n_535), .B(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g665 ( .A(n_535), .B(n_655), .Y(n_665) );
AOI21xp5_ASAP7_75t_L g717 ( .A1(n_535), .A2(n_676), .B(n_718), .Y(n_717) );
AND2x2_ASAP7_75t_L g535 ( .A(n_536), .B(n_537), .Y(n_535) );
AND2x2_ASAP7_75t_L g578 ( .A(n_536), .B(n_579), .Y(n_578) );
BUFx2_ASAP7_75t_L g603 ( .A(n_536), .Y(n_603) );
INVx1_ASAP7_75t_L g627 ( .A(n_536), .Y(n_627) );
OR2x2_ASAP7_75t_L g691 ( .A(n_537), .B(n_550), .Y(n_691) );
NOR2xp67_ASAP7_75t_L g699 ( .A(n_537), .B(n_700), .Y(n_699) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
AND2x2_ASAP7_75t_L g604 ( .A(n_538), .B(n_605), .Y(n_604) );
BUFx2_ASAP7_75t_L g611 ( .A(n_538), .Y(n_611) );
OAI22xp5_ASAP7_75t_L g542 ( .A1(n_543), .A2(n_545), .B1(n_552), .B2(n_554), .Y(n_542) );
OR2x2_ASAP7_75t_L g621 ( .A(n_543), .B(n_571), .Y(n_621) );
INVx1_ASAP7_75t_SL g543 ( .A(n_544), .Y(n_543) );
AOI222xp33_ASAP7_75t_L g662 ( .A1(n_544), .A2(n_663), .B1(n_665), .B2(n_666), .C1(n_667), .C2(n_670), .Y(n_662) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_547), .B(n_551), .Y(n_546) );
INVx1_ASAP7_75t_SL g547 ( .A(n_548), .Y(n_547) );
OR2x2_ASAP7_75t_L g609 ( .A(n_548), .B(n_610), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_549), .B(n_550), .Y(n_548) );
AND2x2_ASAP7_75t_SL g563 ( .A(n_550), .B(n_564), .Y(n_563) );
HB1xp67_ASAP7_75t_L g634 ( .A(n_550), .Y(n_634) );
AND2x2_ASAP7_75t_L g682 ( .A(n_550), .B(n_551), .Y(n_682) );
INVx1_ASAP7_75t_L g700 ( .A(n_550), .Y(n_700) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g666 ( .A(n_553), .B(n_592), .Y(n_666) );
AND2x2_ASAP7_75t_L g708 ( .A(n_553), .B(n_584), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_555), .B(n_558), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_555), .B(n_603), .Y(n_690) );
INVx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
NAND2xp5_ASAP7_75t_SL g587 ( .A(n_556), .B(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g583 ( .A(n_560), .B(n_584), .Y(n_583) );
INVx3_ASAP7_75t_L g651 ( .A(n_560), .Y(n_651) );
O2A1O1Ixp33_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_565), .B(n_569), .C(n_574), .Y(n_561) );
INVxp67_ASAP7_75t_L g575 ( .A(n_562), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_563), .B(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_563), .B(n_610), .Y(n_705) );
BUFx3_ASAP7_75t_L g669 ( .A(n_564), .Y(n_669) );
INVx1_ASAP7_75t_L g576 ( .A(n_565), .Y(n_576) );
AND2x2_ASAP7_75t_L g565 ( .A(n_566), .B(n_568), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g595 ( .A(n_567), .B(n_589), .Y(n_595) );
INVx1_ASAP7_75t_SL g635 ( .A(n_568), .Y(n_635) );
NOR2xp33_ASAP7_75t_L g569 ( .A(n_570), .B(n_571), .Y(n_569) );
INVx1_ASAP7_75t_L g625 ( .A(n_570), .Y(n_625) );
AND2x2_ASAP7_75t_L g648 ( .A(n_570), .B(n_631), .Y(n_648) );
INVx1_ASAP7_75t_SL g619 ( .A(n_571), .Y(n_619) );
INVx1_ASAP7_75t_L g646 ( .A(n_572), .Y(n_646) );
AOI31xp33_ASAP7_75t_L g574 ( .A1(n_575), .A2(n_576), .A3(n_577), .B(n_580), .Y(n_574) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g667 ( .A(n_578), .B(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g641 ( .A(n_579), .Y(n_641) );
BUFx2_ASAP7_75t_L g655 ( .A(n_579), .Y(n_655) );
AND2x2_ASAP7_75t_L g683 ( .A(n_579), .B(n_604), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_581), .B(n_583), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx1_ASAP7_75t_SL g656 ( .A(n_583), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_584), .B(n_651), .Y(n_697) );
AND2x2_ASAP7_75t_L g704 ( .A(n_584), .B(n_630), .Y(n_704) );
AOI211xp5_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_590), .B(n_593), .C(n_608), .Y(n_585) );
INVxp67_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
AOI221xp5_ASAP7_75t_L g616 ( .A1(n_590), .A2(n_617), .B1(n_618), .B2(n_619), .C(n_620), .Y(n_616) );
AND2x2_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
AND2x2_ASAP7_75t_L g624 ( .A(n_591), .B(n_625), .Y(n_624) );
INVx2_ASAP7_75t_L g661 ( .A(n_592), .Y(n_661) );
OAI32xp33_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_596), .A3(n_599), .B1(n_601), .B2(n_606), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
O2A1O1Ixp33_ASAP7_75t_L g647 ( .A1(n_595), .A2(n_648), .B(n_649), .C(n_652), .Y(n_647) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g602 ( .A(n_603), .B(n_604), .Y(n_602) );
OAI21xp5_ASAP7_75t_SL g711 ( .A1(n_603), .A2(n_712), .B(n_713), .Y(n_711) );
INVx1_ASAP7_75t_L g672 ( .A(n_604), .Y(n_672) );
INVxp67_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
NOR2xp33_ASAP7_75t_L g608 ( .A(n_609), .B(n_612), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_610), .B(n_641), .Y(n_640) );
AND2x2_ASAP7_75t_L g658 ( .A(n_610), .B(n_659), .Y(n_658) );
INVx2_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g675 ( .A(n_612), .Y(n_675) );
OR2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
NAND4xp25_ASAP7_75t_SL g615 ( .A(n_616), .B(n_628), .C(n_647), .D(n_662), .Y(n_615) );
AND2x2_ASAP7_75t_L g654 ( .A(n_617), .B(n_655), .Y(n_654) );
AND2x4_ASAP7_75t_L g676 ( .A(n_617), .B(n_669), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_619), .B(n_651), .Y(n_650) );
OAI22xp5_ASAP7_75t_L g620 ( .A1(n_621), .A2(n_622), .B1(n_623), .B2(n_626), .Y(n_620) );
OAI22xp5_ASAP7_75t_L g702 ( .A1(n_621), .A2(n_672), .B1(n_703), .B2(n_705), .Y(n_702) );
O2A1O1Ixp33_ASAP7_75t_L g709 ( .A1(n_621), .A2(n_710), .B(n_711), .C(n_714), .Y(n_709) );
INVx2_ASAP7_75t_L g680 ( .A(n_622), .Y(n_680) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
AOI222xp33_ASAP7_75t_L g674 ( .A1(n_624), .A2(n_658), .B1(n_675), .B2(n_676), .C1(n_677), .C2(n_680), .Y(n_674) );
O2A1O1Ixp33_ASAP7_75t_L g628 ( .A1(n_629), .A2(n_631), .B(n_632), .C(n_636), .Y(n_628) );
INVx1_ASAP7_75t_L g694 ( .A(n_629), .Y(n_694) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
OAI22xp33_ASAP7_75t_L g636 ( .A1(n_633), .A2(n_637), .B1(n_640), .B2(n_642), .Y(n_636) );
OR2x2_ASAP7_75t_L g633 ( .A(n_634), .B(n_635), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_638), .B(n_639), .Y(n_637) );
OR2x2_ASAP7_75t_L g642 ( .A(n_643), .B(n_644), .Y(n_642) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
AND2x2_ASAP7_75t_L g663 ( .A(n_645), .B(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g721 ( .A(n_648), .Y(n_721) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
OAI22xp33_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_656), .B1(n_657), .B2(n_660), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_655), .B(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g712 ( .A(n_660), .Y(n_712) );
INVx1_ASAP7_75t_L g693 ( .A(n_664), .Y(n_693) );
CKINVDCx16_ASAP7_75t_R g720 ( .A(n_666), .Y(n_720) );
INVxp67_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
NAND5xp2_ASAP7_75t_L g673 ( .A(n_674), .B(n_681), .C(n_695), .D(n_701), .E(n_706), .Y(n_673) );
INVx1_ASAP7_75t_SL g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
O2A1O1Ixp33_ASAP7_75t_L g681 ( .A1(n_682), .A2(n_683), .B(n_684), .C(n_687), .Y(n_681) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
AOI31xp33_ASAP7_75t_L g687 ( .A1(n_688), .A2(n_690), .A3(n_691), .B(n_692), .Y(n_687) );
INVx1_ASAP7_75t_L g713 ( .A(n_689), .Y(n_713) );
OR2x2_ASAP7_75t_L g692 ( .A(n_693), .B(n_694), .Y(n_692) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
OAI222xp33_ASAP7_75t_L g716 ( .A1(n_703), .A2(n_705), .B1(n_717), .B2(n_720), .C1(n_721), .C2(n_722), .Y(n_716) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx2_ASAP7_75t_SL g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx2_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx2_ASAP7_75t_SL g731 ( .A(n_732), .Y(n_731) );
CKINVDCx20_ASAP7_75t_R g735 ( .A(n_736), .Y(n_735) );
CKINVDCx14_ASAP7_75t_R g741 ( .A(n_737), .Y(n_741) );
INVx1_ASAP7_75t_SL g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_SL g745 ( .A(n_746), .Y(n_745) );
endmodule