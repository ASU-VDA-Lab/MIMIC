module real_jpeg_6161_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_393;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_14;
wire n_205;
wire n_361;
wire n_261;
wire n_324;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_1),
.A2(n_68),
.B1(n_69),
.B2(n_73),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_1),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_1),
.A2(n_68),
.B1(n_138),
.B2(n_141),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_1),
.A2(n_68),
.B1(n_163),
.B2(n_166),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_1),
.A2(n_68),
.B1(n_180),
.B2(n_194),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_2),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_3),
.A2(n_38),
.B1(n_42),
.B2(n_43),
.Y(n_37)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_3),
.A2(n_42),
.B1(n_108),
.B2(n_111),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_3),
.A2(n_42),
.B1(n_235),
.B2(n_238),
.Y(n_234)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_4),
.Y(n_120)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_5),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_5),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_6),
.Y(n_85)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_6),
.Y(n_96)
);

BUFx5_ASAP7_75t_L g226 ( 
.A(n_6),
.Y(n_226)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_7),
.Y(n_93)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_8),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_8),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_8),
.Y(n_100)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_8),
.Y(n_103)
);

BUFx5_ASAP7_75t_L g180 ( 
.A(n_8),
.Y(n_180)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_8),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_8),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_9),
.Y(n_54)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_9),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_9),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_10),
.A2(n_30),
.B1(n_33),
.B2(n_34),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_10),
.A2(n_33),
.B1(n_123),
.B2(n_147),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_10),
.A2(n_33),
.B1(n_173),
.B2(n_174),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_10),
.B(n_90),
.Y(n_249)
);

O2A1O1Ixp33_ASAP7_75t_L g308 ( 
.A1(n_10),
.A2(n_309),
.B(n_311),
.C(n_319),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_10),
.B(n_335),
.C(n_337),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_10),
.B(n_115),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_10),
.B(n_244),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_10),
.B(n_61),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_11),
.A2(n_180),
.B1(n_181),
.B2(n_182),
.Y(n_179)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_11),
.Y(n_181)
);

OAI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_11),
.A2(n_138),
.B1(n_141),
.B2(n_181),
.Y(n_217)
);

OAI22xp33_ASAP7_75t_SL g325 ( 
.A1(n_11),
.A2(n_148),
.B1(n_181),
.B2(n_315),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_L g344 ( 
.A1(n_11),
.A2(n_181),
.B1(n_345),
.B2(n_349),
.Y(n_344)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);

OAI22xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_205),
.B1(n_401),
.B2(n_402),
.Y(n_13)
);

CKINVDCx14_ASAP7_75t_R g401 ( 
.A(n_14),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_203),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_186),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_16),
.B(n_186),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_104),
.C(n_153),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_17),
.A2(n_104),
.B1(n_105),
.B2(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_17),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_19),
.B1(n_74),
.B2(n_75),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_18),
.A2(n_76),
.B(n_78),
.Y(n_202)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_36),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_20),
.A2(n_76),
.B1(n_77),
.B2(n_78),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_20),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_20),
.A2(n_36),
.B1(n_76),
.B2(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_20),
.B(n_308),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_20),
.A2(n_76),
.B1(n_308),
.B2(n_384),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_27),
.B(n_29),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_21),
.B(n_162),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_21),
.B(n_29),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_21),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_21),
.B(n_344),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_24),
.Y(n_21)
);

INVx3_ASAP7_75t_L g367 ( 
.A(n_22),
.Y(n_367)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_23),
.Y(n_348)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_27),
.Y(n_158)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_29),
.Y(n_159)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_32),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_32),
.Y(n_166)
);

BUFx5_ASAP7_75t_L g337 ( 
.A(n_32),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_33),
.A2(n_100),
.B(n_101),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_33),
.B(n_102),
.Y(n_101)
);

OAI21xp33_ASAP7_75t_L g311 ( 
.A1(n_33),
.A2(n_312),
.B(n_315),
.Y(n_311)
);

AO22x1_ASAP7_75t_SL g61 ( 
.A1(n_34),
.A2(n_54),
.B1(n_62),
.B2(n_64),
.Y(n_61)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_36),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_48),
.B(n_66),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_37),
.A2(n_149),
.B(n_151),
.Y(n_167)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_39),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_40),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_41),
.Y(n_318)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_47),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_47),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_48),
.A2(n_145),
.B(n_149),
.Y(n_198)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_49),
.B(n_67),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_49),
.B(n_146),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_49),
.B(n_325),
.Y(n_324)
);

NOR2x1_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_61),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_53),
.B1(n_55),
.B2(n_58),
.Y(n_50)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g336 ( 
.A(n_57),
.Y(n_336)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_61),
.B(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_61),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_61),
.B(n_325),
.Y(n_339)
);

INVx4_ASAP7_75t_L g349 ( 
.A(n_62),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_63),
.Y(n_237)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_63),
.Y(n_241)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

AND2x2_ASAP7_75t_SL g260 ( 
.A(n_66),
.B(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_66),
.B(n_324),
.Y(n_351)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx6_ASAP7_75t_L g333 ( 
.A(n_72),
.Y(n_333)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_97),
.B(n_98),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_80),
.B(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_80),
.B(n_99),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_80),
.B(n_193),
.Y(n_280)
);

NOR2x1_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_90),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_84),
.B1(n_86),
.B2(n_88),
.Y(n_81)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_85),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_85),
.Y(n_91)
);

NAND2xp33_ASAP7_75t_SL g231 ( 
.A(n_86),
.B(n_232),
.Y(n_231)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_90),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_90),
.B(n_99),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_90),
.B(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_90),
.B(n_179),
.Y(n_212)
);

AO22x1_ASAP7_75t_SL g90 ( 
.A1(n_91),
.A2(n_92),
.B1(n_94),
.B2(n_96),
.Y(n_90)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_92),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_93),
.Y(n_95)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_93),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_93),
.Y(n_140)
);

BUFx5_ASAP7_75t_L g142 ( 
.A(n_93),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_95),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_95),
.Y(n_133)
);

BUFx5_ASAP7_75t_L g224 ( 
.A(n_95),
.Y(n_224)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVxp33_ASAP7_75t_L g230 ( 
.A(n_101),
.Y(n_230)
);

INVx5_ASAP7_75t_L g194 ( 
.A(n_102),
.Y(n_194)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_143),
.B(n_152),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_106),
.B(n_143),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_115),
.B(n_127),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_107),
.A2(n_171),
.B(n_200),
.Y(n_199)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_112),
.A2(n_130),
.B1(n_132),
.B2(n_134),
.Y(n_129)
);

INVx4_ASAP7_75t_SL g112 ( 
.A(n_113),
.Y(n_112)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_115),
.B(n_137),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_115),
.B(n_217),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_115),
.A2(n_171),
.B(n_172),
.Y(n_278)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_116),
.B(n_129),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_116),
.B(n_269),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_121),
.B1(n_124),
.B2(n_125),
.Y(n_116)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx4_ASAP7_75t_L g314 ( 
.A(n_119),
.Y(n_314)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_120),
.Y(n_126)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_120),
.Y(n_131)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_120),
.Y(n_135)
);

INVx3_ASAP7_75t_SL g121 ( 
.A(n_122),
.Y(n_121)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_127),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_128),
.B(n_136),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_128),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_131),
.Y(n_310)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_140),
.Y(n_175)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_140),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_142),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_150),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_144),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_145),
.B(n_149),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVxp67_ASAP7_75t_SL g150 ( 
.A(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_151),
.B(n_339),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_152),
.A2(n_188),
.B1(n_189),
.B2(n_201),
.Y(n_187)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_152),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_153),
.B(n_293),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_168),
.C(n_176),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_154),
.A2(n_155),
.B1(n_287),
.B2(n_288),
.Y(n_286)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_167),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_156),
.B(n_167),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_160),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_157),
.B(n_342),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_159),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_160),
.B(n_360),
.Y(n_359)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_161),
.A2(n_234),
.B(n_242),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_162),
.B(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_168),
.B(n_176),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_169),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_169),
.B(n_247),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_170),
.B(n_216),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_171),
.B(n_217),
.Y(n_247)
);

INVxp67_ASAP7_75t_SL g269 ( 
.A(n_172),
.Y(n_269)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_178),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_178),
.B(n_192),
.Y(n_265)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_202),
.Y(n_186)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_191),
.B1(n_196),
.B2(n_197),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_195),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_195),
.B(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_198),
.A2(n_214),
.B1(n_218),
.B2(n_219),
.Y(n_213)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_198),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_198),
.B(n_211),
.C(n_214),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_205),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_393),
.Y(n_205)
);

NAND3xp33_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_283),
.C(n_298),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_270),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_255),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_209),
.B(n_255),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_220),
.C(n_245),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_210),
.B(n_301),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_211),
.B(n_213),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_212),
.B(n_280),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_214),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_220),
.A2(n_221),
.B1(n_245),
.B2(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_233),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_222),
.B(n_233),
.Y(n_263)
);

AOI32xp33_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_225),
.A3(n_227),
.B1(n_230),
.B2(n_231),
.Y(n_222)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx8_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx8_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_234),
.A2(n_252),
.B(n_259),
.Y(n_258)
);

INVx6_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_244),
.Y(n_362)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_245),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_248),
.C(n_250),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_246),
.B(n_305),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_247),
.B(n_267),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_248),
.A2(n_249),
.B1(n_250),
.B2(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_250),
.Y(n_306)
);

OR2x2_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_251),
.B(n_361),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_SL g371 ( 
.A(n_252),
.B(n_343),
.Y(n_371)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_255),
.B(n_271),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_255),
.B(n_271),
.Y(n_397)
);

FAx1_ASAP7_75t_SL g255 ( 
.A(n_256),
.B(n_257),
.CI(n_262),
.CON(n_255),
.SN(n_255)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_260),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_258),
.B(n_260),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_261),
.B(n_339),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_263),
.B(n_265),
.C(n_266),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g395 ( 
.A1(n_270),
.A2(n_396),
.B(n_397),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_272),
.B(n_274),
.C(n_275),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_279),
.C(n_281),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_281),
.B2(n_282),
.Y(n_277)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_278),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_279),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_295),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_284),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_292),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_285),
.B(n_292),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_289),
.C(n_291),
.Y(n_285)
);

FAx1_ASAP7_75t_SL g296 ( 
.A(n_286),
.B(n_289),
.CI(n_291),
.CON(n_296),
.SN(n_296)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_295),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_296),
.B(n_297),
.Y(n_398)
);

BUFx24_ASAP7_75t_SL g404 ( 
.A(n_296),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_326),
.B(n_392),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_300),
.B(n_303),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_300),
.B(n_303),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_307),
.C(n_321),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_304),
.B(n_388),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_307),
.A2(n_321),
.B1(n_322),
.B2(n_389),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_307),
.Y(n_389)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_308),
.Y(n_384)
);

BUFx3_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx4_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx8_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx4_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_327),
.A2(n_386),
.B(n_391),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_328),
.A2(n_376),
.B(n_385),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_329),
.A2(n_355),
.B(n_375),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_340),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_330),
.B(n_340),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_338),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_331),
.A2(n_332),
.B1(n_338),
.B2(n_358),
.Y(n_357)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_332),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_334),
.Y(n_332)
);

INVx4_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_338),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_350),
.Y(n_340)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_341),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_344),
.B(n_362),
.Y(n_361)
);

BUFx2_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_351),
.A2(n_352),
.B1(n_353),
.B2(n_354),
.Y(n_350)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_351),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_352),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_352),
.B(n_353),
.C(n_378),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_SL g355 ( 
.A1(n_356),
.A2(n_363),
.B(n_374),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_SL g356 ( 
.A(n_357),
.B(n_359),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_357),
.B(n_359),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_364),
.A2(n_370),
.B(n_373),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_369),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_368),
.Y(n_365)
);

INVx1_ASAP7_75t_SL g366 ( 
.A(n_367),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_371),
.B(n_372),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_371),
.B(n_372),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_379),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_377),
.B(n_379),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_383),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_382),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_381),
.B(n_382),
.C(n_383),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_387),
.B(n_390),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_387),
.B(n_390),
.Y(n_391)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g393 ( 
.A1(n_394),
.A2(n_395),
.B(n_398),
.C(n_399),
.D(n_400),
.Y(n_393)
);


endmodule