module real_jpeg_4569_n_27 (n_17, n_8, n_0, n_157, n_21, n_2, n_10, n_9, n_12, n_154, n_156, n_152, n_24, n_6, n_159, n_153, n_151, n_23, n_11, n_14, n_160, n_25, n_7, n_22, n_18, n_3, n_5, n_4, n_1, n_26, n_20, n_19, n_158, n_16, n_15, n_13, n_155, n_27);

input n_17;
input n_8;
input n_0;
input n_157;
input n_21;
input n_2;
input n_10;
input n_9;
input n_12;
input n_154;
input n_156;
input n_152;
input n_24;
input n_6;
input n_159;
input n_153;
input n_151;
input n_23;
input n_11;
input n_14;
input n_160;
input n_25;
input n_7;
input n_22;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_26;
input n_20;
input n_19;
input n_158;
input n_16;
input n_15;
input n_13;
input n_155;

output n_27;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_104;
wire n_64;
wire n_47;
wire n_131;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_141;
wire n_139;
wire n_33;
wire n_65;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_147;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_50;
wire n_143;
wire n_69;
wire n_137;
wire n_31;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_30;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

INVx5_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_0),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_0),
.B(n_85),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_0),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_0),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_1),
.B(n_64),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_1),
.B(n_64),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_2),
.B(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_2),
.B(n_100),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_3),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_4),
.B(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_4),
.B(n_114),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_5),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_6),
.B(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_6),
.B(n_137),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_7),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_8),
.B(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_8),
.B(n_84),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_9),
.B(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_9),
.B(n_142),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_11),
.Y(n_115)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_12),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_13),
.Y(n_120)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_14),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_15),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_16),
.B(n_76),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_17),
.B(n_40),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_17),
.B(n_40),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_18),
.B(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_18),
.B(n_123),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_19),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_20),
.B(n_34),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_20),
.B(n_34),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_21),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_21),
.B(n_45),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_22),
.Y(n_129)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_23),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_24),
.B(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_24),
.B(n_51),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_25),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_26),
.B(n_61),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_26),
.B(n_61),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_140),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_SL g28 ( 
.A1(n_29),
.A2(n_136),
.B(n_139),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_SL g30 ( 
.A1(n_31),
.A2(n_116),
.B(n_130),
.Y(n_30)
);

A2O1A1Ixp33_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_56),
.B(n_104),
.C(n_113),
.Y(n_31)
);

NOR4xp25_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_39),
.C(n_44),
.D(n_50),
.Y(n_32)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_33),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_36),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_62),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_36),
.B(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_36),
.B(n_115),
.Y(n_114)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx11_ASAP7_75t_L g125 ( 
.A(n_38),
.Y(n_125)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_39),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_42),
.Y(n_40)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_44),
.A2(n_108),
.B(n_109),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_47),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g102 ( 
.A(n_47),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_47),
.B(n_128),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_47),
.B(n_138),
.Y(n_137)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_77),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_53),
.Y(n_51)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_55),
.B(n_80),
.Y(n_79)
);

OAI21x1_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_99),
.B(n_103),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_91),
.B(n_98),
.Y(n_57)
);

AO221x1_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_66),
.B1(n_88),
.B2(n_89),
.C(n_90),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_63),
.Y(n_59)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

AO21x1_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_73),
.B(n_87),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_68),
.B(n_72),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_72),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_70),
.Y(n_68)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_83),
.B(n_86),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_78),
.B(n_82),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_79),
.B(n_81),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_79),
.B(n_81),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_92),
.B(n_97),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_92),
.B(n_97),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_94),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_94),
.B(n_120),
.Y(n_119)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_102),
.Y(n_100)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

A2O1A1O1Ixp25_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_107),
.B(n_110),
.C(n_111),
.D(n_112),
.Y(n_105)
);

NAND3xp33_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_121),
.C(n_126),
.Y(n_116)
);

A2O1A1O1Ixp25_ASAP7_75t_L g130 ( 
.A1(n_117),
.A2(n_126),
.B(n_131),
.C(n_134),
.D(n_135),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_119),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_118),
.B(n_119),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_122),
.A2(n_132),
.B(n_133),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_125),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_127),
.B(n_129),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_127),
.B(n_129),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_148),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_144),
.Y(n_142)
);

INVx8_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

BUFx12f_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVxp33_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_151),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_152),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_153),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_154),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_155),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_156),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_157),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_158),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_159),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_160),
.Y(n_101)
);


endmodule