module fake_jpeg_25239_n_409 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_409);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_409;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx11_ASAP7_75t_SL g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx8_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx11_ASAP7_75t_SL g26 ( 
.A(n_6),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx11_ASAP7_75t_SL g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_3),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_18),
.B(n_15),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_46),
.B(n_55),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_47),
.B(n_52),
.Y(n_90)
);

BUFx8_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

INVx3_ASAP7_75t_SL g101 ( 
.A(n_48),
.Y(n_101)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_50),
.Y(n_125)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_18),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_20),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_53),
.B(n_63),
.Y(n_92)
);

BUFx4f_ASAP7_75t_SL g54 ( 
.A(n_19),
.Y(n_54)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_54),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_20),
.B(n_15),
.Y(n_55)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_56),
.Y(n_115)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_58),
.Y(n_103)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_59),
.Y(n_104)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_60),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_61),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_62),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_19),
.B(n_15),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_29),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_64),
.B(n_67),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_65),
.Y(n_129)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_66),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_29),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_68),
.Y(n_106)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_69),
.B(n_70),
.Y(n_99)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_32),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_71),
.B(n_72),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_25),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_27),
.Y(n_73)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_73),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_27),
.Y(n_74)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_74),
.Y(n_122)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_75),
.B(n_76),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_32),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_23),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_77),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_17),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_78),
.B(n_80),
.Y(n_120)
);

BUFx16f_ASAP7_75t_L g79 ( 
.A(n_25),
.Y(n_79)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_79),
.Y(n_126)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_38),
.B(n_0),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_81),
.B(n_82),
.Y(n_85)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_16),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_25),
.Y(n_83)
);

AOI21xp33_ASAP7_75t_SL g107 ( 
.A1(n_83),
.A2(n_84),
.B(n_17),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_17),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_81),
.B(n_38),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_86),
.B(n_110),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_69),
.A2(n_34),
.B1(n_41),
.B2(n_44),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_89),
.A2(n_95),
.B1(n_112),
.B2(n_117),
.Y(n_150)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_94),
.B(n_109),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_75),
.A2(n_34),
.B1(n_44),
.B2(n_36),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_80),
.A2(n_34),
.B1(n_43),
.B2(n_16),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_100),
.A2(n_130),
.B1(n_28),
.B2(n_21),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_107),
.A2(n_83),
.B(n_79),
.Y(n_169)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_46),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_82),
.B(n_38),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_45),
.B(n_38),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_111),
.B(n_30),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_66),
.A2(n_43),
.B1(n_22),
.B2(n_36),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_77),
.A2(n_41),
.B1(n_37),
.B2(n_35),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_114),
.A2(n_59),
.B1(n_51),
.B2(n_30),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_57),
.A2(n_22),
.B1(n_21),
.B2(n_33),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_52),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_118),
.B(n_119),
.Y(n_162)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_53),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_58),
.A2(n_60),
.B1(n_49),
.B2(n_70),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_121),
.A2(n_127),
.B1(n_47),
.B2(n_23),
.Y(n_153)
);

OAI22xp33_ASAP7_75t_L g127 ( 
.A1(n_73),
.A2(n_37),
.B1(n_35),
.B2(n_33),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_64),
.A2(n_37),
.B1(n_35),
.B2(n_33),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_108),
.A2(n_76),
.B1(n_71),
.B2(n_67),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_131),
.A2(n_143),
.B1(n_154),
.B2(n_155),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_96),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_132),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_122),
.Y(n_133)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_133),
.Y(n_186)
);

OAI22xp33_ASAP7_75t_L g135 ( 
.A1(n_122),
.A2(n_74),
.B1(n_54),
.B2(n_84),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_135),
.A2(n_101),
.B1(n_87),
.B2(n_104),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_85),
.B(n_93),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_136),
.B(n_160),
.Y(n_182)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_123),
.Y(n_137)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_137),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_113),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_138),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_86),
.B(n_54),
.C(n_50),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_139),
.B(n_142),
.C(n_124),
.Y(n_202)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_99),
.Y(n_140)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_140),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_85),
.B(n_65),
.C(n_61),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_121),
.Y(n_144)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_144),
.Y(n_197)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_111),
.Y(n_145)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_145),
.Y(n_203)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_91),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_146),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_102),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_147),
.B(n_161),
.Y(n_176)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_123),
.Y(n_148)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_148),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_149),
.B(n_152),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_108),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_151),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_110),
.B(n_30),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_153),
.A2(n_158),
.B1(n_168),
.B2(n_129),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_87),
.A2(n_14),
.B1(n_21),
.B2(n_23),
.Y(n_154)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_100),
.Y(n_156)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_156),
.Y(n_205)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_88),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_157),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_92),
.A2(n_130),
.B1(n_127),
.B2(n_88),
.Y(n_158)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_115),
.Y(n_159)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_159),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_90),
.B(n_72),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_120),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_97),
.B(n_68),
.Y(n_163)
);

OR2x2_ASAP7_75t_L g188 ( 
.A(n_163),
.B(n_105),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_115),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_164),
.B(n_166),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_116),
.Y(n_165)
);

NAND3xp33_ASAP7_75t_L g196 ( 
.A(n_165),
.B(n_101),
.C(n_106),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_97),
.B(n_79),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_103),
.Y(n_167)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_167),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_103),
.A2(n_28),
.B1(n_62),
.B2(n_2),
.Y(n_168)
);

MAJx2_ASAP7_75t_L g179 ( 
.A(n_169),
.B(n_125),
.C(n_106),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_98),
.B(n_28),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_170),
.B(n_171),
.Y(n_193)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_98),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_116),
.Y(n_172)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_172),
.Y(n_210)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_105),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_173),
.B(n_174),
.Y(n_194)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_91),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_175),
.A2(n_190),
.B1(n_192),
.B2(n_207),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_179),
.B(n_211),
.C(n_4),
.Y(n_248)
);

FAx1_ASAP7_75t_SL g180 ( 
.A(n_134),
.B(n_104),
.CI(n_128),
.CON(n_180),
.SN(n_180)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_180),
.B(n_188),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_144),
.A2(n_125),
.B1(n_128),
.B2(n_129),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_191),
.A2(n_135),
.B1(n_133),
.B2(n_151),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_156),
.A2(n_155),
.B1(n_145),
.B2(n_142),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_196),
.A2(n_174),
.B1(n_173),
.B2(n_138),
.Y(n_219)
);

INVx5_ASAP7_75t_L g198 ( 
.A(n_146),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_198),
.B(n_199),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_162),
.B(n_126),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_134),
.B(n_124),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_201),
.B(n_202),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_149),
.A2(n_126),
.B1(n_48),
.B2(n_105),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_132),
.B(n_0),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_208),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_139),
.B(n_48),
.C(n_1),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_150),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_212),
.A2(n_161),
.B1(n_172),
.B2(n_167),
.Y(n_232)
);

AO22x1_ASAP7_75t_L g213 ( 
.A1(n_153),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_213)
);

O2A1O1Ixp33_ASAP7_75t_L g245 ( 
.A1(n_213),
.A2(n_4),
.B(n_5),
.C(n_6),
.Y(n_245)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_163),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_214),
.B(n_141),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_183),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_215),
.Y(n_259)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_194),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_216),
.B(n_217),
.Y(n_265)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_190),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_219),
.A2(n_223),
.B(n_233),
.Y(n_250)
);

OR2x2_ASAP7_75t_L g221 ( 
.A(n_188),
.B(n_152),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_221),
.A2(n_6),
.B(n_11),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_183),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_222),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_205),
.A2(n_169),
.B(n_165),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_192),
.A2(n_205),
.B1(n_197),
.B2(n_191),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_225),
.A2(n_230),
.B1(n_232),
.B2(n_234),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_177),
.B(n_147),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_226),
.B(n_227),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_177),
.B(n_160),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_228),
.B(n_229),
.Y(n_274)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_193),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_197),
.A2(n_159),
.B1(n_164),
.B2(n_140),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_207),
.A2(n_214),
.B1(n_181),
.B2(n_203),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_202),
.A2(n_157),
.B1(n_148),
.B2(n_137),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_189),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_235),
.B(n_238),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_201),
.B(n_171),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_236),
.B(n_203),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_237),
.A2(n_246),
.B1(n_178),
.B2(n_186),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_182),
.B(n_3),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_200),
.Y(n_239)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_239),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_185),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_240),
.Y(n_263)
);

CKINVDCx14_ASAP7_75t_R g241 ( 
.A(n_176),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_241),
.B(n_243),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_185),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_242),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_184),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_245),
.A2(n_4),
.B(n_6),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_212),
.A2(n_133),
.B1(n_151),
.B2(n_7),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_180),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_247),
.B(n_249),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_248),
.B(n_179),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_175),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_254),
.B(n_278),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_255),
.B(n_261),
.C(n_248),
.Y(n_281)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_236),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_256),
.B(n_257),
.Y(n_292)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_230),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_258),
.A2(n_266),
.B1(n_271),
.B2(n_273),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_220),
.B(n_211),
.C(n_180),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_243),
.A2(n_198),
.B1(n_178),
.B2(n_186),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_237),
.A2(n_213),
.B1(n_210),
.B2(n_187),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_267),
.A2(n_218),
.B1(n_233),
.B2(n_221),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_231),
.A2(n_187),
.B(n_213),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_268),
.A2(n_269),
.B(n_272),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_231),
.A2(n_210),
.B(n_209),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_L g271 ( 
.A1(n_249),
.A2(n_204),
.B1(n_195),
.B2(n_209),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_247),
.A2(n_204),
.B(n_195),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_239),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_273),
.B(n_244),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_215),
.B(n_200),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_275),
.B(n_222),
.Y(n_300)
);

AO22x1_ASAP7_75t_SL g276 ( 
.A1(n_225),
.A2(n_184),
.B1(n_206),
.B2(n_9),
.Y(n_276)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_276),
.Y(n_282)
);

CKINVDCx14_ASAP7_75t_R g283 ( 
.A(n_277),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_226),
.B(n_206),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_280),
.B(n_245),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_281),
.B(n_289),
.C(n_290),
.Y(n_312)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_275),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_284),
.B(n_291),
.Y(n_320)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_259),
.Y(n_286)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_286),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_287),
.A2(n_294),
.B1(n_295),
.B2(n_301),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_257),
.A2(n_232),
.B1(n_217),
.B2(n_234),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_288),
.A2(n_267),
.B1(n_256),
.B2(n_258),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_255),
.B(n_220),
.C(n_248),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_261),
.B(n_227),
.C(n_223),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_278),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_253),
.A2(n_233),
.B1(n_218),
.B2(n_221),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_264),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_296),
.B(n_299),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_259),
.B(n_240),
.Y(n_297)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_297),
.Y(n_308)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_298),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_300),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_253),
.A2(n_219),
.B1(n_229),
.B2(n_241),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_250),
.A2(n_246),
.B1(n_242),
.B2(n_235),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_302),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_260),
.Y(n_303)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_303),
.Y(n_327)
);

INVx1_ASAP7_75t_SL g304 ( 
.A(n_254),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_304),
.Y(n_309)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_264),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_305),
.Y(n_311)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_265),
.Y(n_306)
);

INVx2_ASAP7_75t_SL g321 ( 
.A(n_306),
.Y(n_321)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_265),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_307),
.B(n_274),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_281),
.B(n_261),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_SL g346 ( 
.A(n_310),
.B(n_318),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_290),
.B(n_250),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_313),
.B(n_315),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_289),
.B(n_285),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_317),
.A2(n_324),
.B1(n_330),
.B2(n_294),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_285),
.B(n_252),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_282),
.A2(n_270),
.B1(n_252),
.B2(n_272),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_301),
.B(n_269),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_326),
.B(n_312),
.C(n_310),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_295),
.A2(n_270),
.B1(n_279),
.B2(n_260),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_328),
.A2(n_288),
.B1(n_305),
.B2(n_296),
.Y(n_339)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_329),
.Y(n_344)
);

AO22x2_ASAP7_75t_L g330 ( 
.A1(n_282),
.A2(n_276),
.B1(n_271),
.B2(n_277),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_319),
.A2(n_283),
.B(n_302),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g360 ( 
.A(n_331),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_319),
.A2(n_287),
.B1(n_306),
.B2(n_307),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_332),
.A2(n_334),
.B1(n_340),
.B2(n_349),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_325),
.B(n_297),
.Y(n_333)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_333),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_308),
.B(n_303),
.Y(n_335)
);

NAND3xp33_ASAP7_75t_L g361 ( 
.A(n_335),
.B(n_338),
.C(n_343),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_320),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_336),
.A2(n_316),
.B1(n_321),
.B2(n_330),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_337),
.B(n_324),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_323),
.B(n_263),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_339),
.B(n_342),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_314),
.A2(n_274),
.B1(n_292),
.B2(n_300),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g342 ( 
.A(n_330),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_311),
.B(n_263),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_312),
.B(n_315),
.C(n_313),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_345),
.B(n_318),
.C(n_326),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_327),
.B(n_279),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_347),
.A2(n_348),
.B1(n_321),
.B2(n_298),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_309),
.B(n_286),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_322),
.B(n_293),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_350),
.B(n_352),
.C(n_354),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_337),
.B(n_291),
.C(n_328),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_334),
.A2(n_314),
.B1(n_330),
.B2(n_292),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_356),
.A2(n_276),
.B1(n_245),
.B2(n_251),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_345),
.B(n_293),
.C(n_284),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_357),
.B(n_358),
.C(n_346),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_341),
.B(n_317),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_SL g372 ( 
.A1(n_359),
.A2(n_299),
.B(n_251),
.Y(n_372)
);

FAx1_ASAP7_75t_SL g362 ( 
.A(n_349),
.B(n_262),
.CI(n_304),
.CON(n_362),
.SN(n_362)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_362),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_SL g363 ( 
.A(n_341),
.B(n_346),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_363),
.A2(n_224),
.B1(n_280),
.B2(n_228),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_364),
.B(n_344),
.Y(n_366)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_366),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_367),
.B(n_375),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_352),
.B(n_333),
.C(n_332),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_368),
.B(n_354),
.C(n_350),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_355),
.B(n_262),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_369),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_351),
.A2(n_333),
.B1(n_336),
.B2(n_331),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_370),
.A2(n_374),
.B1(n_355),
.B2(n_362),
.Y(n_380)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_372),
.Y(n_379)
);

OAI21xp33_ASAP7_75t_L g373 ( 
.A1(n_353),
.A2(n_268),
.B(n_216),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_373),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_SL g376 ( 
.A(n_357),
.B(n_238),
.Y(n_376)
);

FAx1_ASAP7_75t_SL g387 ( 
.A(n_376),
.B(n_363),
.CI(n_276),
.CON(n_387),
.SN(n_387)
);

OAI21xp5_ASAP7_75t_SL g377 ( 
.A1(n_371),
.A2(n_359),
.B(n_360),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_SL g393 ( 
.A1(n_377),
.A2(n_386),
.B(n_11),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_380),
.A2(n_373),
.B1(n_375),
.B2(n_266),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_365),
.B(n_358),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_383),
.B(n_387),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_385),
.B(n_365),
.C(n_368),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_SL g386 ( 
.A1(n_370),
.A2(n_361),
.B(n_244),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_388),
.B(n_390),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_378),
.B(n_367),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_391),
.A2(n_393),
.B1(n_387),
.B2(n_385),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_380),
.B(n_384),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_392),
.B(n_394),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_386),
.B(n_11),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_379),
.A2(n_12),
.B1(n_13),
.B2(n_382),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_395),
.Y(n_397)
);

A2O1A1O1Ixp25_ASAP7_75t_L g396 ( 
.A1(n_393),
.A2(n_377),
.B(n_387),
.C(n_381),
.D(n_379),
.Y(n_396)
);

NOR4xp25_ASAP7_75t_L g403 ( 
.A(n_396),
.B(n_389),
.C(n_383),
.D(n_13),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_400),
.B(n_381),
.Y(n_402)
);

NOR2xp67_ASAP7_75t_L g401 ( 
.A(n_398),
.B(n_388),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_401),
.B(n_402),
.C(n_403),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_402),
.B(n_399),
.C(n_397),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_405),
.B(n_12),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_406),
.B(n_404),
.Y(n_407)
);

BUFx24_ASAP7_75t_SL g408 ( 
.A(n_407),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_408),
.B(n_12),
.Y(n_409)
);


endmodule