module real_aes_17201_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_857, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_857;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_841;
wire n_318;
wire n_718;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_537;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_693;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_527;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_552;
wire n_402;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_288;
wire n_147;
wire n_150;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_854;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
AND2x4_ASAP7_75t_L g852 ( .A(n_0), .B(n_853), .Y(n_852) );
AOI22xp33_ASAP7_75t_L g183 ( .A1(n_1), .A2(n_34), .B1(n_148), .B2(n_184), .Y(n_183) );
AOI22xp5_ASAP7_75t_L g214 ( .A1(n_2), .A2(n_10), .B1(n_138), .B2(n_215), .Y(n_214) );
INVx1_ASAP7_75t_L g853 ( .A(n_3), .Y(n_853) );
AOI22xp5_ASAP7_75t_L g104 ( .A1(n_4), .A2(n_105), .B1(n_848), .B2(n_854), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g168 ( .A(n_5), .Y(n_168) );
AOI22xp5_ASAP7_75t_L g196 ( .A1(n_6), .A2(n_11), .B1(n_197), .B2(n_200), .Y(n_196) );
OR2x2_ASAP7_75t_L g114 ( .A(n_7), .B(n_30), .Y(n_114) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_8), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g219 ( .A(n_9), .Y(n_219) );
NAND2xp5_ASAP7_75t_SL g500 ( .A(n_12), .B(n_139), .Y(n_500) );
AOI22xp5_ASAP7_75t_L g137 ( .A1(n_13), .A2(n_101), .B1(n_138), .B2(n_141), .Y(n_137) );
AOI22xp33_ASAP7_75t_L g211 ( .A1(n_14), .A2(n_31), .B1(n_173), .B2(n_212), .Y(n_211) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_15), .B(n_139), .Y(n_170) );
OAI21x1_ASAP7_75t_L g156 ( .A1(n_16), .A2(n_45), .B(n_157), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_17), .B(n_542), .Y(n_541) );
CKINVDCx5p33_ASAP7_75t_R g159 ( .A(n_18), .Y(n_159) );
AOI22xp5_ASAP7_75t_L g826 ( .A1(n_19), .A2(n_89), .B1(n_806), .B2(n_827), .Y(n_826) );
INVx1_ASAP7_75t_L g827 ( .A(n_19), .Y(n_827) );
AOI22xp33_ASAP7_75t_L g185 ( .A1(n_20), .A2(n_38), .B1(n_186), .B2(n_187), .Y(n_185) );
CKINVDCx5p33_ASAP7_75t_R g479 ( .A(n_21), .Y(n_479) );
XOR2x2_ASAP7_75t_L g116 ( .A(n_22), .B(n_117), .Y(n_116) );
AOI22xp33_ASAP7_75t_L g266 ( .A1(n_23), .A2(n_43), .B1(n_138), .B2(n_187), .Y(n_266) );
CKINVDCx5p33_ASAP7_75t_R g232 ( .A(n_24), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_25), .B(n_173), .Y(n_172) );
CKINVDCx5p33_ASAP7_75t_R g249 ( .A(n_26), .Y(n_249) );
NAND2xp5_ASAP7_75t_SL g540 ( .A(n_27), .B(n_198), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_28), .B(n_179), .Y(n_490) );
CKINVDCx5p33_ASAP7_75t_R g562 ( .A(n_29), .Y(n_562) );
AOI22xp5_ASAP7_75t_L g224 ( .A1(n_32), .A2(n_83), .B1(n_148), .B2(n_225), .Y(n_224) );
AOI22xp33_ASAP7_75t_L g201 ( .A1(n_33), .A2(n_37), .B1(n_148), .B2(n_169), .Y(n_201) );
AOI22xp33_ASAP7_75t_L g146 ( .A1(n_35), .A2(n_48), .B1(n_138), .B2(n_147), .Y(n_146) );
CKINVDCx5p33_ASAP7_75t_R g484 ( .A(n_36), .Y(n_484) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_39), .B(n_139), .Y(n_527) );
INVx2_ASAP7_75t_L g109 ( .A(n_40), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_41), .B(n_144), .Y(n_537) );
BUFx3_ASAP7_75t_L g112 ( .A(n_42), .Y(n_112) );
INVx1_ASAP7_75t_L g823 ( .A(n_42), .Y(n_823) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_44), .B(n_487), .Y(n_544) );
AND2x2_ASAP7_75t_L g486 ( .A(n_46), .B(n_487), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_47), .B(n_213), .Y(n_591) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_49), .B(n_198), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_50), .B(n_186), .Y(n_566) );
AOI22xp5_ASAP7_75t_L g117 ( .A1(n_51), .A2(n_90), .B1(n_118), .B2(n_119), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_51), .Y(n_119) );
AOI22xp33_ASAP7_75t_L g839 ( .A1(n_52), .A2(n_835), .B1(n_840), .B2(n_841), .Y(n_839) );
AOI22xp33_ASAP7_75t_L g265 ( .A1(n_53), .A2(n_71), .B1(n_147), .B2(n_186), .Y(n_265) );
AOI22xp33_ASAP7_75t_L g247 ( .A1(n_54), .A2(n_74), .B1(n_148), .B2(n_169), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_55), .B(n_513), .Y(n_512) );
A2O1A1Ixp33_ASAP7_75t_L g477 ( .A1(n_56), .A2(n_228), .B(n_478), .C(n_480), .Y(n_477) );
AOI22xp5_ASAP7_75t_L g246 ( .A1(n_57), .A2(n_98), .B1(n_138), .B2(n_200), .Y(n_246) );
AND2x4_ASAP7_75t_L g134 ( .A(n_58), .B(n_135), .Y(n_134) );
INVx1_ASAP7_75t_L g157 ( .A(n_59), .Y(n_157) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_60), .A2(n_61), .B1(n_187), .B2(n_216), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_62), .B(n_179), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_63), .B(n_487), .Y(n_593) );
CKINVDCx5p33_ASAP7_75t_R g485 ( .A(n_64), .Y(n_485) );
NAND2xp5_ASAP7_75t_SL g530 ( .A(n_65), .B(n_187), .Y(n_530) );
INVx1_ASAP7_75t_L g135 ( .A(n_66), .Y(n_135) );
INVx1_ASAP7_75t_L g817 ( .A(n_67), .Y(n_817) );
OAI22xp5_ASAP7_75t_L g825 ( .A1(n_68), .A2(n_826), .B1(n_828), .B2(n_829), .Y(n_825) );
CKINVDCx14_ASAP7_75t_R g828 ( .A(n_68), .Y(n_828) );
CKINVDCx5p33_ASAP7_75t_R g552 ( .A(n_69), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_70), .B(n_179), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_72), .B(n_148), .Y(n_508) );
NAND3xp33_ASAP7_75t_L g538 ( .A(n_73), .B(n_144), .C(n_184), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_75), .B(n_148), .Y(n_493) );
INVx2_ASAP7_75t_L g145 ( .A(n_76), .Y(n_145) );
NAND2xp5_ASAP7_75t_SL g565 ( .A(n_77), .B(n_139), .Y(n_565) );
NAND2xp5_ASAP7_75t_SL g588 ( .A(n_78), .B(n_203), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_79), .B(n_497), .Y(n_496) );
AOI22xp33_ASAP7_75t_L g227 ( .A1(n_80), .A2(n_97), .B1(n_187), .B2(n_228), .Y(n_227) );
CKINVDCx5p33_ASAP7_75t_R g268 ( .A(n_81), .Y(n_268) );
CKINVDCx5p33_ASAP7_75t_R g190 ( .A(n_82), .Y(n_190) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_84), .A2(n_92), .B1(n_198), .B2(n_549), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_85), .B(n_139), .Y(n_563) );
NAND2xp33_ASAP7_75t_SL g592 ( .A(n_86), .B(n_174), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_87), .B(n_142), .Y(n_526) );
CKINVDCx5p33_ASAP7_75t_R g836 ( .A(n_88), .Y(n_836) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_89), .B(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g806 ( .A(n_89), .Y(n_806) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_90), .Y(n_118) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_91), .B(n_179), .Y(n_178) );
CKINVDCx5p33_ASAP7_75t_R g207 ( .A(n_93), .Y(n_207) );
INVx1_ASAP7_75t_L g463 ( .A(n_94), .Y(n_463) );
NOR2xp33_ASAP7_75t_L g821 ( .A(n_94), .B(n_822), .Y(n_821) );
NAND2xp33_ASAP7_75t_L g175 ( .A(n_95), .B(n_139), .Y(n_175) );
NAND2xp33_ASAP7_75t_L g494 ( .A(n_96), .B(n_174), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_99), .B(n_487), .Y(n_515) );
NAND3xp33_ASAP7_75t_L g589 ( .A(n_100), .B(n_174), .C(n_203), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_102), .B(n_148), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g511 ( .A(n_103), .B(n_198), .Y(n_511) );
AO21x2_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_115), .B(n_810), .Y(n_105) );
BUFx6f_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
AND2x6_ASAP7_75t_SL g107 ( .A(n_108), .B(n_110), .Y(n_107) );
BUFx3_ASAP7_75t_L g840 ( .A(n_108), .Y(n_840) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx3_ASAP7_75t_L g815 ( .A(n_109), .Y(n_815) );
NOR2xp33_ASAP7_75t_L g844 ( .A(n_109), .B(n_845), .Y(n_844) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_111), .B(n_113), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
NOR2x1_ASAP7_75t_L g847 ( .A(n_112), .B(n_114), .Y(n_847) );
AND2x6_ASAP7_75t_SL g820 ( .A(n_113), .B(n_821), .Y(n_820) );
INVx1_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
XNOR2xp5_ASAP7_75t_L g115 ( .A(n_116), .B(n_120), .Y(n_115) );
AND2x2_ASAP7_75t_L g120 ( .A(n_121), .B(n_464), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g121 ( .A(n_122), .B(n_461), .Y(n_121) );
OR2x2_ASAP7_75t_L g122 ( .A(n_123), .B(n_364), .Y(n_122) );
NAND4xp25_ASAP7_75t_L g123 ( .A(n_124), .B(n_288), .C(n_319), .D(n_348), .Y(n_123) );
NOR2xp33_ASAP7_75t_L g124 ( .A(n_125), .B(n_255), .Y(n_124) );
OAI322xp33_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_191), .A3(n_220), .B1(n_233), .B2(n_241), .C1(n_250), .C2(n_252), .Y(n_125) );
INVxp67_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_127), .B(n_445), .Y(n_444) );
AND2x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_161), .Y(n_127) );
AND2x2_ASAP7_75t_L g285 ( .A(n_128), .B(n_286), .Y(n_285) );
INVx4_ASAP7_75t_L g321 ( .A(n_128), .Y(n_321) );
INVx3_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
AND2x2_ASAP7_75t_L g296 ( .A(n_129), .B(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g299 ( .A(n_129), .B(n_193), .Y(n_299) );
AND2x2_ASAP7_75t_L g316 ( .A(n_129), .B(n_209), .Y(n_316) );
AND2x2_ASAP7_75t_L g414 ( .A(n_129), .B(n_415), .Y(n_414) );
INVx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx2_ASAP7_75t_L g237 ( .A(n_130), .Y(n_237) );
AND2x4_ASAP7_75t_L g420 ( .A(n_130), .B(n_415), .Y(n_420) );
AO31x2_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_136), .A3(n_152), .B(n_158), .Y(n_130) );
AO31x2_ASAP7_75t_L g244 ( .A1(n_131), .A2(n_204), .A3(n_245), .B(n_248), .Y(n_244) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
NOR2xp67_ASAP7_75t_SL g475 ( .A(n_132), .B(n_153), .Y(n_475) );
INVx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
AO31x2_ASAP7_75t_L g181 ( .A1(n_133), .A2(n_182), .A3(n_188), .B(n_189), .Y(n_181) );
AO31x2_ASAP7_75t_L g194 ( .A1(n_133), .A2(n_195), .A3(n_204), .B(n_206), .Y(n_194) );
AO31x2_ASAP7_75t_L g209 ( .A1(n_133), .A2(n_210), .A3(n_217), .B(n_218), .Y(n_209) );
AO31x2_ASAP7_75t_L g546 ( .A1(n_133), .A2(n_154), .A3(n_547), .B(n_551), .Y(n_546) );
BUFx10_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g177 ( .A(n_134), .Y(n_177) );
BUFx10_ASAP7_75t_L g502 ( .A(n_134), .Y(n_502) );
OAI22xp5_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_143), .B1(n_146), .B2(n_149), .Y(n_136) );
INVx3_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx1_ASAP7_75t_L g542 ( .A(n_139), .Y(n_542) );
OAI21xp5_ASAP7_75t_L g587 ( .A1(n_139), .A2(n_588), .B(n_589), .Y(n_587) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx1_ASAP7_75t_L g142 ( .A(n_140), .Y(n_142) );
INVx3_ASAP7_75t_L g148 ( .A(n_140), .Y(n_148) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_140), .Y(n_174) );
BUFx6f_ASAP7_75t_L g184 ( .A(n_140), .Y(n_184) );
BUFx6f_ASAP7_75t_L g187 ( .A(n_140), .Y(n_187) );
INVx1_ASAP7_75t_L g199 ( .A(n_140), .Y(n_199) );
INVx1_ASAP7_75t_L g213 ( .A(n_140), .Y(n_213) );
INVx1_ASAP7_75t_L g216 ( .A(n_140), .Y(n_216) );
INVx2_ASAP7_75t_L g226 ( .A(n_140), .Y(n_226) );
INVx1_ASAP7_75t_L g228 ( .A(n_140), .Y(n_228) );
O2A1O1Ixp5_ASAP7_75t_L g561 ( .A1(n_141), .A2(n_144), .B(n_562), .C(n_563), .Y(n_561) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
AOI21xp5_ASAP7_75t_L g171 ( .A1(n_143), .A2(n_172), .B(n_175), .Y(n_171) );
OAI22xp5_ASAP7_75t_L g182 ( .A1(n_143), .A2(n_149), .B1(n_183), .B2(n_185), .Y(n_182) );
OAI22xp5_ASAP7_75t_L g195 ( .A1(n_143), .A2(n_196), .B1(n_201), .B2(n_202), .Y(n_195) );
OAI22xp5_ASAP7_75t_L g210 ( .A1(n_143), .A2(n_149), .B1(n_211), .B2(n_214), .Y(n_210) );
OAI22xp5_ASAP7_75t_L g223 ( .A1(n_143), .A2(n_224), .B1(n_227), .B2(n_229), .Y(n_223) );
OAI22xp5_ASAP7_75t_L g245 ( .A1(n_143), .A2(n_202), .B1(n_246), .B2(n_247), .Y(n_245) );
OAI22xp5_ASAP7_75t_L g264 ( .A1(n_143), .A2(n_149), .B1(n_265), .B2(n_266), .Y(n_264) );
OAI22xp5_ASAP7_75t_L g547 ( .A1(n_143), .A2(n_149), .B1(n_548), .B2(n_550), .Y(n_547) );
INVx6_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
O2A1O1Ixp5_ASAP7_75t_L g167 ( .A1(n_144), .A2(n_168), .B(n_169), .C(n_170), .Y(n_167) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_144), .A2(n_529), .B(n_530), .Y(n_528) );
BUFx8_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g151 ( .A(n_145), .Y(n_151) );
INVx1_ASAP7_75t_L g203 ( .A(n_145), .Y(n_203) );
INVx1_ASAP7_75t_L g481 ( .A(n_145), .Y(n_481) );
INVx1_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx4_ASAP7_75t_L g169 ( .A(n_148), .Y(n_169) );
INVx1_ASAP7_75t_L g200 ( .A(n_148), .Y(n_200) );
OAI22xp33_ASAP7_75t_L g483 ( .A1(n_148), .A2(n_187), .B1(n_484), .B2(n_485), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_149), .B(n_483), .Y(n_482) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx2_ASAP7_75t_L g514 ( .A(n_150), .Y(n_514) );
BUFx3_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g498 ( .A(n_151), .Y(n_498) );
AO31x2_ASAP7_75t_L g263 ( .A1(n_152), .A2(n_230), .A3(n_264), .B(n_267), .Y(n_263) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
NOR2xp33_ASAP7_75t_SL g206 ( .A(n_154), .B(n_207), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_154), .B(n_232), .Y(n_231) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx2_ASAP7_75t_L g160 ( .A(n_155), .Y(n_160) );
INVx2_ASAP7_75t_L g205 ( .A(n_155), .Y(n_205) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_156), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g158 ( .A(n_159), .B(n_160), .Y(n_158) );
NOR2xp33_ASAP7_75t_L g267 ( .A(n_160), .B(n_268), .Y(n_267) );
INVx2_ASAP7_75t_L g487 ( .A(n_160), .Y(n_487) );
INVx2_ASAP7_75t_L g505 ( .A(n_160), .Y(n_505) );
AND2x4_ASAP7_75t_L g425 ( .A(n_161), .B(n_326), .Y(n_425) );
INVx1_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx1_ASAP7_75t_L g254 ( .A(n_162), .Y(n_254) );
INVxp67_ASAP7_75t_SL g412 ( .A(n_162), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_163), .B(n_180), .Y(n_162) );
AND2x2_ASAP7_75t_L g242 ( .A(n_163), .B(n_181), .Y(n_242) );
INVx1_ASAP7_75t_L g283 ( .A(n_163), .Y(n_283) );
OAI21x1_ASAP7_75t_L g163 ( .A1(n_164), .A2(n_166), .B(n_178), .Y(n_163) );
OAI21x1_ASAP7_75t_L g278 ( .A1(n_164), .A2(n_166), .B(n_178), .Y(n_278) );
INVx2_ASAP7_75t_SL g164 ( .A(n_165), .Y(n_164) );
INVx4_ASAP7_75t_L g179 ( .A(n_165), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_165), .B(n_190), .Y(n_189) );
BUFx3_ASAP7_75t_L g217 ( .A(n_165), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_165), .B(n_219), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_165), .B(n_249), .Y(n_248) );
AND2x4_ASAP7_75t_SL g501 ( .A(n_165), .B(n_502), .Y(n_501) );
INVx2_ASAP7_75t_L g523 ( .A(n_165), .Y(n_523) );
INVx1_ASAP7_75t_SL g585 ( .A(n_165), .Y(n_585) );
OAI21x1_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_171), .B(n_176), .Y(n_166) );
INVx1_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx2_ASAP7_75t_L g186 ( .A(n_174), .Y(n_186) );
INVx2_ASAP7_75t_SL g176 ( .A(n_177), .Y(n_176) );
INVx2_ASAP7_75t_SL g230 ( .A(n_177), .Y(n_230) );
INVx2_ASAP7_75t_L g188 ( .A(n_179), .Y(n_188) );
INVx2_ASAP7_75t_L g274 ( .A(n_180), .Y(n_274) );
AND2x2_ASAP7_75t_L g338 ( .A(n_180), .B(n_277), .Y(n_338) );
INVx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx1_ASAP7_75t_L g292 ( .A(n_181), .Y(n_292) );
HB1xp67_ASAP7_75t_L g345 ( .A(n_181), .Y(n_345) );
OR2x2_ASAP7_75t_L g416 ( .A(n_181), .B(n_222), .Y(n_416) );
INVx2_ASAP7_75t_L g513 ( .A(n_184), .Y(n_513) );
OAI21xp5_ASAP7_75t_L g536 ( .A1(n_187), .A2(n_537), .B(n_538), .Y(n_536) );
INVx2_ASAP7_75t_L g549 ( .A(n_187), .Y(n_549) );
NAND4xp25_ASAP7_75t_L g294 ( .A(n_191), .B(n_295), .C(n_298), .D(n_300), .Y(n_294) );
INVx1_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
AND2x2_ASAP7_75t_L g432 ( .A(n_192), .B(n_420), .Y(n_432) );
AND2x2_ASAP7_75t_L g192 ( .A(n_193), .B(n_208), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_193), .B(n_261), .Y(n_260) );
AND2x4_ASAP7_75t_L g286 ( .A(n_193), .B(n_287), .Y(n_286) );
INVx2_ASAP7_75t_L g306 ( .A(n_193), .Y(n_306) );
INVx1_ASAP7_75t_L g323 ( .A(n_193), .Y(n_323) );
INVx1_ASAP7_75t_L g331 ( .A(n_193), .Y(n_331) );
HB1xp67_ASAP7_75t_L g445 ( .A(n_193), .Y(n_445) );
INVx4_ASAP7_75t_SL g193 ( .A(n_194), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_194), .B(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_L g363 ( .A(n_194), .B(n_263), .Y(n_363) );
AND2x2_ASAP7_75t_L g371 ( .A(n_194), .B(n_209), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_194), .B(n_394), .Y(n_393) );
BUFx2_ASAP7_75t_L g436 ( .A(n_194), .Y(n_436) );
INVx1_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx1_ASAP7_75t_SL g202 ( .A(n_203), .Y(n_202) );
INVx1_ASAP7_75t_L g229 ( .A(n_203), .Y(n_229) );
INVx1_ASAP7_75t_L g543 ( .A(n_203), .Y(n_543) );
BUFx2_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g551 ( .A(n_205), .B(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx1_ASAP7_75t_L g240 ( .A(n_209), .Y(n_240) );
OR2x2_ASAP7_75t_L g301 ( .A(n_209), .B(n_263), .Y(n_301) );
INVx2_ASAP7_75t_L g308 ( .A(n_209), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_209), .B(n_261), .Y(n_332) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_209), .Y(n_419) );
INVx1_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
INVx1_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
AO31x2_ASAP7_75t_L g222 ( .A1(n_217), .A2(n_223), .A3(n_230), .B(n_231), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g390 ( .A(n_220), .B(n_391), .Y(n_390) );
BUFx2_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
AND2x2_ASAP7_75t_L g243 ( .A(n_222), .B(n_244), .Y(n_243) );
BUFx2_ASAP7_75t_L g253 ( .A(n_222), .Y(n_253) );
INVx2_ASAP7_75t_L g271 ( .A(n_222), .Y(n_271) );
AND2x4_ASAP7_75t_L g303 ( .A(n_222), .B(n_275), .Y(n_303) );
OR2x2_ASAP7_75t_L g383 ( .A(n_222), .B(n_283), .Y(n_383) );
INVx2_ASAP7_75t_SL g225 ( .A(n_226), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g478 ( .A(n_226), .B(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g499 ( .A(n_228), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_234), .B(n_238), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_235), .B(n_251), .Y(n_250) );
OR2x2_ASAP7_75t_L g300 ( .A(n_235), .B(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_235), .B(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_236), .B(n_306), .Y(n_314) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
INVx2_ASAP7_75t_L g259 ( .A(n_237), .Y(n_259) );
OR2x2_ASAP7_75t_L g352 ( .A(n_237), .B(n_262), .Y(n_352) );
INVx1_ASAP7_75t_L g279 ( .A(n_238), .Y(n_279) );
INVx1_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
INVx1_ASAP7_75t_L g251 ( .A(n_239), .Y(n_251) );
INVx1_ASAP7_75t_L g287 ( .A(n_240), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_242), .B(n_243), .Y(n_241) );
OAI322xp33_ASAP7_75t_L g255 ( .A1(n_242), .A2(n_256), .A3(n_269), .B1(n_272), .B2(n_279), .C1(n_280), .C2(n_284), .Y(n_255) );
AND2x4_ASAP7_75t_L g302 ( .A(n_242), .B(n_303), .Y(n_302) );
AOI211xp5_ASAP7_75t_SL g333 ( .A1(n_242), .A2(n_334), .B(n_335), .C(n_339), .Y(n_333) );
AND2x2_ASAP7_75t_L g353 ( .A(n_242), .B(n_243), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_242), .B(n_270), .Y(n_359) );
AND2x4_ASAP7_75t_SL g281 ( .A(n_243), .B(n_282), .Y(n_281) );
NAND3xp33_ASAP7_75t_L g372 ( .A(n_243), .B(n_299), .C(n_327), .Y(n_372) );
AND2x2_ASAP7_75t_L g403 ( .A(n_243), .B(n_404), .Y(n_403) );
AND2x2_ASAP7_75t_L g270 ( .A(n_244), .B(n_271), .Y(n_270) );
INVx3_ASAP7_75t_L g275 ( .A(n_244), .Y(n_275) );
BUFx2_ASAP7_75t_L g343 ( .A(n_244), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_253), .B(n_254), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_253), .B(n_277), .Y(n_276) );
NAND2x1_ASAP7_75t_L g317 ( .A(n_253), .B(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g336 ( .A(n_253), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_254), .B(n_270), .Y(n_401) );
OR2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_260), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
INVx3_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g344 ( .A(n_259), .B(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
HB1xp67_ASAP7_75t_L g297 ( .A(n_263), .Y(n_297) );
AND2x4_ASAP7_75t_L g307 ( .A(n_263), .B(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g394 ( .A(n_263), .Y(n_394) );
INVx2_ASAP7_75t_L g415 ( .A(n_263), .Y(n_415) );
OAI22xp33_ASAP7_75t_L g427 ( .A1(n_269), .A2(n_428), .B1(n_430), .B2(n_431), .Y(n_427) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g339 ( .A(n_270), .B(n_340), .Y(n_339) );
AND2x4_ASAP7_75t_L g293 ( .A(n_271), .B(n_277), .Y(n_293) );
OR2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_276), .Y(n_272) );
INVx1_ASAP7_75t_L g312 ( .A(n_273), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
AND2x4_ASAP7_75t_L g282 ( .A(n_274), .B(n_283), .Y(n_282) );
INVx1_ASAP7_75t_L g404 ( .A(n_274), .Y(n_404) );
INVx2_ASAP7_75t_L g290 ( .A(n_275), .Y(n_290) );
AND2x2_ASAP7_75t_L g318 ( .A(n_275), .B(n_277), .Y(n_318) );
INVx3_ASAP7_75t_L g326 ( .A(n_275), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_275), .B(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g311 ( .A(n_276), .Y(n_311) );
INVx2_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
BUFx2_ASAP7_75t_L g327 ( .A(n_278), .Y(n_327) );
OAI222xp33_ASAP7_75t_L g450 ( .A1(n_280), .A2(n_440), .B1(n_451), .B2(n_454), .C1(n_456), .C2(n_458), .Y(n_450) );
INVx3_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVx1_ASAP7_75t_L g391 ( .A(n_282), .Y(n_391) );
AND2x2_ASAP7_75t_L g455 ( .A(n_282), .B(n_325), .Y(n_455) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_285), .B(n_376), .Y(n_375) );
AOI221xp5_ASAP7_75t_L g288 ( .A1(n_289), .A2(n_294), .B1(n_302), .B2(n_304), .C(n_309), .Y(n_288) );
AND2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
INVx1_ASAP7_75t_L g377 ( .A(n_290), .Y(n_377) );
INVx2_ASAP7_75t_L g439 ( .A(n_291), .Y(n_439) );
AND2x4_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
INVx2_ASAP7_75t_L g340 ( .A(n_292), .Y(n_340) );
AND2x2_ASAP7_75t_L g376 ( .A(n_292), .B(n_377), .Y(n_376) );
AND2x4_ASAP7_75t_L g342 ( .A(n_293), .B(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g368 ( .A(n_293), .B(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g457 ( .A(n_293), .Y(n_457) );
INVx2_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g406 ( .A(n_297), .Y(n_406) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g429 ( .A(n_299), .B(n_307), .Y(n_429) );
AND2x2_ASAP7_75t_L g452 ( .A(n_299), .B(n_453), .Y(n_452) );
OR2x2_ASAP7_75t_L g313 ( .A(n_301), .B(n_314), .Y(n_313) );
INVx2_ASAP7_75t_L g448 ( .A(n_301), .Y(n_448) );
AOI22xp5_ASAP7_75t_L g389 ( .A1(n_302), .A2(n_356), .B1(n_390), .B2(n_392), .Y(n_389) );
OAI21xp5_ASAP7_75t_L g417 ( .A1(n_302), .A2(n_418), .B(n_421), .Y(n_417) );
INVxp67_ASAP7_75t_L g334 ( .A(n_303), .Y(n_334) );
INVx2_ASAP7_75t_SL g438 ( .A(n_303), .Y(n_438) );
AND2x4_ASAP7_75t_L g304 ( .A(n_305), .B(n_307), .Y(n_304) );
OR2x2_ASAP7_75t_L g351 ( .A(n_305), .B(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g449 ( .A(n_305), .B(n_448), .Y(n_449) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g322 ( .A(n_307), .B(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_307), .B(n_331), .Y(n_347) );
INVx2_ASAP7_75t_L g374 ( .A(n_307), .Y(n_374) );
OAI22xp33_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_313), .B1(n_315), .B2(n_317), .Y(n_309) );
NOR2xp33_ASAP7_75t_SL g310 ( .A(n_311), .B(n_312), .Y(n_310) );
AOI22xp5_ASAP7_75t_L g397 ( .A1(n_311), .A2(n_385), .B1(n_398), .B2(n_400), .Y(n_397) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g407 ( .A(n_316), .B(n_408), .Y(n_407) );
AOI21xp5_ASAP7_75t_L g319 ( .A1(n_320), .A2(n_324), .B(n_328), .Y(n_319) );
AND2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
INVx1_ASAP7_75t_L g388 ( .A(n_321), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_321), .B(n_371), .Y(n_399) );
INVx1_ASAP7_75t_L g357 ( .A(n_323), .Y(n_357) );
AND2x2_ASAP7_75t_L g324 ( .A(n_325), .B(n_327), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_325), .B(n_338), .Y(n_430) );
INVx2_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
OAI21xp33_ASAP7_75t_L g443 ( .A1(n_326), .A2(n_444), .B(n_446), .Y(n_443) );
OAI21xp5_ASAP7_75t_SL g328 ( .A1(n_329), .A2(n_333), .B(n_341), .Y(n_328) );
BUFx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
OR2x2_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
INVx1_ASAP7_75t_L g387 ( .A(n_332), .Y(n_387) );
INVx1_ASAP7_75t_L g453 ( .A(n_332), .Y(n_453) );
NOR2xp33_ASAP7_75t_L g335 ( .A(n_336), .B(n_337), .Y(n_335) );
INVx1_ASAP7_75t_L g426 ( .A(n_336), .Y(n_426) );
OR2x2_ASAP7_75t_L g437 ( .A(n_337), .B(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
NAND3xp33_ASAP7_75t_L g341 ( .A(n_342), .B(n_344), .C(n_346), .Y(n_341) );
AOI22xp5_ASAP7_75t_L g402 ( .A1(n_342), .A2(n_403), .B1(n_405), .B2(n_407), .Y(n_402) );
INVx1_ASAP7_75t_L g369 ( .A(n_343), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_344), .B(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g382 ( .A(n_345), .Y(n_382) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_347), .B(n_351), .Y(n_350) );
OAI221xp5_ASAP7_75t_L g409 ( .A1(n_347), .A2(n_410), .B1(n_413), .B2(n_416), .C(n_417), .Y(n_409) );
AOI21xp5_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_353), .B(n_354), .Y(n_348) );
HB1xp67_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx2_ASAP7_75t_L g358 ( .A(n_352), .Y(n_358) );
OAI22xp5_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_359), .B1(n_360), .B2(n_857), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
AND2x4_ASAP7_75t_L g356 ( .A(n_357), .B(n_358), .Y(n_356) );
INVxp67_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx2_ASAP7_75t_SL g361 ( .A(n_362), .Y(n_361) );
AND2x4_ASAP7_75t_L g441 ( .A(n_363), .B(n_419), .Y(n_441) );
NAND4xp25_ASAP7_75t_L g364 ( .A(n_365), .B(n_395), .C(n_422), .D(n_442), .Y(n_364) );
NOR2xp33_ASAP7_75t_L g365 ( .A(n_366), .B(n_378), .Y(n_365) );
OAI221xp5_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_370), .B1(n_372), .B2(n_373), .C(n_375), .Y(n_366) );
AOI22xp33_ASAP7_75t_L g446 ( .A1(n_368), .A2(n_425), .B1(n_447), .B2(n_449), .Y(n_446) );
INVx1_ASAP7_75t_L g421 ( .A(n_370), .Y(n_421) );
INVx2_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g405 ( .A(n_371), .B(n_406), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_371), .B(n_414), .Y(n_413) );
NAND2x1_ASAP7_75t_L g458 ( .A(n_371), .B(n_459), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g434 ( .A(n_373), .B(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g380 ( .A(n_377), .B(n_381), .Y(n_380) );
OAI21xp33_ASAP7_75t_SL g378 ( .A1(n_379), .A2(n_384), .B(n_389), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
NOR2x1_ASAP7_75t_L g381 ( .A(n_382), .B(n_383), .Y(n_381) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_387), .B(n_388), .Y(n_386) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g408 ( .A(n_394), .Y(n_408) );
AOI211xp5_ASAP7_75t_L g422 ( .A1(n_394), .A2(n_423), .B(n_427), .C(n_433), .Y(n_422) );
NOR2xp33_ASAP7_75t_L g395 ( .A(n_396), .B(n_409), .Y(n_395) );
NAND2xp5_ASAP7_75t_SL g396 ( .A(n_397), .B(n_402), .Y(n_396) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
OR2x2_ASAP7_75t_L g456 ( .A(n_404), .B(n_457), .Y(n_456) );
HB1xp67_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
AND2x4_ASAP7_75t_L g418 ( .A(n_419), .B(n_420), .Y(n_418) );
INVx3_ASAP7_75t_L g460 ( .A(n_420), .Y(n_460) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
NAND2x1p5_ASAP7_75t_L g424 ( .A(n_425), .B(n_426), .Y(n_424) );
INVx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
OAI22xp33_ASAP7_75t_R g433 ( .A1(n_434), .A2(n_437), .B1(n_439), .B2(n_440), .Y(n_433) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
AND2x4_ASAP7_75t_L g447 ( .A(n_436), .B(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
NOR2xp33_ASAP7_75t_L g442 ( .A(n_443), .B(n_450), .Y(n_442) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
BUFx8_ASAP7_75t_SL g461 ( .A(n_462), .Y(n_461) );
CKINVDCx5p33_ASAP7_75t_R g809 ( .A(n_462), .Y(n_809) );
AND2x2_ASAP7_75t_L g846 ( .A(n_462), .B(n_847), .Y(n_846) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
NAND2xp5_ASAP7_75t_SL g464 ( .A(n_465), .B(n_805), .Y(n_464) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
AOI21xp5_ASAP7_75t_L g805 ( .A1(n_467), .A2(n_806), .B(n_807), .Y(n_805) );
XNOR2xp5_ASAP7_75t_L g824 ( .A(n_467), .B(n_825), .Y(n_824) );
AND2x4_ASAP7_75t_L g467 ( .A(n_468), .B(n_693), .Y(n_467) );
NOR4xp75_ASAP7_75t_L g468 ( .A(n_469), .B(n_632), .C(n_656), .D(n_675), .Y(n_468) );
NAND3x1_ASAP7_75t_L g469 ( .A(n_470), .B(n_573), .C(n_623), .Y(n_469) );
AOI22xp5_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_516), .B1(n_553), .B2(n_569), .Y(n_470) );
AND2x2_ASAP7_75t_L g754 ( .A(n_471), .B(n_629), .Y(n_754) );
AND2x2_ASAP7_75t_L g471 ( .A(n_472), .B(n_488), .Y(n_471) );
AND2x2_ASAP7_75t_L g704 ( .A(n_472), .B(n_705), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_472), .B(n_709), .Y(n_708) );
INVx2_ASAP7_75t_L g731 ( .A(n_472), .Y(n_731) );
INVx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g577 ( .A(n_473), .Y(n_577) );
INVx2_ASAP7_75t_L g598 ( .A(n_473), .Y(n_598) );
AND2x2_ASAP7_75t_L g692 ( .A(n_473), .B(n_655), .Y(n_692) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g572 ( .A(n_474), .Y(n_572) );
AND2x2_ASAP7_75t_L g671 ( .A(n_474), .B(n_584), .Y(n_671) );
AOI21x1_ASAP7_75t_L g474 ( .A1(n_475), .A2(n_476), .B(n_486), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_477), .B(n_482), .Y(n_476) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_480), .A2(n_493), .B(n_494), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_480), .A2(n_508), .B(n_509), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_480), .A2(n_526), .B(n_527), .Y(n_525) );
AOI21xp5_ASAP7_75t_L g590 ( .A1(n_480), .A2(n_591), .B(n_592), .Y(n_590) );
BUFx4f_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
AND2x2_ASAP7_75t_L g624 ( .A(n_488), .B(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g739 ( .A(n_488), .Y(n_739) );
AND2x2_ASAP7_75t_L g745 ( .A(n_488), .B(n_609), .Y(n_745) );
AND2x2_ASAP7_75t_L g488 ( .A(n_489), .B(n_503), .Y(n_488) );
INVx1_ASAP7_75t_L g582 ( .A(n_489), .Y(n_582) );
INVx4_ASAP7_75t_L g602 ( .A(n_489), .Y(n_602) );
OR2x2_ASAP7_75t_L g651 ( .A(n_489), .B(n_631), .Y(n_651) );
BUFx2_ASAP7_75t_L g720 ( .A(n_489), .Y(n_720) );
AND2x4_ASAP7_75t_L g489 ( .A(n_490), .B(n_491), .Y(n_489) );
OAI21x1_ASAP7_75t_L g491 ( .A1(n_492), .A2(n_495), .B(n_501), .Y(n_491) );
OAI22xp5_ASAP7_75t_L g495 ( .A1(n_496), .A2(n_498), .B1(n_499), .B2(n_500), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g564 ( .A1(n_497), .A2(n_565), .B(n_566), .Y(n_564) );
INVx2_ASAP7_75t_SL g497 ( .A(n_498), .Y(n_497) );
OAI21x1_ASAP7_75t_L g506 ( .A1(n_502), .A2(n_507), .B(n_510), .Y(n_506) );
OAI21x1_ASAP7_75t_L g524 ( .A1(n_502), .A2(n_525), .B(n_528), .Y(n_524) );
OAI21x1_ASAP7_75t_L g535 ( .A1(n_502), .A2(n_536), .B(n_539), .Y(n_535) );
OAI21x1_ASAP7_75t_L g560 ( .A1(n_502), .A2(n_561), .B(n_564), .Y(n_560) );
OAI21x1_ASAP7_75t_L g586 ( .A1(n_502), .A2(n_587), .B(n_590), .Y(n_586) );
AND2x2_ASAP7_75t_L g571 ( .A(n_503), .B(n_572), .Y(n_571) );
INVx2_ASAP7_75t_L g673 ( .A(n_503), .Y(n_673) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g597 ( .A(n_504), .Y(n_597) );
OAI21x1_ASAP7_75t_L g504 ( .A1(n_505), .A2(n_506), .B(n_515), .Y(n_504) );
OAI21xp5_ASAP7_75t_L g559 ( .A1(n_505), .A2(n_560), .B(n_567), .Y(n_559) );
OAI21xp33_ASAP7_75t_SL g611 ( .A1(n_505), .A2(n_506), .B(n_515), .Y(n_611) );
OAI21x1_ASAP7_75t_L g622 ( .A1(n_505), .A2(n_560), .B(n_567), .Y(n_622) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_511), .A2(n_512), .B(n_514), .Y(n_510) );
INVx2_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
NAND2x1_ASAP7_75t_L g742 ( .A(n_518), .B(n_682), .Y(n_742) );
AND2x4_ASAP7_75t_L g518 ( .A(n_519), .B(n_532), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
OR2x2_ASAP7_75t_L g627 ( .A(n_520), .B(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g647 ( .A(n_520), .B(n_648), .Y(n_647) );
HB1xp67_ASAP7_75t_L g681 ( .A(n_520), .Y(n_681) );
INVx3_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
AND2x2_ASAP7_75t_L g637 ( .A(n_521), .B(n_534), .Y(n_637) );
NOR2xp67_ASAP7_75t_L g792 ( .A(n_521), .B(n_533), .Y(n_792) );
BUFx3_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g714 ( .A(n_522), .Y(n_714) );
OAI21x1_ASAP7_75t_L g522 ( .A1(n_523), .A2(n_524), .B(n_531), .Y(n_522) );
OAI21x1_ASAP7_75t_L g534 ( .A1(n_523), .A2(n_535), .B(n_544), .Y(n_534) );
OAI21x1_ASAP7_75t_L g557 ( .A1(n_523), .A2(n_524), .B(n_531), .Y(n_557) );
OA21x2_ASAP7_75t_L g568 ( .A1(n_523), .A2(n_535), .B(n_544), .Y(n_568) );
INVx2_ASAP7_75t_L g735 ( .A(n_532), .Y(n_735) );
AND2x4_ASAP7_75t_L g773 ( .A(n_532), .B(n_712), .Y(n_773) );
AND2x4_ASAP7_75t_L g532 ( .A(n_533), .B(n_545), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g613 ( .A(n_534), .Y(n_613) );
AND2x2_ASAP7_75t_L g648 ( .A(n_534), .B(n_546), .Y(n_648) );
AND2x2_ASAP7_75t_L g771 ( .A(n_534), .B(n_621), .Y(n_771) );
AND2x2_ASAP7_75t_L g782 ( .A(n_534), .B(n_559), .Y(n_782) );
AOI21x1_ASAP7_75t_L g539 ( .A1(n_540), .A2(n_541), .B(n_543), .Y(n_539) );
AND2x2_ASAP7_75t_L g640 ( .A(n_545), .B(n_557), .Y(n_640) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
OR2x2_ASAP7_75t_L g556 ( .A(n_546), .B(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g614 ( .A(n_546), .B(n_557), .Y(n_614) );
OR2x2_ASAP7_75t_L g628 ( .A(n_546), .B(n_568), .Y(n_628) );
AND2x2_ASAP7_75t_L g713 ( .A(n_546), .B(n_714), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_546), .B(n_568), .Y(n_724) );
HB1xp67_ASAP7_75t_L g766 ( .A(n_546), .Y(n_766) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_555), .B(n_558), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g662 ( .A(n_556), .Y(n_662) );
NAND3xp33_ASAP7_75t_L g769 ( .A(n_556), .B(n_770), .C(n_772), .Y(n_769) );
INVx1_ASAP7_75t_L g606 ( .A(n_557), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_558), .B(n_614), .Y(n_736) );
AND2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_568), .Y(n_558) );
INVx1_ASAP7_75t_L g580 ( .A(n_559), .Y(n_580) );
AND2x2_ASAP7_75t_L g785 ( .A(n_568), .B(n_621), .Y(n_785) );
INVx1_ASAP7_75t_L g788 ( .A(n_569), .Y(n_788) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
OR2x2_ASAP7_75t_L g767 ( .A(n_570), .B(n_600), .Y(n_767) );
OR2x2_ASAP7_75t_L g778 ( .A(n_570), .B(n_651), .Y(n_778) );
INVx2_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g654 ( .A(n_571), .B(n_655), .Y(n_654) );
AND2x2_ASAP7_75t_L g802 ( .A(n_571), .B(n_581), .Y(n_802) );
AND2x2_ASAP7_75t_L g610 ( .A(n_572), .B(n_611), .Y(n_610) );
A2O1A1O1Ixp25_ASAP7_75t_L g573 ( .A1(n_574), .A2(n_578), .B(n_594), .C(n_603), .D(n_607), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g688 ( .A(n_576), .B(n_689), .Y(n_688) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g625 ( .A(n_577), .Y(n_625) );
INVx1_ASAP7_75t_L g660 ( .A(n_578), .Y(n_660) );
AND2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_581), .Y(n_578) );
AND2x2_ASAP7_75t_L g639 ( .A(n_579), .B(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
OR2x2_ASAP7_75t_L g630 ( .A(n_580), .B(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g659 ( .A(n_581), .Y(n_659) );
AND2x2_ASAP7_75t_L g730 ( .A(n_581), .B(n_731), .Y(n_730) );
AND2x2_ASAP7_75t_L g776 ( .A(n_581), .B(n_610), .Y(n_776) );
AND2x2_ASAP7_75t_L g581 ( .A(n_582), .B(n_583), .Y(n_581) );
INVx1_ASAP7_75t_L g601 ( .A(n_583), .Y(n_601) );
HB1xp67_ASAP7_75t_L g609 ( .A(n_583), .Y(n_609) );
INVx2_ASAP7_75t_L g655 ( .A(n_583), .Y(n_655) );
INVx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g631 ( .A(n_584), .Y(n_631) );
OAI21x1_ASAP7_75t_L g584 ( .A1(n_585), .A2(n_586), .B(n_593), .Y(n_584) );
INVx1_ASAP7_75t_L g726 ( .A(n_594), .Y(n_726) );
AND2x2_ASAP7_75t_L g594 ( .A(n_595), .B(n_599), .Y(n_594) );
OAI21xp33_ASAP7_75t_L g650 ( .A1(n_595), .A2(n_600), .B(n_651), .Y(n_650) );
AND2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_598), .Y(n_595) );
AND2x2_ASAP7_75t_L g616 ( .A(n_596), .B(n_617), .Y(n_616) );
AND2x2_ASAP7_75t_L g721 ( .A(n_596), .B(n_671), .Y(n_721) );
INVx2_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g653 ( .A(n_597), .B(n_631), .Y(n_653) );
AND2x2_ASAP7_75t_L g677 ( .A(n_598), .B(n_602), .Y(n_677) );
NAND2xp5_ASAP7_75t_SL g761 ( .A(n_598), .B(n_617), .Y(n_761) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx1_ASAP7_75t_SL g705 ( .A(n_600), .Y(n_705) );
OR2x2_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
INVx2_ASAP7_75t_L g617 ( .A(n_602), .Y(n_617) );
NAND2x1_ASAP7_75t_L g672 ( .A(n_602), .B(n_673), .Y(n_672) );
OAI32xp33_ASAP7_75t_L g793 ( .A1(n_603), .A2(n_669), .A3(n_777), .B1(n_794), .B2(n_795), .Y(n_793) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
HB1xp67_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g667 ( .A(n_605), .Y(n_667) );
AND2x2_ASAP7_75t_L g690 ( .A(n_605), .B(n_648), .Y(n_690) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g687 ( .A(n_606), .B(n_621), .Y(n_687) );
OAI22xp33_ASAP7_75t_SL g607 ( .A1(n_608), .A2(n_612), .B1(n_615), .B2(n_618), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_609), .B(n_610), .Y(n_608) );
AND2x2_ASAP7_75t_L g644 ( .A(n_610), .B(n_645), .Y(n_644) );
BUFx2_ASAP7_75t_L g663 ( .A(n_611), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
INVx2_ASAP7_75t_L g777 ( .A(n_613), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_614), .B(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g756 ( .A(n_614), .Y(n_756) );
AND2x2_ASAP7_75t_L g784 ( .A(n_614), .B(n_785), .Y(n_784) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
AND2x4_ASAP7_75t_L g691 ( .A(n_616), .B(n_692), .Y(n_691) );
O2A1O1Ixp33_ASAP7_75t_L g740 ( .A1(n_616), .A2(n_671), .B(n_741), .C(n_743), .Y(n_740) );
INVx1_ASAP7_75t_L g645 ( .A(n_617), .Y(n_645) );
AND2x2_ASAP7_75t_L g689 ( .A(n_617), .B(n_655), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_619), .B(n_640), .Y(n_658) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVxp67_ASAP7_75t_SL g636 ( .A(n_621), .Y(n_636) );
INVxp67_ASAP7_75t_SL g683 ( .A(n_621), .Y(n_683) );
INVx1_ASAP7_75t_L g712 ( .A(n_621), .Y(n_712) );
BUFx3_ASAP7_75t_L g725 ( .A(n_621), .Y(n_725) );
INVx3_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
NAND3xp33_ASAP7_75t_L g623 ( .A(n_624), .B(n_626), .C(n_629), .Y(n_623) );
INVx1_ASAP7_75t_L g747 ( .A(n_624), .Y(n_747) );
OR2x2_ASAP7_75t_L g674 ( .A(n_625), .B(n_659), .Y(n_674) );
OR2x2_ASAP7_75t_L g638 ( .A(n_626), .B(n_639), .Y(n_638) );
INVx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
OAI22xp33_ASAP7_75t_L g664 ( .A1(n_627), .A2(n_665), .B1(n_669), .B2(n_674), .Y(n_664) );
INVx2_ASAP7_75t_L g668 ( .A(n_628), .Y(n_668) );
HB1xp67_ASAP7_75t_L g680 ( .A(n_628), .Y(n_680) );
INVx1_ASAP7_75t_L g699 ( .A(n_628), .Y(n_699) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVxp67_ASAP7_75t_L g643 ( .A(n_631), .Y(n_643) );
HB1xp67_ASAP7_75t_L g738 ( .A(n_631), .Y(n_738) );
OAI22xp5_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_641), .B1(n_646), .B2(n_649), .Y(n_632) );
NOR2x1_ASAP7_75t_L g633 ( .A(n_634), .B(n_638), .Y(n_633) );
BUFx2_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
AND2x4_ASAP7_75t_L g635 ( .A(n_636), .B(n_637), .Y(n_635) );
HB1xp67_ASAP7_75t_L g718 ( .A(n_640), .Y(n_718) );
NAND2x1p5_ASAP7_75t_L g641 ( .A(n_642), .B(n_644), .Y(n_641) );
INVx1_ASAP7_75t_L g709 ( .A(n_642), .Y(n_709) );
BUFx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
AOI221x1_ASAP7_75t_L g695 ( .A1(n_644), .A2(n_696), .B1(n_700), .B2(n_702), .C(n_706), .Y(n_695) );
BUFx2_ASAP7_75t_L g798 ( .A(n_645), .Y(n_798) );
INVx2_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_648), .B(n_687), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_648), .B(n_725), .Y(n_750) );
AND2x2_ASAP7_75t_L g804 ( .A(n_648), .B(n_683), .Y(n_804) );
AOI21xp5_ASAP7_75t_L g649 ( .A1(n_650), .A2(n_652), .B(n_654), .Y(n_649) );
AOI211xp5_ASAP7_75t_L g786 ( .A1(n_651), .A2(n_787), .B(n_793), .C(n_796), .Y(n_786) );
OAI222xp33_ASAP7_75t_L g774 ( .A1(n_652), .A2(n_775), .B1(n_777), .B2(n_778), .C1(n_779), .C2(n_783), .Y(n_774) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
AO21x1_ASAP7_75t_L g656 ( .A1(n_657), .A2(n_663), .B(n_664), .Y(n_656) );
OAI22xp5_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_659), .B1(n_660), .B2(n_661), .Y(n_657) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx2_ASAP7_75t_L g800 ( .A(n_663), .Y(n_800) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
AND2x4_ASAP7_75t_L g666 ( .A(n_667), .B(n_668), .Y(n_666) );
AND2x2_ASAP7_75t_L g701 ( .A(n_668), .B(n_687), .Y(n_701) );
INVx1_ASAP7_75t_L g727 ( .A(n_668), .Y(n_727) );
OAI22xp5_ASAP7_75t_L g722 ( .A1(n_669), .A2(n_723), .B1(n_726), .B2(n_727), .Y(n_722) );
INVx1_ASAP7_75t_L g753 ( .A(n_669), .Y(n_753) );
OR2x6_ASAP7_75t_L g669 ( .A(n_670), .B(n_672), .Y(n_669) );
INVx1_ASAP7_75t_L g799 ( .A(n_670), .Y(n_799) );
INVx2_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_SL g760 ( .A(n_673), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_673), .B(n_689), .Y(n_794) );
OAI21xp33_ASAP7_75t_SL g675 ( .A1(n_676), .A2(n_678), .B(n_684), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx2_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
NOR3x1_ASAP7_75t_L g679 ( .A(n_680), .B(n_681), .C(n_682), .Y(n_679) );
BUFx2_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
AOI22xp5_ASAP7_75t_L g684 ( .A1(n_685), .A2(n_688), .B1(n_690), .B2(n_691), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_687), .B(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g772 ( .A(n_687), .Y(n_772) );
INVx2_ASAP7_75t_L g746 ( .A(n_690), .Y(n_746) );
INVx3_ASAP7_75t_L g707 ( .A(n_691), .Y(n_707) );
NOR2x1_ASAP7_75t_L g693 ( .A(n_694), .B(n_751), .Y(n_693) );
NAND3xp33_ASAP7_75t_L g694 ( .A(n_695), .B(n_715), .C(n_740), .Y(n_694) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
HB1xp67_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx2_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
AOI21xp5_ASAP7_75t_L g706 ( .A1(n_707), .A2(n_708), .B(n_710), .Y(n_706) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
AND2x2_ASAP7_75t_L g711 ( .A(n_712), .B(n_713), .Y(n_711) );
INVx1_ASAP7_75t_L g763 ( .A(n_712), .Y(n_763) );
BUFx2_ASAP7_75t_L g734 ( .A(n_714), .Y(n_734) );
AOI211xp5_ASAP7_75t_L g715 ( .A1(n_716), .A2(n_719), .B(n_722), .C(n_728), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
AND2x4_ASAP7_75t_L g719 ( .A(n_720), .B(n_721), .Y(n_719) );
OR2x2_ASAP7_75t_L g723 ( .A(n_724), .B(n_725), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g791 ( .A(n_725), .B(n_792), .Y(n_791) );
OAI22xp33_ASAP7_75t_L g728 ( .A1(n_729), .A2(n_732), .B1(n_736), .B2(n_737), .Y(n_728) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
OR2x2_ASAP7_75t_L g732 ( .A(n_733), .B(n_735), .Y(n_732) );
AND2x2_ASAP7_75t_L g780 ( .A(n_733), .B(n_771), .Y(n_780) );
INVx2_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
AND2x2_ASAP7_75t_L g781 ( .A(n_734), .B(n_782), .Y(n_781) );
OR2x2_ASAP7_75t_L g737 ( .A(n_738), .B(n_739), .Y(n_737) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
OAI22xp5_ASAP7_75t_L g743 ( .A1(n_744), .A2(n_746), .B1(n_747), .B2(n_748), .Y(n_743) );
INVx3_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVxp67_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
NAND3xp33_ASAP7_75t_L g751 ( .A(n_752), .B(n_757), .C(n_786), .Y(n_751) );
OAI21xp33_ASAP7_75t_L g752 ( .A1(n_753), .A2(n_754), .B(n_755), .Y(n_752) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
NOR2xp33_ASAP7_75t_L g757 ( .A(n_758), .B(n_774), .Y(n_757) );
OAI22xp33_ASAP7_75t_L g758 ( .A1(n_759), .A2(n_762), .B1(n_767), .B2(n_768), .Y(n_758) );
OR2x2_ASAP7_75t_L g759 ( .A(n_760), .B(n_761), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_763), .B(n_764), .Y(n_762) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
NOR2xp67_ASAP7_75t_L g768 ( .A(n_769), .B(n_773), .Y(n_768) );
INVx2_ASAP7_75t_SL g770 ( .A(n_771), .Y(n_770) );
INVx2_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
NOR2xp33_ASAP7_75t_SL g779 ( .A(n_780), .B(n_781), .Y(n_779) );
INVx2_ASAP7_75t_L g795 ( .A(n_781), .Y(n_795) );
INVx2_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
NOR2xp33_ASAP7_75t_L g787 ( .A(n_788), .B(n_789), .Y(n_787) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
INVx1_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
AOI21xp33_ASAP7_75t_L g796 ( .A1(n_797), .A2(n_801), .B(n_803), .Y(n_796) );
NAND3x2_ASAP7_75t_L g797 ( .A(n_798), .B(n_799), .C(n_800), .Y(n_797) );
INVx1_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
INVxp67_ASAP7_75t_SL g803 ( .A(n_804), .Y(n_803) );
INVx4_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
BUFx12f_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
OAI21xp5_ASAP7_75t_L g810 ( .A1(n_811), .A2(n_816), .B(n_839), .Y(n_810) );
INVx4_ASAP7_75t_SL g811 ( .A(n_812), .Y(n_811) );
BUFx6f_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
CKINVDCx11_ASAP7_75t_R g813 ( .A(n_814), .Y(n_813) );
BUFx6f_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
AOI21xp5_ASAP7_75t_L g816 ( .A1(n_817), .A2(n_818), .B(n_830), .Y(n_816) );
OAI31xp33_ASAP7_75t_SL g830 ( .A1(n_817), .A2(n_824), .A3(n_831), .B(n_834), .Y(n_830) );
AND2x2_ASAP7_75t_L g818 ( .A(n_819), .B(n_824), .Y(n_818) );
CKINVDCx5p33_ASAP7_75t_R g819 ( .A(n_820), .Y(n_819) );
INVx5_ASAP7_75t_L g833 ( .A(n_820), .Y(n_833) );
INVx4_ASAP7_75t_L g838 ( .A(n_820), .Y(n_838) );
INVx1_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
INVx1_ASAP7_75t_L g829 ( .A(n_826), .Y(n_829) );
INVx1_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
BUFx2_ASAP7_75t_SL g832 ( .A(n_833), .Y(n_832) );
INVxp67_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
NOR2xp33_ASAP7_75t_L g835 ( .A(n_836), .B(n_837), .Y(n_835) );
BUFx12f_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
INVx2_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
INVx1_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
BUFx10_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
INVx1_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
AND2x6_ASAP7_75t_L g851 ( .A(n_846), .B(n_852), .Y(n_851) );
BUFx6f_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
CKINVDCx5p33_ASAP7_75t_R g849 ( .A(n_850), .Y(n_849) );
INVx5_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
BUFx5_ASAP7_75t_L g855 ( .A(n_851), .Y(n_855) );
CKINVDCx11_ASAP7_75t_R g854 ( .A(n_855), .Y(n_854) );
endmodule