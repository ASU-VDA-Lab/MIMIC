module fake_jpeg_15435_n_313 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_313);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_313;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx24_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_20),
.B(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_20),
.B(n_0),
.Y(n_38)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_26),
.B(n_1),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_22),
.Y(n_51)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_17),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_17),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_40),
.A2(n_35),
.B(n_38),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_44),
.A2(n_46),
.B1(n_55),
.B2(n_39),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_43),
.A2(n_20),
.B1(n_21),
.B2(n_32),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_45),
.B(n_51),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_40),
.A2(n_38),
.B1(n_35),
.B2(n_37),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_61),
.Y(n_72)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

BUFx4f_ASAP7_75t_SL g74 ( 
.A(n_48),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_43),
.A2(n_21),
.B1(n_23),
.B2(n_32),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_50),
.A2(n_63),
.B1(n_67),
.B2(n_41),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_26),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_54),
.B(n_56),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_37),
.A2(n_27),
.B1(n_31),
.B2(n_30),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_26),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_57),
.Y(n_96)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_58),
.B(n_60),
.Y(n_92)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_23),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_36),
.A2(n_25),
.B1(n_31),
.B2(n_30),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_26),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_66),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_27),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_39),
.A2(n_25),
.B1(n_41),
.B2(n_18),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_66),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_69),
.B(n_70),
.Y(n_102)
);

INVx6_ASAP7_75t_SL g70 ( 
.A(n_49),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_71),
.B(n_73),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_56),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_33),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_75),
.B(n_80),
.Y(n_110)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_76),
.Y(n_101)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_77),
.Y(n_123)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_78),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_46),
.B(n_39),
.Y(n_80)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_81),
.Y(n_105)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_83),
.Y(n_122)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

AND2x2_ASAP7_75t_SL g85 ( 
.A(n_51),
.B(n_64),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_85),
.A2(n_44),
.B(n_68),
.Y(n_100)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_86),
.B(n_89),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_L g88 ( 
.A1(n_54),
.A2(n_39),
.B1(n_24),
.B2(n_29),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_88),
.A2(n_94),
.B1(n_53),
.B2(n_58),
.Y(n_111)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_57),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_90),
.B(n_95),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_91),
.B(n_2),
.Y(n_106)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_93),
.Y(n_113)
);

OA22x2_ASAP7_75t_L g94 ( 
.A1(n_53),
.A2(n_33),
.B1(n_24),
.B2(n_29),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_65),
.B(n_33),
.Y(n_95)
);

INVx2_ASAP7_75t_R g98 ( 
.A(n_93),
.Y(n_98)
);

OAI21xp33_ASAP7_75t_SL g129 ( 
.A1(n_98),
.A2(n_111),
.B(n_94),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_92),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_99),
.B(n_109),
.Y(n_134)
);

MAJx2_ASAP7_75t_L g143 ( 
.A(n_100),
.B(n_117),
.C(n_98),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_68),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_103),
.B(n_69),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_106),
.A2(n_107),
.B(n_117),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_87),
.B(n_2),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_84),
.Y(n_108)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_108),
.Y(n_127)
);

INVx13_ASAP7_75t_L g109 ( 
.A(n_74),
.Y(n_109)
);

INVx13_ASAP7_75t_L g114 ( 
.A(n_74),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_118),
.Y(n_139)
);

AND2x6_ASAP7_75t_L g116 ( 
.A(n_91),
.B(n_2),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_116),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_82),
.A2(n_60),
.B(n_33),
.Y(n_117)
);

INVx13_ASAP7_75t_L g118 ( 
.A(n_74),
.Y(n_118)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_78),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_119),
.B(n_122),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_79),
.B(n_73),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_120),
.A2(n_94),
.B(n_83),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_85),
.B(n_48),
.C(n_57),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_124),
.B(n_75),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_101),
.A2(n_80),
.B1(n_79),
.B2(n_82),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_125),
.A2(n_138),
.B1(n_137),
.B2(n_135),
.Y(n_175)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_126),
.B(n_152),
.Y(n_179)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_104),
.Y(n_128)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_128),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_129),
.A2(n_101),
.B1(n_113),
.B2(n_106),
.Y(n_155)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_104),
.Y(n_131)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_131),
.Y(n_184)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_97),
.Y(n_132)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_132),
.Y(n_157)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_97),
.Y(n_133)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_133),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_135),
.B(n_136),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_103),
.B(n_82),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_120),
.B(n_85),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_137),
.B(n_138),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_120),
.B(n_85),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_108),
.Y(n_140)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_140),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_141),
.B(n_113),
.C(n_111),
.Y(n_156)
);

XNOR2x1_ASAP7_75t_L g185 ( 
.A(n_143),
.B(n_22),
.Y(n_185)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_144),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_121),
.B(n_72),
.Y(n_145)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_145),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_102),
.B(n_72),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_146),
.B(n_148),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_110),
.B(n_71),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_147),
.B(n_150),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_110),
.B(n_94),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_149),
.A2(n_22),
.B(n_74),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_100),
.B(n_124),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_112),
.B(n_98),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_151),
.B(n_28),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_115),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_122),
.Y(n_153)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_153),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_107),
.B(n_86),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_154),
.A2(n_109),
.B(n_114),
.Y(n_181)
);

AO21x1_ASAP7_75t_L g210 ( 
.A1(n_155),
.A2(n_165),
.B(n_181),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_156),
.B(n_141),
.C(n_130),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_150),
.A2(n_106),
.B1(n_116),
.B2(n_107),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_159),
.A2(n_163),
.B1(n_168),
.B2(n_171),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_127),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_160),
.B(n_170),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_136),
.A2(n_99),
.B1(n_123),
.B2(n_77),
.Y(n_163)
);

BUFx12f_ASAP7_75t_L g167 ( 
.A(n_127),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_167),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_149),
.A2(n_123),
.B1(n_119),
.B2(n_90),
.Y(n_168)
);

XOR2x2_ASAP7_75t_L g169 ( 
.A(n_143),
.B(n_19),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_169),
.A2(n_172),
.B(n_178),
.Y(n_198)
);

INVx13_ASAP7_75t_L g170 ( 
.A(n_139),
.Y(n_170)
);

AO21x2_ASAP7_75t_SL g171 ( 
.A1(n_143),
.A2(n_147),
.B(n_151),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_142),
.A2(n_70),
.B1(n_96),
.B2(n_109),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_173),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_175),
.B(n_176),
.Y(n_202)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_153),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_142),
.A2(n_148),
.B(n_130),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_185),
.B(n_134),
.Y(n_211)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_183),
.Y(n_187)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_187),
.Y(n_227)
);

BUFx24_ASAP7_75t_SL g189 ( 
.A(n_180),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_189),
.B(n_194),
.Y(n_220)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_183),
.Y(n_191)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_191),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_157),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_193),
.B(n_197),
.Y(n_215)
);

BUFx24_ASAP7_75t_SL g194 ( 
.A(n_158),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_167),
.Y(n_195)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_195),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_162),
.B(n_125),
.Y(n_196)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_196),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_162),
.B(n_128),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_167),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_199),
.B(n_200),
.Y(n_230)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_164),
.Y(n_200)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_179),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_201),
.Y(n_223)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_174),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_203),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_204),
.B(n_156),
.C(n_182),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_170),
.B(n_152),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_205),
.Y(n_219)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_161),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_206),
.Y(n_234)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_161),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_207),
.B(n_209),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_185),
.B(n_154),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_208),
.A2(n_202),
.B(n_188),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_166),
.B(n_131),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_211),
.B(n_118),
.Y(n_233)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_184),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_212),
.A2(n_176),
.B1(n_184),
.B2(n_177),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_213),
.B(n_214),
.C(n_216),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_204),
.B(n_169),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_198),
.B(n_178),
.Y(n_216)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_218),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_211),
.B(n_175),
.C(n_171),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_221),
.B(n_224),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_198),
.B(n_171),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_190),
.A2(n_171),
.B1(n_173),
.B2(n_155),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_225),
.B(n_208),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_196),
.B(n_159),
.C(n_181),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_226),
.B(n_231),
.Y(n_247)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_228),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_188),
.B(n_163),
.C(n_172),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_233),
.B(n_236),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_197),
.B(n_140),
.C(n_133),
.Y(n_236)
);

AOI22x1_ASAP7_75t_L g237 ( 
.A1(n_210),
.A2(n_126),
.B1(n_105),
.B2(n_24),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_237),
.A2(n_201),
.B1(n_192),
.B2(n_132),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_216),
.A2(n_190),
.B(n_208),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_238),
.A2(n_243),
.B(n_256),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_220),
.B(n_209),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_239),
.B(n_251),
.Y(n_262)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_223),
.Y(n_241)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_241),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_224),
.B(n_210),
.Y(n_243)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_230),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_246),
.B(n_250),
.Y(n_258)
);

OR2x2_ASAP7_75t_L g259 ( 
.A(n_248),
.B(n_253),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_249),
.A2(n_236),
.B1(n_221),
.B2(n_213),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_223),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_222),
.B(n_186),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_219),
.B(n_186),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_252),
.B(n_253),
.Y(n_263)
);

BUFx12_ASAP7_75t_L g253 ( 
.A(n_237),
.Y(n_253)
);

AO21x1_ASAP7_75t_L g254 ( 
.A1(n_235),
.A2(n_29),
.B(n_34),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_254),
.B(n_255),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_217),
.B(n_18),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_215),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_259),
.B(n_268),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_243),
.A2(n_226),
.B1(n_231),
.B2(n_234),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_261),
.B(n_267),
.Y(n_277)
);

INVxp67_ASAP7_75t_SL g266 ( 
.A(n_250),
.Y(n_266)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_266),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_242),
.A2(n_232),
.B1(n_229),
.B2(n_227),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_245),
.B(n_214),
.C(n_233),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_269),
.B(n_270),
.C(n_271),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_245),
.B(n_105),
.C(n_48),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_257),
.B(n_48),
.C(n_34),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_257),
.B(n_34),
.C(n_28),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_272),
.B(n_253),
.Y(n_282)
);

NAND3xp33_ASAP7_75t_L g273 ( 
.A(n_262),
.B(n_244),
.C(n_238),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_273),
.B(n_285),
.Y(n_296)
);

BUFx24_ASAP7_75t_SL g274 ( 
.A(n_258),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_280),
.Y(n_287)
);

OAI21xp33_ASAP7_75t_L g278 ( 
.A1(n_260),
.A2(n_240),
.B(n_244),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_278),
.A2(n_281),
.B(n_282),
.Y(n_294)
);

NOR2xp67_ASAP7_75t_L g279 ( 
.A(n_270),
.B(n_254),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_279),
.B(n_28),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_263),
.A2(n_247),
.B(n_248),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_247),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_265),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_284),
.B(n_89),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_266),
.A2(n_3),
.B(n_4),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_283),
.B(n_264),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_286),
.B(n_289),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_275),
.A2(n_259),
.B1(n_271),
.B2(n_272),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_288),
.B(n_292),
.Y(n_300)
);

AO21x1_ASAP7_75t_L g290 ( 
.A1(n_278),
.A2(n_3),
.B(n_4),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_290),
.B(n_295),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_291),
.A2(n_7),
.B(n_8),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_277),
.B(n_96),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_276),
.A2(n_281),
.B1(n_4),
.B2(n_6),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_276),
.B(n_18),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_296),
.B(n_81),
.C(n_6),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_297),
.B(n_298),
.C(n_301),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_293),
.B(n_6),
.C(n_7),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_299),
.B(n_9),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_294),
.B(n_8),
.C(n_9),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_304),
.A2(n_306),
.B1(n_307),
.B2(n_308),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_302),
.B(n_287),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_300),
.A2(n_303),
.B(n_288),
.Y(n_307)
);

AOI322xp5_ASAP7_75t_L g308 ( 
.A1(n_300),
.A2(n_9),
.A3(n_10),
.B1(n_11),
.B2(n_13),
.C1(n_14),
.C2(n_15),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_305),
.A2(n_10),
.B1(n_13),
.B2(n_14),
.Y(n_310)
);

OA21x2_ASAP7_75t_L g311 ( 
.A1(n_310),
.A2(n_10),
.B(n_15),
.Y(n_311)
);

BUFx24_ASAP7_75t_SL g312 ( 
.A(n_311),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_312),
.B(n_309),
.Y(n_313)
);


endmodule