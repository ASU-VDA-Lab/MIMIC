module fake_jpeg_17068_n_313 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_313);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_313;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_145;
wire n_20;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

BUFx4f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx8_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx4f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_15),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_27),
.Y(n_37)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_29),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_17),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_51),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_49),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_32),
.B(n_31),
.Y(n_51)
);

A2O1A1Ixp33_ASAP7_75t_L g52 ( 
.A1(n_37),
.A2(n_30),
.B(n_29),
.C(n_21),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_52),
.B(n_21),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_35),
.A2(n_30),
.B1(n_26),
.B2(n_27),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_53),
.A2(n_35),
.B1(n_30),
.B2(n_34),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_56),
.A2(n_33),
.B1(n_39),
.B2(n_25),
.Y(n_94)
);

AND2x2_ASAP7_75t_SL g57 ( 
.A(n_42),
.B(n_51),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_57),
.B(n_65),
.C(n_69),
.Y(n_89)
);

INVx2_ASAP7_75t_R g58 ( 
.A(n_52),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_58),
.A2(n_76),
.B(n_80),
.Y(n_91)
);

CKINVDCx12_ASAP7_75t_R g59 ( 
.A(n_55),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_59),
.B(n_63),
.Y(n_101)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_43),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_44),
.A2(n_35),
.B1(n_34),
.B2(n_32),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_64),
.A2(n_83),
.B1(n_48),
.B2(n_39),
.Y(n_93)
);

AND2x2_ASAP7_75t_SL g65 ( 
.A(n_46),
.B(n_54),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_66),
.Y(n_92)
);

AND2x2_ASAP7_75t_SL g69 ( 
.A(n_44),
.B(n_37),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_70),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_49),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_72),
.B(n_81),
.Y(n_98)
);

BUFx12_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_73),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_37),
.Y(n_75)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_75),
.Y(n_100)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx4_ASAP7_75t_SL g85 ( 
.A(n_77),
.Y(n_85)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_78),
.Y(n_104)
);

INVx13_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

INVx4_ASAP7_75t_SL g96 ( 
.A(n_79),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_41),
.A2(n_34),
.B1(n_35),
.B2(n_28),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_45),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_48),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_41),
.A2(n_33),
.B1(n_39),
.B2(n_28),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_50),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_84),
.B(n_102),
.Y(n_130)
);

AND2x2_ASAP7_75t_SL g86 ( 
.A(n_58),
.B(n_40),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_86),
.A2(n_69),
.B(n_65),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_61),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_90),
.B(n_97),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_93),
.A2(n_94),
.B1(n_95),
.B2(n_78),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_67),
.A2(n_39),
.B1(n_40),
.B2(n_38),
.Y(n_95)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_74),
.Y(n_99)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_99),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_57),
.B(n_36),
.C(n_40),
.Y(n_102)
);

INVx2_ASAP7_75t_SL g103 ( 
.A(n_63),
.Y(n_103)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_103),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_67),
.B(n_50),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_110),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_66),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_107),
.B(n_77),
.Y(n_118)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_60),
.Y(n_108)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_108),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_67),
.B(n_40),
.Y(n_110)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_68),
.Y(n_111)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_111),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_113),
.A2(n_115),
.B(n_117),
.Y(n_161)
);

BUFx12_ASAP7_75t_L g114 ( 
.A(n_106),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_114),
.B(n_122),
.Y(n_140)
);

AND2x2_ASAP7_75t_SL g115 ( 
.A(n_84),
.B(n_58),
.Y(n_115)
);

AO22x1_ASAP7_75t_L g116 ( 
.A1(n_86),
.A2(n_62),
.B1(n_65),
.B2(n_69),
.Y(n_116)
);

AO21x2_ASAP7_75t_SL g150 ( 
.A1(n_116),
.A2(n_102),
.B(n_38),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_91),
.A2(n_76),
.B(n_72),
.Y(n_117)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_118),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_86),
.A2(n_62),
.B(n_71),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_119),
.A2(n_121),
.B(n_23),
.Y(n_165)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_106),
.Y(n_120)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_120),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_91),
.A2(n_71),
.B(n_80),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_104),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_123),
.B(n_136),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_99),
.A2(n_74),
.B1(n_33),
.B2(n_81),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_125),
.A2(n_103),
.B1(n_85),
.B2(n_111),
.Y(n_157)
);

INVx13_ASAP7_75t_L g126 ( 
.A(n_96),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_126),
.B(n_36),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_105),
.A2(n_64),
.B1(n_33),
.B2(n_70),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_129),
.A2(n_95),
.B1(n_110),
.B2(n_93),
.Y(n_145)
);

BUFx2_ASAP7_75t_SL g131 ( 
.A(n_96),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_131),
.Y(n_142)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_108),
.Y(n_132)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_132),
.Y(n_141)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_97),
.Y(n_133)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_133),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_135),
.A2(n_127),
.B1(n_113),
.B2(n_139),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_98),
.B(n_73),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_100),
.B(n_73),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_137),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_101),
.B(n_73),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_138),
.Y(n_159)
);

INVx2_ASAP7_75t_SL g139 ( 
.A(n_107),
.Y(n_139)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_139),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_145),
.B(n_124),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_146),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_115),
.B(n_89),
.Y(n_147)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_147),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_130),
.B(n_89),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_149),
.B(n_152),
.C(n_166),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_150),
.A2(n_160),
.B1(n_163),
.B2(n_126),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_115),
.B(n_134),
.Y(n_151)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_151),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_130),
.B(n_87),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_135),
.A2(n_87),
.B1(n_109),
.B2(n_88),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_154),
.A2(n_156),
.B1(n_157),
.B2(n_162),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_134),
.A2(n_121),
.B1(n_129),
.B2(n_116),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_114),
.B(n_103),
.Y(n_158)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_158),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_117),
.A2(n_85),
.B1(n_109),
.B2(n_25),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_119),
.A2(n_92),
.B1(n_20),
.B2(n_24),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_165),
.B(n_172),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_116),
.B(n_36),
.C(n_38),
.Y(n_166)
);

INVx2_ASAP7_75t_SL g167 ( 
.A(n_128),
.Y(n_167)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_167),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_133),
.B(n_19),
.Y(n_168)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_168),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_122),
.B(n_112),
.Y(n_169)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_169),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_112),
.B(n_36),
.C(n_38),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_170),
.B(n_68),
.C(n_22),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_127),
.A2(n_20),
.B1(n_24),
.B2(n_18),
.Y(n_171)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_171),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_120),
.A2(n_22),
.B(n_19),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_153),
.B(n_114),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_173),
.B(n_182),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_140),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_174),
.B(n_179),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_175),
.A2(n_164),
.B1(n_165),
.B2(n_170),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_151),
.B(n_139),
.Y(n_176)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_176),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_169),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_141),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_155),
.B(n_114),
.Y(n_184)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_184),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_148),
.B(n_124),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_187),
.B(n_190),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_159),
.B(n_132),
.Y(n_190)
);

NAND3xp33_ASAP7_75t_L g192 ( 
.A(n_147),
.B(n_18),
.C(n_22),
.Y(n_192)
);

NAND3xp33_ASAP7_75t_L g220 ( 
.A(n_192),
.B(n_12),
.C(n_14),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_144),
.B(n_128),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_193),
.B(n_164),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_194),
.A2(n_160),
.B1(n_166),
.B2(n_150),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_149),
.B(n_152),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_195),
.B(n_197),
.C(n_199),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_143),
.B(n_22),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_196),
.B(n_203),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_156),
.B(n_18),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_167),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_200),
.Y(n_210)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_167),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_201),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_161),
.B(n_68),
.C(n_18),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_202),
.B(n_172),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_143),
.B(n_0),
.Y(n_203)
);

OAI32xp33_ASAP7_75t_L g204 ( 
.A1(n_176),
.A2(n_150),
.A3(n_161),
.B1(n_145),
.B2(n_154),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_204),
.B(n_216),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_183),
.B(n_150),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_206),
.A2(n_212),
.B(n_226),
.Y(n_247)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_207),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_188),
.B(n_168),
.Y(n_209)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_209),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_185),
.Y(n_214)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_214),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_215),
.B(n_23),
.C(n_7),
.Y(n_245)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_185),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_189),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_217),
.B(n_220),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_221),
.A2(n_178),
.B1(n_202),
.B2(n_191),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_195),
.B(n_191),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_222),
.B(n_196),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_223),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_188),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_225),
.A2(n_203),
.B(n_186),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_180),
.B(n_141),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_226),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_194),
.A2(n_142),
.B1(n_79),
.B2(n_0),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_227),
.A2(n_198),
.B1(n_186),
.B2(n_181),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_228),
.A2(n_242),
.B1(n_207),
.B2(n_7),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_222),
.B(n_199),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_229),
.B(n_235),
.Y(n_262)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_230),
.Y(n_261)
);

MAJx2_ASAP7_75t_L g231 ( 
.A(n_204),
.B(n_178),
.C(n_183),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_231),
.B(n_237),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_232),
.A2(n_208),
.B1(n_227),
.B2(n_205),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_224),
.B(n_197),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_236),
.B(n_239),
.C(n_241),
.Y(n_252)
);

XNOR2x1_ASAP7_75t_SL g237 ( 
.A(n_206),
.B(n_180),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_224),
.B(n_177),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_215),
.B(n_15),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_206),
.A2(n_7),
.B(n_14),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_245),
.B(n_213),
.C(n_205),
.Y(n_253)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_247),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_240),
.B(n_210),
.Y(n_248)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_248),
.Y(n_266)
);

BUFx24_ASAP7_75t_SL g249 ( 
.A(n_239),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_249),
.B(n_253),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_246),
.B(n_218),
.Y(n_250)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_250),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_238),
.B(n_211),
.Y(n_251)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_251),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_234),
.A2(n_217),
.B1(n_209),
.B2(n_216),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_254),
.A2(n_257),
.B1(n_241),
.B2(n_236),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_233),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_256),
.B(n_258),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_244),
.A2(n_237),
.B1(n_231),
.B2(n_247),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_243),
.B(n_219),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_259),
.B(n_242),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_260),
.B(n_245),
.C(n_228),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_262),
.B(n_235),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_265),
.B(n_272),
.Y(n_282)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_269),
.Y(n_279)
);

OR2x2_ASAP7_75t_L g284 ( 
.A(n_270),
.B(n_271),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_261),
.B(n_253),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_254),
.B(n_229),
.Y(n_273)
);

OR2x2_ASAP7_75t_L g288 ( 
.A(n_273),
.B(n_252),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_263),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_274),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_23),
.C(n_1),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_275),
.B(n_276),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_252),
.B(n_2),
.C(n_3),
.Y(n_276)
);

BUFx24_ASAP7_75t_SL g278 ( 
.A(n_266),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_278),
.B(n_286),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_277),
.B(n_257),
.Y(n_280)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_280),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_281),
.A2(n_272),
.B1(n_276),
.B2(n_275),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_267),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_283),
.B(n_287),
.Y(n_291)
);

BUFx24_ASAP7_75t_SL g286 ( 
.A(n_268),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_270),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_288),
.B(n_255),
.Y(n_294)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_290),
.Y(n_299)
);

NOR2xp67_ASAP7_75t_L g292 ( 
.A(n_284),
.B(n_255),
.Y(n_292)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_292),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_282),
.B(n_264),
.C(n_265),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_293),
.B(n_295),
.Y(n_298)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_294),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_279),
.A2(n_4),
.B(n_5),
.Y(n_295)
);

NOR2xp67_ASAP7_75t_SL g296 ( 
.A(n_285),
.B(n_6),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_296),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_300),
.B(n_291),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g303 ( 
.A(n_289),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_303),
.B(n_302),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_304),
.A2(n_305),
.B1(n_306),
.B2(n_299),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_301),
.A2(n_292),
.B(n_297),
.Y(n_306)
);

NAND3xp33_ASAP7_75t_L g308 ( 
.A(n_307),
.B(n_298),
.C(n_303),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_308),
.A2(n_8),
.B(n_11),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_309),
.B(n_13),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_310),
.B(n_11),
.C(n_12),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_311),
.B(n_12),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_312),
.B(n_13),
.Y(n_313)
);


endmodule