module fake_jpeg_24439_n_281 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_281);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_281;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx5_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx24_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

BUFx24_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_32),
.Y(n_49)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_35),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_18),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_37),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_18),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_38),
.A2(n_14),
.B1(n_29),
.B2(n_15),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_36),
.B(n_25),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_48),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_36),
.B(n_24),
.Y(n_45)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_38),
.A2(n_23),
.B1(n_29),
.B2(n_15),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_46),
.A2(n_33),
.B1(n_19),
.B2(n_28),
.Y(n_74)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_25),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_50),
.B(n_37),
.Y(n_75)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_30),
.A2(n_22),
.B1(n_14),
.B2(n_20),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_53),
.A2(n_56),
.B1(n_33),
.B2(n_34),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_30),
.A2(n_22),
.B1(n_20),
.B2(n_29),
.Y(n_56)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

INVxp33_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_37),
.B(n_27),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_59),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_55),
.A2(n_30),
.B1(n_19),
.B2(n_28),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_61),
.B(n_69),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_40),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_63),
.B(n_67),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_66),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_38),
.Y(n_67)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_73),
.Y(n_88)
);

OA22x2_ASAP7_75t_L g72 ( 
.A1(n_49),
.A2(n_32),
.B1(n_31),
.B2(n_34),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_72),
.A2(n_74),
.B1(n_76),
.B2(n_79),
.Y(n_82)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_47),
.A2(n_27),
.B1(n_26),
.B2(n_24),
.Y(n_76)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_47),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_41),
.A2(n_21),
.B1(n_16),
.B2(n_26),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_81),
.A2(n_56),
.B1(n_53),
.B2(n_55),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_48),
.C(n_49),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_83),
.B(n_89),
.C(n_98),
.Y(n_109)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_85),
.B(n_95),
.Y(n_114)
);

AND2x4_ASAP7_75t_SL g86 ( 
.A(n_75),
.B(n_51),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_86),
.A2(n_102),
.B(n_72),
.Y(n_115)
);

MAJx2_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_35),
.C(n_39),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_91),
.A2(n_103),
.B1(n_71),
.B2(n_54),
.Y(n_112)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_67),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_92),
.B(n_94),
.Y(n_111)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_93),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_68),
.B(n_52),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_66),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_68),
.B(n_62),
.Y(n_97)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_79),
.B(n_35),
.C(n_39),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_62),
.B(n_59),
.Y(n_99)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_99),
.Y(n_110)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_74),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_104),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_72),
.B(n_55),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_61),
.A2(n_44),
.B1(n_45),
.B2(n_58),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_100),
.A2(n_64),
.B1(n_70),
.B2(n_81),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_106),
.A2(n_99),
.B1(n_102),
.B2(n_44),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_95),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_107),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_112),
.A2(n_98),
.B1(n_89),
.B2(n_82),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_93),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_113),
.B(n_116),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_115),
.A2(n_120),
.B(n_122),
.Y(n_134)
);

INVx2_ASAP7_75t_SL g116 ( 
.A(n_85),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_88),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_117),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_88),
.Y(n_118)
);

BUFx24_ASAP7_75t_SL g137 ( 
.A(n_118),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_94),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_119),
.Y(n_141)
);

A2O1A1Ixp33_ASAP7_75t_SL g120 ( 
.A1(n_91),
.A2(n_72),
.B(n_31),
.C(n_34),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_84),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_121),
.B(n_123),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_86),
.A2(n_44),
.B(n_72),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_84),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_70),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_124),
.B(n_35),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_103),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_126),
.Y(n_132)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_101),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_127),
.B(n_104),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_114),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_128),
.B(n_140),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_109),
.B(n_83),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_129),
.B(n_130),
.C(n_133),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_109),
.B(n_86),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_127),
.B(n_87),
.C(n_92),
.Y(n_133)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_116),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_135),
.B(n_144),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_124),
.B(n_86),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_138),
.B(n_110),
.C(n_105),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_120),
.A2(n_90),
.B1(n_87),
.B2(n_97),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_139),
.A2(n_146),
.B1(n_105),
.B2(n_110),
.Y(n_161)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_125),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_142),
.A2(n_120),
.B1(n_122),
.B2(n_121),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_107),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_112),
.A2(n_89),
.B1(n_82),
.B2(n_102),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_145),
.A2(n_120),
.B1(n_123),
.B2(n_108),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_117),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_147),
.B(n_149),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_119),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_150),
.B(n_111),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_151),
.B(n_77),
.Y(n_162)
);

AO21x1_ASAP7_75t_L g154 ( 
.A1(n_139),
.A2(n_115),
.B(n_108),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_154),
.B(n_155),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_143),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_156),
.B(n_158),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_157),
.A2(n_168),
.B1(n_148),
.B2(n_128),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_159),
.B(n_169),
.C(n_173),
.Y(n_176)
);

XNOR2x1_ASAP7_75t_L g160 ( 
.A(n_130),
.B(n_120),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_160),
.B(n_163),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_161),
.A2(n_136),
.B1(n_54),
.B2(n_65),
.Y(n_194)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_162),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_129),
.B(n_39),
.Y(n_163)
);

OR2x2_ASAP7_75t_L g164 ( 
.A(n_141),
.B(n_116),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_164),
.B(n_171),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_140),
.B(n_96),
.Y(n_165)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_165),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_135),
.Y(n_166)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_166),
.Y(n_185)
);

A2O1A1Ixp33_ASAP7_75t_L g167 ( 
.A1(n_146),
.A2(n_16),
.B(n_21),
.C(n_77),
.Y(n_167)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_167),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_132),
.A2(n_96),
.B1(n_54),
.B2(n_73),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_138),
.B(n_80),
.Y(n_169)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_148),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_133),
.B(n_54),
.C(n_77),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_132),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_174),
.B(n_131),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_137),
.B(n_12),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_175),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_152),
.B(n_142),
.C(n_134),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_180),
.B(n_193),
.C(n_176),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_183),
.A2(n_187),
.B1(n_167),
.B2(n_153),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_172),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_186),
.B(n_197),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_157),
.A2(n_160),
.B1(n_134),
.B2(n_154),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_164),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_189),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_170),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_190),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_191),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_152),
.B(n_150),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_192),
.B(n_163),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_169),
.B(n_151),
.C(n_145),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_194),
.A2(n_195),
.B1(n_57),
.B2(n_43),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_174),
.A2(n_78),
.B1(n_65),
.B2(n_57),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_155),
.B(n_21),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_198),
.B(n_200),
.C(n_202),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_192),
.B(n_159),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_199),
.B(n_207),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_182),
.B(n_158),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_182),
.B(n_173),
.Y(n_202)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_203),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_180),
.B(n_65),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_204),
.B(n_179),
.C(n_181),
.Y(n_229)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_206),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_191),
.B(n_8),
.Y(n_209)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_209),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_181),
.B(n_16),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_211),
.B(n_212),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_176),
.B(n_31),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_194),
.B(n_195),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_213),
.B(n_186),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_183),
.A2(n_7),
.B1(n_13),
.B2(n_12),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_214),
.B(n_197),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_184),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_215),
.A2(n_196),
.B1(n_201),
.B2(n_178),
.Y(n_221)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_218),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_205),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_219),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_208),
.A2(n_184),
.B(n_188),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_220),
.B(n_222),
.Y(n_235)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_221),
.Y(n_241)
);

FAx1_ASAP7_75t_SL g222 ( 
.A(n_211),
.B(n_193),
.CI(n_187),
.CON(n_222),
.SN(n_222)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_210),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_226),
.B(n_227),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_204),
.B(n_185),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_228),
.B(n_202),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_229),
.B(n_231),
.C(n_6),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_198),
.B(n_188),
.C(n_178),
.Y(n_231)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_233),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_224),
.B(n_185),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_234),
.B(n_221),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_223),
.A2(n_207),
.B1(n_200),
.B2(n_199),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_236),
.A2(n_217),
.B1(n_225),
.B2(n_216),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_230),
.B(n_177),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_237),
.B(n_238),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_229),
.B(n_7),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_231),
.B(n_6),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_239),
.B(n_13),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_242),
.B(n_244),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_230),
.B(n_9),
.Y(n_244)
);

NOR2xp67_ASAP7_75t_SL g245 ( 
.A(n_222),
.B(n_9),
.Y(n_245)
);

MAJx2_ASAP7_75t_L g247 ( 
.A(n_245),
.B(n_13),
.C(n_12),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_243),
.B(n_220),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_246),
.B(n_249),
.Y(n_259)
);

OAI21xp33_ASAP7_75t_L g258 ( 
.A1(n_247),
.A2(n_10),
.B(n_1),
.Y(n_258)
);

BUFx24_ASAP7_75t_SL g248 ( 
.A(n_244),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_248),
.B(n_238),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_250),
.B(n_251),
.Y(n_257)
);

INVx11_ASAP7_75t_L g251 ( 
.A(n_239),
.Y(n_251)
);

OR2x2_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_222),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_253),
.B(n_241),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_256),
.B(n_57),
.C(n_1),
.Y(n_265)
);

OA21x2_ASAP7_75t_SL g269 ( 
.A1(n_258),
.A2(n_259),
.B(n_1),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_SL g260 ( 
.A(n_246),
.B(n_242),
.Y(n_260)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_260),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_255),
.A2(n_232),
.B(n_240),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_261),
.A2(n_253),
.B(n_254),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_262),
.B(n_0),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_263),
.A2(n_257),
.B(n_259),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_252),
.B(n_217),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_264),
.B(n_265),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_266),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_268),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_269),
.B(n_270),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_267),
.B(n_57),
.C(n_3),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_273),
.B(n_274),
.Y(n_276)
);

A2O1A1O1Ixp25_ASAP7_75t_L g277 ( 
.A1(n_272),
.A2(n_271),
.B(n_3),
.C(n_4),
.D(n_2),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_277),
.A2(n_275),
.B1(n_273),
.B2(n_4),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_278),
.B(n_276),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_279),
.B(n_3),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_280),
.B(n_4),
.Y(n_281)
);


endmodule