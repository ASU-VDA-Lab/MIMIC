module fake_jpeg_3500_n_437 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_437);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_437;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

INVx6_ASAP7_75t_SL g29 ( 
.A(n_5),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_12),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx16f_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_44),
.Y(n_109)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx4_ASAP7_75t_SL g92 ( 
.A(n_45),
.Y(n_92)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_47),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx4_ASAP7_75t_SL g96 ( 
.A(n_48),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_49),
.Y(n_107)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_51),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_52),
.Y(n_119)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_53),
.Y(n_128)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g124 ( 
.A(n_54),
.Y(n_124)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_55),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_21),
.B(n_0),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_56),
.B(n_59),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_57),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_58),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_23),
.B(n_0),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_60),
.Y(n_103)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_61),
.B(n_83),
.Y(n_87)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_62),
.Y(n_121)
);

BUFx24_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_64),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_65),
.Y(n_133)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_66),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_67),
.Y(n_102)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_17),
.Y(n_68)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_68),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_69),
.Y(n_122)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_17),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g130 ( 
.A(n_70),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_71),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g129 ( 
.A(n_72),
.Y(n_129)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_73),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_74),
.Y(n_120)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_75),
.Y(n_126)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_76),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_24),
.B(n_32),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_77),
.B(n_79),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_78),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_24),
.B(n_1),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_38),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_80),
.B(n_81),
.Y(n_90)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_41),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_82),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_25),
.B(n_32),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_43),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_84),
.B(n_17),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_38),
.Y(n_85)
);

AOI21xp33_ASAP7_75t_SL g99 ( 
.A1(n_85),
.A2(n_18),
.B(n_42),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_49),
.A2(n_40),
.B1(n_39),
.B2(n_43),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_88),
.A2(n_95),
.B1(n_98),
.B2(n_112),
.Y(n_156)
);

INVxp33_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_89),
.Y(n_164)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_94),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_47),
.A2(n_42),
.B1(n_37),
.B2(n_40),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_48),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_97),
.B(n_117),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_51),
.A2(n_40),
.B1(n_43),
.B2(n_27),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_99),
.A2(n_63),
.B(n_18),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_44),
.A2(n_42),
.B1(n_37),
.B2(n_40),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_48),
.A2(n_42),
.B1(n_37),
.B2(n_43),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_116),
.A2(n_96),
.B1(n_46),
.B2(n_76),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_73),
.B(n_31),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_75),
.B(n_31),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_118),
.B(n_67),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_78),
.B(n_25),
.C(n_26),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_131),
.B(n_37),
.Y(n_135)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_132),
.Y(n_134)
);

BUFx2_ASAP7_75t_L g189 ( 
.A(n_134),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_135),
.B(n_154),
.Y(n_185)
);

OAI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_98),
.A2(n_88),
.B1(n_95),
.B2(n_112),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_136),
.A2(n_140),
.B1(n_146),
.B2(n_168),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_90),
.B(n_81),
.Y(n_137)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_137),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g138 ( 
.A(n_124),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_138),
.Y(n_192)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_89),
.Y(n_139)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_139),
.Y(n_182)
);

OAI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_116),
.A2(n_55),
.B1(n_70),
.B2(n_85),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_90),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_141),
.B(n_143),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_142),
.B(n_122),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_86),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_128),
.Y(n_144)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_144),
.Y(n_193)
);

BUFx2_ASAP7_75t_L g145 ( 
.A(n_101),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_145),
.Y(n_191)
);

OAI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_110),
.A2(n_82),
.B1(n_74),
.B2(n_72),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_111),
.B(n_26),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_147),
.B(n_151),
.Y(n_187)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_91),
.Y(n_148)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_148),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_86),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_149),
.B(n_169),
.Y(n_204)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_107),
.Y(n_150)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_150),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_114),
.A2(n_33),
.B1(n_36),
.B2(n_20),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_151),
.A2(n_175),
.B(n_36),
.Y(n_184)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_103),
.Y(n_152)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_152),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_124),
.B(n_67),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_107),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_155),
.Y(n_206)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_113),
.Y(n_157)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_157),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_102),
.Y(n_158)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_158),
.Y(n_203)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_105),
.Y(n_159)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_159),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_126),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_160),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_108),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_162),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_105),
.B(n_68),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_163),
.B(n_167),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_87),
.A2(n_33),
.B1(n_27),
.B2(n_15),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_165),
.A2(n_166),
.B1(n_170),
.B2(n_178),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_93),
.A2(n_58),
.B1(n_71),
.B2(n_69),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_121),
.Y(n_167)
);

INVx11_ASAP7_75t_L g168 ( 
.A(n_104),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_115),
.Y(n_169)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_109),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_171),
.B(n_172),
.Y(n_180)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_109),
.Y(n_172)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_104),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_173),
.B(n_174),
.Y(n_196)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_93),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_96),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_176),
.B(n_50),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_100),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_177),
.B(n_37),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_120),
.A2(n_16),
.B1(n_20),
.B2(n_28),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_156),
.A2(n_123),
.B1(n_52),
.B2(n_57),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_181),
.A2(n_215),
.B1(n_162),
.B2(n_155),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_184),
.A2(n_1),
.B(n_2),
.Y(n_249)
);

AOI32xp33_ASAP7_75t_L g186 ( 
.A1(n_175),
.A2(n_92),
.A3(n_123),
.B1(n_35),
.B2(n_16),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_186),
.B(n_209),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_187),
.B(n_154),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_135),
.B(n_92),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_188),
.B(n_201),
.C(n_220),
.Y(n_225)
);

A2O1A1O1Ixp25_ASAP7_75t_L g194 ( 
.A1(n_135),
.A2(n_35),
.B(n_28),
.C(n_15),
.D(n_27),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_194),
.A2(n_198),
.B(n_148),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_153),
.B(n_133),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_195),
.B(n_211),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_139),
.A2(n_15),
.B(n_130),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_144),
.B(n_122),
.C(n_125),
.Y(n_201)
);

INVxp33_ASAP7_75t_L g255 ( 
.A(n_207),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_208),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_161),
.B(n_37),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_166),
.A2(n_66),
.B1(n_64),
.B2(n_65),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_210),
.A2(n_218),
.B1(n_221),
.B2(n_164),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_147),
.B(n_133),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_152),
.B(n_127),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_212),
.B(n_14),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_137),
.A2(n_108),
.B1(n_125),
.B2(n_119),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_216),
.B(n_176),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_137),
.A2(n_127),
.B1(n_106),
.B2(n_119),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_167),
.B(n_129),
.C(n_104),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_174),
.A2(n_106),
.B1(n_129),
.B2(n_42),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_187),
.B(n_169),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_222),
.B(n_231),
.Y(n_261)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_193),
.Y(n_224)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_224),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_226),
.A2(n_228),
.B1(n_238),
.B2(n_251),
.Y(n_271)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_227),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_181),
.A2(n_134),
.B1(n_163),
.B2(n_154),
.Y(n_228)
);

INVx3_ASAP7_75t_SL g229 ( 
.A(n_219),
.Y(n_229)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_229),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_204),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_232),
.B(n_247),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_188),
.B(n_163),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_233),
.B(n_242),
.C(n_246),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_214),
.Y(n_234)
);

INVx4_ASAP7_75t_L g262 ( 
.A(n_234),
.Y(n_262)
);

FAx1_ASAP7_75t_SL g235 ( 
.A(n_185),
.B(n_164),
.CI(n_145),
.CON(n_235),
.SN(n_235)
);

A2O1A1Ixp33_ASAP7_75t_L g293 ( 
.A1(n_235),
.A2(n_199),
.B(n_203),
.C(n_206),
.Y(n_293)
);

INVxp33_ASAP7_75t_L g279 ( 
.A(n_236),
.Y(n_279)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_193),
.Y(n_237)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_237),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_202),
.A2(n_185),
.B1(n_211),
.B2(n_210),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_219),
.Y(n_239)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_239),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_195),
.B(n_157),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_240),
.B(n_243),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_185),
.A2(n_171),
.B1(n_172),
.B2(n_173),
.Y(n_241)
);

AO21x1_ASAP7_75t_L g284 ( 
.A1(n_241),
.A2(n_200),
.B(n_196),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_217),
.B(n_168),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_179),
.B(n_158),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_216),
.B(n_150),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_244),
.B(n_252),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_245),
.A2(n_248),
.B(n_249),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_217),
.B(n_129),
.C(n_42),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_212),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_190),
.A2(n_18),
.B1(n_2),
.B2(n_3),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_214),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_250),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_213),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_183),
.B(n_2),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_254),
.B(n_205),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_189),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_256),
.B(n_259),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_184),
.A2(n_3),
.B(n_4),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_257),
.A2(n_194),
.B(n_198),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_190),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_258),
.A2(n_200),
.B1(n_221),
.B2(n_182),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_192),
.B(n_6),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_260),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_232),
.B(n_192),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_266),
.B(n_267),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_253),
.B(n_231),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_245),
.A2(n_186),
.B(n_180),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_269),
.A2(n_270),
.B(n_246),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_257),
.A2(n_182),
.B(n_183),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_272),
.A2(n_284),
.B(n_235),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_275),
.B(n_277),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_241),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_276),
.B(n_289),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_247),
.B(n_197),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_238),
.A2(n_218),
.B1(n_201),
.B2(n_215),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_283),
.A2(n_228),
.B1(n_227),
.B2(n_255),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_233),
.B(n_220),
.C(n_200),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_285),
.B(n_286),
.C(n_287),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_225),
.B(n_242),
.C(n_230),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_225),
.B(n_197),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_230),
.B(n_205),
.C(n_199),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_288),
.B(n_203),
.C(n_189),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_234),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_250),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_290),
.B(n_294),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_293),
.A2(n_249),
.B(n_255),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_254),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_295),
.A2(n_300),
.B1(n_302),
.B2(n_308),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_298),
.Y(n_334)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_273),
.Y(n_299)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_299),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_280),
.A2(n_226),
.B1(n_223),
.B2(n_251),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_280),
.A2(n_253),
.B1(n_224),
.B2(n_237),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_304),
.A2(n_311),
.B(n_293),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_277),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_305),
.B(n_306),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_268),
.B(n_275),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_268),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_307),
.B(n_310),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_283),
.A2(n_256),
.B1(n_206),
.B2(n_229),
.Y(n_308)
);

BUFx2_ASAP7_75t_L g310 ( 
.A(n_291),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_281),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_312),
.B(n_318),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_313),
.B(n_264),
.Y(n_327)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_273),
.Y(n_314)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_314),
.Y(n_341)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_282),
.Y(n_316)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_316),
.Y(n_344)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_282),
.Y(n_317)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_317),
.Y(n_346)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_288),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_287),
.B(n_235),
.C(n_189),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_319),
.B(n_322),
.C(n_260),
.Y(n_326)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_291),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_320),
.B(n_265),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_271),
.A2(n_229),
.B1(n_239),
.B2(n_191),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_321),
.A2(n_323),
.B1(n_281),
.B2(n_290),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_286),
.B(n_191),
.C(n_7),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_271),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_318),
.B(n_279),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_324),
.B(n_343),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_326),
.B(n_328),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_327),
.B(n_328),
.C(n_330),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_301),
.B(n_264),
.C(n_285),
.Y(n_328)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_329),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_301),
.B(n_261),
.C(n_294),
.Y(n_330)
);

AND2x6_ASAP7_75t_L g331 ( 
.A(n_309),
.B(n_269),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_331),
.A2(n_332),
.B1(n_342),
.B2(n_345),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_295),
.A2(n_276),
.B1(n_278),
.B2(n_261),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_319),
.B(n_304),
.C(n_313),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_335),
.B(n_337),
.C(n_348),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_336),
.B(n_296),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_322),
.B(n_263),
.C(n_270),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_297),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_305),
.A2(n_263),
.B1(n_274),
.B2(n_278),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_312),
.B(n_274),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_347),
.B(n_325),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_303),
.B(n_292),
.C(n_272),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_303),
.B(n_292),
.C(n_289),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_349),
.B(n_316),
.C(n_314),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_333),
.A2(n_307),
.B1(n_315),
.B2(n_297),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_350),
.A2(n_357),
.B1(n_310),
.B2(n_262),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_351),
.B(n_367),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_L g354 ( 
.A1(n_334),
.A2(n_315),
.B(n_311),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_SL g378 ( 
.A1(n_354),
.A2(n_355),
.B(n_336),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_L g355 ( 
.A1(n_332),
.A2(n_298),
.B(n_302),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_333),
.A2(n_308),
.B1(n_306),
.B2(n_300),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_338),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_SL g384 ( 
.A(n_358),
.B(n_265),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_345),
.A2(n_296),
.B1(n_321),
.B2(n_317),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_359),
.A2(n_370),
.B1(n_344),
.B2(n_341),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g360 ( 
.A(n_349),
.Y(n_360)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_360),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_361),
.B(n_363),
.Y(n_387)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_362),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_327),
.B(n_284),
.Y(n_363)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_339),
.Y(n_366)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_366),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_330),
.B(n_284),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g374 ( 
.A(n_368),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_335),
.B(n_340),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_369),
.B(n_326),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_342),
.A2(n_299),
.B1(n_323),
.B2(n_320),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_356),
.B(n_346),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_371),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_372),
.B(n_373),
.Y(n_398)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_370),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g376 ( 
.A1(n_354),
.A2(n_355),
.B(n_365),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_L g397 ( 
.A1(n_376),
.A2(n_364),
.B(n_352),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_378),
.B(n_361),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_379),
.A2(n_373),
.B1(n_376),
.B2(n_374),
.Y(n_394)
);

NAND4xp25_ASAP7_75t_L g380 ( 
.A(n_350),
.B(n_331),
.C(n_348),
.D(n_337),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_380),
.A2(n_357),
.B(n_368),
.Y(n_388)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_353),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_381),
.A2(n_384),
.B1(n_385),
.B2(n_359),
.Y(n_392)
);

AOI21x1_ASAP7_75t_L g386 ( 
.A1(n_367),
.A2(n_310),
.B(n_262),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_386),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_388),
.B(n_389),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_387),
.B(n_369),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_390),
.B(n_377),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_375),
.B(n_363),
.Y(n_391)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_391),
.Y(n_406)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_392),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_SL g393 ( 
.A1(n_380),
.A2(n_352),
.B(n_364),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_393),
.B(n_400),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_394),
.A2(n_397),
.B1(n_387),
.B2(n_383),
.Y(n_408)
);

BUFx24_ASAP7_75t_SL g395 ( 
.A(n_382),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_SL g402 ( 
.A(n_395),
.B(n_381),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_377),
.B(n_351),
.C(n_10),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_SL g421 ( 
.A(n_402),
.B(n_12),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_399),
.A2(n_379),
.B1(n_385),
.B2(n_378),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_403),
.B(n_408),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g404 ( 
.A(n_400),
.Y(n_404)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_404),
.Y(n_414)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_389),
.A2(n_371),
.B(n_386),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_L g419 ( 
.A1(n_405),
.A2(n_409),
.B(n_390),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_407),
.B(n_411),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g409 ( 
.A1(n_398),
.A2(n_9),
.B(n_10),
.Y(n_409)
);

INVx11_ASAP7_75t_L g411 ( 
.A(n_396),
.Y(n_411)
);

INVx6_ASAP7_75t_L g415 ( 
.A(n_410),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_415),
.B(n_407),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_406),
.B(n_396),
.Y(n_416)
);

OR2x2_ASAP7_75t_L g427 ( 
.A(n_416),
.B(n_417),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_412),
.B(n_391),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_419),
.Y(n_426)
);

OAI21xp33_ASAP7_75t_L g420 ( 
.A1(n_408),
.A2(n_11),
.B(n_12),
.Y(n_420)
);

A2O1A1Ixp33_ASAP7_75t_SL g428 ( 
.A1(n_420),
.A2(n_13),
.B(n_415),
.C(n_413),
.Y(n_428)
);

INVx11_ASAP7_75t_L g425 ( 
.A(n_421),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_418),
.A2(n_401),
.B1(n_411),
.B2(n_405),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_422),
.B(n_424),
.Y(n_430)
);

NOR3xp33_ASAP7_75t_L g431 ( 
.A(n_423),
.B(n_428),
.C(n_13),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_414),
.B(n_403),
.C(n_409),
.Y(n_424)
);

NAND2xp33_ASAP7_75t_SL g429 ( 
.A(n_426),
.B(n_420),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_SL g434 ( 
.A1(n_429),
.A2(n_432),
.B(n_425),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_431),
.B(n_422),
.C(n_428),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_427),
.B(n_13),
.Y(n_432)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_433),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_435),
.B(n_430),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_436),
.B(n_434),
.Y(n_437)
);


endmodule