module real_jpeg_15915_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_131;
wire n_47;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_13;
wire n_113;
wire n_155;
wire n_120;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_0),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_1),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_2),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_3),
.Y(n_60)
);

AND2x2_ASAP7_75t_SL g19 ( 
.A(n_4),
.B(n_20),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_4),
.B(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_4),
.B(n_59),
.Y(n_58)
);

AND2x4_ASAP7_75t_SL g62 ( 
.A(n_4),
.B(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_4),
.B(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_4),
.Y(n_119)
);

AND2x2_ASAP7_75t_SL g156 ( 
.A(n_4),
.B(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_5),
.B(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_6),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_6),
.Y(n_88)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_7),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_7),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_8),
.B(n_30),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_8),
.B(n_46),
.Y(n_45)
);

AND2x4_ASAP7_75t_SL g54 ( 
.A(n_8),
.B(n_55),
.Y(n_54)
);

AND2x4_ASAP7_75t_L g75 ( 
.A(n_8),
.B(n_76),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_8),
.B(n_88),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_8),
.B(n_27),
.Y(n_103)
);

NAND2x1p5_ASAP7_75t_L g123 ( 
.A(n_8),
.B(n_124),
.Y(n_123)
);

NAND2x1_ASAP7_75t_L g167 ( 
.A(n_8),
.B(n_168),
.Y(n_167)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_9),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g25 ( 
.A(n_10),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_10),
.B(n_72),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_10),
.B(n_91),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_10),
.B(n_133),
.Y(n_132)
);

BUFx8_ASAP7_75t_L g168 ( 
.A(n_11),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_143),
.Y(n_12)
);

HB1xp67_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_112),
.B(n_142),
.Y(n_14)
);

OAI21xp5_ASAP7_75t_SL g15 ( 
.A1(n_16),
.A2(n_84),
.B(n_111),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_49),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_17),
.B(n_49),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_34),
.C(n_42),
.Y(n_17)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_18),
.B(n_96),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_22),
.B1(n_32),
.B2(n_33),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_19),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_19),
.A2(n_32),
.B1(n_131),
.B2(n_135),
.Y(n_130)
);

O2A1O1Ixp33_ASAP7_75t_L g151 ( 
.A1(n_19),
.A2(n_94),
.B(n_103),
.C(n_132),
.Y(n_151)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_28),
.B2(n_29),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_24),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_24),
.B(n_28),
.C(n_32),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_26),
.Y(n_24)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_25),
.B(n_40),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g173 ( 
.A(n_25),
.B(n_174),
.Y(n_173)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_31),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_34),
.A2(n_42),
.B1(n_43),
.B2(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_34),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_34),
.A2(n_35),
.B(n_38),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_38),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_35),
.A2(n_44),
.B1(n_45),
.B2(n_48),
.Y(n_43)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_38),
.A2(n_39),
.B1(n_53),
.B2(n_54),
.Y(n_141)
);

INVx2_ASAP7_75t_SL g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g44 ( 
.A(n_45),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g64 ( 
.A1(n_45),
.A2(n_54),
.B(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_54),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_45),
.B(n_90),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_46),
.Y(n_172)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

XOR2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_68),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_50),
.B(n_69),
.C(n_83),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_61),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_52),
.A2(n_100),
.B(n_104),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_52),
.A2(n_62),
.B(n_67),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_58),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_58),
.A2(n_90),
.B1(n_92),
.B2(n_93),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_64),
.B1(n_66),
.B2(n_67),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_62),
.Y(n_66)
);

O2A1O1Ixp33_ASAP7_75t_SL g86 ( 
.A1(n_62),
.A2(n_87),
.B(n_89),
.C(n_94),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_62),
.B(n_87),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_62),
.A2(n_66),
.B1(n_87),
.B2(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_64),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_65),
.B(n_117),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_65),
.B(n_118),
.C(n_123),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_69),
.A2(n_70),
.B1(n_82),
.B2(n_83),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_73),
.B1(n_74),
.B2(n_81),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_71),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_71),
.B(n_75),
.C(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_78),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_77),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_77),
.Y(n_176)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_78),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_78),
.A2(n_139),
.B1(n_155),
.B2(n_161),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_98),
.B(n_110),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_95),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_95),
.Y(n_110)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_87),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_87),
.B(n_102),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_89),
.B(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_90),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_90),
.A2(n_92),
.B1(n_156),
.B2(n_160),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_97),
.B(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_97),
.B(n_106),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_105),
.B(n_109),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_101),
.B(n_102),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_101),
.B(n_102),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_102),
.A2(n_103),
.B1(n_132),
.B2(n_134),
.Y(n_131)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_114),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_113),
.B(n_114),
.Y(n_142)
);

XOR2x2_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_129),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_128),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_116),
.B(n_128),
.C(n_129),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_122),
.B1(n_123),
.B2(n_127),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_118),
.Y(n_127)
);

OR2x6_ASAP7_75t_SL g118 ( 
.A(n_119),
.B(n_120),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_SL g122 ( 
.A(n_123),
.Y(n_122)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_136),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_137),
.C(n_141),
.Y(n_148)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_131),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_132),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_138),
.B1(n_140),
.B2(n_141),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_179),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_145),
.B(n_146),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_162),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_149),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_154),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_155),
.Y(n_161)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_156),
.Y(n_160)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_163),
.B(n_178),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_170),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_166),
.B1(n_167),
.B2(n_169),
.Y(n_164)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_165),
.Y(n_169)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_173),
.B(n_177),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_171),
.B(n_173),
.Y(n_177)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);


endmodule