module fake_ariane_879_n_750 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_143, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_136, n_28, n_80, n_97, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_750);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_136;
input n_28;
input n_80;
input n_97;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_750;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_698;
wire n_695;
wire n_160;
wire n_180;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_176;
wire n_691;
wire n_404;
wire n_172;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_564;
wire n_610;
wire n_205;
wire n_341;
wire n_245;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_690;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_286;
wire n_443;
wire n_586;
wire n_686;
wire n_605;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_524;
wire n_391;
wire n_349;
wire n_634;
wire n_466;
wire n_346;
wire n_214;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_162;
wire n_264;
wire n_737;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_372;
wire n_377;
wire n_396;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_363;
wire n_720;
wire n_354;
wire n_725;
wire n_419;
wire n_151;
wire n_146;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_154;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_145;
wire n_193;
wire n_733;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_668;
wire n_339;
wire n_738;
wire n_672;
wire n_487;
wire n_740;
wire n_167;
wire n_422;
wire n_153;
wire n_648;
wire n_269;
wire n_597;
wire n_158;
wire n_259;
wire n_446;
wire n_553;
wire n_566;
wire n_578;
wire n_701;
wire n_625;
wire n_152;
wire n_405;
wire n_557;
wire n_169;
wire n_173;
wire n_242;
wire n_645;
wire n_309;
wire n_320;
wire n_331;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_166;
wire n_253;
wire n_561;
wire n_218;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_247;
wire n_569;
wire n_567;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_510;
wire n_256;
wire n_326;
wire n_681;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_689;
wire n_694;
wire n_282;
wire n_328;
wire n_368;
wire n_699;
wire n_590;
wire n_727;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_644;
wire n_536;
wire n_293;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_303;
wire n_671;
wire n_442;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_661;
wire n_488;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_163;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_149;
wire n_383;
wire n_623;
wire n_237;
wire n_175;
wire n_711;
wire n_453;
wire n_734;
wire n_491;
wire n_181;
wire n_723;
wire n_616;
wire n_617;
wire n_705;
wire n_630;
wire n_658;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_371;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_178;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_710;
wire n_249;
wire n_534;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_148;
wire n_652;
wire n_451;
wire n_745;
wire n_613;
wire n_475;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_716;
wire n_742;
wire n_182;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_577;
wire n_407;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_280;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_161;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_655;
wire n_540;
wire n_216;
wire n_544;
wire n_692;
wire n_599;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_389;
wire n_657;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_150;
wire n_375;
wire n_324;
wire n_585;
wire n_669;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_697;
wire n_622;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_156;
wire n_292;
wire n_174;
wire n_275;
wire n_704;
wire n_147;
wire n_204;
wire n_615;
wire n_521;
wire n_496;
wire n_739;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_428;
wire n_159;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_165;
wire n_317;
wire n_243;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_749;
wire n_289;
wire n_548;
wire n_542;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_157;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_425;
wire n_431;
wire n_508;
wire n_624;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_353;
wire n_736;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_558;
wire n_592;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_155;
wire n_573;
wire n_531;
wire n_675;

INVx1_ASAP7_75t_L g145 ( 
.A(n_4),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_133),
.Y(n_146)
);

INVx1_ASAP7_75t_SL g147 ( 
.A(n_102),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_67),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_6),
.Y(n_149)
);

INVx2_ASAP7_75t_SL g150 ( 
.A(n_141),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_24),
.Y(n_151)
);

INVx1_ASAP7_75t_SL g152 ( 
.A(n_66),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_106),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_3),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_70),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_131),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_135),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_39),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_127),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_49),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_89),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_108),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_63),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_105),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_33),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_4),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_103),
.Y(n_167)
);

OR2x2_ASAP7_75t_L g168 ( 
.A(n_76),
.B(n_12),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_130),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_14),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_114),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_60),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_136),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_129),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_54),
.Y(n_175)
);

BUFx10_ASAP7_75t_L g176 ( 
.A(n_10),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_43),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_93),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_26),
.Y(n_179)
);

BUFx2_ASAP7_75t_L g180 ( 
.A(n_71),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_74),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_132),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_47),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_92),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_17),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_53),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_137),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_35),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_113),
.Y(n_189)
);

NOR2xp67_ASAP7_75t_L g190 ( 
.A(n_25),
.B(n_88),
.Y(n_190)
);

INVx2_ASAP7_75t_SL g191 ( 
.A(n_128),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_101),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_144),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_134),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_96),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_3),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_176),
.B(n_0),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_196),
.Y(n_198)
);

AND2x6_ASAP7_75t_L g199 ( 
.A(n_192),
.B(n_18),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_180),
.B(n_0),
.Y(n_200)
);

BUFx2_ASAP7_75t_L g201 ( 
.A(n_185),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_173),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_173),
.Y(n_203)
);

OAI22x1_ASAP7_75t_R g204 ( 
.A1(n_154),
.A2(n_1),
.B1(n_2),
.B2(n_5),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_146),
.B(n_1),
.Y(n_205)
);

INVx2_ASAP7_75t_SL g206 ( 
.A(n_176),
.Y(n_206)
);

AOI22x1_ASAP7_75t_SL g207 ( 
.A1(n_154),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_151),
.B(n_7),
.Y(n_208)
);

INVx5_ASAP7_75t_L g209 ( 
.A(n_173),
.Y(n_209)
);

BUFx12f_ASAP7_75t_L g210 ( 
.A(n_150),
.Y(n_210)
);

OAI22x1_ASAP7_75t_L g211 ( 
.A1(n_145),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_211)
);

BUFx12f_ASAP7_75t_L g212 ( 
.A(n_191),
.Y(n_212)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_196),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_149),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_163),
.B(n_8),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_167),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_166),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_173),
.Y(n_218)
);

INVxp67_ASAP7_75t_SL g219 ( 
.A(n_196),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_194),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_148),
.B(n_11),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_196),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_170),
.Y(n_223)
);

OA21x2_ASAP7_75t_L g224 ( 
.A1(n_155),
.A2(n_12),
.B(n_13),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g225 ( 
.A(n_170),
.Y(n_225)
);

AND2x4_ASAP7_75t_L g226 ( 
.A(n_148),
.B(n_13),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_156),
.Y(n_227)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_186),
.Y(n_228)
);

BUFx12f_ASAP7_75t_L g229 ( 
.A(n_153),
.Y(n_229)
);

AND2x4_ASAP7_75t_L g230 ( 
.A(n_186),
.B(n_14),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_192),
.Y(n_231)
);

INVx5_ASAP7_75t_L g232 ( 
.A(n_190),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_167),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_157),
.Y(n_234)
);

INVx5_ASAP7_75t_L g235 ( 
.A(n_159),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_158),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_216),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_213),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_216),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_219),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_214),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_228),
.B(n_169),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_234),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_233),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_229),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_234),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_R g247 ( 
.A(n_229),
.B(n_195),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_210),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_210),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_223),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_217),
.Y(n_251)
);

OAI21x1_ASAP7_75t_L g252 ( 
.A1(n_227),
.A2(n_175),
.B(n_189),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_212),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_212),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_201),
.Y(n_255)
);

INVx5_ASAP7_75t_L g256 ( 
.A(n_199),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_202),
.Y(n_257)
);

NAND2xp33_ASAP7_75t_R g258 ( 
.A(n_225),
.B(n_160),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_235),
.Y(n_259)
);

INVxp67_ASAP7_75t_SL g260 ( 
.A(n_228),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_235),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_206),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_202),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_235),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_206),
.B(n_147),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_213),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_235),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_213),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_235),
.Y(n_269)
);

OAI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_215),
.A2(n_220),
.B1(n_200),
.B2(n_208),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_R g271 ( 
.A(n_221),
.B(n_161),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_232),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_232),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_232),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_232),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_197),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_236),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_232),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_236),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_236),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_236),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_202),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_255),
.B(n_226),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_270),
.B(n_226),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_241),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_251),
.Y(n_286)
);

AO221x1_ASAP7_75t_L g287 ( 
.A1(n_276),
.A2(n_211),
.B1(n_204),
.B2(n_215),
.C(n_207),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_271),
.B(n_226),
.Y(n_288)
);

AND2x4_ASAP7_75t_L g289 ( 
.A(n_265),
.B(n_230),
.Y(n_289)
);

NOR2xp67_ASAP7_75t_L g290 ( 
.A(n_243),
.B(n_209),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_240),
.B(n_230),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_279),
.B(n_230),
.Y(n_292)
);

NOR2xp67_ASAP7_75t_L g293 ( 
.A(n_246),
.B(n_209),
.Y(n_293)
);

BUFx2_ASAP7_75t_L g294 ( 
.A(n_239),
.Y(n_294)
);

BUFx6f_ASAP7_75t_SL g295 ( 
.A(n_245),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_266),
.Y(n_296)
);

NOR2xp67_ASAP7_75t_L g297 ( 
.A(n_248),
.B(n_249),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_238),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_262),
.B(n_200),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_268),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_242),
.B(n_205),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_272),
.B(n_231),
.Y(n_302)
);

NOR3xp33_ASAP7_75t_L g303 ( 
.A(n_277),
.B(n_168),
.C(n_177),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_273),
.B(n_231),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_274),
.B(n_231),
.Y(n_305)
);

NAND3xp33_ASAP7_75t_L g306 ( 
.A(n_258),
.B(n_231),
.C(n_224),
.Y(n_306)
);

NAND2xp33_ASAP7_75t_L g307 ( 
.A(n_256),
.B(n_199),
.Y(n_307)
);

NAND2xp33_ASAP7_75t_L g308 ( 
.A(n_256),
.B(n_199),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_253),
.B(n_198),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_275),
.B(n_198),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_278),
.B(n_280),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_281),
.B(n_222),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_252),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_257),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_257),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_257),
.Y(n_316)
);

AO221x1_ASAP7_75t_L g317 ( 
.A1(n_257),
.A2(n_211),
.B1(n_172),
.B2(n_174),
.C(n_171),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_282),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_259),
.B(n_222),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_263),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_263),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_263),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_261),
.B(n_209),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_264),
.B(n_209),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_267),
.B(n_209),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_263),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_254),
.B(n_224),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_269),
.B(n_152),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_282),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_256),
.B(n_202),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_282),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_256),
.B(n_162),
.Y(n_332)
);

NOR2xp67_ASAP7_75t_L g333 ( 
.A(n_282),
.B(n_164),
.Y(n_333)
);

INVx4_ASAP7_75t_L g334 ( 
.A(n_247),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_244),
.B(n_203),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_250),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_237),
.B(n_203),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_241),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_260),
.B(n_203),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_241),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_238),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_260),
.B(n_203),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_260),
.B(n_218),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_241),
.Y(n_344)
);

BUFx6f_ASAP7_75t_SL g345 ( 
.A(n_245),
.Y(n_345)
);

HB1xp67_ASAP7_75t_L g346 ( 
.A(n_289),
.Y(n_346)
);

BUFx3_ASAP7_75t_L g347 ( 
.A(n_294),
.Y(n_347)
);

INVx4_ASAP7_75t_L g348 ( 
.A(n_334),
.Y(n_348)
);

OAI22xp33_ASAP7_75t_L g349 ( 
.A1(n_284),
.A2(n_224),
.B1(n_183),
.B2(n_193),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_284),
.A2(n_182),
.B1(n_178),
.B2(n_188),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_289),
.B(n_283),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_285),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_286),
.Y(n_353)
);

OAI21xp33_ASAP7_75t_L g354 ( 
.A1(n_301),
.A2(n_187),
.B(n_184),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_300),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_301),
.B(n_165),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_288),
.B(n_179),
.Y(n_357)
);

AND2x6_ASAP7_75t_SL g358 ( 
.A(n_336),
.B(n_299),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_337),
.B(n_181),
.Y(n_359)
);

OR2x2_ASAP7_75t_L g360 ( 
.A(n_335),
.B(n_15),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_288),
.B(n_334),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_313),
.A2(n_199),
.B(n_218),
.Y(n_362)
);

AND2x4_ASAP7_75t_L g363 ( 
.A(n_309),
.B(n_199),
.Y(n_363)
);

INVx2_ASAP7_75t_SL g364 ( 
.A(n_327),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_338),
.Y(n_365)
);

AND2x4_ASAP7_75t_L g366 ( 
.A(n_297),
.B(n_340),
.Y(n_366)
);

OR2x2_ASAP7_75t_L g367 ( 
.A(n_344),
.B(n_15),
.Y(n_367)
);

INVxp67_ASAP7_75t_SL g368 ( 
.A(n_315),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_296),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_345),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_303),
.A2(n_292),
.B1(n_291),
.B2(n_293),
.Y(n_371)
);

AND2x6_ASAP7_75t_SL g372 ( 
.A(n_287),
.B(n_16),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_303),
.A2(n_16),
.B1(n_17),
.B2(n_218),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_328),
.B(n_199),
.Y(n_374)
);

INVx3_ASAP7_75t_L g375 ( 
.A(n_318),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_290),
.A2(n_218),
.B1(n_20),
.B2(n_21),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_R g377 ( 
.A(n_295),
.B(n_345),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_311),
.B(n_143),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_341),
.B(n_19),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_339),
.A2(n_22),
.B(n_23),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_298),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_312),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_311),
.B(n_142),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_319),
.B(n_27),
.Y(n_384)
);

AOI22xp33_ASAP7_75t_L g385 ( 
.A1(n_317),
.A2(n_306),
.B1(n_302),
.B2(n_319),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_333),
.B(n_28),
.Y(n_386)
);

A2O1A1Ixp33_ASAP7_75t_L g387 ( 
.A1(n_342),
.A2(n_29),
.B(n_30),
.C(n_31),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_302),
.A2(n_32),
.B1(n_34),
.B2(n_36),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_343),
.B(n_37),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_L g390 ( 
.A1(n_323),
.A2(n_38),
.B(n_40),
.Y(n_390)
);

INVx4_ASAP7_75t_L g391 ( 
.A(n_295),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_310),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_304),
.B(n_41),
.Y(n_393)
);

NAND2x1_ASAP7_75t_L g394 ( 
.A(n_318),
.B(n_42),
.Y(n_394)
);

BUFx2_ASAP7_75t_L g395 ( 
.A(n_305),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_316),
.Y(n_396)
);

BUFx12f_ASAP7_75t_L g397 ( 
.A(n_315),
.Y(n_397)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_315),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_314),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g400 ( 
.A1(n_326),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_400)
);

INVx2_ASAP7_75t_SL g401 ( 
.A(n_320),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_329),
.B(n_48),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_321),
.B(n_50),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_331),
.B(n_307),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_330),
.Y(n_405)
);

INVx2_ASAP7_75t_SL g406 ( 
.A(n_315),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_332),
.B(n_51),
.Y(n_407)
);

BUFx2_ASAP7_75t_L g408 ( 
.A(n_322),
.Y(n_408)
);

OR2x2_ASAP7_75t_L g409 ( 
.A(n_322),
.B(n_140),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_307),
.B(n_52),
.Y(n_410)
);

INVx3_ASAP7_75t_L g411 ( 
.A(n_322),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_351),
.B(n_348),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_352),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_373),
.A2(n_332),
.B1(n_322),
.B2(n_308),
.Y(n_414)
);

BUFx2_ASAP7_75t_L g415 ( 
.A(n_347),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g416 ( 
.A1(n_374),
.A2(n_308),
.B(n_325),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_346),
.B(n_324),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_353),
.Y(n_418)
);

A2O1A1Ixp33_ASAP7_75t_L g419 ( 
.A1(n_378),
.A2(n_55),
.B(n_56),
.C(n_57),
.Y(n_419)
);

INVx2_ASAP7_75t_SL g420 ( 
.A(n_366),
.Y(n_420)
);

AOI221xp5_ASAP7_75t_L g421 ( 
.A1(n_373),
.A2(n_58),
.B1(n_59),
.B2(n_61),
.C(n_62),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_348),
.B(n_64),
.Y(n_422)
);

INVx6_ASAP7_75t_L g423 ( 
.A(n_391),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_365),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_356),
.B(n_65),
.Y(n_425)
);

INVx4_ASAP7_75t_L g426 ( 
.A(n_397),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_392),
.B(n_68),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_371),
.B(n_69),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_369),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_377),
.Y(n_430)
);

NOR2xp67_ASAP7_75t_SL g431 ( 
.A(n_367),
.B(n_391),
.Y(n_431)
);

O2A1O1Ixp33_ASAP7_75t_L g432 ( 
.A1(n_354),
.A2(n_72),
.B(n_73),
.C(n_75),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_361),
.B(n_395),
.Y(n_433)
);

INVx5_ASAP7_75t_L g434 ( 
.A(n_358),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_366),
.B(n_77),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_383),
.A2(n_78),
.B1(n_79),
.B2(n_80),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g437 ( 
.A1(n_404),
.A2(n_81),
.B(n_82),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_357),
.B(n_360),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_372),
.A2(n_83),
.B1(n_84),
.B2(n_85),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_359),
.B(n_86),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_370),
.B(n_87),
.Y(n_441)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_381),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_355),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g444 ( 
.A(n_364),
.B(n_90),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_350),
.B(n_91),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_382),
.Y(n_446)
);

INVxp67_ASAP7_75t_SL g447 ( 
.A(n_406),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_SL g448 ( 
.A(n_400),
.B(n_94),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_405),
.B(n_139),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_363),
.B(n_95),
.Y(n_450)
);

OAI21x1_ASAP7_75t_L g451 ( 
.A1(n_362),
.A2(n_97),
.B(n_98),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_408),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_396),
.Y(n_453)
);

INVx4_ASAP7_75t_L g454 ( 
.A(n_398),
.Y(n_454)
);

O2A1O1Ixp5_ASAP7_75t_L g455 ( 
.A1(n_384),
.A2(n_99),
.B(n_100),
.C(n_104),
.Y(n_455)
);

INVx2_ASAP7_75t_SL g456 ( 
.A(n_363),
.Y(n_456)
);

AOI21xp5_ASAP7_75t_L g457 ( 
.A1(n_404),
.A2(n_389),
.B(n_362),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_385),
.B(n_107),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_L g459 ( 
.A1(n_368),
.A2(n_109),
.B(n_110),
.Y(n_459)
);

AOI21xp5_ASAP7_75t_L g460 ( 
.A1(n_410),
.A2(n_111),
.B(n_112),
.Y(n_460)
);

HB1xp67_ASAP7_75t_L g461 ( 
.A(n_401),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_399),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_398),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_L g464 ( 
.A1(n_410),
.A2(n_115),
.B(n_116),
.Y(n_464)
);

O2A1O1Ixp33_ASAP7_75t_L g465 ( 
.A1(n_349),
.A2(n_400),
.B(n_375),
.C(n_407),
.Y(n_465)
);

AND2x4_ASAP7_75t_L g466 ( 
.A(n_411),
.B(n_117),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_443),
.Y(n_467)
);

INVx3_ASAP7_75t_L g468 ( 
.A(n_454),
.Y(n_468)
);

BUFx3_ASAP7_75t_L g469 ( 
.A(n_415),
.Y(n_469)
);

INVx2_ASAP7_75t_SL g470 ( 
.A(n_423),
.Y(n_470)
);

OR2x6_ASAP7_75t_L g471 ( 
.A(n_426),
.B(n_409),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_413),
.Y(n_472)
);

BUFx3_ASAP7_75t_L g473 ( 
.A(n_430),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_L g474 ( 
.A1(n_457),
.A2(n_402),
.B(n_393),
.Y(n_474)
);

BUFx2_ASAP7_75t_R g475 ( 
.A(n_452),
.Y(n_475)
);

BUFx3_ASAP7_75t_L g476 ( 
.A(n_423),
.Y(n_476)
);

AO21x2_ASAP7_75t_L g477 ( 
.A1(n_425),
.A2(n_402),
.B(n_403),
.Y(n_477)
);

INVxp33_ASAP7_75t_L g478 ( 
.A(n_433),
.Y(n_478)
);

CKINVDCx16_ASAP7_75t_R g479 ( 
.A(n_426),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_456),
.Y(n_480)
);

AND2x2_ASAP7_75t_SL g481 ( 
.A(n_448),
.B(n_388),
.Y(n_481)
);

OA21x2_ASAP7_75t_L g482 ( 
.A1(n_451),
.A2(n_403),
.B(n_379),
.Y(n_482)
);

BUFx12f_ASAP7_75t_L g483 ( 
.A(n_434),
.Y(n_483)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_454),
.Y(n_484)
);

INVx5_ASAP7_75t_L g485 ( 
.A(n_463),
.Y(n_485)
);

INVx3_ASAP7_75t_SL g486 ( 
.A(n_434),
.Y(n_486)
);

OAI21x1_ASAP7_75t_L g487 ( 
.A1(n_416),
.A2(n_394),
.B(n_390),
.Y(n_487)
);

NAND2x1p5_ASAP7_75t_L g488 ( 
.A(n_463),
.B(n_375),
.Y(n_488)
);

INVxp67_ASAP7_75t_L g489 ( 
.A(n_412),
.Y(n_489)
);

BUFx8_ASAP7_75t_L g490 ( 
.A(n_420),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_418),
.Y(n_491)
);

OA21x2_ASAP7_75t_L g492 ( 
.A1(n_437),
.A2(n_380),
.B(n_387),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_446),
.B(n_386),
.Y(n_493)
);

INVx2_ASAP7_75t_SL g494 ( 
.A(n_450),
.Y(n_494)
);

BUFx2_ASAP7_75t_L g495 ( 
.A(n_461),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_453),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_463),
.Y(n_497)
);

OAI21xp5_ASAP7_75t_L g498 ( 
.A1(n_465),
.A2(n_428),
.B(n_449),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_424),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_429),
.B(n_376),
.Y(n_500)
);

BUFx10_ASAP7_75t_L g501 ( 
.A(n_422),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_466),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_462),
.Y(n_503)
);

OR2x6_ASAP7_75t_L g504 ( 
.A(n_442),
.B(n_138),
.Y(n_504)
);

INVx2_ASAP7_75t_SL g505 ( 
.A(n_434),
.Y(n_505)
);

OAI21x1_ASAP7_75t_L g506 ( 
.A1(n_460),
.A2(n_118),
.B(n_119),
.Y(n_506)
);

AND2x4_ASAP7_75t_L g507 ( 
.A(n_466),
.B(n_120),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_438),
.B(n_121),
.Y(n_508)
);

BUFx12f_ASAP7_75t_L g509 ( 
.A(n_441),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_427),
.Y(n_510)
);

INVx3_ASAP7_75t_SL g511 ( 
.A(n_435),
.Y(n_511)
);

INVx2_ASAP7_75t_SL g512 ( 
.A(n_417),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_496),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_472),
.Y(n_514)
);

AOI21xp5_ASAP7_75t_L g515 ( 
.A1(n_481),
.A2(n_498),
.B(n_474),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_467),
.Y(n_516)
);

HB1xp67_ASAP7_75t_L g517 ( 
.A(n_495),
.Y(n_517)
);

HB1xp67_ASAP7_75t_L g518 ( 
.A(n_469),
.Y(n_518)
);

AO21x2_ASAP7_75t_L g519 ( 
.A1(n_477),
.A2(n_440),
.B(n_458),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_L g520 ( 
.A1(n_481),
.A2(n_414),
.B1(n_445),
.B2(n_439),
.Y(n_520)
);

INVx2_ASAP7_75t_SL g521 ( 
.A(n_476),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_467),
.Y(n_522)
);

OAI22xp33_ASAP7_75t_L g523 ( 
.A1(n_478),
.A2(n_448),
.B1(n_421),
.B2(n_436),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_496),
.Y(n_524)
);

CKINVDCx11_ASAP7_75t_R g525 ( 
.A(n_486),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_491),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_503),
.Y(n_527)
);

INVx3_ASAP7_75t_L g528 ( 
.A(n_507),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_499),
.Y(n_529)
);

AOI21x1_ASAP7_75t_L g530 ( 
.A1(n_482),
.A2(n_487),
.B(n_492),
.Y(n_530)
);

AOI22xp33_ASAP7_75t_SL g531 ( 
.A1(n_509),
.A2(n_439),
.B1(n_414),
.B2(n_444),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_502),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_493),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_507),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_489),
.A2(n_431),
.B1(n_447),
.B2(n_436),
.Y(n_535)
);

INVx1_ASAP7_75t_SL g536 ( 
.A(n_475),
.Y(n_536)
);

AOI22xp33_ASAP7_75t_L g537 ( 
.A1(n_509),
.A2(n_464),
.B1(n_459),
.B2(n_432),
.Y(n_537)
);

BUFx2_ASAP7_75t_L g538 ( 
.A(n_469),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_512),
.Y(n_539)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_507),
.Y(n_540)
);

BUFx4f_ASAP7_75t_SL g541 ( 
.A(n_483),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_502),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_500),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_510),
.Y(n_544)
);

INVx2_ASAP7_75t_SL g545 ( 
.A(n_476),
.Y(n_545)
);

CKINVDCx11_ASAP7_75t_R g546 ( 
.A(n_486),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_488),
.Y(n_547)
);

HB1xp67_ASAP7_75t_L g548 ( 
.A(n_480),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_488),
.Y(n_549)
);

AOI22xp33_ASAP7_75t_L g550 ( 
.A1(n_511),
.A2(n_419),
.B1(n_455),
.B2(n_124),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_506),
.Y(n_551)
);

AND2x4_ASAP7_75t_L g552 ( 
.A(n_485),
.B(n_122),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_506),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_538),
.B(n_478),
.Y(n_554)
);

AOI22xp33_ASAP7_75t_L g555 ( 
.A1(n_520),
.A2(n_511),
.B1(n_504),
.B2(n_501),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_527),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_538),
.B(n_489),
.Y(n_557)
);

BUFx2_ASAP7_75t_L g558 ( 
.A(n_518),
.Y(n_558)
);

AOI22xp33_ASAP7_75t_L g559 ( 
.A1(n_531),
.A2(n_504),
.B1(n_501),
.B2(n_494),
.Y(n_559)
);

NAND2xp33_ASAP7_75t_SL g560 ( 
.A(n_528),
.B(n_494),
.Y(n_560)
);

AO31x2_ASAP7_75t_L g561 ( 
.A1(n_515),
.A2(n_508),
.A3(n_477),
.B(n_482),
.Y(n_561)
);

CKINVDCx8_ASAP7_75t_R g562 ( 
.A(n_552),
.Y(n_562)
);

OR2x2_ASAP7_75t_L g563 ( 
.A(n_527),
.B(n_517),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_548),
.B(n_545),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_514),
.Y(n_565)
);

OAI21x1_ASAP7_75t_L g566 ( 
.A1(n_530),
.A2(n_487),
.B(n_492),
.Y(n_566)
);

AO31x2_ASAP7_75t_L g567 ( 
.A1(n_551),
.A2(n_492),
.A3(n_501),
.B(n_504),
.Y(n_567)
);

HB1xp67_ASAP7_75t_L g568 ( 
.A(n_551),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_526),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_513),
.Y(n_570)
);

HB1xp67_ASAP7_75t_L g571 ( 
.A(n_530),
.Y(n_571)
);

NOR3xp33_ASAP7_75t_SL g572 ( 
.A(n_523),
.B(n_479),
.C(n_473),
.Y(n_572)
);

NAND2xp33_ASAP7_75t_R g573 ( 
.A(n_552),
.B(n_471),
.Y(n_573)
);

CKINVDCx12_ASAP7_75t_R g574 ( 
.A(n_541),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_526),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_529),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_529),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_535),
.B(n_497),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_521),
.B(n_480),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_521),
.B(n_470),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_545),
.B(n_470),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_525),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_513),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_524),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_543),
.B(n_533),
.Y(n_585)
);

OR2x2_ASAP7_75t_L g586 ( 
.A(n_524),
.B(n_473),
.Y(n_586)
);

OR2x6_ASAP7_75t_L g587 ( 
.A(n_528),
.B(n_471),
.Y(n_587)
);

OAI22xp5_ASAP7_75t_L g588 ( 
.A1(n_528),
.A2(n_471),
.B1(n_484),
.B2(n_468),
.Y(n_588)
);

NAND2xp33_ASAP7_75t_R g589 ( 
.A(n_540),
.B(n_484),
.Y(n_589)
);

NOR3xp33_ASAP7_75t_SL g590 ( 
.A(n_534),
.B(n_483),
.C(n_490),
.Y(n_590)
);

INVxp67_ASAP7_75t_L g591 ( 
.A(n_543),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_546),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_544),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_544),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_539),
.B(n_505),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_516),
.Y(n_596)
);

NAND2xp33_ASAP7_75t_L g597 ( 
.A(n_540),
.B(n_468),
.Y(n_597)
);

BUFx10_ASAP7_75t_L g598 ( 
.A(n_552),
.Y(n_598)
);

INVx8_ASAP7_75t_L g599 ( 
.A(n_540),
.Y(n_599)
);

BUFx2_ASAP7_75t_L g600 ( 
.A(n_567),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_583),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_569),
.Y(n_602)
);

HB1xp67_ASAP7_75t_L g603 ( 
.A(n_563),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_584),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_575),
.B(n_519),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_570),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_576),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_577),
.B(n_593),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_594),
.Y(n_609)
);

BUFx6f_ASAP7_75t_L g610 ( 
.A(n_562),
.Y(n_610)
);

AOI21xp5_ASAP7_75t_SL g611 ( 
.A1(n_587),
.A2(n_519),
.B(n_578),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_565),
.B(n_542),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_596),
.Y(n_613)
);

OR2x2_ASAP7_75t_L g614 ( 
.A(n_591),
.B(n_533),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_557),
.B(n_542),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_568),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_568),
.Y(n_617)
);

INVxp67_ASAP7_75t_SL g618 ( 
.A(n_589),
.Y(n_618)
);

OR2x2_ASAP7_75t_L g619 ( 
.A(n_591),
.B(n_585),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_556),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_554),
.B(n_532),
.Y(n_621)
);

AND2x4_ASAP7_75t_L g622 ( 
.A(n_567),
.B(n_549),
.Y(n_622)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_567),
.B(n_564),
.Y(n_623)
);

BUFx6f_ASAP7_75t_L g624 ( 
.A(n_598),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_567),
.B(n_532),
.Y(n_625)
);

INVx3_ASAP7_75t_L g626 ( 
.A(n_599),
.Y(n_626)
);

AND2x4_ASAP7_75t_L g627 ( 
.A(n_585),
.B(n_547),
.Y(n_627)
);

BUFx2_ASAP7_75t_L g628 ( 
.A(n_571),
.Y(n_628)
);

OR2x2_ASAP7_75t_L g629 ( 
.A(n_558),
.B(n_522),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_574),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_571),
.B(n_547),
.Y(n_631)
);

INVx3_ASAP7_75t_SL g632 ( 
.A(n_582),
.Y(n_632)
);

AND2x4_ASAP7_75t_L g633 ( 
.A(n_572),
.B(n_522),
.Y(n_633)
);

INVx1_ASAP7_75t_SL g634 ( 
.A(n_586),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_623),
.B(n_561),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_606),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_603),
.B(n_579),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_601),
.Y(n_638)
);

OA21x2_ASAP7_75t_L g639 ( 
.A1(n_600),
.A2(n_566),
.B(n_553),
.Y(n_639)
);

OR2x2_ASAP7_75t_L g640 ( 
.A(n_623),
.B(n_619),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_610),
.B(n_572),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_631),
.B(n_561),
.Y(n_642)
);

HB1xp67_ASAP7_75t_L g643 ( 
.A(n_619),
.Y(n_643)
);

NAND2x1_ASAP7_75t_L g644 ( 
.A(n_616),
.B(n_553),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_615),
.B(n_581),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_615),
.B(n_614),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_608),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_606),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_608),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_601),
.Y(n_650)
);

AND2x4_ASAP7_75t_SL g651 ( 
.A(n_610),
.B(n_598),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_614),
.B(n_580),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_629),
.B(n_555),
.Y(n_653)
);

OAI221xp5_ASAP7_75t_SL g654 ( 
.A1(n_618),
.A2(n_555),
.B1(n_559),
.B2(n_537),
.C(n_550),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_602),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_631),
.B(n_561),
.Y(n_656)
);

BUFx2_ASAP7_75t_L g657 ( 
.A(n_628),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_604),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_604),
.Y(n_659)
);

BUFx2_ASAP7_75t_L g660 ( 
.A(n_628),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_629),
.B(n_634),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_643),
.B(n_617),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_638),
.Y(n_663)
);

BUFx3_ASAP7_75t_L g664 ( 
.A(n_657),
.Y(n_664)
);

OR2x2_ASAP7_75t_L g665 ( 
.A(n_640),
.B(n_616),
.Y(n_665)
);

HB1xp67_ASAP7_75t_L g666 ( 
.A(n_657),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_647),
.B(n_617),
.Y(n_667)
);

OR2x2_ASAP7_75t_L g668 ( 
.A(n_640),
.B(n_621),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_649),
.B(n_607),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_650),
.Y(n_670)
);

INVxp67_ASAP7_75t_SL g671 ( 
.A(n_660),
.Y(n_671)
);

INVx3_ASAP7_75t_L g672 ( 
.A(n_644),
.Y(n_672)
);

NAND4xp25_ASAP7_75t_L g673 ( 
.A(n_660),
.B(n_559),
.C(n_609),
.D(n_595),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_635),
.B(n_605),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_635),
.B(n_605),
.Y(n_675)
);

AND2x4_ASAP7_75t_L g676 ( 
.A(n_642),
.B(n_625),
.Y(n_676)
);

OR2x2_ASAP7_75t_L g677 ( 
.A(n_646),
.B(n_625),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_663),
.Y(n_678)
);

NAND4xp75_ASAP7_75t_L g679 ( 
.A(n_674),
.B(n_641),
.C(n_653),
.D(n_642),
.Y(n_679)
);

NOR2x1_ASAP7_75t_L g680 ( 
.A(n_664),
.B(n_637),
.Y(n_680)
);

OAI31xp33_ASAP7_75t_L g681 ( 
.A1(n_673),
.A2(n_654),
.A3(n_656),
.B(n_600),
.Y(n_681)
);

OAI32xp33_ASAP7_75t_L g682 ( 
.A1(n_665),
.A2(n_652),
.A3(n_645),
.B1(n_589),
.B2(n_655),
.Y(n_682)
);

INVx1_ASAP7_75t_SL g683 ( 
.A(n_668),
.Y(n_683)
);

INVx1_ASAP7_75t_SL g684 ( 
.A(n_662),
.Y(n_684)
);

AO221x1_ASAP7_75t_L g685 ( 
.A1(n_672),
.A2(n_610),
.B1(n_624),
.B2(n_638),
.C(n_659),
.Y(n_685)
);

OAI33xp33_ASAP7_75t_L g686 ( 
.A1(n_677),
.A2(n_661),
.A3(n_659),
.B1(n_630),
.B2(n_592),
.B3(n_670),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_664),
.B(n_656),
.Y(n_687)
);

NAND3xp33_ASAP7_75t_L g688 ( 
.A(n_666),
.B(n_671),
.C(n_672),
.Y(n_688)
);

AOI22xp5_ASAP7_75t_L g689 ( 
.A1(n_679),
.A2(n_676),
.B1(n_573),
.B2(n_675),
.Y(n_689)
);

INVx1_ASAP7_75t_SL g690 ( 
.A(n_684),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_687),
.B(n_667),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_686),
.B(n_632),
.Y(n_692)
);

OAI21xp33_ASAP7_75t_L g693 ( 
.A1(n_680),
.A2(n_688),
.B(n_682),
.Y(n_693)
);

OAI22xp33_ASAP7_75t_L g694 ( 
.A1(n_689),
.A2(n_681),
.B1(n_677),
.B2(n_683),
.Y(n_694)
);

AOI21xp5_ASAP7_75t_L g695 ( 
.A1(n_693),
.A2(n_681),
.B(n_685),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_690),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_691),
.Y(n_697)
);

OR2x2_ASAP7_75t_L g698 ( 
.A(n_692),
.B(n_678),
.Y(n_698)
);

AOI21xp5_ASAP7_75t_L g699 ( 
.A1(n_695),
.A2(n_694),
.B(n_698),
.Y(n_699)
);

OAI211xp5_ASAP7_75t_L g700 ( 
.A1(n_696),
.A2(n_630),
.B(n_536),
.C(n_672),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_697),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_696),
.B(n_669),
.Y(n_702)
);

AOI22xp5_ASAP7_75t_L g703 ( 
.A1(n_699),
.A2(n_676),
.B1(n_612),
.B2(n_675),
.Y(n_703)
);

OAI21xp33_ASAP7_75t_L g704 ( 
.A1(n_701),
.A2(n_702),
.B(n_700),
.Y(n_704)
);

OAI211xp5_ASAP7_75t_SL g705 ( 
.A1(n_699),
.A2(n_590),
.B(n_632),
.C(n_626),
.Y(n_705)
);

AOI22xp5_ASAP7_75t_L g706 ( 
.A1(n_703),
.A2(n_676),
.B1(n_612),
.B2(n_633),
.Y(n_706)
);

AOI321xp33_ASAP7_75t_L g707 ( 
.A1(n_704),
.A2(n_633),
.A3(n_627),
.B1(n_674),
.B2(n_622),
.C(n_588),
.Y(n_707)
);

AOI21xp5_ASAP7_75t_L g708 ( 
.A1(n_705),
.A2(n_644),
.B(n_669),
.Y(n_708)
);

OAI211xp5_ASAP7_75t_L g709 ( 
.A1(n_704),
.A2(n_626),
.B(n_590),
.C(n_667),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_709),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_707),
.Y(n_711)
);

NOR2x1_ASAP7_75t_L g712 ( 
.A(n_708),
.B(n_626),
.Y(n_712)
);

NOR2x1_ASAP7_75t_L g713 ( 
.A(n_706),
.B(n_610),
.Y(n_713)
);

NOR2x1_ASAP7_75t_L g714 ( 
.A(n_709),
.B(n_610),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_709),
.B(n_651),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_709),
.Y(n_716)
);

AOI22xp5_ASAP7_75t_L g717 ( 
.A1(n_709),
.A2(n_633),
.B1(n_560),
.B2(n_651),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_710),
.Y(n_718)
);

NOR2x1_ASAP7_75t_L g719 ( 
.A(n_716),
.B(n_497),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_711),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_715),
.B(n_712),
.Y(n_721)
);

AND2x2_ASAP7_75t_SL g722 ( 
.A(n_717),
.B(n_624),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_714),
.Y(n_723)
);

NAND3xp33_ASAP7_75t_L g724 ( 
.A(n_713),
.B(n_490),
.C(n_485),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_710),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_725),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_718),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_718),
.Y(n_728)
);

OAI31xp33_ASAP7_75t_SL g729 ( 
.A1(n_721),
.A2(n_490),
.A3(n_627),
.B(n_670),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_720),
.Y(n_730)
);

XNOR2xp5_ASAP7_75t_L g731 ( 
.A(n_723),
.B(n_719),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_722),
.Y(n_732)
);

AOI22xp5_ASAP7_75t_L g733 ( 
.A1(n_730),
.A2(n_724),
.B1(n_624),
.B2(n_597),
.Y(n_733)
);

AO22x2_ASAP7_75t_L g734 ( 
.A1(n_727),
.A2(n_658),
.B1(n_650),
.B2(n_627),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_730),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_728),
.Y(n_736)
);

OAI22xp5_ASAP7_75t_L g737 ( 
.A1(n_726),
.A2(n_624),
.B1(n_639),
.B2(n_658),
.Y(n_737)
);

OAI22xp5_ASAP7_75t_L g738 ( 
.A1(n_735),
.A2(n_732),
.B1(n_731),
.B2(n_729),
.Y(n_738)
);

OAI22xp33_ASAP7_75t_L g739 ( 
.A1(n_733),
.A2(n_736),
.B1(n_737),
.B2(n_734),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_735),
.B(n_639),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_735),
.B(n_624),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_740),
.Y(n_742)
);

AOI22xp5_ASAP7_75t_L g743 ( 
.A1(n_738),
.A2(n_639),
.B1(n_622),
.B2(n_599),
.Y(n_743)
);

AO211x2_ASAP7_75t_L g744 ( 
.A1(n_739),
.A2(n_620),
.B(n_485),
.C(n_611),
.Y(n_744)
);

AOI211xp5_ASAP7_75t_L g745 ( 
.A1(n_742),
.A2(n_741),
.B(n_497),
.C(n_611),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_743),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_746),
.B(n_744),
.Y(n_747)
);

AOI22xp5_ASAP7_75t_L g748 ( 
.A1(n_747),
.A2(n_745),
.B1(n_485),
.B2(n_622),
.Y(n_748)
);

AOI221xp5_ASAP7_75t_L g749 ( 
.A1(n_748),
.A2(n_648),
.B1(n_636),
.B2(n_599),
.C(n_613),
.Y(n_749)
);

AOI211xp5_ASAP7_75t_L g750 ( 
.A1(n_749),
.A2(n_123),
.B(n_125),
.C(n_126),
.Y(n_750)
);


endmodule