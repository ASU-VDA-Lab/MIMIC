module real_aes_8281_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_421;
wire n_555;
wire n_319;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_659;
wire n_547;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_417;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_505;
wire n_434;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g260 ( .A1(n_0), .A2(n_261), .B(n_262), .C(n_265), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_1), .B(n_249), .Y(n_266) );
INVx1_ASAP7_75t_L g105 ( .A(n_2), .Y(n_105) );
NAND2xp5_ASAP7_75t_SL g176 ( .A(n_3), .B(n_177), .Y(n_176) );
A2O1A1Ixp33_ASAP7_75t_L g539 ( .A1(n_4), .A2(n_138), .B(n_141), .C(n_540), .Y(n_539) );
AOI21xp5_ASAP7_75t_L g563 ( .A1(n_5), .A2(n_133), .B(n_564), .Y(n_563) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_6), .A2(n_133), .B(n_243), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_7), .B(n_249), .Y(n_570) );
AO21x2_ASAP7_75t_L g204 ( .A1(n_8), .A2(n_168), .B(n_205), .Y(n_204) );
AND2x6_ASAP7_75t_L g138 ( .A(n_9), .B(n_139), .Y(n_138) );
A2O1A1Ixp33_ASAP7_75t_L g221 ( .A1(n_10), .A2(n_138), .B(n_141), .C(n_222), .Y(n_221) );
INVx1_ASAP7_75t_L g508 ( .A(n_11), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_12), .B(n_111), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_12), .B(n_40), .Y(n_456) );
NAND2xp5_ASAP7_75t_SL g542 ( .A(n_13), .B(n_225), .Y(n_542) );
INVx1_ASAP7_75t_L g159 ( .A(n_14), .Y(n_159) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_15), .B(n_177), .Y(n_211) );
A2O1A1Ixp33_ASAP7_75t_L g525 ( .A1(n_16), .A2(n_178), .B(n_526), .C(n_528), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_17), .B(n_249), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_18), .B(n_153), .Y(n_499) );
A2O1A1Ixp33_ASAP7_75t_L g140 ( .A1(n_19), .A2(n_141), .B(n_144), .C(n_152), .Y(n_140) );
A2O1A1Ixp33_ASAP7_75t_L g515 ( .A1(n_20), .A2(n_213), .B(n_264), .C(n_516), .Y(n_515) );
NAND2xp5_ASAP7_75t_SL g559 ( .A(n_21), .B(n_225), .Y(n_559) );
AOI22xp5_ASAP7_75t_L g119 ( .A1(n_22), .A2(n_120), .B1(n_121), .B2(n_449), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g449 ( .A(n_22), .Y(n_449) );
NAND2xp5_ASAP7_75t_SL g481 ( .A(n_23), .B(n_225), .Y(n_481) );
CKINVDCx16_ASAP7_75t_R g555 ( .A(n_24), .Y(n_555) );
INVx1_ASAP7_75t_L g480 ( .A(n_25), .Y(n_480) );
A2O1A1Ixp33_ASAP7_75t_L g207 ( .A1(n_26), .A2(n_141), .B(n_152), .C(n_208), .Y(n_207) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_27), .Y(n_137) );
CKINVDCx20_ASAP7_75t_R g538 ( .A(n_28), .Y(n_538) );
INVx1_ASAP7_75t_L g496 ( .A(n_29), .Y(n_496) );
NAND2xp5_ASAP7_75t_SL g457 ( .A(n_30), .B(n_458), .Y(n_457) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_31), .A2(n_133), .B(n_258), .Y(n_257) );
INVx2_ASAP7_75t_L g136 ( .A(n_32), .Y(n_136) );
A2O1A1Ixp33_ASAP7_75t_L g189 ( .A1(n_33), .A2(n_181), .B(n_190), .C(n_192), .Y(n_189) );
CKINVDCx20_ASAP7_75t_R g545 ( .A(n_34), .Y(n_545) );
A2O1A1Ixp33_ASAP7_75t_L g566 ( .A1(n_35), .A2(n_264), .B(n_567), .C(n_569), .Y(n_566) );
INVxp67_ASAP7_75t_L g497 ( .A(n_36), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_37), .B(n_210), .Y(n_209) );
A2O1A1Ixp33_ASAP7_75t_L g478 ( .A1(n_38), .A2(n_141), .B(n_152), .C(n_479), .Y(n_478) );
CKINVDCx14_ASAP7_75t_R g565 ( .A(n_39), .Y(n_565) );
INVx1_ASAP7_75t_L g111 ( .A(n_40), .Y(n_111) );
A2O1A1Ixp33_ASAP7_75t_L g505 ( .A1(n_41), .A2(n_265), .B(n_506), .C(n_507), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_42), .B(n_132), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g227 ( .A(n_43), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_44), .B(n_177), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_45), .B(n_133), .Y(n_206) );
CKINVDCx20_ASAP7_75t_R g483 ( .A(n_46), .Y(n_483) );
CKINVDCx20_ASAP7_75t_R g493 ( .A(n_47), .Y(n_493) );
A2O1A1Ixp33_ASAP7_75t_L g233 ( .A1(n_48), .A2(n_181), .B(n_190), .C(n_234), .Y(n_233) );
INVx1_ASAP7_75t_L g263 ( .A(n_49), .Y(n_263) );
OAI22xp5_ASAP7_75t_L g121 ( .A1(n_50), .A2(n_122), .B1(n_123), .B2(n_448), .Y(n_121) );
CKINVDCx16_ASAP7_75t_R g122 ( .A(n_50), .Y(n_122) );
INVx1_ASAP7_75t_L g235 ( .A(n_51), .Y(n_235) );
INVx1_ASAP7_75t_L g514 ( .A(n_52), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_53), .B(n_133), .Y(n_232) );
CKINVDCx20_ASAP7_75t_R g161 ( .A(n_54), .Y(n_161) );
CKINVDCx14_ASAP7_75t_R g504 ( .A(n_55), .Y(n_504) );
INVx1_ASAP7_75t_L g139 ( .A(n_56), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_57), .B(n_133), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_58), .B(n_249), .Y(n_248) );
A2O1A1Ixp33_ASAP7_75t_L g245 ( .A1(n_59), .A2(n_151), .B(n_174), .C(n_246), .Y(n_245) );
INVx1_ASAP7_75t_L g158 ( .A(n_60), .Y(n_158) );
OAI22xp5_ASAP7_75t_L g461 ( .A1(n_61), .A2(n_100), .B1(n_462), .B2(n_463), .Y(n_461) );
CKINVDCx20_ASAP7_75t_R g463 ( .A(n_61), .Y(n_463) );
INVx1_ASAP7_75t_SL g568 ( .A(n_62), .Y(n_568) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_63), .Y(n_117) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_64), .B(n_177), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_65), .B(n_249), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_66), .B(n_178), .Y(n_223) );
INVx1_ASAP7_75t_L g558 ( .A(n_67), .Y(n_558) );
CKINVDCx16_ASAP7_75t_R g259 ( .A(n_68), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_69), .B(n_146), .Y(n_145) );
A2O1A1Ixp33_ASAP7_75t_L g171 ( .A1(n_70), .A2(n_141), .B(n_172), .C(n_181), .Y(n_171) );
CKINVDCx16_ASAP7_75t_R g244 ( .A(n_71), .Y(n_244) );
INVx1_ASAP7_75t_L g109 ( .A(n_72), .Y(n_109) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_73), .A2(n_133), .B(n_503), .Y(n_502) );
CKINVDCx20_ASAP7_75t_R g561 ( .A(n_74), .Y(n_561) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_75), .A2(n_133), .B(n_523), .Y(n_522) );
AOI222xp33_ASAP7_75t_SL g460 ( .A1(n_76), .A2(n_461), .B1(n_464), .B2(n_743), .C1(n_744), .C2(n_748), .Y(n_460) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_77), .A2(n_132), .B(n_492), .Y(n_491) );
CKINVDCx16_ASAP7_75t_R g477 ( .A(n_78), .Y(n_477) );
INVx1_ASAP7_75t_L g524 ( .A(n_79), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g148 ( .A(n_80), .B(n_149), .Y(n_148) );
AOI22xp5_ASAP7_75t_L g101 ( .A1(n_81), .A2(n_102), .B1(n_112), .B2(n_752), .Y(n_101) );
CKINVDCx20_ASAP7_75t_R g198 ( .A(n_82), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_83), .A2(n_133), .B(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g527 ( .A(n_84), .Y(n_527) );
INVx2_ASAP7_75t_L g156 ( .A(n_85), .Y(n_156) );
INVx1_ASAP7_75t_L g541 ( .A(n_86), .Y(n_541) );
CKINVDCx20_ASAP7_75t_R g185 ( .A(n_87), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_88), .B(n_225), .Y(n_224) );
INVx2_ASAP7_75t_L g106 ( .A(n_89), .Y(n_106) );
OR2x2_ASAP7_75t_L g453 ( .A(n_89), .B(n_454), .Y(n_453) );
OR2x2_ASAP7_75t_L g467 ( .A(n_89), .B(n_455), .Y(n_467) );
A2O1A1Ixp33_ASAP7_75t_L g556 ( .A1(n_90), .A2(n_141), .B(n_181), .C(n_557), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_91), .B(n_133), .Y(n_188) );
INVx1_ASAP7_75t_L g193 ( .A(n_92), .Y(n_193) );
INVxp67_ASAP7_75t_L g247 ( .A(n_93), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_94), .B(n_168), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_95), .B(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g173 ( .A(n_96), .Y(n_173) );
INVx1_ASAP7_75t_L g219 ( .A(n_97), .Y(n_219) );
INVx2_ASAP7_75t_L g517 ( .A(n_98), .Y(n_517) );
AND2x2_ASAP7_75t_L g237 ( .A(n_99), .B(n_155), .Y(n_237) );
CKINVDCx20_ASAP7_75t_R g462 ( .A(n_100), .Y(n_462) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
HB1xp67_ASAP7_75t_L g752 ( .A(n_103), .Y(n_752) );
OR2x2_ASAP7_75t_L g103 ( .A(n_104), .B(n_110), .Y(n_103) );
NAND3xp33_ASAP7_75t_SL g104 ( .A(n_105), .B(n_106), .C(n_107), .Y(n_104) );
AND2x2_ASAP7_75t_L g455 ( .A(n_105), .B(n_456), .Y(n_455) );
OR2x2_ASAP7_75t_L g468 ( .A(n_106), .B(n_455), .Y(n_468) );
NOR2x2_ASAP7_75t_L g750 ( .A(n_106), .B(n_454), .Y(n_750) );
INVx1_ASAP7_75t_SL g107 ( .A(n_108), .Y(n_107) );
OA21x2_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_118), .B(n_459), .Y(n_112) );
INVx1_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
INVx1_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
BUFx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx1_ASAP7_75t_L g751 ( .A(n_117), .Y(n_751) );
OAI21xp5_ASAP7_75t_SL g118 ( .A1(n_119), .A2(n_450), .B(n_457), .Y(n_118) );
INVxp67_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
OAI22xp5_ASAP7_75t_SL g744 ( .A1(n_123), .A2(n_470), .B1(n_745), .B2(n_746), .Y(n_744) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
BUFx2_ASAP7_75t_L g448 ( .A(n_124), .Y(n_448) );
AND3x1_ASAP7_75t_L g124 ( .A(n_125), .B(n_352), .C(n_409), .Y(n_124) );
NOR3xp33_ASAP7_75t_L g125 ( .A(n_126), .B(n_297), .C(n_333), .Y(n_125) );
OAI211xp5_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_199), .B(n_251), .C(n_284), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_128), .B(n_163), .Y(n_127) );
HB1xp67_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
AND2x4_ASAP7_75t_L g254 ( .A(n_129), .B(n_255), .Y(n_254) );
INVx5_ASAP7_75t_L g283 ( .A(n_129), .Y(n_283) );
AND2x2_ASAP7_75t_L g356 ( .A(n_129), .B(n_272), .Y(n_356) );
AND2x2_ASAP7_75t_L g394 ( .A(n_129), .B(n_300), .Y(n_394) );
AND2x2_ASAP7_75t_L g414 ( .A(n_129), .B(n_256), .Y(n_414) );
OR2x6_ASAP7_75t_L g129 ( .A(n_130), .B(n_160), .Y(n_129) );
AOI21xp5_ASAP7_75t_SL g130 ( .A1(n_131), .A2(n_140), .B(n_153), .Y(n_130) );
BUFx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
AND2x4_ASAP7_75t_L g133 ( .A(n_134), .B(n_138), .Y(n_133) );
NAND2x1p5_ASAP7_75t_L g220 ( .A(n_134), .B(n_138), .Y(n_220) );
AND2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_137), .Y(n_134) );
INVx1_ASAP7_75t_L g151 ( .A(n_135), .Y(n_151) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx2_ASAP7_75t_L g142 ( .A(n_136), .Y(n_142) );
INVx1_ASAP7_75t_L g214 ( .A(n_136), .Y(n_214) );
INVx1_ASAP7_75t_L g143 ( .A(n_137), .Y(n_143) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_137), .Y(n_147) );
INVx3_ASAP7_75t_L g178 ( .A(n_137), .Y(n_178) );
INVx1_ASAP7_75t_L g210 ( .A(n_137), .Y(n_210) );
BUFx6f_ASAP7_75t_L g225 ( .A(n_137), .Y(n_225) );
BUFx3_ASAP7_75t_L g152 ( .A(n_138), .Y(n_152) );
INVx4_ASAP7_75t_SL g182 ( .A(n_138), .Y(n_182) );
INVx5_ASAP7_75t_L g191 ( .A(n_141), .Y(n_191) );
AND2x6_ASAP7_75t_L g141 ( .A(n_142), .B(n_143), .Y(n_141) );
BUFx6f_ASAP7_75t_L g180 ( .A(n_142), .Y(n_180) );
BUFx3_ASAP7_75t_L g196 ( .A(n_142), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_148), .B(n_150), .Y(n_144) );
INVx2_ASAP7_75t_L g149 ( .A(n_146), .Y(n_149) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx4_ASAP7_75t_L g175 ( .A(n_147), .Y(n_175) );
O2A1O1Ixp33_ASAP7_75t_L g192 ( .A1(n_149), .A2(n_193), .B(n_194), .C(n_195), .Y(n_192) );
O2A1O1Ixp33_ASAP7_75t_L g234 ( .A1(n_149), .A2(n_195), .B(n_235), .C(n_236), .Y(n_234) );
O2A1O1Ixp5_ASAP7_75t_L g540 ( .A1(n_149), .A2(n_541), .B(n_542), .C(n_543), .Y(n_540) );
O2A1O1Ixp33_ASAP7_75t_L g557 ( .A1(n_149), .A2(n_543), .B(n_558), .C(n_559), .Y(n_557) );
O2A1O1Ixp33_ASAP7_75t_L g479 ( .A1(n_150), .A2(n_177), .B(n_480), .C(n_481), .Y(n_479) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
NAND2xp5_ASAP7_75t_SL g494 ( .A(n_151), .B(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
NOR2xp33_ASAP7_75t_L g560 ( .A(n_154), .B(n_561), .Y(n_560) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx1_ASAP7_75t_L g162 ( .A(n_155), .Y(n_162) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_155), .A2(n_188), .B(n_189), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_155), .A2(n_232), .B(n_233), .Y(n_231) );
O2A1O1Ixp33_ASAP7_75t_L g476 ( .A1(n_155), .A2(n_220), .B(n_477), .C(n_478), .Y(n_476) );
OA21x2_ASAP7_75t_L g501 ( .A1(n_155), .A2(n_502), .B(n_509), .Y(n_501) );
AND2x2_ASAP7_75t_SL g155 ( .A(n_156), .B(n_157), .Y(n_155) );
AND2x2_ASAP7_75t_L g169 ( .A(n_156), .B(n_157), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_158), .B(n_159), .Y(n_157) );
NOR2xp33_ASAP7_75t_L g160 ( .A(n_161), .B(n_162), .Y(n_160) );
AO21x2_ASAP7_75t_L g536 ( .A1(n_162), .A2(n_537), .B(n_544), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_163), .B(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g163 ( .A(n_164), .B(n_186), .Y(n_163) );
HB1xp67_ASAP7_75t_L g295 ( .A(n_164), .Y(n_295) );
AND2x2_ASAP7_75t_L g309 ( .A(n_164), .B(n_255), .Y(n_309) );
INVx1_ASAP7_75t_L g332 ( .A(n_164), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_164), .B(n_283), .Y(n_371) );
OR2x2_ASAP7_75t_L g408 ( .A(n_164), .B(n_253), .Y(n_408) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
HB1xp67_ASAP7_75t_L g344 ( .A(n_165), .Y(n_344) );
AND2x2_ASAP7_75t_L g351 ( .A(n_165), .B(n_256), .Y(n_351) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
AND2x2_ASAP7_75t_L g272 ( .A(n_166), .B(n_256), .Y(n_272) );
BUFx2_ASAP7_75t_L g300 ( .A(n_166), .Y(n_300) );
AO21x2_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_170), .B(n_184), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g184 ( .A(n_167), .B(n_185), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_167), .B(n_198), .Y(n_197) );
AO21x2_ASAP7_75t_L g217 ( .A1(n_167), .A2(n_218), .B(n_226), .Y(n_217) );
INVx3_ASAP7_75t_L g249 ( .A(n_167), .Y(n_249) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_167), .B(n_483), .Y(n_482) );
NOR2xp33_ASAP7_75t_L g544 ( .A(n_167), .B(n_545), .Y(n_544) );
AO21x2_ASAP7_75t_L g553 ( .A1(n_167), .A2(n_554), .B(n_560), .Y(n_553) );
INVx4_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_168), .A2(n_206), .B(n_207), .Y(n_205) );
HB1xp67_ASAP7_75t_L g241 ( .A(n_168), .Y(n_241) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx1_ASAP7_75t_L g228 ( .A(n_169), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_171), .B(n_183), .Y(n_170) );
O2A1O1Ixp33_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_174), .B(n_176), .C(n_179), .Y(n_172) );
INVx1_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
OAI22xp33_ASAP7_75t_L g495 ( .A1(n_175), .A2(n_177), .B1(n_496), .B2(n_497), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_175), .B(n_517), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_175), .B(n_527), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_177), .B(n_247), .Y(n_246) );
INVx2_ASAP7_75t_L g261 ( .A(n_177), .Y(n_261) );
INVx5_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g507 ( .A(n_178), .B(n_508), .Y(n_507) );
HB1xp67_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx3_ASAP7_75t_L g569 ( .A(n_180), .Y(n_569) );
INVx1_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
O2A1O1Ixp33_ASAP7_75t_L g243 ( .A1(n_182), .A2(n_191), .B(n_244), .C(n_245), .Y(n_243) );
O2A1O1Ixp33_ASAP7_75t_SL g258 ( .A1(n_182), .A2(n_191), .B(n_259), .C(n_260), .Y(n_258) );
O2A1O1Ixp33_ASAP7_75t_SL g492 ( .A1(n_182), .A2(n_191), .B(n_493), .C(n_494), .Y(n_492) );
O2A1O1Ixp33_ASAP7_75t_SL g503 ( .A1(n_182), .A2(n_191), .B(n_504), .C(n_505), .Y(n_503) );
O2A1O1Ixp33_ASAP7_75t_SL g513 ( .A1(n_182), .A2(n_191), .B(n_514), .C(n_515), .Y(n_513) );
O2A1O1Ixp33_ASAP7_75t_SL g523 ( .A1(n_182), .A2(n_191), .B(n_524), .C(n_525), .Y(n_523) );
O2A1O1Ixp33_ASAP7_75t_L g564 ( .A1(n_182), .A2(n_191), .B(n_565), .C(n_566), .Y(n_564) );
INVx5_ASAP7_75t_L g253 ( .A(n_186), .Y(n_253) );
BUFx2_ASAP7_75t_L g276 ( .A(n_186), .Y(n_276) );
AND2x2_ASAP7_75t_L g433 ( .A(n_186), .B(n_287), .Y(n_433) );
OR2x6_ASAP7_75t_L g186 ( .A(n_187), .B(n_197), .Y(n_186) );
INVx2_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
HB1xp67_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
INVx2_ASAP7_75t_L g265 ( .A(n_196), .Y(n_265) );
INVx1_ASAP7_75t_L g528 ( .A(n_196), .Y(n_528) );
INVx1_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
NAND2xp33_ASAP7_75t_L g200 ( .A(n_201), .B(n_238), .Y(n_200) );
OAI221xp5_ASAP7_75t_L g333 ( .A1(n_201), .A2(n_334), .B1(n_341), .B2(n_342), .C(n_345), .Y(n_333) );
OR2x2_ASAP7_75t_L g201 ( .A(n_202), .B(n_215), .Y(n_201) );
AND2x2_ASAP7_75t_L g239 ( .A(n_202), .B(n_240), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_202), .B(n_328), .Y(n_327) );
INVx1_ASAP7_75t_SL g202 ( .A(n_203), .Y(n_202) );
AND2x2_ASAP7_75t_L g268 ( .A(n_203), .B(n_216), .Y(n_268) );
NAND2xp5_ASAP7_75t_SL g278 ( .A(n_203), .B(n_217), .Y(n_278) );
OR2x2_ASAP7_75t_L g289 ( .A(n_203), .B(n_240), .Y(n_289) );
AND2x2_ASAP7_75t_L g292 ( .A(n_203), .B(n_280), .Y(n_292) );
AND2x2_ASAP7_75t_L g308 ( .A(n_203), .B(n_229), .Y(n_308) );
OR2x2_ASAP7_75t_L g324 ( .A(n_203), .B(n_217), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_203), .B(n_240), .Y(n_386) );
INVx2_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_204), .B(n_229), .Y(n_378) );
AND2x2_ASAP7_75t_L g381 ( .A(n_204), .B(n_217), .Y(n_381) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_209), .A2(n_211), .B(n_212), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_212), .A2(n_223), .B(n_224), .Y(n_222) );
INVx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
INVx3_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
OR2x2_ASAP7_75t_L g302 ( .A(n_215), .B(n_289), .Y(n_302) );
INVx2_ASAP7_75t_L g328 ( .A(n_215), .Y(n_328) );
OR2x2_ASAP7_75t_L g215 ( .A(n_216), .B(n_229), .Y(n_215) );
AND2x2_ASAP7_75t_L g250 ( .A(n_216), .B(n_230), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_216), .B(n_240), .Y(n_307) );
OR2x2_ASAP7_75t_L g318 ( .A(n_216), .B(n_230), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_216), .B(n_280), .Y(n_377) );
OAI221xp5_ASAP7_75t_L g410 ( .A1(n_216), .A2(n_411), .B1(n_413), .B2(n_415), .C(n_418), .Y(n_410) );
INVx5_ASAP7_75t_SL g216 ( .A(n_217), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_217), .B(n_240), .Y(n_349) );
OAI21xp5_ASAP7_75t_L g218 ( .A1(n_219), .A2(n_220), .B(n_221), .Y(n_218) );
OAI21xp5_ASAP7_75t_L g537 ( .A1(n_220), .A2(n_538), .B(n_539), .Y(n_537) );
OAI21xp5_ASAP7_75t_L g554 ( .A1(n_220), .A2(n_555), .B(n_556), .Y(n_554) );
INVx4_ASAP7_75t_L g264 ( .A(n_225), .Y(n_264) );
INVx2_ASAP7_75t_L g506 ( .A(n_225), .Y(n_506) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_227), .B(n_228), .Y(n_226) );
INVx2_ASAP7_75t_L g489 ( .A(n_228), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_229), .B(n_280), .Y(n_279) );
NOR2xp33_ASAP7_75t_L g290 ( .A(n_229), .B(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g296 ( .A(n_229), .B(n_268), .Y(n_296) );
OR2x2_ASAP7_75t_L g340 ( .A(n_229), .B(n_240), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_229), .B(n_292), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_229), .B(n_385), .Y(n_384) );
AND2x2_ASAP7_75t_L g405 ( .A(n_229), .B(n_406), .Y(n_405) );
INVx5_ASAP7_75t_SL g229 ( .A(n_230), .Y(n_229) );
AND2x2_ASAP7_75t_SL g269 ( .A(n_230), .B(n_239), .Y(n_269) );
O2A1O1Ixp33_ASAP7_75t_SL g273 ( .A1(n_230), .A2(n_274), .B(n_277), .C(n_281), .Y(n_273) );
OR2x2_ASAP7_75t_L g311 ( .A(n_230), .B(n_307), .Y(n_311) );
OR2x2_ASAP7_75t_L g347 ( .A(n_230), .B(n_289), .Y(n_347) );
OAI311xp33_ASAP7_75t_L g353 ( .A1(n_230), .A2(n_292), .A3(n_354), .B1(n_357), .C1(n_364), .Y(n_353) );
AND2x2_ASAP7_75t_L g404 ( .A(n_230), .B(n_240), .Y(n_404) );
AND2x2_ASAP7_75t_L g412 ( .A(n_230), .B(n_267), .Y(n_412) );
HB1xp67_ASAP7_75t_L g430 ( .A(n_230), .Y(n_430) );
AND2x2_ASAP7_75t_L g447 ( .A(n_230), .B(n_268), .Y(n_447) );
OR2x6_ASAP7_75t_L g230 ( .A(n_231), .B(n_237), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_239), .B(n_250), .Y(n_238) );
AND2x2_ASAP7_75t_L g275 ( .A(n_239), .B(n_276), .Y(n_275) );
INVx2_ASAP7_75t_L g431 ( .A(n_239), .Y(n_431) );
AND2x2_ASAP7_75t_L g267 ( .A(n_240), .B(n_268), .Y(n_267) );
INVx3_ASAP7_75t_L g280 ( .A(n_240), .Y(n_280) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_240), .Y(n_323) );
INVxp67_ASAP7_75t_L g362 ( .A(n_240), .Y(n_362) );
OA21x2_ASAP7_75t_L g240 ( .A1(n_241), .A2(n_242), .B(n_248), .Y(n_240) );
OA21x2_ASAP7_75t_L g511 ( .A1(n_241), .A2(n_512), .B(n_518), .Y(n_511) );
OA21x2_ASAP7_75t_L g521 ( .A1(n_241), .A2(n_522), .B(n_529), .Y(n_521) );
OA21x2_ASAP7_75t_L g562 ( .A1(n_241), .A2(n_563), .B(n_570), .Y(n_562) );
OA21x2_ASAP7_75t_L g256 ( .A1(n_249), .A2(n_257), .B(n_266), .Y(n_256) );
AND2x2_ASAP7_75t_L g440 ( .A(n_250), .B(n_288), .Y(n_440) );
AOI221xp5_ASAP7_75t_L g251 ( .A1(n_252), .A2(n_267), .B1(n_269), .B2(n_270), .C(n_273), .Y(n_251) );
AND2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_254), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_253), .B(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g293 ( .A(n_253), .B(n_283), .Y(n_293) );
AND2x2_ASAP7_75t_L g301 ( .A(n_253), .B(n_255), .Y(n_301) );
OR2x2_ASAP7_75t_L g313 ( .A(n_253), .B(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g331 ( .A(n_253), .B(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g355 ( .A(n_253), .B(n_356), .Y(n_355) );
HB1xp67_ASAP7_75t_L g375 ( .A(n_253), .Y(n_375) );
AND2x2_ASAP7_75t_L g427 ( .A(n_253), .B(n_351), .Y(n_427) );
OAI31xp33_ASAP7_75t_L g435 ( .A1(n_253), .A2(n_304), .A3(n_403), .B(n_436), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_254), .B(n_331), .Y(n_330) );
INVx1_ASAP7_75t_SL g399 ( .A(n_254), .Y(n_399) );
NOR2xp33_ASAP7_75t_L g407 ( .A(n_254), .B(n_408), .Y(n_407) );
AND2x4_ASAP7_75t_L g287 ( .A(n_255), .B(n_283), .Y(n_287) );
INVx1_ASAP7_75t_L g374 ( .A(n_255), .Y(n_374) );
INVx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g424 ( .A(n_256), .B(n_283), .Y(n_424) );
NOR2xp33_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
NOR2xp33_ASAP7_75t_L g567 ( .A(n_264), .B(n_568), .Y(n_567) );
INVx2_ASAP7_75t_L g543 ( .A(n_265), .Y(n_543) );
INVx1_ASAP7_75t_SL g434 ( .A(n_267), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_268), .B(n_339), .Y(n_338) );
AOI22xp5_ASAP7_75t_L g418 ( .A1(n_269), .A2(n_381), .B1(n_419), .B2(n_422), .Y(n_418) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g282 ( .A(n_272), .B(n_283), .Y(n_282) );
INVx1_ASAP7_75t_L g341 ( .A(n_272), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_272), .B(n_293), .Y(n_446) );
INVx1_ASAP7_75t_SL g274 ( .A(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g416 ( .A(n_275), .B(n_417), .Y(n_416) );
AOI21xp5_ASAP7_75t_L g334 ( .A1(n_276), .A2(n_335), .B(n_337), .Y(n_334) );
OR2x2_ASAP7_75t_L g342 ( .A(n_276), .B(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g363 ( .A(n_276), .B(n_351), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_276), .B(n_374), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_276), .B(n_414), .Y(n_413) );
OAI221xp5_ASAP7_75t_SL g390 ( .A1(n_277), .A2(n_391), .B1(n_396), .B2(n_399), .C(n_400), .Y(n_390) );
OR2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
OR2x2_ASAP7_75t_L g367 ( .A(n_278), .B(n_340), .Y(n_367) );
INVx1_ASAP7_75t_L g406 ( .A(n_278), .Y(n_406) );
INVx2_ASAP7_75t_L g382 ( .A(n_279), .Y(n_382) );
INVx1_ASAP7_75t_L g316 ( .A(n_280), .Y(n_316) );
INVx1_ASAP7_75t_SL g281 ( .A(n_282), .Y(n_281) );
INVx2_ASAP7_75t_L g321 ( .A(n_283), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_283), .B(n_344), .Y(n_343) );
AND2x2_ASAP7_75t_L g350 ( .A(n_283), .B(n_351), .Y(n_350) );
OR2x2_ASAP7_75t_L g438 ( .A(n_283), .B(n_408), .Y(n_438) );
AOI222xp33_ASAP7_75t_L g284 ( .A1(n_285), .A2(n_288), .B1(n_290), .B2(n_293), .C1(n_294), .C2(n_296), .Y(n_284) );
INVxp67_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g294 ( .A(n_287), .B(n_295), .Y(n_294) );
AOI22xp33_ASAP7_75t_L g364 ( .A1(n_287), .A2(n_337), .B1(n_365), .B2(n_366), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_287), .B(n_421), .Y(n_420) );
INVx1_ASAP7_75t_SL g288 ( .A(n_289), .Y(n_288) );
INVx1_ASAP7_75t_SL g291 ( .A(n_292), .Y(n_291) );
OAI21xp33_ASAP7_75t_SL g325 ( .A1(n_296), .A2(n_326), .B(n_329), .Y(n_325) );
OAI211xp5_ASAP7_75t_SL g297 ( .A1(n_298), .A2(n_302), .B(n_303), .C(n_325), .Y(n_297) );
INVxp67_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
AOI221xp5_ASAP7_75t_L g303 ( .A1(n_301), .A2(n_304), .B1(n_309), .B2(n_310), .C(n_312), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_301), .B(n_389), .Y(n_388) );
INVxp67_ASAP7_75t_L g395 ( .A(n_301), .Y(n_395) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_306), .B(n_308), .Y(n_305) );
AND2x2_ASAP7_75t_L g397 ( .A(n_306), .B(n_398), .Y(n_397) );
INVx1_ASAP7_75t_SL g306 ( .A(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g314 ( .A(n_309), .Y(n_314) );
AND2x2_ASAP7_75t_L g320 ( .A(n_309), .B(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
OAI22xp5_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_315), .B1(n_319), .B2(n_322), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_316), .B(n_328), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_317), .B(n_362), .Y(n_361) );
INVx1_ASAP7_75t_SL g317 ( .A(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g417 ( .A(n_321), .Y(n_417) );
AND2x2_ASAP7_75t_L g436 ( .A(n_321), .B(n_351), .Y(n_436) );
OR2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_328), .B(n_385), .Y(n_444) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
NOR2xp33_ASAP7_75t_L g442 ( .A(n_331), .B(n_399), .Y(n_442) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g365 ( .A(n_343), .Y(n_365) );
BUFx2_ASAP7_75t_L g389 ( .A(n_344), .Y(n_389) );
OAI21xp5_ASAP7_75t_SL g345 ( .A1(n_346), .A2(n_348), .B(n_350), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
NOR3xp33_ASAP7_75t_L g352 ( .A(n_353), .B(n_368), .C(n_390), .Y(n_352) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
OAI21xp5_ASAP7_75t_L g357 ( .A1(n_358), .A2(n_360), .B(n_363), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_SL g366 ( .A(n_367), .Y(n_366) );
A2O1A1Ixp33_ASAP7_75t_SL g368 ( .A1(n_369), .A2(n_372), .B(n_376), .C(n_379), .Y(n_368) );
NAND2xp5_ASAP7_75t_SL g401 ( .A(n_369), .B(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
NOR2xp67_ASAP7_75t_SL g373 ( .A(n_374), .B(n_375), .Y(n_373) );
OR2x2_ASAP7_75t_L g376 ( .A(n_377), .B(n_378), .Y(n_376) );
INVx1_ASAP7_75t_SL g398 ( .A(n_378), .Y(n_398) );
OAI21xp5_ASAP7_75t_L g379 ( .A1(n_380), .A2(n_383), .B(n_387), .Y(n_379) );
AND2x4_ASAP7_75t_L g380 ( .A(n_381), .B(n_382), .Y(n_380) );
AND2x2_ASAP7_75t_L g403 ( .A(n_381), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_SL g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
NOR2xp33_ASAP7_75t_L g392 ( .A(n_393), .B(n_395), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
AOI22xp33_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_403), .B1(n_405), .B2(n_407), .Y(n_400) );
INVx2_ASAP7_75t_SL g421 ( .A(n_408), .Y(n_421) );
NOR3xp33_ASAP7_75t_L g409 ( .A(n_410), .B(n_425), .C(n_437), .Y(n_409) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVxp67_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVxp67_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_421), .B(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
OAI221xp5_ASAP7_75t_L g425 ( .A1(n_426), .A2(n_428), .B1(n_432), .B2(n_434), .C(n_435), .Y(n_425) );
A2O1A1Ixp33_ASAP7_75t_L g437 ( .A1(n_426), .A2(n_438), .B(n_439), .C(n_441), .Y(n_437) );
INVx1_ASAP7_75t_SL g426 ( .A(n_427), .Y(n_426) );
INVxp67_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
NOR2xp33_ASAP7_75t_L g429 ( .A(n_430), .B(n_431), .Y(n_429) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
AOI22xp5_ASAP7_75t_L g441 ( .A1(n_442), .A2(n_443), .B1(n_445), .B2(n_447), .Y(n_441) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
OAI22xp5_ASAP7_75t_L g464 ( .A1(n_448), .A2(n_465), .B1(n_468), .B2(n_469), .Y(n_464) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_SL g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_SL g452 ( .A(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g458 ( .A(n_453), .Y(n_458) );
INVx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
NAND3xp33_ASAP7_75t_L g459 ( .A(n_457), .B(n_460), .C(n_751), .Y(n_459) );
INVx1_ASAP7_75t_L g743 ( .A(n_461), .Y(n_743) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g745 ( .A(n_466), .Y(n_745) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g747 ( .A(n_468), .Y(n_747) );
INVx1_ASAP7_75t_SL g469 ( .A(n_470), .Y(n_469) );
OR5x1_ASAP7_75t_L g470 ( .A(n_471), .B(n_637), .C(n_701), .D(n_717), .E(n_732), .Y(n_470) );
NAND4xp25_ASAP7_75t_L g471 ( .A(n_472), .B(n_571), .C(n_598), .D(n_621), .Y(n_471) );
AOI21xp5_ASAP7_75t_L g472 ( .A1(n_473), .A2(n_519), .B(n_530), .Y(n_472) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_474), .B(n_484), .Y(n_473) );
HB1xp67_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx3_ASAP7_75t_SL g550 ( .A(n_475), .Y(n_550) );
AND2x4_ASAP7_75t_L g584 ( .A(n_475), .B(n_573), .Y(n_584) );
OR2x2_ASAP7_75t_L g594 ( .A(n_475), .B(n_552), .Y(n_594) );
OR2x2_ASAP7_75t_L g640 ( .A(n_475), .B(n_487), .Y(n_640) );
AND2x2_ASAP7_75t_L g654 ( .A(n_475), .B(n_551), .Y(n_654) );
AND2x2_ASAP7_75t_L g697 ( .A(n_475), .B(n_587), .Y(n_697) );
AND2x2_ASAP7_75t_L g704 ( .A(n_475), .B(n_562), .Y(n_704) );
AND2x2_ASAP7_75t_L g723 ( .A(n_475), .B(n_613), .Y(n_723) );
AND2x2_ASAP7_75t_L g741 ( .A(n_475), .B(n_583), .Y(n_741) );
OR2x6_ASAP7_75t_L g475 ( .A(n_476), .B(n_482), .Y(n_475) );
INVx1_ASAP7_75t_L g706 ( .A(n_484), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_485), .B(n_500), .Y(n_484) );
AND2x2_ASAP7_75t_L g616 ( .A(n_485), .B(n_551), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_485), .B(n_636), .Y(n_635) );
AOI32xp33_ASAP7_75t_L g649 ( .A1(n_485), .A2(n_650), .A3(n_653), .B1(n_655), .B2(n_659), .Y(n_649) );
AND2x2_ASAP7_75t_L g719 ( .A(n_485), .B(n_613), .Y(n_719) );
INVx2_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_SL g486 ( .A(n_487), .Y(n_486) );
AND2x2_ASAP7_75t_L g583 ( .A(n_487), .B(n_552), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_487), .B(n_593), .Y(n_592) );
AND2x2_ASAP7_75t_L g625 ( .A(n_487), .B(n_572), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_487), .B(n_704), .Y(n_703) );
AO21x2_ASAP7_75t_L g487 ( .A1(n_488), .A2(n_490), .B(n_498), .Y(n_487) );
INVx1_ASAP7_75t_L g588 ( .A(n_488), .Y(n_588) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
OA21x2_ASAP7_75t_L g587 ( .A1(n_491), .A2(n_499), .B(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
AND2x2_ASAP7_75t_L g590 ( .A(n_500), .B(n_534), .Y(n_590) );
AND2x2_ASAP7_75t_L g666 ( .A(n_500), .B(n_667), .Y(n_666) );
INVx1_ASAP7_75t_SL g738 ( .A(n_500), .Y(n_738) );
AND2x2_ASAP7_75t_L g500 ( .A(n_501), .B(n_510), .Y(n_500) );
OR2x2_ASAP7_75t_L g533 ( .A(n_501), .B(n_511), .Y(n_533) );
AND2x2_ASAP7_75t_L g547 ( .A(n_501), .B(n_548), .Y(n_547) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_501), .B(n_576), .Y(n_575) );
INVx2_ASAP7_75t_L g597 ( .A(n_501), .Y(n_597) );
AND2x2_ASAP7_75t_L g624 ( .A(n_501), .B(n_511), .Y(n_624) );
BUFx3_ASAP7_75t_L g627 ( .A(n_501), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_501), .B(n_602), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_501), .B(n_721), .Y(n_720) );
INVx2_ASAP7_75t_L g578 ( .A(n_510), .Y(n_578) );
AND2x2_ASAP7_75t_L g596 ( .A(n_510), .B(n_576), .Y(n_596) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
AND2x2_ASAP7_75t_L g607 ( .A(n_511), .B(n_521), .Y(n_607) );
HB1xp67_ASAP7_75t_L g620 ( .A(n_511), .Y(n_620) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_520), .B(n_627), .Y(n_677) );
HB1xp67_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx1_ASAP7_75t_SL g548 ( .A(n_521), .Y(n_548) );
NAND3xp33_ASAP7_75t_L g595 ( .A(n_521), .B(n_596), .C(n_597), .Y(n_595) );
OR2x2_ASAP7_75t_L g603 ( .A(n_521), .B(n_576), .Y(n_603) );
AND2x2_ASAP7_75t_L g623 ( .A(n_521), .B(n_576), .Y(n_623) );
AND2x2_ASAP7_75t_L g667 ( .A(n_521), .B(n_536), .Y(n_667) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_531), .A2(n_546), .B(n_549), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g531 ( .A(n_532), .B(n_534), .Y(n_531) );
AND2x2_ASAP7_75t_L g742 ( .A(n_532), .B(n_667), .Y(n_742) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
OAI22xp5_ASAP7_75t_L g681 ( .A1(n_533), .A2(n_640), .B1(n_682), .B2(n_684), .Y(n_681) );
OR2x2_ASAP7_75t_L g688 ( .A(n_533), .B(n_603), .Y(n_688) );
OR2x2_ASAP7_75t_L g712 ( .A(n_533), .B(n_713), .Y(n_712) );
NOR2xp33_ASAP7_75t_L g725 ( .A(n_533), .B(n_632), .Y(n_725) );
AND2x2_ASAP7_75t_L g618 ( .A(n_534), .B(n_619), .Y(n_618) );
AOI21xp5_ASAP7_75t_L g705 ( .A1(n_534), .A2(n_691), .B(n_706), .Y(n_705) );
AOI32xp33_ASAP7_75t_L g726 ( .A1(n_534), .A2(n_616), .A3(n_727), .B1(n_729), .B2(n_730), .Y(n_726) );
OR2x2_ASAP7_75t_L g737 ( .A(n_534), .B(n_738), .Y(n_737) );
CKINVDCx16_ASAP7_75t_R g534 ( .A(n_535), .Y(n_534) );
OR2x2_ASAP7_75t_L g605 ( .A(n_535), .B(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_535), .B(n_619), .Y(n_684) );
BUFx3_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx4_ASAP7_75t_L g576 ( .A(n_536), .Y(n_576) );
AND2x2_ASAP7_75t_L g642 ( .A(n_536), .B(n_607), .Y(n_642) );
AND3x2_ASAP7_75t_L g651 ( .A(n_536), .B(n_547), .C(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g577 ( .A(n_548), .B(n_578), .Y(n_577) );
HB1xp67_ASAP7_75t_L g632 ( .A(n_548), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_548), .B(n_576), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_550), .B(n_551), .Y(n_549) );
AND2x2_ASAP7_75t_L g572 ( .A(n_550), .B(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g612 ( .A(n_550), .B(n_613), .Y(n_612) );
AND2x2_ASAP7_75t_L g630 ( .A(n_550), .B(n_562), .Y(n_630) );
AND2x2_ASAP7_75t_L g648 ( .A(n_550), .B(n_552), .Y(n_648) );
OR2x2_ASAP7_75t_L g662 ( .A(n_550), .B(n_663), .Y(n_662) );
AND2x2_ASAP7_75t_L g708 ( .A(n_550), .B(n_636), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_551), .B(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g551 ( .A(n_552), .B(n_562), .Y(n_551) );
AND2x2_ASAP7_75t_L g609 ( .A(n_552), .B(n_587), .Y(n_609) );
OR2x2_ASAP7_75t_L g663 ( .A(n_552), .B(n_587), .Y(n_663) );
AND2x2_ASAP7_75t_L g716 ( .A(n_552), .B(n_573), .Y(n_716) );
INVx2_ASAP7_75t_SL g552 ( .A(n_553), .Y(n_552) );
BUFx2_ASAP7_75t_L g614 ( .A(n_553), .Y(n_614) );
AND2x2_ASAP7_75t_L g636 ( .A(n_553), .B(n_562), .Y(n_636) );
INVx2_ASAP7_75t_L g573 ( .A(n_562), .Y(n_573) );
INVx1_ASAP7_75t_L g593 ( .A(n_562), .Y(n_593) );
AOI211xp5_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_574), .B(n_579), .C(n_591), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_572), .B(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g735 ( .A(n_572), .Y(n_735) );
AND2x2_ASAP7_75t_L g613 ( .A(n_573), .B(n_614), .Y(n_613) );
AND2x2_ASAP7_75t_L g574 ( .A(n_575), .B(n_577), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_576), .B(n_577), .Y(n_585) );
INVx1_ASAP7_75t_L g670 ( .A(n_576), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_576), .B(n_597), .Y(n_694) );
AND2x2_ASAP7_75t_L g710 ( .A(n_576), .B(n_624), .Y(n_710) );
NAND2xp5_ASAP7_75t_SL g692 ( .A(n_577), .B(n_693), .Y(n_692) );
INVx2_ASAP7_75t_L g601 ( .A(n_578), .Y(n_601) );
OAI22xp5_ASAP7_75t_L g579 ( .A1(n_580), .A2(n_585), .B1(n_586), .B2(n_589), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
NOR2xp33_ASAP7_75t_L g581 ( .A(n_582), .B(n_584), .Y(n_581) );
NOR2xp33_ASAP7_75t_L g734 ( .A(n_582), .B(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_583), .B(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g608 ( .A(n_584), .B(n_609), .Y(n_608) );
AOI221xp5_ASAP7_75t_SL g673 ( .A1(n_584), .A2(n_626), .B1(n_674), .B2(n_679), .C(n_681), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_584), .B(n_647), .Y(n_680) );
INVx1_ASAP7_75t_L g740 ( .A(n_586), .Y(n_740) );
BUFx3_ASAP7_75t_L g647 ( .A(n_587), .Y(n_647) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
AOI21xp33_ASAP7_75t_SL g591 ( .A1(n_592), .A2(n_594), .B(n_595), .Y(n_591) );
INVx1_ASAP7_75t_L g656 ( .A(n_593), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_593), .B(n_647), .Y(n_700) );
INVx1_ASAP7_75t_L g657 ( .A(n_594), .Y(n_657) );
NAND2xp5_ASAP7_75t_SL g658 ( .A(n_594), .B(n_647), .Y(n_658) );
INVxp67_ASAP7_75t_L g678 ( .A(n_596), .Y(n_678) );
AND2x2_ASAP7_75t_L g619 ( .A(n_597), .B(n_620), .Y(n_619) );
O2A1O1Ixp33_ASAP7_75t_L g598 ( .A1(n_599), .A2(n_604), .B(n_608), .C(n_610), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
INVx1_ASAP7_75t_SL g633 ( .A(n_601), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_602), .B(n_633), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_602), .B(n_624), .Y(n_675) );
INVx2_ASAP7_75t_SL g602 ( .A(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
OAI22xp5_ASAP7_75t_L g610 ( .A1(n_605), .A2(n_611), .B1(n_615), .B2(n_617), .Y(n_610) );
INVx1_ASAP7_75t_SL g606 ( .A(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g626 ( .A(n_607), .B(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g671 ( .A(n_607), .B(n_672), .Y(n_671) );
OAI21xp33_ASAP7_75t_L g674 ( .A1(n_609), .A2(n_675), .B(n_676), .Y(n_674) );
INVx1_ASAP7_75t_SL g611 ( .A(n_612), .Y(n_611) );
AOI221xp5_ASAP7_75t_L g621 ( .A1(n_613), .A2(n_622), .B1(n_625), .B2(n_626), .C(n_628), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_613), .B(n_647), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_613), .B(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g729 ( .A(n_619), .Y(n_729) );
INVxp67_ASAP7_75t_L g652 ( .A(n_620), .Y(n_652) );
INVx1_ASAP7_75t_L g659 ( .A(n_622), .Y(n_659) );
AND2x2_ASAP7_75t_L g622 ( .A(n_623), .B(n_624), .Y(n_622) );
AND2x2_ASAP7_75t_L g698 ( .A(n_623), .B(n_627), .Y(n_698) );
INVx1_ASAP7_75t_L g672 ( .A(n_627), .Y(n_672) );
NAND2xp5_ASAP7_75t_SL g702 ( .A(n_627), .B(n_642), .Y(n_702) );
OAI32xp33_ASAP7_75t_L g628 ( .A1(n_629), .A2(n_631), .A3(n_633), .B1(n_634), .B2(n_635), .Y(n_628) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
INVx2_ASAP7_75t_SL g641 ( .A(n_636), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_636), .B(n_668), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_636), .B(n_697), .Y(n_728) );
NAND2x1p5_ASAP7_75t_L g736 ( .A(n_636), .B(n_647), .Y(n_736) );
NAND5xp2_ASAP7_75t_L g637 ( .A(n_638), .B(n_660), .C(n_673), .D(n_685), .E(n_686), .Y(n_637) );
AOI221xp5_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_642), .B1(n_643), .B2(n_645), .C(n_649), .Y(n_638) );
NOR2xp33_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .Y(n_639) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
NAND2xp33_ASAP7_75t_SL g664 ( .A(n_644), .B(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_647), .B(n_648), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_647), .B(n_716), .Y(n_715) );
AOI22xp33_ASAP7_75t_L g660 ( .A1(n_648), .A2(n_661), .B1(n_664), .B2(n_668), .Y(n_660) );
INVx2_ASAP7_75t_SL g650 ( .A(n_651), .Y(n_650) );
OAI211xp5_ASAP7_75t_SL g655 ( .A1(n_651), .A2(n_656), .B(n_657), .C(n_658), .Y(n_655) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_SL g683 ( .A(n_663), .Y(n_683) );
INVx1_ASAP7_75t_SL g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_SL g668 ( .A(n_669), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_670), .B(n_671), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_672), .B(n_721), .Y(n_731) );
OR2x2_ASAP7_75t_L g676 ( .A(n_677), .B(n_678), .Y(n_676) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
AOI222xp33_ASAP7_75t_L g686 ( .A1(n_687), .A2(n_689), .B1(n_691), .B2(n_695), .C1(n_698), .C2(n_699), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
OAI221xp5_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_703), .B1(n_705), .B2(n_707), .C(n_709), .Y(n_701) );
INVx1_ASAP7_75t_SL g707 ( .A(n_708), .Y(n_707) );
OAI21xp33_ASAP7_75t_L g709 ( .A1(n_710), .A2(n_711), .B(n_714), .Y(n_709) );
INVx2_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g721 ( .A(n_713), .Y(n_721) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
OAI221xp5_ASAP7_75t_L g717 ( .A1(n_718), .A2(n_720), .B1(n_722), .B2(n_724), .C(n_726), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_SL g722 ( .A(n_723), .Y(n_722) );
INVxp67_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
A2O1A1Ixp33_ASAP7_75t_L g732 ( .A1(n_733), .A2(n_736), .B(n_737), .C(n_739), .Y(n_732) );
INVxp67_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
OAI21xp33_ASAP7_75t_L g739 ( .A1(n_740), .A2(n_741), .B(n_742), .Y(n_739) );
INVx2_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_SL g748 ( .A(n_749), .Y(n_748) );
INVx3_ASAP7_75t_SL g749 ( .A(n_750), .Y(n_749) );
endmodule