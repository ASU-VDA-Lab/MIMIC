module real_jpeg_17175_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_202;
wire n_128;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_516;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_15;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

OAI21xp5_ASAP7_75t_L g14 ( 
.A1(n_0),
.A2(n_15),
.B(n_16),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_0),
.B(n_17),
.Y(n_16)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_1),
.A2(n_110),
.B1(n_115),
.B2(n_119),
.Y(n_109)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_1),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_1),
.A2(n_119),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_1),
.A2(n_119),
.B1(n_252),
.B2(n_254),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_1),
.A2(n_119),
.B1(n_337),
.B2(n_340),
.Y(n_336)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_2),
.Y(n_126)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_2),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_2),
.Y(n_134)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_2),
.Y(n_138)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_3),
.Y(n_80)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_3),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_3),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_3),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_4),
.A2(n_227),
.B1(n_228),
.B2(n_229),
.Y(n_226)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_4),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_4),
.A2(n_228),
.B1(n_284),
.B2(n_286),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_4),
.A2(n_228),
.B1(n_310),
.B2(n_327),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_L g395 ( 
.A1(n_4),
.A2(n_228),
.B1(n_396),
.B2(n_399),
.Y(n_395)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_5),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_5),
.Y(n_181)
);

CKINVDCx14_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

INVx2_ASAP7_75t_SL g23 ( 
.A(n_7),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_7),
.A2(n_23),
.B1(n_102),
.B2(n_104),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_7),
.A2(n_23),
.B1(n_184),
.B2(n_188),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_7),
.B(n_219),
.Y(n_218)
);

OAI32xp33_ASAP7_75t_L g369 ( 
.A1(n_7),
.A2(n_370),
.A3(n_373),
.B1(n_376),
.B2(n_380),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_7),
.B(n_132),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_7),
.B(n_416),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_7),
.B(n_78),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_8),
.Y(n_93)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_8),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_8),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_8),
.Y(n_107)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_8),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_8),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g311 ( 
.A(n_8),
.Y(n_311)
);

BUFx5_ASAP7_75t_L g328 ( 
.A(n_8),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_9),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_55)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_9),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_L g140 ( 
.A1(n_9),
.A2(n_57),
.B1(n_141),
.B2(n_144),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_9),
.A2(n_57),
.B1(n_156),
.B2(n_159),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g211 ( 
.A(n_9),
.B(n_212),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_10),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_10),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_11),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_12),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_12),
.Y(n_177)
);

BUFx4f_ASAP7_75t_L g187 ( 
.A(n_12),
.Y(n_187)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_12),
.Y(n_191)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_13),
.Y(n_231)
);

BUFx8_ASAP7_75t_L g258 ( 
.A(n_13),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_517),
.Y(n_17)
);

OAI221xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_61),
.B1(n_65),
.B2(n_275),
.C(n_511),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_19),
.B(n_61),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_20),
.B(n_274),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_20),
.B(n_274),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_41),
.Y(n_20)
);

NAND2xp33_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_32),
.Y(n_21)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_22),
.B(n_43),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B(n_28),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_23),
.B(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_23),
.B(n_221),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_R g300 ( 
.A(n_23),
.B(n_33),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_23),
.B(n_345),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_23),
.B(n_377),
.Y(n_376)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_27),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_28),
.A2(n_344),
.B1(n_347),
.B2(n_356),
.Y(n_343)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_32),
.B(n_55),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_32),
.B(n_226),
.Y(n_359)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_44),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_33),
.A2(n_63),
.B(n_64),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_33),
.A2(n_63),
.B1(n_64),
.B2(n_225),
.Y(n_224)
);

OAI21xp33_ASAP7_75t_SL g250 ( 
.A1(n_33),
.A2(n_41),
.B(n_251),
.Y(n_250)
);

OA22x2_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_36),
.B1(n_38),
.B2(n_40),
.Y(n_33)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_34),
.Y(n_346)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_35),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_35),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_35),
.Y(n_143)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_39),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_42),
.B(n_359),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_55),
.Y(n_42)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_43),
.B(n_226),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_45),
.A2(n_46),
.B1(n_50),
.B2(n_54),
.Y(n_44)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_57),
.B(n_295),
.Y(n_294)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_SL g227 ( 
.A(n_60),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_61),
.A2(n_164),
.B(n_201),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_62),
.A2(n_166),
.B1(n_201),
.B2(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_62),
.Y(n_238)
);

OAI21x1_ASAP7_75t_R g267 ( 
.A1(n_63),
.A2(n_73),
.B(n_251),
.Y(n_267)
);

NAND3xp33_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_262),
.C(n_273),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_239),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_68),
.B(n_202),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_68),
.B(n_202),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_163),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_70),
.A2(n_71),
.B1(n_146),
.B2(n_147),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_71),
.B(n_146),
.C(n_163),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_75),
.Y(n_71)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_72),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_72),
.A2(n_242),
.B1(n_244),
.B2(n_260),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_72),
.B(n_244),
.C(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_74),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_73),
.B(n_463),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_74),
.B(n_359),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_76),
.A2(n_77),
.B1(n_108),
.B2(n_145),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_76),
.A2(n_77),
.B1(n_246),
.B2(n_247),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_76),
.A2(n_77),
.B1(n_361),
.B2(n_362),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_76),
.B(n_358),
.C(n_362),
.Y(n_480)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_R g241 ( 
.A(n_77),
.B(n_108),
.C(n_242),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_77),
.B(n_247),
.C(n_249),
.Y(n_272)
);

OA21x2_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_89),
.B(n_101),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_78),
.B(n_101),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_78),
.B(n_155),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_78),
.B(n_194),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_78),
.B(n_326),
.Y(n_388)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

AND2x2_ASAP7_75t_SL g89 ( 
.A(n_79),
.B(n_90),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_81),
.B1(n_83),
.B2(n_87),
.Y(n_79)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_82),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_82),
.Y(n_340)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_82),
.Y(n_398)
);

OAI22xp33_ASAP7_75t_L g90 ( 
.A1(n_83),
.A2(n_91),
.B1(n_94),
.B2(n_97),
.Y(n_90)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_89),
.B(n_155),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_89),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_89),
.B(n_326),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_89),
.B(n_101),
.Y(n_389)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_93),
.Y(n_158)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_93),
.Y(n_162)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_100),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g321 ( 
.A(n_107),
.Y(n_321)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_108),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_120),
.B(n_139),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_109),
.Y(n_149)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_114),
.Y(n_118)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx8_ASAP7_75t_L g287 ( 
.A(n_118),
.Y(n_287)
);

NOR2x1_ASAP7_75t_L g215 ( 
.A(n_120),
.B(n_216),
.Y(n_215)
);

AOI21x1_ASAP7_75t_L g268 ( 
.A1(n_120),
.A2(n_216),
.B(n_269),
.Y(n_268)
);

INVx2_ASAP7_75t_SL g120 ( 
.A(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_121),
.B(n_140),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_121),
.B(n_283),
.Y(n_282)
);

NOR2x1_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_132),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_125),
.B1(n_127),
.B2(n_130),
.Y(n_122)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_123),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_128),
.Y(n_315)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_128),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_130),
.Y(n_306)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_131),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_132),
.B(n_140),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_132),
.A2(n_149),
.B(n_150),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_132),
.B(n_217),
.Y(n_248)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_132),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_132),
.B(n_283),
.Y(n_363)
);

AO22x2_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_135),
.B1(n_136),
.B2(n_137),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_135),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_139),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_139),
.B(n_282),
.Y(n_281)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_143),
.Y(n_219)
);

INVx6_ASAP7_75t_L g356 ( 
.A(n_144),
.Y(n_356)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

OA21x2_ASAP7_75t_L g232 ( 
.A1(n_147),
.A2(n_148),
.B(n_152),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_152),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_151),
.B(n_248),
.Y(n_247)
);

AND2x4_ASAP7_75t_SL g362 ( 
.A(n_151),
.B(n_363),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_154),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_153),
.Y(n_324)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_154),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_154),
.B(n_440),
.Y(n_439)
);

BUFx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_157),
.Y(n_195)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_164),
.A2(n_165),
.B1(n_236),
.B2(n_237),
.Y(n_235)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_192),
.Y(n_165)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_166),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_166),
.B(n_302),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_166),
.A2(n_201),
.B1(n_302),
.B2(n_445),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_166),
.A2(n_192),
.B1(n_201),
.B2(n_493),
.Y(n_492)
);

OA21x2_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_172),
.B(n_182),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx4_ASAP7_75t_SL g209 ( 
.A(n_169),
.Y(n_209)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_169),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_171),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_173),
.B(n_211),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_173),
.B(n_183),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_173),
.B(n_395),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_SL g470 ( 
.A1(n_173),
.A2(n_336),
.B(n_471),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_178),
.Y(n_173)
);

BUFx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_176),
.Y(n_339)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g375 ( 
.A(n_177),
.Y(n_375)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_178),
.Y(n_393)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_181),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_182),
.A2(n_208),
.B(n_210),
.Y(n_207)
);

AO21x1_ASAP7_75t_L g391 ( 
.A1(n_182),
.A2(n_392),
.B(n_394),
.Y(n_391)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_186),
.Y(n_379)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_187),
.Y(n_212)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_189),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx3_ASAP7_75t_L g414 ( 
.A(n_190),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_191),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g493 ( 
.A(n_192),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_199),
.B(n_200),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_200),
.B(n_325),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_200),
.B(n_389),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_232),
.C(n_233),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_203),
.B(n_502),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_213),
.C(n_223),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_204),
.B(n_495),
.Y(n_494)
);

AOI21x1_ASAP7_75t_SL g204 ( 
.A1(n_205),
.A2(n_206),
.B(n_207),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_205),
.B(n_206),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_207),
.B(n_466),
.Y(n_465)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_210),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_211),
.A2(n_293),
.B(n_296),
.Y(n_292)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_214),
.B(n_224),
.Y(n_495)
);

NOR2xp67_ASAP7_75t_SL g214 ( 
.A(n_215),
.B(n_222),
.Y(n_214)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_215),
.Y(n_443)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_220),
.Y(n_217)
);

OAI32xp33_ASAP7_75t_L g302 ( 
.A1(n_220),
.A2(n_303),
.A3(n_307),
.B1(n_312),
.B2(n_316),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx5_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

BUFx12f_ASAP7_75t_L g253 ( 
.A(n_231),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g502 ( 
.A1(n_232),
.A2(n_234),
.B1(n_235),
.B2(n_503),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_232),
.Y(n_503)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g512 ( 
.A1(n_239),
.A2(n_513),
.B(n_514),
.Y(n_512)
);

NOR2xp67_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_261),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_240),
.B(n_261),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_243),
.Y(n_240)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_241),
.Y(n_264)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_244),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_245),
.A2(n_249),
.B1(n_250),
.B2(n_259),
.Y(n_244)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_245),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_247),
.Y(n_246)
);

AND2x4_ASAP7_75t_SL g460 ( 
.A(n_248),
.B(n_282),
.Y(n_460)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g511 ( 
.A1(n_262),
.A2(n_273),
.B(n_512),
.C(n_515),
.D(n_516),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_263),
.B(n_265),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_263),
.B(n_265),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_272),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_267),
.A2(n_268),
.B1(n_270),
.B2(n_271),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_267),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_267),
.B(n_271),
.C(n_272),
.Y(n_274)
);

INVx2_ASAP7_75t_SL g271 ( 
.A(n_268),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_268),
.A2(n_271),
.B1(n_473),
.B2(n_474),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_271),
.B(n_468),
.C(n_474),
.Y(n_490)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

AO221x1_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_454),
.B1(n_504),
.B2(n_509),
.C(n_510),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_364),
.B(n_453),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_329),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_279),
.B(n_329),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_301),
.C(n_322),
.Y(n_279)
);

XOR2x1_ASAP7_75t_L g448 ( 
.A(n_280),
.B(n_449),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_281),
.B(n_288),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_281),
.B(n_289),
.C(n_300),
.Y(n_332)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_289),
.A2(n_290),
.B1(n_299),
.B2(n_300),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g418 ( 
.A(n_291),
.B(n_419),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_SL g424 ( 
.A(n_292),
.B(n_394),
.Y(n_424)
);

INVxp67_ASAP7_75t_L g471 ( 
.A(n_292),
.Y(n_471)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx6_ASAP7_75t_L g341 ( 
.A(n_298),
.Y(n_341)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_301),
.A2(n_322),
.B1(n_323),
.B2(n_450),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_301),
.Y(n_450)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_302),
.Y(n_445)
);

INVx1_ASAP7_75t_SL g303 ( 
.A(n_304),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_310),
.Y(n_372)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_320),
.Y(n_316)
);

HB1xp67_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_325),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_357),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_331),
.A2(n_332),
.B1(n_333),
.B2(n_334),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_331),
.B(n_334),
.C(n_357),
.Y(n_483)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_343),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_335),
.B(n_343),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_336),
.A2(n_341),
.B(n_342),
.Y(n_335)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

HB1xp67_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_342),
.B(n_429),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_352),
.Y(n_347)
);

INVx2_ASAP7_75t_SL g348 ( 
.A(n_349),
.Y(n_348)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx4_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx3_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_360),
.Y(n_357)
);

CKINVDCx16_ASAP7_75t_R g361 ( 
.A(n_362),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_363),
.B(n_443),
.Y(n_442)
);

AOI21x1_ASAP7_75t_SL g364 ( 
.A1(n_365),
.A2(n_447),
.B(n_452),
.Y(n_364)
);

OAI21x1_ASAP7_75t_L g365 ( 
.A1(n_366),
.A2(n_433),
.B(n_446),
.Y(n_365)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_367),
.A2(n_408),
.B(n_432),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_390),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_368),
.B(n_390),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_387),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_369),
.B(n_387),
.Y(n_430)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

BUFx3_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

BUFx3_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_384),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx5_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

BUFx2_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_389),
.Y(n_387)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_388),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_403),
.Y(n_390)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_391),
.Y(n_435)
);

BUFx2_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_395),
.B(n_420),
.Y(n_419)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_404),
.A2(n_405),
.B1(n_406),
.B2(n_407),
.Y(n_403)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_404),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_405),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_405),
.B(n_406),
.C(n_435),
.Y(n_434)
);

OAI21xp5_ASAP7_75t_L g408 ( 
.A1(n_409),
.A2(n_427),
.B(n_431),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_L g409 ( 
.A1(n_410),
.A2(n_423),
.B(n_426),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_418),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_415),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_419),
.Y(n_429)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

HB1xp67_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_424),
.B(n_425),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_424),
.B(n_425),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_430),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_428),
.B(n_430),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_436),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_434),
.B(n_436),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_444),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_438),
.A2(n_439),
.B1(n_441),
.B2(n_442),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_438),
.B(n_442),
.C(n_444),
.Y(n_451)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_448),
.B(n_451),
.Y(n_447)
);

NOR2xp67_ASAP7_75t_L g452 ( 
.A(n_448),
.B(n_451),
.Y(n_452)
);

NOR3xp33_ASAP7_75t_L g454 ( 
.A(n_455),
.B(n_486),
.C(n_498),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_456),
.B(n_482),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_456),
.B(n_507),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_457),
.B(n_475),
.Y(n_456)
);

OR2x2_ASAP7_75t_L g505 ( 
.A(n_457),
.B(n_475),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_458),
.B(n_464),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_458),
.B(n_465),
.C(n_488),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_460),
.C(n_461),
.Y(n_458)
);

XOR2x1_ASAP7_75t_SL g477 ( 
.A(n_459),
.B(n_478),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_460),
.A2(n_461),
.B1(n_462),
.B2(n_479),
.Y(n_478)
);

CKINVDCx16_ASAP7_75t_R g479 ( 
.A(n_460),
.Y(n_479)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_467),
.Y(n_464)
);

HB1xp67_ASAP7_75t_L g488 ( 
.A(n_467),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_468),
.B(n_472),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_470),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_469),
.B(n_470),
.Y(n_481)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_473),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_480),
.C(n_481),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_477),
.B(n_485),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_480),
.B(n_481),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_483),
.B(n_484),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_483),
.B(n_484),
.Y(n_507)
);

A2O1A1Ixp33_ASAP7_75t_L g504 ( 
.A1(n_486),
.A2(n_505),
.B(n_506),
.C(n_508),
.Y(n_504)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_487),
.B(n_489),
.Y(n_486)
);

OR2x2_ASAP7_75t_L g508 ( 
.A(n_487),
.B(n_489),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_490),
.B(n_491),
.Y(n_489)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_490),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_L g491 ( 
.A1(n_492),
.A2(n_494),
.B1(n_496),
.B2(n_497),
.Y(n_491)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_492),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_492),
.B(n_496),
.C(n_500),
.Y(n_499)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_494),
.Y(n_496)
);

INVxp67_ASAP7_75t_L g509 ( 
.A(n_498),
.Y(n_509)
);

NOR2x1_ASAP7_75t_L g498 ( 
.A(n_499),
.B(n_501),
.Y(n_498)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_499),
.B(n_501),
.Y(n_510)
);


endmodule