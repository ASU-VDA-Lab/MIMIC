module fake_jpeg_240_n_70 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_70);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_70;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_15;
wire n_66;

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_7),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_7),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_8),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_5),
.B(n_0),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_3),
.B(n_0),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

AOI22xp33_ASAP7_75t_SL g19 ( 
.A1(n_16),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_19),
.A2(n_22),
.B1(n_11),
.B2(n_9),
.Y(n_31)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_13),
.B(n_1),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_21),
.B(n_24),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g22 ( 
.A1(n_14),
.A2(n_5),
.B1(n_6),
.B2(n_16),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_13),
.B(n_6),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_17),
.B(n_10),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_25),
.B(n_18),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_25),
.B(n_17),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_28),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_21),
.B(n_11),
.Y(n_30)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_24),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_31),
.A2(n_23),
.B1(n_9),
.B2(n_19),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_20),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_32),
.Y(n_38)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_33),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_41),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_SL g50 ( 
.A1(n_39),
.A2(n_15),
.B(n_26),
.Y(n_50)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_12),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_31),
.A2(n_23),
.B1(n_12),
.B2(n_15),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_42),
.B(n_32),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_43),
.B(n_47),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_46),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_38),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_30),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_48),
.B(n_26),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_50),
.A2(n_42),
.B(n_34),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g57 ( 
.A(n_53),
.B(n_50),
.Y(n_57)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_56),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_55),
.B(n_44),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_49),
.B(n_37),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_57),
.B(n_53),
.C(n_52),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_58),
.B(n_59),
.Y(n_63)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_61),
.B(n_62),
.Y(n_64)
);

BUFx24_ASAP7_75t_SL g62 ( 
.A(n_60),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_63),
.B(n_45),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_65),
.B(n_45),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_66),
.B(n_67),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_64),
.B(n_57),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_68),
.B(n_43),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_69),
.B(n_40),
.Y(n_70)
);


endmodule