module fake_jpeg_21890_n_232 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_232);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_232;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_4),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_17),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_36),
.Y(n_44)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g36 ( 
.A(n_17),
.B(n_0),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_37),
.A2(n_31),
.B1(n_22),
.B2(n_21),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_19),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_40),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_23),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_30),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_42),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_2),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_16),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_48),
.A2(n_35),
.B1(n_40),
.B2(n_20),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_41),
.A2(n_31),
.B1(n_22),
.B2(n_16),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_49),
.A2(n_55),
.B1(n_58),
.B2(n_59),
.Y(n_83)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx3_ASAP7_75t_SL g79 ( 
.A(n_50),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_53),
.B(n_39),
.Y(n_76)
);

CKINVDCx9p33_ASAP7_75t_R g54 ( 
.A(n_42),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_37),
.A2(n_22),
.B1(n_16),
.B2(n_21),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_36),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_37),
.A2(n_21),
.B1(n_18),
.B2(n_20),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_37),
.A2(n_23),
.B1(n_30),
.B2(n_28),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

A2O1A1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_43),
.A2(n_30),
.B(n_28),
.C(n_32),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_61),
.B(n_56),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_62),
.B(n_80),
.Y(n_91)
);

NAND3xp33_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_41),
.C(n_42),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_63),
.B(n_69),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_36),
.Y(n_64)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_64),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_34),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_65),
.B(n_66),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_47),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

BUFx24_ASAP7_75t_L g92 ( 
.A(n_67),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_68),
.A2(n_71),
.B1(n_45),
.B2(n_46),
.Y(n_93)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_61),
.A2(n_40),
.B1(n_35),
.B2(n_38),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_36),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_72),
.B(n_75),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_73),
.A2(n_77),
.B(n_24),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_52),
.B(n_38),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_76),
.B(n_78),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_61),
.A2(n_18),
.B1(n_27),
.B2(n_26),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_58),
.B(n_55),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_51),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_45),
.B(n_34),
.Y(n_82)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_45),
.B(n_29),
.Y(n_84)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_51),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_26),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_87),
.B(n_90),
.Y(n_117)
);

O2A1O1Ixp33_ASAP7_75t_L g88 ( 
.A1(n_78),
.A2(n_48),
.B(n_59),
.C(n_50),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_88),
.A2(n_97),
.B1(n_101),
.B2(n_60),
.Y(n_135)
);

OAI21xp33_ASAP7_75t_L g115 ( 
.A1(n_89),
.A2(n_105),
.B(n_108),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_76),
.B(n_52),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_93),
.A2(n_83),
.B1(n_72),
.B2(n_62),
.Y(n_119)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_96),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_77),
.B(n_19),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_100),
.B(n_106),
.Y(n_114)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_101),
.B(n_102),
.Y(n_134)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_67),
.Y(n_102)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_67),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_104),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_76),
.B(n_46),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_65),
.B(n_29),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_65),
.B(n_27),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_107),
.B(n_87),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_66),
.A2(n_24),
.B(n_25),
.Y(n_108)
);

CKINVDCx5p33_ASAP7_75t_R g110 ( 
.A(n_86),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_110),
.Y(n_120)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_80),
.Y(n_111)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_111),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_96),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_116),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_109),
.A2(n_73),
.B(n_83),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_118),
.A2(n_122),
.B(n_128),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_119),
.A2(n_126),
.B1(n_97),
.B2(n_94),
.Y(n_141)
);

OAI21xp33_ASAP7_75t_L g122 ( 
.A1(n_105),
.A2(n_63),
.B(n_75),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_109),
.B(n_76),
.C(n_46),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_131),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_92),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_124),
.Y(n_152)
);

AND2x6_ASAP7_75t_L g125 ( 
.A(n_95),
.B(n_50),
.Y(n_125)
);

NAND3xp33_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_103),
.C(n_98),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_93),
.A2(n_60),
.B1(n_81),
.B2(n_85),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_127),
.B(n_129),
.Y(n_156)
);

O2A1O1Ixp33_ASAP7_75t_L g128 ( 
.A1(n_90),
.A2(n_99),
.B(n_91),
.C(n_103),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_92),
.Y(n_129)
);

OA21x2_ASAP7_75t_L g130 ( 
.A1(n_88),
.A2(n_39),
.B(n_54),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_130),
.A2(n_70),
.B(n_84),
.Y(n_151)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_111),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_91),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_108),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_110),
.Y(n_133)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_133),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_135),
.A2(n_81),
.B1(n_70),
.B2(n_69),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_118),
.A2(n_89),
.B1(n_99),
.B2(n_100),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_138),
.A2(n_148),
.B1(n_153),
.B2(n_133),
.Y(n_164)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_134),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_140),
.B(n_149),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_141),
.A2(n_147),
.B1(n_112),
.B2(n_120),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_142),
.B(n_155),
.Y(n_165)
);

NAND3xp33_ASAP7_75t_L g143 ( 
.A(n_132),
.B(n_98),
.C(n_94),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_143),
.B(n_146),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_119),
.B(n_107),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_144),
.B(n_114),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_145),
.B(n_154),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_113),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_126),
.A2(n_128),
.B1(n_130),
.B2(n_123),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_135),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_151),
.A2(n_157),
.B(n_158),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_125),
.A2(n_106),
.B1(n_74),
.B2(n_87),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_117),
.B(n_74),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_121),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_121),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_117),
.B(n_92),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_137),
.B(n_115),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_159),
.B(n_166),
.C(n_168),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_137),
.A2(n_130),
.B(n_116),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_160),
.A2(n_169),
.B(n_171),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_138),
.B(n_127),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_161),
.B(n_163),
.Y(n_185)
);

AOI221xp5_ASAP7_75t_L g188 ( 
.A1(n_162),
.A2(n_158),
.B1(n_150),
.B2(n_157),
.C(n_28),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_164),
.A2(n_141),
.B1(n_154),
.B2(n_158),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_136),
.B(n_112),
.C(n_131),
.Y(n_166)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_146),
.Y(n_167)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_167),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_136),
.B(n_129),
.C(n_124),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_139),
.B(n_120),
.Y(n_169)
);

CKINVDCx14_ASAP7_75t_R g170 ( 
.A(n_156),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_170),
.B(n_173),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_139),
.A2(n_151),
.B(n_152),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_145),
.B(n_114),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_147),
.A2(n_113),
.B(n_25),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_175),
.A2(n_150),
.B(n_92),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_168),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_178),
.B(n_179),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_162),
.A2(n_153),
.B1(n_152),
.B2(n_155),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_180),
.B(n_187),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_164),
.A2(n_171),
.B1(n_174),
.B2(n_160),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_181),
.A2(n_182),
.B(n_30),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_159),
.B(n_144),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_186),
.B(n_188),
.Y(n_196)
);

BUFx12_ASAP7_75t_L g187 ( 
.A(n_169),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_165),
.A2(n_172),
.B1(n_176),
.B2(n_166),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_189),
.B(n_192),
.Y(n_197)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_169),
.Y(n_192)
);

OAI21x1_ASAP7_75t_L g194 ( 
.A1(n_180),
.A2(n_177),
.B(n_175),
.Y(n_194)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_194),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_190),
.A2(n_172),
.B(n_176),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_195),
.A2(n_200),
.B1(n_202),
.B2(n_203),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_184),
.B(n_161),
.C(n_163),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_198),
.B(n_199),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_184),
.B(n_104),
.C(n_102),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_178),
.A2(n_79),
.B(n_15),
.Y(n_202)
);

NOR2x1_ASAP7_75t_L g203 ( 
.A(n_183),
.B(n_79),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_198),
.B(n_185),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_205),
.B(n_208),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_197),
.A2(n_190),
.B1(n_191),
.B2(n_189),
.Y(n_206)
);

AOI322xp5_ASAP7_75t_L g214 ( 
.A1(n_206),
.A2(n_203),
.A3(n_187),
.B1(n_15),
.B2(n_28),
.C1(n_79),
.C2(n_8),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_196),
.B(n_185),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_201),
.B(n_182),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_210),
.B(n_211),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_196),
.B(n_186),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_199),
.B(n_187),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_212),
.B(n_13),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_209),
.A2(n_193),
.B(n_195),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_213),
.A2(n_211),
.B(n_204),
.Y(n_220)
);

AOI31xp33_ASAP7_75t_L g221 ( 
.A1(n_214),
.A2(n_219),
.A3(n_5),
.B(n_6),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_216),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_207),
.A2(n_2),
.B(n_4),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_217),
.A2(n_7),
.B(n_9),
.Y(n_223)
);

AOI322xp5_ASAP7_75t_L g219 ( 
.A1(n_208),
.A2(n_4),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_9),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_220),
.A2(n_219),
.B(n_10),
.Y(n_226)
);

OAI21x1_ASAP7_75t_L g228 ( 
.A1(n_221),
.A2(n_7),
.B(n_10),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_215),
.A2(n_204),
.B(n_205),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_222),
.B(n_223),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_224),
.B(n_218),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_225),
.B(n_226),
.Y(n_230)
);

AOI322xp5_ASAP7_75t_L g229 ( 
.A1(n_228),
.A2(n_10),
.A3(n_11),
.B1(n_12),
.B2(n_221),
.C1(n_100),
.C2(n_115),
.Y(n_229)
);

MAJx2_ASAP7_75t_L g231 ( 
.A(n_229),
.B(n_227),
.C(n_11),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_231),
.B(n_230),
.Y(n_232)
);


endmodule