module real_jpeg_9063_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_282, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_282;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_238;
wire n_76;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_268;
wire n_42;
wire n_112;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_277;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_187;
wire n_75;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_216;
wire n_128;
wire n_202;
wire n_179;
wire n_167;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_273;
wire n_269;
wire n_89;

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_1),
.A2(n_30),
.B1(n_31),
.B2(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_1),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_1),
.A2(n_44),
.B1(n_45),
.B2(n_50),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_1),
.A2(n_50),
.B1(n_56),
.B2(n_57),
.Y(n_92)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_2),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_2),
.A2(n_27),
.B1(n_30),
.B2(n_31),
.Y(n_29)
);

AOI21xp33_ASAP7_75t_L g198 ( 
.A1(n_2),
.A2(n_11),
.B(n_31),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_3),
.A2(n_26),
.B1(n_33),
.B2(n_34),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_3),
.A2(n_30),
.B1(n_31),
.B2(n_34),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_3),
.A2(n_34),
.B1(n_56),
.B2(n_57),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_3),
.A2(n_34),
.B1(n_44),
.B2(n_45),
.Y(n_212)
);

BUFx10_ASAP7_75t_L g73 ( 
.A(n_4),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_5),
.Y(n_57)
);

A2O1A1Ixp33_ASAP7_75t_SL g53 ( 
.A1(n_6),
.A2(n_44),
.B(n_54),
.C(n_55),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_6),
.B(n_44),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_6),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_55)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_6),
.Y(n_58)
);

BUFx6f_ASAP7_75t_SL g41 ( 
.A(n_7),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_9),
.A2(n_44),
.B1(n_45),
.B2(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_9),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_9),
.A2(n_56),
.B1(n_57),
.B2(n_60),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_10),
.A2(n_26),
.B1(n_33),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_10),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_10),
.A2(n_30),
.B1(n_31),
.B2(n_36),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_10),
.A2(n_36),
.B1(n_44),
.B2(n_45),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_10),
.A2(n_36),
.B1(n_56),
.B2(n_57),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_11),
.A2(n_44),
.B(n_122),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_11),
.B(n_44),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_11),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_11),
.A2(n_71),
.B1(n_74),
.B2(n_133),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_11),
.A2(n_30),
.B(n_158),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_11),
.B(n_30),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_11),
.B(n_179),
.Y(n_178)
);

OAI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_11),
.A2(n_26),
.B1(n_33),
.B2(n_135),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_12),
.A2(n_44),
.B1(n_45),
.B2(n_124),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_12),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_12),
.A2(n_56),
.B1(n_57),
.B2(n_124),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_12),
.A2(n_30),
.B1(n_31),
.B2(n_124),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_12),
.A2(n_26),
.B1(n_33),
.B2(n_124),
.Y(n_220)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_14),
.A2(n_30),
.B1(n_31),
.B2(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_14),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_14),
.A2(n_44),
.B1(n_45),
.B2(n_48),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_14),
.A2(n_48),
.B1(n_56),
.B2(n_57),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_15),
.A2(n_26),
.B1(n_33),
.B2(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_15),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_15),
.A2(n_56),
.B1(n_57),
.B2(n_98),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_15),
.A2(n_44),
.B1(n_45),
.B2(n_98),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_15),
.A2(n_30),
.B1(n_31),
.B2(n_98),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_16),
.A2(n_26),
.B1(n_33),
.B2(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_16),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_16),
.A2(n_56),
.B1(n_57),
.B2(n_81),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_16),
.A2(n_44),
.B1(n_45),
.B2(n_81),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_16),
.A2(n_30),
.B1(n_31),
.B2(n_81),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_17),
.A2(n_56),
.B1(n_57),
.B2(n_115),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_17),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_17),
.A2(n_44),
.B1(n_45),
.B2(n_115),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_17),
.A2(n_30),
.B1(n_31),
.B2(n_115),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_17),
.A2(n_26),
.B1(n_33),
.B2(n_115),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_104),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_102),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_82),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_21),
.B(n_82),
.Y(n_103)
);

BUFx24_ASAP7_75t_SL g281 ( 
.A(n_21),
.Y(n_281)
);

FAx1_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_62),
.CI(n_67),
.CON(n_21),
.SN(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_37),
.B2(n_38),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_29),
.B1(n_32),
.B2(n_35),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_25),
.A2(n_29),
.B1(n_32),
.B2(n_80),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_25),
.A2(n_29),
.B1(n_80),
.B2(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_25),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_25),
.A2(n_29),
.B1(n_231),
.B2(n_232),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_25),
.A2(n_29),
.B1(n_97),
.B2(n_232),
.Y(n_249)
);

A2O1A1Ixp33_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B(n_28),
.C(n_29),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_26),
.B(n_27),
.Y(n_28)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

A2O1A1Ixp33_ASAP7_75t_L g197 ( 
.A1(n_26),
.A2(n_27),
.B(n_135),
.C(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_29),
.Y(n_179)
);

A2O1A1Ixp33_ASAP7_75t_L g40 ( 
.A1(n_30),
.A2(n_41),
.B(n_42),
.C(n_43),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_41),
.Y(n_42)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_51),
.B1(n_52),
.B2(n_61),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_39),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_40),
.A2(n_43),
.B1(n_47),
.B2(n_49),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_40),
.A2(n_43),
.B1(n_47),
.B2(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_40),
.A2(n_43),
.B1(n_64),
.B2(n_101),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_40),
.A2(n_43),
.B1(n_157),
.B2(n_159),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_40),
.A2(n_43),
.B1(n_159),
.B2(n_175),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_40),
.A2(n_43),
.B1(n_175),
.B2(n_216),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_40),
.A2(n_43),
.B1(n_216),
.B2(n_228),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_40),
.A2(n_43),
.B1(n_101),
.B2(n_228),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_41),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_41),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_42),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_43),
.B(n_135),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_44),
.B(n_46),
.Y(n_163)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_45),
.A2(n_162),
.B1(n_163),
.B2(n_164),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_53),
.A2(n_55),
.B(n_59),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_53),
.A2(n_55),
.B1(n_59),
.B2(n_66),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_53),
.A2(n_55),
.B1(n_66),
.B2(n_77),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_53),
.A2(n_55),
.B1(n_77),
.B2(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_53),
.A2(n_55),
.B1(n_121),
.B2(n_123),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_53),
.A2(n_55),
.B1(n_123),
.B2(n_148),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_53),
.A2(n_55),
.B1(n_148),
.B2(n_155),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_53),
.A2(n_55),
.B1(n_155),
.B2(n_187),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_53),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_53),
.A2(n_55),
.B1(n_94),
.B2(n_238),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_54),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_55),
.B(n_135),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_55),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_73),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_56),
.B(n_58),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_56),
.B(n_139),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_57),
.A2(n_126),
.B1(n_127),
.B2(n_128),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_62),
.A2(n_63),
.B(n_65),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_65),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_78),
.B(n_79),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_68),
.A2(n_69),
.B1(n_84),
.B2(n_85),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_76),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_70),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_70),
.A2(n_78),
.B1(n_79),
.B2(n_86),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_70),
.A2(n_76),
.B1(n_78),
.B2(n_263),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_74),
.B(n_75),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_71),
.A2(n_74),
.B1(n_75),
.B2(n_92),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_71),
.A2(n_74),
.B1(n_114),
.B2(n_133),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_71),
.A2(n_74),
.B1(n_117),
.B2(n_150),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_71),
.A2(n_74),
.B1(n_150),
.B2(n_166),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_71),
.A2(n_74),
.B1(n_201),
.B2(n_202),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_71),
.A2(n_74),
.B1(n_92),
.B2(n_202),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_72),
.A2(n_73),
.B1(n_113),
.B2(n_116),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_72),
.A2(n_73),
.B1(n_167),
.B2(n_181),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_73),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_74),
.B(n_135),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_76),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_79),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_87),
.C(n_88),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_83),
.B(n_87),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_88),
.A2(n_89),
.B1(n_266),
.B2(n_267),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_95),
.C(n_99),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_90),
.B(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_93),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_91),
.B(n_93),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_95),
.A2(n_96),
.B1(n_99),
.B2(n_100),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

AOI321xp33_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_257),
.A3(n_268),
.B1(n_274),
.B2(n_279),
.C(n_282),
.Y(n_104)
);

NOR3xp33_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_222),
.C(n_253),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_191),
.B(n_221),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_108),
.A2(n_169),
.B(n_190),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_152),
.B(n_168),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_110),
.A2(n_142),
.B(n_151),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_130),
.B(n_141),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_118),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_112),
.B(n_118),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_119),
.A2(n_120),
.B1(n_125),
.B2(n_129),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_119),
.B(n_129),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_122),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_125),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_136),
.B(n_140),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_134),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_132),
.B(n_134),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_137),
.B(n_138),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_144),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_143),
.B(n_144),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_145),
.B(n_153),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_145),
.B(n_153),
.Y(n_168)
);

FAx1_ASAP7_75t_SL g145 ( 
.A(n_146),
.B(n_147),
.CI(n_149),
.CON(n_145),
.SN(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_153),
.Y(n_170)
);

FAx1_ASAP7_75t_SL g153 ( 
.A(n_154),
.B(n_156),
.CI(n_160),
.CON(n_153),
.SN(n_153)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_158),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_165),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_161),
.B(n_165),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_170),
.B(n_171),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_173),
.B1(n_183),
.B2(n_184),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_172),
.B(n_186),
.C(n_188),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_176),
.B1(n_177),
.B2(n_182),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_174),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_180),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_178),
.B(n_180),
.C(n_182),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_179),
.A2(n_218),
.B1(n_219),
.B2(n_220),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_181),
.Y(n_201)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_185),
.A2(n_186),
.B1(n_188),
.B2(n_189),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_185),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_186),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_187),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_192),
.B(n_193),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_206),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_203),
.B1(n_204),
.B2(n_205),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_195),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_195),
.B(n_205),
.C(n_206),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_197),
.B1(n_199),
.B2(n_200),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_196),
.B(n_200),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_197),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_200),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_203),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_217),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_209),
.B1(n_214),
.B2(n_215),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_209),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_209),
.B(n_214),
.C(n_217),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_211),
.B1(n_212),
.B2(n_213),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_212),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_215),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_220),
.Y(n_231)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

AOI21xp33_ASAP7_75t_L g275 ( 
.A1(n_223),
.A2(n_276),
.B(n_277),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_240),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_224),
.B(n_240),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_235),
.C(n_239),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_225),
.B(n_256),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_226),
.B(n_234),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_227),
.A2(n_229),
.B1(n_230),
.B2(n_233),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_227),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_SL g251 ( 
.A(n_229),
.B(n_233),
.C(n_234),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_230),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_235),
.B(n_239),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_236),
.B(n_237),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_241),
.A2(n_242),
.B1(n_251),
.B2(n_252),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_242),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_243),
.B(n_244),
.C(n_252),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_245),
.B(n_248),
.C(n_250),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_247),
.A2(n_248),
.B1(n_249),
.B2(n_250),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_247),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_249),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_251),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_254),
.B(n_255),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_265),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_258),
.B(n_265),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_262),
.C(n_264),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_259),
.A2(n_260),
.B1(n_262),
.B2(n_273),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_260),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_262),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_264),
.B(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_269),
.A2(n_275),
.B(n_278),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_270),
.B(n_271),
.Y(n_278)
);


endmodule