module fake_netlist_5_1059_n_70 (n_16, n_0, n_12, n_9, n_18, n_1, n_8, n_10, n_4, n_11, n_17, n_19, n_7, n_15, n_20, n_5, n_14, n_2, n_13, n_3, n_6, n_70);

input n_16;
input n_0;
input n_12;
input n_9;
input n_18;
input n_1;
input n_8;
input n_10;
input n_4;
input n_11;
input n_17;
input n_19;
input n_7;
input n_15;
input n_20;
input n_5;
input n_14;
input n_2;
input n_13;
input n_3;
input n_6;

output n_70;

wire n_54;
wire n_29;
wire n_43;
wire n_47;
wire n_58;
wire n_67;
wire n_69;
wire n_36;
wire n_25;
wire n_53;
wire n_27;
wire n_42;
wire n_64;
wire n_22;
wire n_45;
wire n_24;
wire n_46;
wire n_28;
wire n_21;
wire n_44;
wire n_40;
wire n_34;
wire n_62;
wire n_38;
wire n_61;
wire n_68;
wire n_32;
wire n_41;
wire n_35;
wire n_65;
wire n_56;
wire n_51;
wire n_63;
wire n_57;
wire n_37;
wire n_59;
wire n_26;
wire n_30;
wire n_33;
wire n_55;
wire n_48;
wire n_31;
wire n_23;
wire n_50;
wire n_66;
wire n_49;
wire n_52;
wire n_60;
wire n_39;

BUFx3_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_19),
.Y(n_23)
);

CKINVDCx5p33_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

AND2x4_ASAP7_75t_L g25 ( 
.A(n_14),
.B(n_13),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

OA21x2_ASAP7_75t_L g28 ( 
.A1(n_3),
.A2(n_18),
.B(n_7),
.Y(n_28)
);

AND2x4_ASAP7_75t_L g29 ( 
.A(n_4),
.B(n_12),
.Y(n_29)
);

CKINVDCx5p33_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

OA21x2_ASAP7_75t_L g31 ( 
.A1(n_0),
.A2(n_10),
.B(n_1),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_2),
.B(n_1),
.Y(n_34)
);

NOR3xp33_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_15),
.C(n_17),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_21),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_21),
.B(n_27),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_34),
.A2(n_29),
.B1(n_25),
.B2(n_23),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_32),
.B(n_33),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

AND2x4_ASAP7_75t_L g41 ( 
.A(n_25),
.B(n_29),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

NOR2xp67_ASAP7_75t_L g44 ( 
.A(n_42),
.B(n_32),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_30),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_45),
.B(n_38),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_51),
.B(n_37),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_48),
.Y(n_53)
);

AND2x4_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_35),
.Y(n_54)
);

AND2x4_ASAP7_75t_SL g55 ( 
.A(n_50),
.B(n_23),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

NOR2xp67_ASAP7_75t_L g57 ( 
.A(n_53),
.B(n_36),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_52),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_56),
.Y(n_59)
);

OAI221xp5_ASAP7_75t_L g60 ( 
.A1(n_57),
.A2(n_53),
.B1(n_56),
.B2(n_39),
.C(n_30),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_60),
.Y(n_61)
);

NOR3xp33_ASAP7_75t_L g62 ( 
.A(n_60),
.B(n_58),
.C(n_54),
.Y(n_62)
);

NAND4xp75_ASAP7_75t_L g63 ( 
.A(n_61),
.B(n_31),
.C(n_28),
.D(n_44),
.Y(n_63)
);

NOR2x1_ASAP7_75t_L g64 ( 
.A(n_62),
.B(n_59),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_64),
.A2(n_55),
.B1(n_54),
.B2(n_63),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_64),
.B(n_59),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_66),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_65),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_67),
.B(n_31),
.Y(n_69)
);

OR2x6_ASAP7_75t_L g70 ( 
.A(n_69),
.B(n_68),
.Y(n_70)
);


endmodule