module fake_jpeg_9220_n_62 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_62);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_62;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_27;
wire n_55;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_36;
wire n_31;
wire n_25;
wire n_56;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_32;

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx24_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_15),
.B(n_5),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_7),
.A2(n_3),
.B1(n_5),
.B2(n_21),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_26),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_37),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_29),
.A2(n_23),
.B1(n_10),
.B2(n_11),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_33),
.A2(n_30),
.B1(n_14),
.B2(n_17),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_27),
.B(n_0),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_2),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_24),
.B(n_1),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_4),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_1),
.Y(n_36)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_25),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_41),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_2),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_28),
.Y(n_42)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_46),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_4),
.Y(n_44)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_45),
.A2(n_6),
.B1(n_19),
.B2(n_20),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g47 ( 
.A1(n_35),
.A2(n_25),
.B(n_30),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_47),
.B(n_25),
.C(n_7),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_50),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_L g50 ( 
.A1(n_48),
.A2(n_8),
.B1(n_9),
.B2(n_12),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_53),
.B(n_45),
.C(n_46),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_56),
.B(n_49),
.C(n_52),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_58),
.B(n_54),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_L g60 ( 
.A1(n_59),
.A2(n_38),
.B(n_55),
.Y(n_60)
);

AOI21x1_ASAP7_75t_L g61 ( 
.A1(n_60),
.A2(n_40),
.B(n_57),
.Y(n_61)
);

OAI221xp5_ASAP7_75t_L g62 ( 
.A1(n_61),
.A2(n_47),
.B1(n_50),
.B2(n_39),
.C(n_51),
.Y(n_62)
);


endmodule