module real_aes_17163_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_800;
wire n_778;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_320;
wire n_884;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_889;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_874;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_142;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_649;
wire n_193;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_397;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_653;
wire n_290;
wire n_365;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_623;
wire n_249;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_888;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
AND2x4_ASAP7_75t_L g523 ( .A(n_0), .B(n_524), .Y(n_523) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_1), .A2(n_33), .B1(n_165), .B2(n_185), .Y(n_601) );
AOI22xp5_ASAP7_75t_L g650 ( .A1(n_2), .A2(n_9), .B1(n_562), .B2(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g524 ( .A(n_3), .Y(n_524) );
CKINVDCx5p33_ASAP7_75t_R g619 ( .A(n_4), .Y(n_619) );
AOI22xp5_ASAP7_75t_L g584 ( .A1(n_5), .A2(n_10), .B1(n_585), .B2(n_586), .Y(n_584) );
OR2x2_ASAP7_75t_L g115 ( .A(n_6), .B(n_28), .Y(n_115) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_7), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g653 ( .A(n_8), .Y(n_653) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_11), .B(n_170), .Y(n_196) );
AOI22xp5_ASAP7_75t_L g561 ( .A1(n_12), .A2(n_101), .B1(n_255), .B2(n_562), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g648 ( .A1(n_13), .A2(n_29), .B1(n_623), .B2(n_649), .Y(n_648) );
NAND2xp5_ASAP7_75t_SL g620 ( .A(n_14), .B(n_170), .Y(n_620) );
OAI21x1_ASAP7_75t_L g150 ( .A1(n_15), .A2(n_45), .B(n_151), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_16), .B(n_169), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g877 ( .A(n_17), .B(n_878), .Y(n_877) );
CKINVDCx5p33_ASAP7_75t_R g567 ( .A(n_18), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_19), .A2(n_37), .B1(n_136), .B2(n_261), .Y(n_602) );
CKINVDCx5p33_ASAP7_75t_R g239 ( .A(n_20), .Y(n_239) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_21), .A2(n_43), .B1(n_136), .B2(n_562), .Y(n_572) );
CKINVDCx5p33_ASAP7_75t_R g636 ( .A(n_22), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_23), .B(n_623), .Y(n_622) );
NAND2xp5_ASAP7_75t_SL g167 ( .A(n_24), .B(n_138), .Y(n_167) );
CKINVDCx5p33_ASAP7_75t_R g512 ( .A(n_25), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_26), .B(n_181), .Y(n_180) );
CKINVDCx5p33_ASAP7_75t_R g254 ( .A(n_27), .Y(n_254) );
AOI22xp5_ASAP7_75t_L g631 ( .A1(n_30), .A2(n_83), .B1(n_185), .B2(n_632), .Y(n_631) );
OAI22xp5_ASAP7_75t_L g529 ( .A1(n_31), .A2(n_530), .B1(n_532), .B2(n_533), .Y(n_529) );
INVx1_ASAP7_75t_L g533 ( .A(n_31), .Y(n_533) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_32), .A2(n_36), .B1(n_185), .B2(n_588), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_34), .A2(n_48), .B1(n_562), .B2(n_564), .Y(n_563) );
CKINVDCx5p33_ASAP7_75t_R g243 ( .A(n_35), .Y(n_243) );
XNOR2x2_ASAP7_75t_L g530 ( .A(n_38), .B(n_531), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g275 ( .A(n_39), .B(n_170), .Y(n_275) );
INVx2_ASAP7_75t_L g108 ( .A(n_40), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_41), .B(n_141), .Y(n_163) );
INVx1_ASAP7_75t_L g113 ( .A(n_42), .Y(n_113) );
BUFx3_ASAP7_75t_L g542 ( .A(n_42), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_44), .B(n_175), .Y(n_174) );
AND2x2_ASAP7_75t_L g245 ( .A(n_46), .B(n_175), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_47), .B(n_221), .Y(n_220) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_49), .B(n_138), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_50), .B(n_261), .Y(n_260) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_51), .A2(n_71), .B1(n_261), .B2(n_564), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_52), .A2(n_74), .B1(n_185), .B2(n_588), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_53), .B(n_208), .Y(n_207) );
A2O1A1Ixp33_ASAP7_75t_L g237 ( .A1(n_54), .A2(n_188), .B(n_195), .C(n_238), .Y(n_237) );
OAI22xp5_ASAP7_75t_L g118 ( .A1(n_55), .A2(n_60), .B1(n_119), .B2(n_120), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_55), .Y(n_119) );
AOI22xp5_ASAP7_75t_L g610 ( .A1(n_56), .A2(n_97), .B1(n_562), .B2(n_586), .Y(n_610) );
INVx1_ASAP7_75t_L g151 ( .A(n_57), .Y(n_151) );
AND2x4_ASAP7_75t_L g153 ( .A(n_58), .B(n_154), .Y(n_153) );
AOI22xp33_ASAP7_75t_L g143 ( .A1(n_59), .A2(n_62), .B1(n_136), .B2(n_144), .Y(n_143) );
INVx1_ASAP7_75t_L g120 ( .A(n_60), .Y(n_120) );
OAI22x1_ASAP7_75t_L g122 ( .A1(n_61), .A2(n_92), .B1(n_123), .B2(n_124), .Y(n_122) );
INVx1_ASAP7_75t_L g124 ( .A(n_61), .Y(n_124) );
XOR2xp5_ASAP7_75t_SL g534 ( .A(n_61), .B(n_125), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_63), .B(n_181), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_64), .B(n_175), .Y(n_223) );
CKINVDCx5p33_ASAP7_75t_R g244 ( .A(n_65), .Y(n_244) );
NAND2xp5_ASAP7_75t_SL g278 ( .A(n_66), .B(n_136), .Y(n_278) );
INVx1_ASAP7_75t_L g154 ( .A(n_67), .Y(n_154) );
CKINVDCx5p33_ASAP7_75t_R g156 ( .A(n_68), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_69), .B(n_181), .Y(n_279) );
XNOR2xp5_ASAP7_75t_L g528 ( .A(n_70), .B(n_529), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_72), .B(n_185), .Y(n_203) );
NAND3xp33_ASAP7_75t_L g164 ( .A(n_73), .B(n_141), .C(n_165), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_75), .B(n_185), .Y(n_184) );
INVx2_ASAP7_75t_L g142 ( .A(n_76), .Y(n_142) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_77), .B(n_172), .Y(n_217) );
NAND2xp5_ASAP7_75t_SL g259 ( .A(n_78), .B(n_170), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_79), .B(n_192), .Y(n_191) );
AOI22xp33_ASAP7_75t_L g633 ( .A1(n_80), .A2(n_98), .B1(n_136), .B2(n_195), .Y(n_633) );
CKINVDCx5p33_ASAP7_75t_R g576 ( .A(n_81), .Y(n_576) );
CKINVDCx5p33_ASAP7_75t_R g605 ( .A(n_82), .Y(n_605) );
AOI22xp33_ASAP7_75t_L g134 ( .A1(n_84), .A2(n_91), .B1(n_135), .B2(n_138), .Y(n_134) );
CKINVDCx20_ASAP7_75t_R g519 ( .A(n_85), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_86), .B(n_170), .Y(n_257) );
NAND2xp33_ASAP7_75t_SL g222 ( .A(n_87), .B(n_187), .Y(n_222) );
INVx1_ASAP7_75t_L g531 ( .A(n_88), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_89), .B(n_256), .Y(n_274) );
NAND2xp5_ASAP7_75t_SL g626 ( .A(n_90), .B(n_181), .Y(n_626) );
INVx1_ASAP7_75t_L g123 ( .A(n_92), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g592 ( .A(n_93), .Y(n_592) );
NOR2xp33_ASAP7_75t_L g111 ( .A(n_94), .B(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g539 ( .A(n_94), .Y(n_539) );
NAND2xp33_ASAP7_75t_L g624 ( .A(n_95), .B(n_170), .Y(n_624) );
NAND2xp33_ASAP7_75t_L g186 ( .A(n_96), .B(n_187), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_99), .B(n_175), .Y(n_210) );
NAND3xp33_ASAP7_75t_L g218 ( .A(n_100), .B(n_172), .C(n_187), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_102), .B(n_185), .Y(n_277) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_103), .B(n_138), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_523), .B(n_525), .Y(n_104) );
OAI21x1_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_116), .B(n_514), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
AND2x2_ASAP7_75t_L g107 ( .A(n_108), .B(n_109), .Y(n_107) );
INVx3_ASAP7_75t_L g517 ( .A(n_108), .Y(n_517) );
NOR2xp33_ASAP7_75t_L g889 ( .A(n_108), .B(n_890), .Y(n_889) );
INVx5_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
CKINVDCx8_ASAP7_75t_R g522 ( .A(n_110), .Y(n_522) );
INVx3_ASAP7_75t_L g890 ( .A(n_110), .Y(n_890) );
AND2x6_ASAP7_75t_SL g110 ( .A(n_111), .B(n_114), .Y(n_110) );
INVx1_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
NOR2x1_ASAP7_75t_L g541 ( .A(n_115), .B(n_542), .Y(n_541) );
AOI22xp5_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_511), .B1(n_512), .B2(n_513), .Y(n_116) );
XOR2xp5_ASAP7_75t_L g117 ( .A(n_118), .B(n_121), .Y(n_117) );
XNOR2x1_ASAP7_75t_L g513 ( .A(n_118), .B(n_121), .Y(n_513) );
XNOR2x1_ASAP7_75t_L g121 ( .A(n_122), .B(n_125), .Y(n_121) );
OR2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_399), .Y(n_125) );
NAND4xp25_ASAP7_75t_L g126 ( .A(n_127), .B(n_306), .C(n_347), .D(n_379), .Y(n_126) );
NOR2xp33_ASAP7_75t_SL g127 ( .A(n_128), .B(n_285), .Y(n_127) );
NAND3xp33_ASAP7_75t_SL g128 ( .A(n_129), .B(n_246), .C(n_265), .Y(n_128) );
AOI22xp5_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_177), .B1(n_224), .B2(n_228), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_130), .B(n_292), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_130), .B(n_392), .Y(n_498) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
OR2x2_ASAP7_75t_L g248 ( .A(n_131), .B(n_249), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_132), .B(n_158), .Y(n_131) );
OR2x2_ASAP7_75t_L g227 ( .A(n_132), .B(n_158), .Y(n_227) );
INVx1_ASAP7_75t_L g295 ( .A(n_132), .Y(n_295) );
AND2x2_ASAP7_75t_L g298 ( .A(n_132), .B(n_269), .Y(n_298) );
AND2x2_ASAP7_75t_L g346 ( .A(n_132), .B(n_319), .Y(n_346) );
AND2x2_ASAP7_75t_L g354 ( .A(n_132), .B(n_328), .Y(n_354) );
OR2x2_ASAP7_75t_L g365 ( .A(n_132), .B(n_319), .Y(n_365) );
HB1xp67_ASAP7_75t_L g405 ( .A(n_132), .Y(n_405) );
AO31x2_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_148), .A3(n_152), .B(n_155), .Y(n_132) );
OAI22xp5_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_140), .B1(n_143), .B2(n_145), .Y(n_133) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
OAI21xp5_ASAP7_75t_L g162 ( .A1(n_136), .A2(n_163), .B(n_164), .Y(n_162) );
OAI22xp33_ASAP7_75t_L g242 ( .A1(n_136), .A2(n_185), .B1(n_243), .B2(n_244), .Y(n_242) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx1_ASAP7_75t_L g139 ( .A(n_137), .Y(n_139) );
INVx1_ASAP7_75t_L g144 ( .A(n_137), .Y(n_144) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_137), .Y(n_165) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_137), .Y(n_170) );
INVx3_ASAP7_75t_L g185 ( .A(n_137), .Y(n_185) );
BUFx6f_ASAP7_75t_L g187 ( .A(n_137), .Y(n_187) );
INVx1_ASAP7_75t_L g195 ( .A(n_137), .Y(n_195) );
INVx1_ASAP7_75t_L g221 ( .A(n_137), .Y(n_221) );
INVx2_ASAP7_75t_L g240 ( .A(n_137), .Y(n_240) );
INVx1_ASAP7_75t_L g256 ( .A(n_137), .Y(n_256) );
INVx1_ASAP7_75t_L g585 ( .A(n_138), .Y(n_585) );
INVx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
OAI22xp5_ASAP7_75t_L g560 ( .A1(n_140), .A2(n_145), .B1(n_561), .B2(n_563), .Y(n_560) );
OAI22xp5_ASAP7_75t_L g570 ( .A1(n_140), .A2(n_145), .B1(n_571), .B2(n_572), .Y(n_570) );
OAI22xp5_ASAP7_75t_L g583 ( .A1(n_140), .A2(n_584), .B1(n_587), .B2(n_589), .Y(n_583) );
OAI22xp5_ASAP7_75t_L g600 ( .A1(n_140), .A2(n_145), .B1(n_601), .B2(n_602), .Y(n_600) );
OAI22xp5_ASAP7_75t_L g609 ( .A1(n_140), .A2(n_589), .B1(n_610), .B2(n_611), .Y(n_609) );
AOI21xp5_ASAP7_75t_L g621 ( .A1(n_140), .A2(n_622), .B(n_624), .Y(n_621) );
OAI22xp5_ASAP7_75t_L g630 ( .A1(n_140), .A2(n_631), .B1(n_633), .B2(n_634), .Y(n_630) );
OAI22xp5_ASAP7_75t_L g647 ( .A1(n_140), .A2(n_145), .B1(n_648), .B2(n_650), .Y(n_647) );
INVx6_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
O2A1O1Ixp5_ASAP7_75t_L g253 ( .A1(n_141), .A2(n_254), .B(n_255), .C(n_257), .Y(n_253) );
AOI21xp5_ASAP7_75t_L g276 ( .A1(n_141), .A2(n_277), .B(n_278), .Y(n_276) );
O2A1O1Ixp5_ASAP7_75t_L g618 ( .A1(n_141), .A2(n_588), .B(n_619), .C(n_620), .Y(n_618) );
BUFx8_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx2_ASAP7_75t_L g147 ( .A(n_142), .Y(n_147) );
INVx1_ASAP7_75t_L g172 ( .A(n_142), .Y(n_172) );
INVx1_ASAP7_75t_L g189 ( .A(n_142), .Y(n_189) );
INVx1_ASAP7_75t_L g651 ( .A(n_144), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_145), .B(n_242), .Y(n_241) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g209 ( .A(n_146), .Y(n_209) );
BUFx3_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g193 ( .A(n_147), .Y(n_193) );
INVx2_ASAP7_75t_L g234 ( .A(n_148), .Y(n_234) );
NOR2xp33_ASAP7_75t_SL g591 ( .A(n_148), .B(n_592), .Y(n_591) );
NOR2xp33_ASAP7_75t_L g635 ( .A(n_148), .B(n_636), .Y(n_635) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx2_ASAP7_75t_L g157 ( .A(n_149), .Y(n_157) );
INVx2_ASAP7_75t_L g176 ( .A(n_149), .Y(n_176) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_150), .Y(n_160) );
INVx2_ASAP7_75t_L g235 ( .A(n_152), .Y(n_235) );
AO31x2_ASAP7_75t_L g582 ( .A1(n_152), .A2(n_583), .A3(n_590), .B(n_591), .Y(n_582) );
AO31x2_ASAP7_75t_L g599 ( .A1(n_152), .A2(n_600), .A3(n_603), .B(n_604), .Y(n_599) );
AO31x2_ASAP7_75t_L g646 ( .A1(n_152), .A2(n_629), .A3(n_647), .B(n_652), .Y(n_646) );
BUFx10_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
BUFx10_ASAP7_75t_L g173 ( .A(n_153), .Y(n_173) );
INVx1_ASAP7_75t_L g574 ( .A(n_153), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g155 ( .A(n_156), .B(n_157), .Y(n_155) );
BUFx2_ASAP7_75t_L g590 ( .A(n_157), .Y(n_590) );
AND2x2_ASAP7_75t_L g324 ( .A(n_158), .B(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g353 ( .A(n_158), .B(n_250), .Y(n_353) );
OA21x2_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_161), .B(n_174), .Y(n_158) );
OAI21x1_ASAP7_75t_L g269 ( .A1(n_159), .A2(n_161), .B(n_174), .Y(n_269) );
OAI21x1_ASAP7_75t_L g271 ( .A1(n_159), .A2(n_272), .B(n_279), .Y(n_271) );
OAI21x1_ASAP7_75t_L g319 ( .A1(n_159), .A2(n_272), .B(n_279), .Y(n_319) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx4_ASAP7_75t_L g181 ( .A(n_160), .Y(n_181) );
AND2x4_ASAP7_75t_SL g197 ( .A(n_160), .B(n_173), .Y(n_197) );
INVx1_ASAP7_75t_SL g214 ( .A(n_160), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g604 ( .A(n_160), .B(n_605), .Y(n_604) );
NOR2xp33_ASAP7_75t_L g612 ( .A(n_160), .B(n_512), .Y(n_612) );
INVx2_ASAP7_75t_SL g616 ( .A(n_160), .Y(n_616) );
BUFx3_ASAP7_75t_L g629 ( .A(n_160), .Y(n_629) );
NOR2xp33_ASAP7_75t_L g652 ( .A(n_160), .B(n_653), .Y(n_652) );
OAI21x1_ASAP7_75t_L g161 ( .A1(n_162), .A2(n_166), .B(n_173), .Y(n_161) );
INVx2_ASAP7_75t_L g208 ( .A(n_165), .Y(n_208) );
AOI21x1_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_168), .B(n_171), .Y(n_166) );
INVx1_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
OAI21xp5_ASAP7_75t_L g216 ( .A1(n_170), .A2(n_217), .B(n_218), .Y(n_216) );
INVx3_ASAP7_75t_L g562 ( .A(n_170), .Y(n_562) );
INVx1_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx1_ASAP7_75t_SL g589 ( .A(n_172), .Y(n_589) );
INVx1_ASAP7_75t_L g634 ( .A(n_172), .Y(n_634) );
OAI21x1_ASAP7_75t_L g201 ( .A1(n_173), .A2(n_202), .B(n_205), .Y(n_201) );
OAI21x1_ASAP7_75t_L g215 ( .A1(n_173), .A2(n_216), .B(n_219), .Y(n_215) );
OAI21x1_ASAP7_75t_L g252 ( .A1(n_173), .A2(n_253), .B(n_258), .Y(n_252) );
OAI21x1_ASAP7_75t_L g272 ( .A1(n_173), .A2(n_273), .B(n_276), .Y(n_272) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx2_ASAP7_75t_L g200 ( .A(n_176), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_176), .B(n_567), .Y(n_566) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_176), .B(n_576), .Y(n_575) );
OAI21xp5_ASAP7_75t_L g465 ( .A1(n_177), .A2(n_324), .B(n_460), .Y(n_465) );
AND2x2_ASAP7_75t_L g177 ( .A(n_178), .B(n_211), .Y(n_177) );
AND2x2_ASAP7_75t_L g228 ( .A(n_178), .B(n_229), .Y(n_228) );
AND2x2_ASAP7_75t_L g263 ( .A(n_178), .B(n_264), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_178), .B(n_361), .Y(n_360) );
NAND2xp33_ASAP7_75t_R g395 ( .A(n_178), .B(n_361), .Y(n_395) );
INVx1_ASAP7_75t_L g429 ( .A(n_178), .Y(n_429) );
HB1xp67_ASAP7_75t_L g479 ( .A(n_178), .Y(n_479) );
AND2x2_ASAP7_75t_L g178 ( .A(n_179), .B(n_198), .Y(n_178) );
INVx1_ASAP7_75t_L g282 ( .A(n_179), .Y(n_282) );
INVx4_ASAP7_75t_L g303 ( .A(n_179), .Y(n_303) );
OR2x2_ASAP7_75t_L g386 ( .A(n_179), .B(n_311), .Y(n_386) );
BUFx2_ASAP7_75t_L g455 ( .A(n_179), .Y(n_455) );
AND2x4_ASAP7_75t_L g179 ( .A(n_180), .B(n_182), .Y(n_179) );
INVx2_ASAP7_75t_L g603 ( .A(n_181), .Y(n_603) );
OAI21x1_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_190), .B(n_197), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_184), .A2(n_186), .B(n_188), .Y(n_183) );
INVx1_ASAP7_75t_L g564 ( .A(n_185), .Y(n_564) );
INVx1_ASAP7_75t_L g586 ( .A(n_185), .Y(n_586) );
INVx4_ASAP7_75t_L g588 ( .A(n_185), .Y(n_588) );
INVx2_ASAP7_75t_L g261 ( .A(n_187), .Y(n_261) );
INVx1_ASAP7_75t_L g623 ( .A(n_187), .Y(n_623) );
AOI21xp5_ASAP7_75t_L g202 ( .A1(n_188), .A2(n_203), .B(n_204), .Y(n_202) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_188), .A2(n_220), .B(n_222), .Y(n_219) );
AOI21xp5_ASAP7_75t_L g273 ( .A1(n_188), .A2(n_274), .B(n_275), .Y(n_273) );
BUFx4f_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
OAI22xp5_ASAP7_75t_L g190 ( .A1(n_191), .A2(n_193), .B1(n_194), .B2(n_196), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g258 ( .A1(n_192), .A2(n_259), .B(n_260), .Y(n_258) );
INVx2_ASAP7_75t_SL g192 ( .A(n_193), .Y(n_192) );
INVx1_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
AND2x2_ASAP7_75t_L g283 ( .A(n_198), .B(n_284), .Y(n_283) );
INVx2_ASAP7_75t_L g370 ( .A(n_198), .Y(n_370) );
AND2x2_ASAP7_75t_L g456 ( .A(n_198), .B(n_264), .Y(n_456) );
AND2x2_ASAP7_75t_L g478 ( .A(n_198), .B(n_303), .Y(n_478) );
INVx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx1_ASAP7_75t_L g333 ( .A(n_199), .Y(n_333) );
OAI21x1_ASAP7_75t_L g199 ( .A1(n_200), .A2(n_201), .B(n_210), .Y(n_199) );
OAI21x1_ASAP7_75t_L g251 ( .A1(n_200), .A2(n_252), .B(n_262), .Y(n_251) );
OAI21xp33_ASAP7_75t_SL g315 ( .A1(n_200), .A2(n_201), .B(n_210), .Y(n_315) );
OAI21xp5_ASAP7_75t_L g325 ( .A1(n_200), .A2(n_252), .B(n_262), .Y(n_325) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_206), .A2(n_207), .B(n_209), .Y(n_205) );
HB1xp67_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
AND2x2_ASAP7_75t_L g281 ( .A(n_212), .B(n_282), .Y(n_281) );
INVx2_ASAP7_75t_L g304 ( .A(n_212), .Y(n_304) );
INVx1_ASAP7_75t_L g341 ( .A(n_212), .Y(n_341) );
INVx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
INVx1_ASAP7_75t_L g311 ( .A(n_213), .Y(n_311) );
AND2x2_ASAP7_75t_L g368 ( .A(n_213), .B(n_232), .Y(n_368) );
OAI21x1_ASAP7_75t_L g213 ( .A1(n_214), .A2(n_215), .B(n_223), .Y(n_213) );
INVx1_ASAP7_75t_L g649 ( .A(n_221), .Y(n_649) );
NOR2xp33_ASAP7_75t_SL g363 ( .A(n_224), .B(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
AND2x4_ASAP7_75t_L g410 ( .A(n_226), .B(n_411), .Y(n_410) );
INVx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
OR2x2_ASAP7_75t_L g426 ( .A(n_227), .B(n_292), .Y(n_426) );
INVx1_ASAP7_75t_L g434 ( .A(n_227), .Y(n_434) );
OR2x2_ASAP7_75t_L g355 ( .A(n_229), .B(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
HB1xp67_ASAP7_75t_L g305 ( .A(n_230), .Y(n_305) );
INVx1_ASAP7_75t_L g463 ( .A(n_230), .Y(n_463) );
INVx1_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
INVx2_ASAP7_75t_L g264 ( .A(n_231), .Y(n_264) );
AND2x2_ASAP7_75t_L g361 ( .A(n_231), .B(n_304), .Y(n_361) );
INVx2_ASAP7_75t_L g420 ( .A(n_231), .Y(n_420) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx1_ASAP7_75t_L g284 ( .A(n_232), .Y(n_284) );
AOI21x1_ASAP7_75t_L g232 ( .A1(n_233), .A2(n_236), .B(n_245), .Y(n_232) );
NOR2xp67_ASAP7_75t_SL g233 ( .A(n_234), .B(n_235), .Y(n_233) );
INVx2_ASAP7_75t_L g565 ( .A(n_234), .Y(n_565) );
INVx1_ASAP7_75t_L g559 ( .A(n_235), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_237), .B(n_241), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_239), .B(n_240), .Y(n_238) );
INVx2_ASAP7_75t_SL g632 ( .A(n_240), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_247), .B(n_263), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
INVx2_ASAP7_75t_L g374 ( .A(n_249), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_249), .B(n_298), .Y(n_431) );
NAND2xp5_ASAP7_75t_SL g470 ( .A(n_249), .B(n_364), .Y(n_470) );
AND2x2_ASAP7_75t_L g496 ( .A(n_249), .B(n_354), .Y(n_496) );
BUFx3_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
INVxp67_ASAP7_75t_SL g267 ( .A(n_250), .Y(n_267) );
INVxp67_ASAP7_75t_SL g289 ( .A(n_250), .Y(n_289) );
AND2x2_ASAP7_75t_L g322 ( .A(n_250), .B(n_269), .Y(n_322) );
INVx1_ASAP7_75t_L g393 ( .A(n_250), .Y(n_393) );
INVx1_ASAP7_75t_L g408 ( .A(n_250), .Y(n_408) );
AND2x2_ASAP7_75t_L g460 ( .A(n_250), .B(n_413), .Y(n_460) );
INVx3_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
INVx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g331 ( .A(n_264), .B(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g338 ( .A(n_264), .B(n_339), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_264), .B(n_488), .Y(n_487) );
INVx2_ASAP7_75t_L g507 ( .A(n_264), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_266), .B(n_280), .Y(n_265) );
INVx1_ASAP7_75t_L g336 ( .A(n_266), .Y(n_336) );
AND2x4_ASAP7_75t_L g266 ( .A(n_267), .B(n_268), .Y(n_266) );
NAND2x1_ASAP7_75t_L g510 ( .A(n_267), .B(n_410), .Y(n_510) );
AND2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
INVx1_ASAP7_75t_L g294 ( .A(n_269), .Y(n_294) );
AND2x2_ASAP7_75t_L g359 ( .A(n_269), .B(n_325), .Y(n_359) );
INVx1_ASAP7_75t_L g373 ( .A(n_269), .Y(n_373) );
INVx3_ASAP7_75t_L g292 ( .A(n_270), .Y(n_292) );
BUFx3_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
INVx1_ASAP7_75t_L g328 ( .A(n_271), .Y(n_328) );
AND2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_283), .Y(n_280) );
INVx1_ASAP7_75t_L g356 ( .A(n_281), .Y(n_356) );
AND2x2_ASAP7_75t_L g383 ( .A(n_281), .B(n_314), .Y(n_383) );
AND2x2_ASAP7_75t_L g444 ( .A(n_281), .B(n_445), .Y(n_444) );
AND2x2_ASAP7_75t_L g506 ( .A(n_281), .B(n_507), .Y(n_506) );
INVx2_ASAP7_75t_L g387 ( .A(n_283), .Y(n_387) );
AND2x2_ASAP7_75t_L g415 ( .A(n_283), .B(n_304), .Y(n_415) );
AND2x2_ASAP7_75t_L g314 ( .A(n_284), .B(n_315), .Y(n_314) );
AOI21xp5_ASAP7_75t_L g285 ( .A1(n_286), .A2(n_296), .B(n_299), .Y(n_285) );
OAI22xp5_ASAP7_75t_SL g504 ( .A1(n_286), .A2(n_505), .B1(n_508), .B2(n_510), .Y(n_504) );
NAND2x1p5_ASAP7_75t_L g286 ( .A(n_287), .B(n_290), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
NAND2x1_ASAP7_75t_L g489 ( .A(n_288), .B(n_290), .Y(n_489) );
BUFx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AND2x4_ASAP7_75t_L g290 ( .A(n_291), .B(n_293), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_291), .B(n_353), .Y(n_398) );
INVx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g297 ( .A(n_292), .B(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_292), .B(n_373), .Y(n_372) );
AND2x4_ASAP7_75t_L g450 ( .A(n_293), .B(n_408), .Y(n_450) );
INVx1_ASAP7_75t_L g503 ( .A(n_293), .Y(n_503) );
AND2x4_ASAP7_75t_L g293 ( .A(n_294), .B(n_295), .Y(n_293) );
AND2x2_ASAP7_75t_L g318 ( .A(n_295), .B(n_319), .Y(n_318) );
INVx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_305), .Y(n_300) );
AND2x2_ASAP7_75t_L g301 ( .A(n_302), .B(n_304), .Y(n_301) );
INVx1_ASAP7_75t_L g313 ( .A(n_302), .Y(n_313) );
AND2x2_ASAP7_75t_L g377 ( .A(n_302), .B(n_378), .Y(n_377) );
AND3x2_ASAP7_75t_L g419 ( .A(n_302), .B(n_332), .C(n_420), .Y(n_419) );
NAND2xp5_ASAP7_75t_SL g476 ( .A(n_302), .B(n_420), .Y(n_476) );
INVx2_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
OR2x2_ASAP7_75t_L g340 ( .A(n_303), .B(n_341), .Y(n_340) );
NAND2x1_ASAP7_75t_L g369 ( .A(n_303), .B(n_370), .Y(n_369) );
BUFx2_ASAP7_75t_L g424 ( .A(n_303), .Y(n_424) );
AND2x2_ASAP7_75t_L g485 ( .A(n_303), .B(n_420), .Y(n_485) );
OR2x2_ASAP7_75t_L g464 ( .A(n_304), .B(n_333), .Y(n_464) );
INVx1_ASAP7_75t_L g425 ( .A(n_305), .Y(n_425) );
AOI321xp33_ASAP7_75t_L g306 ( .A1(n_307), .A2(n_316), .A3(n_320), .B1(n_323), .B2(n_329), .C(n_335), .Y(n_306) );
AOI211xp5_ASAP7_75t_SL g347 ( .A1(n_307), .A2(n_348), .B(n_350), .C(n_362), .Y(n_347) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
NAND2x1p5_ASAP7_75t_L g308 ( .A(n_309), .B(n_312), .Y(n_308) );
NOR3xp33_ASAP7_75t_L g473 ( .A(n_309), .B(n_412), .C(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g488 ( .A(n_309), .Y(n_488) );
BUFx2_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVxp67_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g332 ( .A(n_311), .B(n_333), .Y(n_332) );
OR2x2_ASAP7_75t_L g482 ( .A(n_311), .B(n_446), .Y(n_482) );
INVx1_ASAP7_75t_L g334 ( .A(n_312), .Y(n_334) );
AND2x2_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
BUFx2_ASAP7_75t_L g491 ( .A(n_313), .Y(n_491) );
INVx1_ASAP7_75t_L g344 ( .A(n_314), .Y(n_344) );
AND2x2_ASAP7_75t_L g471 ( .A(n_314), .B(n_455), .Y(n_471) );
BUFx2_ASAP7_75t_L g494 ( .A(n_315), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_316), .B(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g413 ( .A(n_319), .Y(n_413) );
OAI321xp33_ASAP7_75t_L g457 ( .A1(n_320), .A2(n_411), .A3(n_458), .B1(n_459), .B2(n_462), .C(n_465), .Y(n_457) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx2_ASAP7_75t_SL g321 ( .A(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g382 ( .A(n_322), .B(n_326), .Y(n_382) );
AND2x2_ASAP7_75t_L g323 ( .A(n_324), .B(n_326), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_324), .B(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g446 ( .A(n_325), .Y(n_446) );
INVx2_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
BUFx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_330), .B(n_334), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g484 ( .A(n_332), .B(n_485), .Y(n_484) );
INVx2_ASAP7_75t_L g378 ( .A(n_333), .Y(n_378) );
OAI22xp5_ASAP7_75t_L g335 ( .A1(n_336), .A2(n_337), .B1(n_342), .B2(n_345), .Y(n_335) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
AOI31xp33_ASAP7_75t_L g422 ( .A1(n_338), .A2(n_374), .A3(n_423), .B(n_425), .Y(n_422) );
INVx1_ASAP7_75t_SL g339 ( .A(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g437 ( .A(n_340), .Y(n_437) );
OR2x2_ASAP7_75t_L g458 ( .A(n_340), .B(n_344), .Y(n_458) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
BUFx2_ASAP7_75t_L g390 ( .A(n_346), .Y(n_390) );
INVx1_ASAP7_75t_L g448 ( .A(n_346), .Y(n_448) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
OAI22xp33_ASAP7_75t_L g350 ( .A1(n_351), .A2(n_355), .B1(n_357), .B2(n_360), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_353), .B(n_354), .Y(n_352) );
INVx2_ASAP7_75t_L g442 ( .A(n_354), .Y(n_442) );
INVx2_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
OAI21xp5_ASAP7_75t_L g388 ( .A1(n_358), .A2(n_389), .B(n_391), .Y(n_388) );
BUFx2_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
NAND2x1_ASAP7_75t_L g447 ( .A(n_359), .B(n_448), .Y(n_447) );
AND2x4_ASAP7_75t_L g376 ( .A(n_361), .B(n_377), .Y(n_376) );
OAI22xp33_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_366), .B1(n_371), .B2(n_375), .Y(n_362) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
OR2x2_ASAP7_75t_L g391 ( .A(n_365), .B(n_392), .Y(n_391) );
OR2x6_ASAP7_75t_L g366 ( .A(n_367), .B(n_369), .Y(n_366) );
NOR2x1_ASAP7_75t_SL g428 ( .A(n_367), .B(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g492 ( .A(n_367), .Y(n_492) );
INVx2_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g397 ( .A(n_368), .B(n_378), .Y(n_397) );
OR2x2_ASAP7_75t_L g371 ( .A(n_372), .B(n_374), .Y(n_371) );
INVx2_ASAP7_75t_L g418 ( .A(n_373), .Y(n_418) );
AOI22xp33_ASAP7_75t_L g475 ( .A1(n_373), .A2(n_418), .B1(n_476), .B2(n_477), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_374), .B(n_434), .Y(n_433) );
INVx3_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
AND2x2_ASAP7_75t_L g436 ( .A(n_378), .B(n_420), .Y(n_436) );
AOI221xp5_ASAP7_75t_L g379 ( .A1(n_380), .A2(n_383), .B1(n_384), .B2(n_388), .C(n_394), .Y(n_379) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_382), .B(n_484), .Y(n_483) );
INVx2_ASAP7_75t_L g502 ( .A(n_383), .Y(n_502) );
INVx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
OR2x2_ASAP7_75t_L g385 ( .A(n_386), .B(n_387), .Y(n_385) );
INVx1_ASAP7_75t_L g440 ( .A(n_387), .Y(n_440) );
INVxp67_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
AOI21xp33_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_396), .B(n_398), .Y(n_394) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_397), .B(n_407), .Y(n_406) );
AND2x4_ASAP7_75t_L g501 ( .A(n_397), .B(n_455), .Y(n_501) );
NAND2xp5_ASAP7_75t_SL g399 ( .A(n_400), .B(n_466), .Y(n_399) );
NOR4xp25_ASAP7_75t_L g400 ( .A(n_401), .B(n_421), .C(n_438), .D(n_457), .Y(n_400) );
OAI221xp5_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_406), .B1(n_409), .B2(n_414), .C(n_416), .Y(n_401) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
AOI22xp33_ASAP7_75t_L g439 ( .A1(n_403), .A2(n_425), .B1(n_440), .B2(n_441), .Y(n_439) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
NAND2xp5_ASAP7_75t_SL g474 ( .A(n_405), .B(n_408), .Y(n_474) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx2_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
OAI221xp5_ASAP7_75t_L g438 ( .A1(n_414), .A2(n_439), .B1(n_443), .B2(n_447), .C(n_449), .Y(n_438) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_417), .B(n_419), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
OAI21xp5_ASAP7_75t_SL g421 ( .A1(n_422), .A2(n_426), .B(n_427), .Y(n_421) );
INVxp67_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
AND2x2_ASAP7_75t_L g509 ( .A(n_424), .B(n_436), .Y(n_509) );
INVx2_ASAP7_75t_L g451 ( .A(n_426), .Y(n_451) );
AOI22xp5_ASAP7_75t_L g427 ( .A1(n_428), .A2(n_430), .B1(n_432), .B2(n_435), .Y(n_427) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g461 ( .A(n_434), .Y(n_461) );
INVx1_ASAP7_75t_L g481 ( .A(n_434), .Y(n_481) );
AND2x2_ASAP7_75t_L g435 ( .A(n_436), .B(n_437), .Y(n_435) );
INVxp67_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
OAI21xp5_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_451), .B(n_452), .Y(n_449) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_454), .B(n_456), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
OR3x2_ASAP7_75t_L g462 ( .A(n_455), .B(n_463), .C(n_464), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_460), .B(n_461), .Y(n_459) );
NOR4xp75_ASAP7_75t_SL g466 ( .A(n_467), .B(n_486), .C(n_499), .D(n_504), .Y(n_466) );
NAND3x1_ASAP7_75t_L g467 ( .A(n_468), .B(n_472), .C(n_483), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_469), .B(n_471), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
AOI22xp5_ASAP7_75t_L g472 ( .A1(n_473), .A2(n_475), .B1(n_479), .B2(n_480), .Y(n_472) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
NOR2x1_ASAP7_75t_SL g480 ( .A(n_481), .B(n_482), .Y(n_480) );
OAI22xp5_ASAP7_75t_L g486 ( .A1(n_487), .A2(n_489), .B1(n_490), .B2(n_495), .Y(n_486) );
NAND3x2_ASAP7_75t_L g490 ( .A(n_491), .B(n_492), .C(n_493), .Y(n_490) );
INVx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g495 ( .A(n_496), .B(n_497), .Y(n_495) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_500), .A2(n_502), .B(n_503), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
CKINVDCx5p33_ASAP7_75t_R g883 ( .A(n_511), .Y(n_883) );
CKINVDCx5p33_ASAP7_75t_R g511 ( .A(n_512), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_515), .B(n_518), .Y(n_514) );
INVxp67_ASAP7_75t_SL g515 ( .A(n_516), .Y(n_515) );
BUFx8_ASAP7_75t_SL g516 ( .A(n_517), .Y(n_516) );
BUFx2_ASAP7_75t_L g882 ( .A(n_517), .Y(n_882) );
NOR2xp33_ASAP7_75t_L g518 ( .A(n_519), .B(n_520), .Y(n_518) );
INVx3_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g880 ( .A(n_521), .B(n_881), .Y(n_880) );
INVx3_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
NAND2xp5_ASAP7_75t_SL g881 ( .A(n_523), .B(n_882), .Y(n_881) );
INVx2_ASAP7_75t_SL g888 ( .A(n_523), .Y(n_888) );
OAI22xp33_ASAP7_75t_L g525 ( .A1(n_526), .A2(n_879), .B1(n_883), .B2(n_884), .Y(n_525) );
AOI21x1_ASAP7_75t_L g526 ( .A1(n_527), .A2(n_535), .B(n_543), .Y(n_526) );
OR2x2_ASAP7_75t_L g527 ( .A(n_528), .B(n_534), .Y(n_527) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_528), .A2(n_534), .B(n_536), .Y(n_535) );
XOR2xp5_ASAP7_75t_L g547 ( .A(n_528), .B(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g532 ( .A(n_530), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_537), .B(n_540), .Y(n_536) );
NOR2x1_ASAP7_75t_R g545 ( .A(n_537), .B(n_546), .Y(n_545) );
CKINVDCx5p33_ASAP7_75t_R g537 ( .A(n_538), .Y(n_537) );
AND2x2_ASAP7_75t_L g878 ( .A(n_538), .B(n_541), .Y(n_878) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVxp67_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
BUFx2_ASAP7_75t_L g546 ( .A(n_541), .Y(n_546) );
OAI21x1_ASAP7_75t_L g543 ( .A1(n_544), .A2(n_547), .B(n_877), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
AND3x4_ASAP7_75t_L g550 ( .A(n_551), .B(n_739), .C(n_793), .Y(n_550) );
NOR2x1_ASAP7_75t_L g551 ( .A(n_552), .B(n_699), .Y(n_551) );
NAND3xp33_ASAP7_75t_L g552 ( .A(n_553), .B(n_637), .C(n_681), .Y(n_552) );
OAI21xp33_ASAP7_75t_L g553 ( .A1(n_554), .A2(n_577), .B(n_594), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
HB1xp67_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
OR2x2_ASAP7_75t_L g731 ( .A(n_556), .B(n_641), .Y(n_731) );
INVx2_ASAP7_75t_L g757 ( .A(n_556), .Y(n_757) );
OR2x2_ASAP7_75t_L g556 ( .A(n_557), .B(n_568), .Y(n_556) );
INVx1_ASAP7_75t_L g656 ( .A(n_557), .Y(n_656) );
INVx2_ASAP7_75t_L g771 ( .A(n_557), .Y(n_771) );
INVx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx2_ASAP7_75t_L g580 ( .A(n_558), .Y(n_580) );
AND2x4_ASAP7_75t_L g714 ( .A(n_558), .B(n_676), .Y(n_714) );
AO31x2_ASAP7_75t_L g558 ( .A1(n_559), .A2(n_560), .A3(n_565), .B(n_566), .Y(n_558) );
AO31x2_ASAP7_75t_L g608 ( .A1(n_559), .A2(n_590), .A3(n_609), .B(n_612), .Y(n_608) );
AO31x2_ASAP7_75t_L g569 ( .A1(n_565), .A2(n_570), .A3(n_573), .B(n_575), .Y(n_569) );
INVx1_ASAP7_75t_L g767 ( .A(n_568), .Y(n_767) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g593 ( .A(n_569), .Y(n_593) );
AND2x4_ASAP7_75t_L g644 ( .A(n_569), .B(n_645), .Y(n_644) );
HB1xp67_ASAP7_75t_L g673 ( .A(n_569), .Y(n_673) );
INVx2_ASAP7_75t_L g676 ( .A(n_569), .Y(n_676) );
OR2x2_ASAP7_75t_L g690 ( .A(n_569), .B(n_646), .Y(n_690) );
AND2x2_ASAP7_75t_L g792 ( .A(n_569), .B(n_582), .Y(n_792) );
AO31x2_ASAP7_75t_L g628 ( .A1(n_573), .A2(n_629), .A3(n_630), .B(n_635), .Y(n_628) );
INVx2_ASAP7_75t_SL g573 ( .A(n_574), .Y(n_573) );
INVx2_ASAP7_75t_SL g625 ( .A(n_574), .Y(n_625) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
NAND2xp5_ASAP7_75t_SL g847 ( .A(n_578), .B(n_848), .Y(n_847) );
OR2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_581), .Y(n_578) );
OR2x2_ASAP7_75t_L g674 ( .A(n_579), .B(n_675), .Y(n_674) );
NAND2xp5_ASAP7_75t_SL g738 ( .A(n_579), .B(n_693), .Y(n_738) );
AND2x2_ASAP7_75t_L g803 ( .A(n_579), .B(n_779), .Y(n_803) );
INVx4_ASAP7_75t_L g837 ( .A(n_579), .Y(n_837) );
INVx3_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g672 ( .A(n_580), .B(n_673), .Y(n_672) );
AND2x2_ASAP7_75t_L g710 ( .A(n_580), .B(n_643), .Y(n_710) );
AND2x2_ASAP7_75t_L g820 ( .A(n_580), .B(n_646), .Y(n_820) );
AND2x2_ASAP7_75t_L g854 ( .A(n_580), .B(n_676), .Y(n_854) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_582), .B(n_593), .Y(n_581) );
INVx4_ASAP7_75t_SL g643 ( .A(n_582), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_582), .B(n_670), .Y(n_669) );
AND2x2_ASAP7_75t_L g755 ( .A(n_582), .B(n_646), .Y(n_755) );
BUFx2_ASAP7_75t_L g773 ( .A(n_582), .Y(n_773) );
AOI222xp33_ASAP7_75t_L g681 ( .A1(n_593), .A2(n_682), .B1(n_687), .B2(n_688), .C1(n_691), .C2(n_695), .Y(n_681) );
INVx1_ASAP7_75t_L g812 ( .A(n_593), .Y(n_812) );
AND2x2_ASAP7_75t_L g594 ( .A(n_595), .B(n_606), .Y(n_594) );
AND2x2_ASAP7_75t_L g849 ( .A(n_595), .B(n_661), .Y(n_849) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_L g870 ( .A(n_596), .B(n_871), .Y(n_870) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
AND2x4_ASAP7_75t_L g679 ( .A(n_597), .B(n_680), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g818 ( .A(n_597), .B(n_662), .Y(n_818) );
INVx2_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_598), .B(n_666), .Y(n_708) );
AND2x2_ASAP7_75t_L g736 ( .A(n_598), .B(n_614), .Y(n_736) );
INVx2_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g665 ( .A(n_599), .B(n_666), .Y(n_665) );
OR2x2_ASAP7_75t_L g698 ( .A(n_599), .B(n_628), .Y(n_698) );
INVx1_ASAP7_75t_L g726 ( .A(n_599), .Y(n_726) );
HB1xp67_ASAP7_75t_L g832 ( .A(n_599), .Y(n_832) );
AOI222xp33_ASAP7_75t_L g781 ( .A1(n_606), .A2(n_724), .B1(n_782), .B2(n_783), .C1(n_785), .C2(n_787), .Y(n_781) );
AND2x4_ASAP7_75t_L g606 ( .A(n_607), .B(n_613), .Y(n_606) );
INVx1_ASAP7_75t_L g716 ( .A(n_607), .Y(n_716) );
BUFx2_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx3_ASAP7_75t_L g662 ( .A(n_608), .Y(n_662) );
AND2x2_ASAP7_75t_L g667 ( .A(n_608), .B(n_628), .Y(n_667) );
AND2x2_ASAP7_75t_L g727 ( .A(n_608), .B(n_627), .Y(n_727) );
AND2x2_ASAP7_75t_L g715 ( .A(n_613), .B(n_716), .Y(n_715) );
AND2x4_ASAP7_75t_L g810 ( .A(n_613), .B(n_726), .Y(n_810) );
NAND2xp5_ASAP7_75t_L g816 ( .A(n_613), .B(n_817), .Y(n_816) );
AND3x1_ASAP7_75t_L g875 ( .A(n_613), .B(n_644), .C(n_876), .Y(n_875) );
AND2x4_ASAP7_75t_L g613 ( .A(n_614), .B(n_627), .Y(n_613) );
AND2x2_ASAP7_75t_L g696 ( .A(n_614), .B(n_662), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g845 ( .A(n_614), .B(n_798), .Y(n_845) );
INVx2_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
BUFx2_ASAP7_75t_L g659 ( .A(n_615), .Y(n_659) );
OAI21x1_ASAP7_75t_L g615 ( .A1(n_616), .A2(n_617), .B(n_626), .Y(n_615) );
OAI21x1_ASAP7_75t_L g666 ( .A1(n_616), .A2(n_617), .B(n_626), .Y(n_666) );
OAI21x1_ASAP7_75t_L g617 ( .A1(n_618), .A2(n_621), .B(n_625), .Y(n_617) );
INVx2_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
AND2x4_ASAP7_75t_L g661 ( .A(n_628), .B(n_662), .Y(n_661) );
OR2x2_ASAP7_75t_L g694 ( .A(n_628), .B(n_680), .Y(n_694) );
INVx1_ASAP7_75t_L g704 ( .A(n_628), .Y(n_704) );
BUFx2_ASAP7_75t_L g798 ( .A(n_628), .Y(n_798) );
AOI21xp5_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_657), .B(n_663), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
NAND2x1_ASAP7_75t_L g639 ( .A(n_640), .B(n_654), .Y(n_639) );
AOI221xp5_ASAP7_75t_SL g721 ( .A1(n_640), .A2(n_722), .B1(n_728), .B2(n_732), .C(n_737), .Y(n_721) );
AND2x4_ASAP7_75t_L g640 ( .A(n_641), .B(n_644), .Y(n_640) );
INVx2_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g842 ( .A(n_642), .B(n_656), .Y(n_842) );
INVx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_643), .B(n_676), .Y(n_675) );
AND2x4_ASAP7_75t_L g684 ( .A(n_643), .B(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g720 ( .A(n_643), .Y(n_720) );
INVx1_ASAP7_75t_L g730 ( .A(n_643), .Y(n_730) );
AND2x2_ASAP7_75t_L g749 ( .A(n_643), .B(n_750), .Y(n_749) );
OR2x2_ASAP7_75t_L g761 ( .A(n_643), .B(n_762), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g874 ( .A(n_643), .B(n_767), .Y(n_874) );
INVx2_ASAP7_75t_L g709 ( .A(n_644), .Y(n_709) );
AND2x2_ASAP7_75t_L g719 ( .A(n_644), .B(n_720), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_644), .B(n_730), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g862 ( .A(n_644), .B(n_863), .Y(n_862) );
INVx2_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g670 ( .A(n_646), .Y(n_670) );
HB1xp67_ASAP7_75t_L g713 ( .A(n_646), .Y(n_713) );
INVx1_ASAP7_75t_L g750 ( .A(n_646), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_646), .B(n_767), .Y(n_766) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
OR2x2_ASAP7_75t_L g689 ( .A(n_655), .B(n_690), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g791 ( .A(n_655), .B(n_792), .Y(n_791) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
HB1xp67_ASAP7_75t_L g748 ( .A(n_656), .Y(n_748) );
NOR2xp33_ASAP7_75t_R g657 ( .A(n_658), .B(n_660), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
NOR3xp33_ASAP7_75t_L g737 ( .A(n_659), .B(n_729), .C(n_738), .Y(n_737) );
AND2x2_ASAP7_75t_L g760 ( .A(n_659), .B(n_667), .Y(n_760) );
AND2x2_ASAP7_75t_L g789 ( .A(n_659), .B(n_759), .Y(n_789) );
OR2x2_ASAP7_75t_L g856 ( .A(n_659), .B(n_857), .Y(n_856) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
AND2x4_ASAP7_75t_L g782 ( .A(n_661), .B(n_665), .Y(n_782) );
INVx2_ASAP7_75t_SL g866 ( .A(n_661), .Y(n_866) );
INVx2_ASAP7_75t_L g693 ( .A(n_662), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_662), .B(n_707), .Y(n_706) );
INVx3_ASAP7_75t_L g735 ( .A(n_662), .Y(n_735) );
HB1xp67_ASAP7_75t_L g808 ( .A(n_662), .Y(n_808) );
OAI32xp33_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_668), .A3(n_671), .B1(n_674), .B2(n_677), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_665), .B(n_667), .Y(n_664) );
AND2x2_ASAP7_75t_L g687 ( .A(n_665), .B(n_667), .Y(n_687) );
AND2x2_ASAP7_75t_L g745 ( .A(n_665), .B(n_727), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_665), .B(n_727), .Y(n_753) );
INVx1_ASAP7_75t_L g680 ( .A(n_666), .Y(n_680) );
AND2x4_ASAP7_75t_SL g678 ( .A(n_667), .B(n_679), .Y(n_678) );
INVx1_ASAP7_75t_SL g822 ( .A(n_667), .Y(n_822) );
INVx2_ASAP7_75t_L g857 ( .A(n_667), .Y(n_857) );
AND2x2_ASAP7_75t_L g869 ( .A(n_667), .B(n_736), .Y(n_869) );
NOR3xp33_ASAP7_75t_L g799 ( .A(n_668), .B(n_790), .C(n_800), .Y(n_799) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g685 ( .A(n_670), .Y(n_685) );
AOI321xp33_ASAP7_75t_L g868 ( .A1(n_671), .A2(n_730), .A3(n_869), .B1(n_870), .B2(n_872), .C(n_875), .Y(n_868) );
INVx2_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g686 ( .A(n_673), .Y(n_686) );
OAI22xp5_ASAP7_75t_L g872 ( .A1(n_675), .A2(n_694), .B1(n_873), .B2(n_874), .Y(n_872) );
INVx3_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
AND2x2_ASAP7_75t_L g775 ( .A(n_679), .B(n_734), .Y(n_775) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
NAND2xp5_ASAP7_75t_SL g683 ( .A(n_684), .B(n_686), .Y(n_683) );
INVx1_ASAP7_75t_L g809 ( .A(n_684), .Y(n_809) );
NAND2x1_ASAP7_75t_L g836 ( .A(n_684), .B(n_837), .Y(n_836) );
NAND2xp5_ASAP7_75t_L g853 ( .A(n_684), .B(n_854), .Y(n_853) );
AND2x2_ASAP7_75t_L g834 ( .A(n_686), .B(n_820), .Y(n_834) );
INVx2_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx2_ASAP7_75t_L g774 ( .A(n_690), .Y(n_774) );
OR2x2_ASAP7_75t_L g841 ( .A(n_690), .B(n_842), .Y(n_841) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
OR2x2_ASAP7_75t_L g692 ( .A(n_693), .B(n_694), .Y(n_692) );
NOR2xp33_ASAP7_75t_L g718 ( .A(n_693), .B(n_694), .Y(n_718) );
NOR2x1p5_ASAP7_75t_L g759 ( .A(n_693), .B(n_698), .Y(n_759) );
INVx1_ASAP7_75t_L g829 ( .A(n_693), .Y(n_829) );
NOR2x1_ASAP7_75t_L g830 ( .A(n_694), .B(n_831), .Y(n_830) );
AND2x2_ASAP7_75t_L g695 ( .A(n_696), .B(n_697), .Y(n_695) );
INVxp67_ASAP7_75t_SL g873 ( .A(n_696), .Y(n_873) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
NAND3xp33_ASAP7_75t_L g699 ( .A(n_700), .B(n_711), .C(n_721), .Y(n_699) );
NAND3xp33_ASAP7_75t_L g700 ( .A(n_701), .B(n_709), .C(n_710), .Y(n_700) );
AND2x4_ASAP7_75t_L g701 ( .A(n_702), .B(n_705), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
BUFx2_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g851 ( .A(n_705), .Y(n_851) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVxp67_ASAP7_75t_SL g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g743 ( .A(n_708), .Y(n_743) );
INVx1_ASAP7_75t_L g779 ( .A(n_708), .Y(n_779) );
NAND2xp33_ASAP7_75t_L g783 ( .A(n_709), .B(n_784), .Y(n_783) );
INVx1_ASAP7_75t_L g787 ( .A(n_709), .Y(n_787) );
INVx1_ASAP7_75t_L g813 ( .A(n_710), .Y(n_813) );
AOI21xp5_ASAP7_75t_L g711 ( .A1(n_712), .A2(n_715), .B(n_717), .Y(n_711) );
AND2x4_ASAP7_75t_L g712 ( .A(n_713), .B(n_714), .Y(n_712) );
INVx3_ASAP7_75t_L g762 ( .A(n_714), .Y(n_762) );
AND2x2_ASAP7_75t_L g717 ( .A(n_718), .B(n_719), .Y(n_717) );
INVxp67_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
AND2x2_ASAP7_75t_L g724 ( .A(n_725), .B(n_727), .Y(n_724) );
INVx2_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
AND2x2_ASAP7_75t_L g839 ( .A(n_726), .B(n_829), .Y(n_839) );
AND2x2_ASAP7_75t_L g742 ( .A(n_727), .B(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g807 ( .A(n_727), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_729), .B(n_731), .Y(n_728) );
OR2x2_ASAP7_75t_L g765 ( .A(n_730), .B(n_766), .Y(n_765) );
INVx2_ASAP7_75t_L g744 ( .A(n_731), .Y(n_744) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_734), .B(n_736), .Y(n_733) );
INVx2_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
AND2x4_ASAP7_75t_L g778 ( .A(n_735), .B(n_779), .Y(n_778) );
INVx1_ASAP7_75t_L g867 ( .A(n_736), .Y(n_867) );
NOR2xp67_ASAP7_75t_L g739 ( .A(n_740), .B(n_776), .Y(n_739) );
NAND3xp33_ASAP7_75t_SL g740 ( .A(n_741), .B(n_751), .C(n_763), .Y(n_740) );
AOI22xp33_ASAP7_75t_L g741 ( .A1(n_742), .A2(n_744), .B1(n_745), .B2(n_746), .Y(n_741) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_748), .B(n_749), .Y(n_747) );
INVx1_ASAP7_75t_L g784 ( .A(n_749), .Y(n_784) );
AND2x2_ASAP7_75t_L g859 ( .A(n_749), .B(n_770), .Y(n_859) );
INVx1_ASAP7_75t_L g806 ( .A(n_750), .Y(n_806) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
OAI32xp33_ASAP7_75t_L g752 ( .A1(n_753), .A2(n_754), .A3(n_756), .B1(n_758), .B2(n_761), .Y(n_752) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx2_ASAP7_75t_L g786 ( .A(n_755), .Y(n_786) );
NAND2x1_ASAP7_75t_L g824 ( .A(n_755), .B(n_825), .Y(n_824) );
HB1xp67_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
AND2x2_ASAP7_75t_L g785 ( .A(n_757), .B(n_786), .Y(n_785) );
NOR2x1_ASAP7_75t_L g758 ( .A(n_759), .B(n_760), .Y(n_758) );
OAI211xp5_ASAP7_75t_SL g811 ( .A1(n_762), .A2(n_805), .B(n_812), .C(n_813), .Y(n_811) );
INVx2_ASAP7_75t_L g825 ( .A(n_762), .Y(n_825) );
OAI21xp5_ASAP7_75t_L g763 ( .A1(n_764), .A2(n_768), .B(n_775), .Y(n_763) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
INVx1_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
HB1xp67_ASAP7_75t_L g780 ( .A(n_769), .Y(n_780) );
NAND2x1_ASAP7_75t_L g769 ( .A(n_770), .B(n_772), .Y(n_769) );
INVx2_ASAP7_75t_L g863 ( .A(n_770), .Y(n_863) );
INVx3_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
AND2x2_ASAP7_75t_L g871 ( .A(n_771), .B(n_806), .Y(n_871) );
AND2x2_ASAP7_75t_L g876 ( .A(n_771), .B(n_832), .Y(n_876) );
AND2x4_ASAP7_75t_L g772 ( .A(n_773), .B(n_774), .Y(n_772) );
INVx1_ASAP7_75t_L g801 ( .A(n_774), .Y(n_801) );
OAI211xp5_ASAP7_75t_L g776 ( .A1(n_777), .A2(n_780), .B(n_781), .C(n_788), .Y(n_776) );
INVxp67_ASAP7_75t_SL g777 ( .A(n_778), .Y(n_777) );
NAND2x1p5_ASAP7_75t_L g795 ( .A(n_778), .B(n_796), .Y(n_795) );
NAND2xp5_ASAP7_75t_L g788 ( .A(n_789), .B(n_790), .Y(n_788) );
INVx2_ASAP7_75t_SL g790 ( .A(n_791), .Y(n_790) );
NOR3xp33_ASAP7_75t_L g793 ( .A(n_794), .B(n_826), .C(n_855), .Y(n_793) );
OAI211xp5_ASAP7_75t_L g794 ( .A1(n_795), .A2(n_799), .B(n_802), .C(n_814), .Y(n_794) );
INVx1_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
AOI22xp5_ASAP7_75t_L g838 ( .A1(n_800), .A2(n_839), .B1(n_840), .B2(n_843), .Y(n_838) );
INVx1_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
AOI22xp5_ASAP7_75t_L g802 ( .A1(n_803), .A2(n_804), .B1(n_810), .B2(n_811), .Y(n_802) );
OAI22xp33_ASAP7_75t_L g804 ( .A1(n_805), .A2(n_807), .B1(n_808), .B2(n_809), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g848 ( .A(n_805), .B(n_837), .Y(n_848) );
INVx1_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
AND2x2_ASAP7_75t_L g819 ( .A(n_812), .B(n_820), .Y(n_819) );
AOI22xp5_ASAP7_75t_L g814 ( .A1(n_815), .A2(n_819), .B1(n_821), .B2(n_823), .Y(n_814) );
INVx1_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
INVx1_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
OR2x2_ASAP7_75t_L g844 ( .A(n_818), .B(n_845), .Y(n_844) );
INVx2_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
INVx1_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
OAI211xp5_ASAP7_75t_SL g826 ( .A1(n_827), .A2(n_833), .B(n_838), .C(n_846), .Y(n_826) );
INVx2_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
AND2x2_ASAP7_75t_L g828 ( .A(n_829), .B(n_830), .Y(n_828) );
INVx1_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
NOR2xp33_ASAP7_75t_L g833 ( .A(n_834), .B(n_835), .Y(n_833) );
INVx2_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
INVx1_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
INVx2_ASAP7_75t_SL g843 ( .A(n_844), .Y(n_843) );
AOI22xp5_ASAP7_75t_L g846 ( .A1(n_847), .A2(n_849), .B1(n_850), .B2(n_852), .Y(n_846) );
INVx1_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
INVx1_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
OAI211xp5_ASAP7_75t_SL g855 ( .A1(n_856), .A2(n_858), .B(n_860), .C(n_868), .Y(n_855) );
INVxp67_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
NAND2xp5_ASAP7_75t_L g860 ( .A(n_861), .B(n_864), .Y(n_860) );
INVx1_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
INVx1_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
OR2x2_ASAP7_75t_L g865 ( .A(n_866), .B(n_867), .Y(n_865) );
INVx1_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
INVx6_ASAP7_75t_SL g884 ( .A(n_885), .Y(n_884) );
BUFx10_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
OR2x4_ASAP7_75t_L g886 ( .A(n_887), .B(n_889), .Y(n_886) );
BUFx2_ASAP7_75t_L g887 ( .A(n_888), .Y(n_887) );
endmodule