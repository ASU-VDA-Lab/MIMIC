module fake_aes_5004_n_558 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_558);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_558;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_540;
wire n_119;
wire n_141;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_554;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_428;
wire n_364;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
BUFx6f_ASAP7_75t_L g79 ( .A(n_42), .Y(n_79) );
CKINVDCx5p33_ASAP7_75t_R g80 ( .A(n_22), .Y(n_80) );
CKINVDCx14_ASAP7_75t_R g81 ( .A(n_15), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_17), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_48), .Y(n_83) );
BUFx3_ASAP7_75t_L g84 ( .A(n_76), .Y(n_84) );
CKINVDCx5p33_ASAP7_75t_R g85 ( .A(n_12), .Y(n_85) );
BUFx2_ASAP7_75t_L g86 ( .A(n_58), .Y(n_86) );
INVxp67_ASAP7_75t_SL g87 ( .A(n_59), .Y(n_87) );
INVx2_ASAP7_75t_L g88 ( .A(n_60), .Y(n_88) );
CKINVDCx20_ASAP7_75t_R g89 ( .A(n_27), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_64), .Y(n_90) );
CKINVDCx20_ASAP7_75t_R g91 ( .A(n_57), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_17), .Y(n_92) );
BUFx2_ASAP7_75t_SL g93 ( .A(n_65), .Y(n_93) );
BUFx3_ASAP7_75t_L g94 ( .A(n_73), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_66), .Y(n_95) );
CKINVDCx20_ASAP7_75t_R g96 ( .A(n_38), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_12), .Y(n_97) );
CKINVDCx16_ASAP7_75t_R g98 ( .A(n_11), .Y(n_98) );
BUFx6f_ASAP7_75t_L g99 ( .A(n_16), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_5), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_26), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_33), .Y(n_102) );
CKINVDCx20_ASAP7_75t_R g103 ( .A(n_39), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_35), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_29), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_37), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_7), .Y(n_107) );
HB1xp67_ASAP7_75t_L g108 ( .A(n_24), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_40), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_55), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_23), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_9), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_13), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_47), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_3), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_30), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_41), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_36), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_16), .Y(n_119) );
BUFx6f_ASAP7_75t_L g120 ( .A(n_79), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_90), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_90), .Y(n_122) );
NOR2xp33_ASAP7_75t_L g123 ( .A(n_86), .B(n_0), .Y(n_123) );
AND2x6_ASAP7_75t_L g124 ( .A(n_84), .B(n_43), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_88), .Y(n_125) );
AND2x2_ASAP7_75t_L g126 ( .A(n_86), .B(n_0), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_116), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_81), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_108), .B(n_1), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_89), .Y(n_130) );
OAI21x1_ASAP7_75t_L g131 ( .A1(n_88), .A2(n_44), .B(n_77), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_91), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g133 ( .A(n_98), .Y(n_133) );
INVx6_ASAP7_75t_L g134 ( .A(n_79), .Y(n_134) );
INVx3_ASAP7_75t_L g135 ( .A(n_99), .Y(n_135) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_79), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_96), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_116), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_85), .B(n_1), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_117), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_117), .Y(n_141) );
AND2x4_ASAP7_75t_L g142 ( .A(n_126), .B(n_119), .Y(n_142) );
NOR2xp33_ASAP7_75t_L g143 ( .A(n_121), .B(n_83), .Y(n_143) );
AND2x6_ASAP7_75t_L g144 ( .A(n_126), .B(n_118), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_130), .Y(n_145) );
INVx4_ASAP7_75t_L g146 ( .A(n_124), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_120), .Y(n_147) );
INVxp67_ASAP7_75t_L g148 ( .A(n_123), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_120), .Y(n_149) );
INVx3_ASAP7_75t_L g150 ( .A(n_125), .Y(n_150) );
BUFx10_ASAP7_75t_L g151 ( .A(n_124), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_135), .Y(n_152) );
AND2x2_ASAP7_75t_L g153 ( .A(n_141), .B(n_80), .Y(n_153) );
NAND2xp5_ASAP7_75t_SL g154 ( .A(n_121), .B(n_80), .Y(n_154) );
INVx5_ASAP7_75t_L g155 ( .A(n_124), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g156 ( .A(n_122), .B(n_95), .Y(n_156) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_120), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_122), .B(n_102), .Y(n_158) );
AND2x2_ASAP7_75t_L g159 ( .A(n_141), .B(n_101), .Y(n_159) );
CKINVDCx5p33_ASAP7_75t_R g160 ( .A(n_132), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_120), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_135), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_120), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_135), .Y(n_164) );
BUFx3_ASAP7_75t_L g165 ( .A(n_124), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_135), .Y(n_166) );
INVxp67_ASAP7_75t_L g167 ( .A(n_153), .Y(n_167) );
AND2x2_ASAP7_75t_L g168 ( .A(n_153), .B(n_129), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_153), .B(n_140), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_159), .B(n_127), .Y(n_170) );
CKINVDCx5p33_ASAP7_75t_R g171 ( .A(n_145), .Y(n_171) );
A2O1A1Ixp33_ASAP7_75t_SL g172 ( .A1(n_148), .A2(n_140), .B(n_138), .C(n_127), .Y(n_172) );
AOI22xp5_ASAP7_75t_L g173 ( .A1(n_144), .A2(n_138), .B1(n_139), .B2(n_124), .Y(n_173) );
NAND2x1p5_ASAP7_75t_L g174 ( .A(n_146), .B(n_131), .Y(n_174) );
NAND2xp33_ASAP7_75t_SL g175 ( .A(n_159), .B(n_103), .Y(n_175) );
CKINVDCx5p33_ASAP7_75t_R g176 ( .A(n_160), .Y(n_176) );
INVx2_ASAP7_75t_SL g177 ( .A(n_159), .Y(n_177) );
BUFx4f_ASAP7_75t_SL g178 ( .A(n_154), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_142), .B(n_101), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_150), .Y(n_180) );
AND2x2_ASAP7_75t_L g181 ( .A(n_142), .B(n_85), .Y(n_181) );
AND2x2_ASAP7_75t_SL g182 ( .A(n_146), .B(n_118), .Y(n_182) );
BUFx3_ASAP7_75t_L g183 ( .A(n_165), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_142), .B(n_106), .Y(n_184) );
BUFx3_ASAP7_75t_L g185 ( .A(n_165), .Y(n_185) );
NAND2x1p5_ASAP7_75t_L g186 ( .A(n_146), .B(n_131), .Y(n_186) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_146), .B(n_106), .Y(n_187) );
INVxp67_ASAP7_75t_SL g188 ( .A(n_165), .Y(n_188) );
AND2x6_ASAP7_75t_SL g189 ( .A(n_142), .B(n_133), .Y(n_189) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_155), .B(n_111), .Y(n_190) );
INVx3_ASAP7_75t_L g191 ( .A(n_150), .Y(n_191) );
INVx2_ASAP7_75t_SL g192 ( .A(n_155), .Y(n_192) );
AOI22xp33_ASAP7_75t_L g193 ( .A1(n_144), .A2(n_148), .B1(n_143), .B2(n_156), .Y(n_193) );
OAI22x1_ASAP7_75t_L g194 ( .A1(n_143), .A2(n_137), .B1(n_107), .B2(n_111), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_150), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_150), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_144), .B(n_158), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_158), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_144), .B(n_124), .Y(n_199) );
BUFx12f_ASAP7_75t_L g200 ( .A(n_189), .Y(n_200) );
A2O1A1Ixp33_ASAP7_75t_L g201 ( .A1(n_198), .A2(n_125), .B(n_112), .C(n_82), .Y(n_201) );
NOR2xp67_ASAP7_75t_SL g202 ( .A(n_183), .B(n_155), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_198), .Y(n_203) );
BUFx2_ASAP7_75t_L g204 ( .A(n_182), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_168), .B(n_144), .Y(n_205) );
BUFx6f_ASAP7_75t_L g206 ( .A(n_183), .Y(n_206) );
BUFx3_ASAP7_75t_L g207 ( .A(n_183), .Y(n_207) );
HB1xp67_ASAP7_75t_L g208 ( .A(n_167), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_180), .Y(n_209) );
BUFx6f_ASAP7_75t_L g210 ( .A(n_185), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_180), .Y(n_211) );
OR2x6_ASAP7_75t_L g212 ( .A(n_177), .B(n_93), .Y(n_212) );
AOI221xp5_ASAP7_75t_L g213 ( .A1(n_168), .A2(n_128), .B1(n_107), .B2(n_92), .C(n_113), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_182), .B(n_155), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_195), .Y(n_215) );
BUFx12f_ASAP7_75t_L g216 ( .A(n_189), .Y(n_216) );
INVx2_ASAP7_75t_SL g217 ( .A(n_185), .Y(n_217) );
AND2x4_ASAP7_75t_L g218 ( .A(n_177), .B(n_169), .Y(n_218) );
INVx2_ASAP7_75t_SL g219 ( .A(n_185), .Y(n_219) );
O2A1O1Ixp33_ASAP7_75t_L g220 ( .A1(n_169), .A2(n_100), .B(n_115), .C(n_97), .Y(n_220) );
BUFx12f_ASAP7_75t_L g221 ( .A(n_171), .Y(n_221) );
AOI22xp33_ASAP7_75t_SL g222 ( .A1(n_182), .A2(n_144), .B1(n_124), .B2(n_114), .Y(n_222) );
INVx4_ASAP7_75t_L g223 ( .A(n_191), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_195), .Y(n_224) );
INVx3_ASAP7_75t_L g225 ( .A(n_191), .Y(n_225) );
OAI22xp5_ASAP7_75t_L g226 ( .A1(n_197), .A2(n_144), .B1(n_155), .B2(n_114), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_196), .Y(n_227) );
AND2x4_ASAP7_75t_L g228 ( .A(n_170), .B(n_144), .Y(n_228) );
INVx4_ASAP7_75t_L g229 ( .A(n_191), .Y(n_229) );
BUFx6f_ASAP7_75t_L g230 ( .A(n_199), .Y(n_230) );
O2A1O1Ixp33_ASAP7_75t_L g231 ( .A1(n_172), .A2(n_110), .B(n_104), .C(n_105), .Y(n_231) );
BUFx6f_ASAP7_75t_L g232 ( .A(n_199), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_211), .Y(n_233) );
INVx3_ASAP7_75t_L g234 ( .A(n_206), .Y(n_234) );
AO32x2_ASAP7_75t_L g235 ( .A1(n_226), .A2(n_174), .A3(n_186), .B1(n_173), .B2(n_193), .Y(n_235) );
OR2x2_ASAP7_75t_L g236 ( .A(n_203), .B(n_181), .Y(n_236) );
INVx2_ASAP7_75t_SL g237 ( .A(n_203), .Y(n_237) );
AND2x4_ASAP7_75t_L g238 ( .A(n_218), .B(n_191), .Y(n_238) );
HB1xp67_ASAP7_75t_L g239 ( .A(n_208), .Y(n_239) );
OAI21x1_ASAP7_75t_L g240 ( .A1(n_231), .A2(n_186), .B(n_174), .Y(n_240) );
AOI22xp33_ASAP7_75t_L g241 ( .A1(n_204), .A2(n_175), .B1(n_181), .B2(n_194), .Y(n_241) );
AOI22xp5_ASAP7_75t_L g242 ( .A1(n_204), .A2(n_173), .B1(n_179), .B2(n_184), .Y(n_242) );
OAI21x1_ASAP7_75t_L g243 ( .A1(n_209), .A2(n_174), .B(n_186), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_205), .B(n_178), .Y(n_244) );
OR2x2_ASAP7_75t_L g245 ( .A(n_218), .B(n_176), .Y(n_245) );
OAI21x1_ASAP7_75t_SL g246 ( .A1(n_223), .A2(n_196), .B(n_109), .Y(n_246) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_209), .A2(n_155), .B(n_187), .Y(n_247) );
AOI22xp33_ASAP7_75t_L g248 ( .A1(n_228), .A2(n_194), .B1(n_155), .B2(n_188), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_218), .B(n_228), .Y(n_249) );
INVxp67_ASAP7_75t_SL g250 ( .A(n_206), .Y(n_250) );
AO21x2_ASAP7_75t_L g251 ( .A1(n_201), .A2(n_87), .B(n_190), .Y(n_251) );
OR2x6_ASAP7_75t_L g252 ( .A(n_212), .B(n_93), .Y(n_252) );
OAI21x1_ASAP7_75t_L g253 ( .A1(n_227), .A2(n_161), .B(n_149), .Y(n_253) );
AOI21xp33_ASAP7_75t_L g254 ( .A1(n_212), .A2(n_220), .B(n_222), .Y(n_254) );
OAI21x1_ASAP7_75t_L g255 ( .A1(n_227), .A2(n_161), .B(n_149), .Y(n_255) );
AO31x2_ASAP7_75t_L g256 ( .A1(n_211), .A2(n_149), .A3(n_163), .B(n_161), .Y(n_256) );
BUFx12f_ASAP7_75t_L g257 ( .A(n_221), .Y(n_257) );
AOI22xp33_ASAP7_75t_SL g258 ( .A1(n_200), .A2(n_84), .B1(n_94), .B2(n_99), .Y(n_258) );
OAI21x1_ASAP7_75t_L g259 ( .A1(n_215), .A2(n_147), .B(n_163), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_215), .Y(n_260) );
AOI22xp33_ASAP7_75t_L g261 ( .A1(n_254), .A2(n_216), .B1(n_200), .B2(n_218), .Y(n_261) );
BUFx6f_ASAP7_75t_L g262 ( .A(n_238), .Y(n_262) );
OAI21x1_ASAP7_75t_L g263 ( .A1(n_243), .A2(n_224), .B(n_225), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_236), .B(n_228), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_236), .B(n_228), .Y(n_265) );
AOI22xp33_ASAP7_75t_L g266 ( .A1(n_241), .A2(n_216), .B1(n_212), .B2(n_213), .Y(n_266) );
OAI221xp5_ASAP7_75t_L g267 ( .A1(n_245), .A2(n_212), .B1(n_214), .B2(n_225), .C(n_224), .Y(n_267) );
OAI22xp5_ASAP7_75t_L g268 ( .A1(n_237), .A2(n_212), .B1(n_207), .B2(n_217), .Y(n_268) );
OAI221xp5_ASAP7_75t_L g269 ( .A1(n_245), .A2(n_225), .B1(n_229), .B2(n_223), .C(n_219), .Y(n_269) );
OR2x2_ASAP7_75t_L g270 ( .A(n_239), .B(n_223), .Y(n_270) );
AOI221xp5_ASAP7_75t_L g271 ( .A1(n_244), .A2(n_99), .B1(n_229), .B2(n_230), .C(n_232), .Y(n_271) );
AOI221xp5_ASAP7_75t_L g272 ( .A1(n_242), .A2(n_99), .B1(n_229), .B2(n_230), .C(n_232), .Y(n_272) );
OAI22xp33_ASAP7_75t_L g273 ( .A1(n_252), .A2(n_221), .B1(n_219), .B2(n_217), .Y(n_273) );
OAI22xp5_ASAP7_75t_L g274 ( .A1(n_237), .A2(n_207), .B1(n_210), .B2(n_206), .Y(n_274) );
BUFx2_ASAP7_75t_L g275 ( .A(n_257), .Y(n_275) );
A2O1A1Ixp33_ASAP7_75t_L g276 ( .A1(n_260), .A2(n_94), .B(n_230), .C(n_232), .Y(n_276) );
A2O1A1Ixp33_ASAP7_75t_L g277 ( .A1(n_242), .A2(n_202), .B(n_230), .C(n_232), .Y(n_277) );
AND2x2_ASAP7_75t_L g278 ( .A(n_238), .B(n_2), .Y(n_278) );
AOI22xp33_ASAP7_75t_L g279 ( .A1(n_252), .A2(n_99), .B1(n_230), .B2(n_232), .Y(n_279) );
OAI22xp33_ASAP7_75t_L g280 ( .A1(n_252), .A2(n_210), .B1(n_206), .B2(n_79), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_260), .B(n_210), .Y(n_281) );
OAI22xp5_ASAP7_75t_L g282 ( .A1(n_252), .A2(n_233), .B1(n_249), .B2(n_238), .Y(n_282) );
OA21x2_ASAP7_75t_L g283 ( .A1(n_240), .A2(n_163), .B(n_147), .Y(n_283) );
AOI22xp33_ASAP7_75t_SL g284 ( .A1(n_257), .A2(n_210), .B1(n_206), .B2(n_79), .Y(n_284) );
INVxp67_ASAP7_75t_L g285 ( .A(n_270), .Y(n_285) );
BUFx6f_ASAP7_75t_L g286 ( .A(n_263), .Y(n_286) );
AND2x2_ASAP7_75t_L g287 ( .A(n_278), .B(n_233), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_281), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_283), .Y(n_289) );
HB1xp67_ASAP7_75t_L g290 ( .A(n_276), .Y(n_290) );
BUFx3_ASAP7_75t_L g291 ( .A(n_262), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_283), .Y(n_292) );
NOR2x1_ASAP7_75t_R g293 ( .A(n_275), .B(n_250), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_283), .Y(n_294) );
INVxp67_ASAP7_75t_SL g295 ( .A(n_282), .Y(n_295) );
BUFx3_ASAP7_75t_L g296 ( .A(n_262), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_262), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_262), .Y(n_298) );
AND2x4_ASAP7_75t_SL g299 ( .A(n_279), .B(n_234), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_264), .Y(n_300) );
BUFx6f_ASAP7_75t_L g301 ( .A(n_265), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_261), .B(n_234), .Y(n_302) );
OR2x2_ASAP7_75t_L g303 ( .A(n_261), .B(n_266), .Y(n_303) );
HB1xp67_ASAP7_75t_L g304 ( .A(n_276), .Y(n_304) );
AND2x2_ASAP7_75t_L g305 ( .A(n_266), .B(n_234), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_277), .B(n_243), .Y(n_306) );
INVx4_ASAP7_75t_R g307 ( .A(n_273), .Y(n_307) );
AOI22xp33_ASAP7_75t_L g308 ( .A1(n_303), .A2(n_267), .B1(n_258), .B2(n_271), .Y(n_308) );
AND2x2_ASAP7_75t_L g309 ( .A(n_289), .B(n_235), .Y(n_309) );
AND2x4_ASAP7_75t_L g310 ( .A(n_302), .B(n_240), .Y(n_310) );
BUFx3_ASAP7_75t_L g311 ( .A(n_291), .Y(n_311) );
OR2x2_ASAP7_75t_L g312 ( .A(n_303), .B(n_268), .Y(n_312) );
INVx1_ASAP7_75t_SL g313 ( .A(n_299), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_294), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_289), .B(n_235), .Y(n_315) );
AND2x2_ASAP7_75t_L g316 ( .A(n_292), .B(n_235), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_292), .Y(n_317) );
AOI33xp33_ASAP7_75t_L g318 ( .A1(n_302), .A2(n_248), .A3(n_279), .B1(n_284), .B2(n_166), .B3(n_164), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_294), .Y(n_319) );
OR2x2_ASAP7_75t_L g320 ( .A(n_285), .B(n_274), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_287), .B(n_235), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_294), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_300), .B(n_272), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_286), .Y(n_324) );
INVx3_ASAP7_75t_L g325 ( .A(n_286), .Y(n_325) );
OR2x2_ASAP7_75t_L g326 ( .A(n_285), .B(n_251), .Y(n_326) );
AOI221xp5_ASAP7_75t_L g327 ( .A1(n_295), .A2(n_246), .B1(n_269), .B2(n_280), .C(n_251), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_286), .Y(n_328) );
BUFx3_ASAP7_75t_L g329 ( .A(n_291), .Y(n_329) );
HB1xp67_ASAP7_75t_L g330 ( .A(n_306), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_288), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_288), .Y(n_332) );
AOI211xp5_ASAP7_75t_L g333 ( .A1(n_293), .A2(n_120), .B(n_136), .C(n_247), .Y(n_333) );
OR2x2_ASAP7_75t_L g334 ( .A(n_300), .B(n_251), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_305), .B(n_235), .Y(n_335) );
OAI321xp33_ASAP7_75t_L g336 ( .A1(n_305), .A2(n_136), .A3(n_3), .B1(n_4), .B2(n_5), .C(n_6), .Y(n_336) );
AND2x2_ASAP7_75t_L g337 ( .A(n_335), .B(n_295), .Y(n_337) );
AND2x2_ASAP7_75t_L g338 ( .A(n_335), .B(n_306), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_331), .B(n_300), .Y(n_339) );
OR2x2_ASAP7_75t_L g340 ( .A(n_312), .B(n_301), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_335), .B(n_290), .Y(n_341) );
HB1xp67_ASAP7_75t_L g342 ( .A(n_320), .Y(n_342) );
AND2x4_ASAP7_75t_L g343 ( .A(n_310), .B(n_286), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_321), .B(n_290), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_331), .B(n_304), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_317), .Y(n_346) );
NOR2xp33_ASAP7_75t_SL g347 ( .A(n_313), .B(n_293), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_321), .B(n_304), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_314), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_317), .Y(n_350) );
HB1xp67_ASAP7_75t_L g351 ( .A(n_320), .Y(n_351) );
OR2x2_ASAP7_75t_L g352 ( .A(n_312), .B(n_301), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_310), .B(n_297), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_310), .B(n_297), .Y(n_354) );
AOI31xp33_ASAP7_75t_SL g355 ( .A1(n_333), .A2(n_307), .A3(n_298), .B(n_297), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_314), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_314), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_310), .B(n_298), .Y(n_358) );
OR2x2_ASAP7_75t_L g359 ( .A(n_326), .B(n_301), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_309), .B(n_298), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_332), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_309), .B(n_301), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_319), .Y(n_363) );
OR2x2_ASAP7_75t_L g364 ( .A(n_326), .B(n_301), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_309), .B(n_301), .Y(n_365) );
INVx3_ASAP7_75t_L g366 ( .A(n_325), .Y(n_366) );
OR2x2_ASAP7_75t_L g367 ( .A(n_319), .B(n_287), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_315), .B(n_286), .Y(n_368) );
HB1xp67_ASAP7_75t_L g369 ( .A(n_322), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_315), .B(n_286), .Y(n_370) );
NAND4xp25_ASAP7_75t_L g371 ( .A(n_308), .B(n_296), .C(n_291), .D(n_307), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_332), .Y(n_372) );
OAI21xp5_ASAP7_75t_L g373 ( .A1(n_336), .A2(n_259), .B(n_255), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_322), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_315), .B(n_296), .Y(n_375) );
INVx1_ASAP7_75t_SL g376 ( .A(n_313), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_334), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_316), .B(n_296), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_316), .B(n_299), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_378), .B(n_311), .Y(n_380) );
OR2x2_ASAP7_75t_L g381 ( .A(n_342), .B(n_334), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_351), .B(n_316), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_346), .Y(n_383) );
AOI22xp33_ASAP7_75t_L g384 ( .A1(n_371), .A2(n_327), .B1(n_330), .B2(n_323), .Y(n_384) );
OR2x2_ASAP7_75t_L g385 ( .A(n_367), .B(n_330), .Y(n_385) );
INVx1_ASAP7_75t_SL g386 ( .A(n_367), .Y(n_386) );
OAI21xp5_ASAP7_75t_L g387 ( .A1(n_347), .A2(n_336), .B(n_333), .Y(n_387) );
INVx1_ASAP7_75t_SL g388 ( .A(n_376), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_337), .B(n_323), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_346), .Y(n_390) );
NAND2x1p5_ASAP7_75t_L g391 ( .A(n_376), .B(n_311), .Y(n_391) );
OR2x2_ASAP7_75t_L g392 ( .A(n_340), .B(n_311), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_337), .B(n_329), .Y(n_393) );
OR2x2_ASAP7_75t_L g394 ( .A(n_340), .B(n_329), .Y(n_394) );
INVx3_ASAP7_75t_L g395 ( .A(n_363), .Y(n_395) );
HB1xp67_ASAP7_75t_L g396 ( .A(n_369), .Y(n_396) );
INVxp67_ASAP7_75t_L g397 ( .A(n_369), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_349), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_378), .B(n_329), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_350), .Y(n_400) );
NOR2xp33_ASAP7_75t_L g401 ( .A(n_371), .B(n_2), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_379), .B(n_325), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_341), .B(n_318), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_379), .B(n_325), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_341), .B(n_327), .Y(n_405) );
NOR2xp33_ASAP7_75t_L g406 ( .A(n_361), .B(n_4), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_344), .B(n_325), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_344), .B(n_328), .Y(n_408) );
CKINVDCx16_ASAP7_75t_R g409 ( .A(n_347), .Y(n_409) );
CKINVDCx20_ASAP7_75t_R g410 ( .A(n_375), .Y(n_410) );
BUFx6f_ASAP7_75t_L g411 ( .A(n_343), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_348), .B(n_328), .Y(n_412) );
INVx3_ASAP7_75t_SL g413 ( .A(n_359), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_348), .B(n_328), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_349), .Y(n_415) );
AND2x4_ASAP7_75t_L g416 ( .A(n_343), .B(n_324), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_338), .B(n_324), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_338), .B(n_324), .Y(n_418) );
NAND2xp5_ASAP7_75t_SL g419 ( .A(n_363), .B(n_299), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_350), .Y(n_420) );
NAND2x1p5_ASAP7_75t_L g421 ( .A(n_374), .B(n_210), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_349), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_361), .B(n_6), .Y(n_423) );
OR2x2_ASAP7_75t_L g424 ( .A(n_352), .B(n_7), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_372), .Y(n_425) );
BUFx3_ASAP7_75t_L g426 ( .A(n_363), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_372), .Y(n_427) );
NAND4xp25_ASAP7_75t_L g428 ( .A(n_345), .B(n_8), .C(n_9), .D(n_10), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_374), .Y(n_429) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_345), .B(n_8), .Y(n_430) );
OR2x6_ASAP7_75t_L g431 ( .A(n_339), .B(n_246), .Y(n_431) );
AOI22xp5_ASAP7_75t_L g432 ( .A1(n_401), .A2(n_353), .B1(n_354), .B2(n_358), .Y(n_432) );
AOI22xp5_ASAP7_75t_L g433 ( .A1(n_401), .A2(n_353), .B1(n_354), .B2(n_358), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_385), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_383), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_426), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_426), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_386), .B(n_377), .Y(n_438) );
AOI21xp33_ASAP7_75t_SL g439 ( .A1(n_409), .A2(n_355), .B(n_339), .Y(n_439) );
OAI31xp33_ASAP7_75t_L g440 ( .A1(n_428), .A2(n_355), .A3(n_377), .B(n_343), .Y(n_440) );
AOI322xp5_ASAP7_75t_L g441 ( .A1(n_430), .A2(n_362), .A3(n_365), .B1(n_375), .B2(n_360), .C1(n_368), .C2(n_370), .Y(n_441) );
AOI322xp5_ASAP7_75t_L g442 ( .A1(n_430), .A2(n_362), .A3(n_365), .B1(n_360), .B2(n_370), .C1(n_368), .C2(n_343), .Y(n_442) );
NOR2xp33_ASAP7_75t_L g443 ( .A(n_410), .B(n_352), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_413), .B(n_364), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_389), .B(n_364), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_382), .B(n_357), .Y(n_446) );
OAI32xp33_ASAP7_75t_L g447 ( .A1(n_410), .A2(n_359), .A3(n_366), .B1(n_357), .B2(n_356), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_405), .B(n_357), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_390), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_400), .Y(n_450) );
OAI32xp33_ASAP7_75t_L g451 ( .A1(n_387), .A2(n_366), .A3(n_356), .B1(n_373), .B2(n_14), .Y(n_451) );
OR2x2_ASAP7_75t_L g452 ( .A(n_413), .B(n_356), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_397), .B(n_366), .Y(n_453) );
INVxp67_ASAP7_75t_SL g454 ( .A(n_396), .Y(n_454) );
NOR3xp33_ASAP7_75t_L g455 ( .A(n_406), .B(n_366), .C(n_373), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_420), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_425), .Y(n_457) );
AOI222xp33_ASAP7_75t_L g458 ( .A1(n_403), .A2(n_136), .B1(n_134), .B2(n_13), .C1(n_14), .C2(n_15), .Y(n_458) );
OAI21xp33_ASAP7_75t_L g459 ( .A1(n_384), .A2(n_136), .B(n_147), .Y(n_459) );
NAND2x1_ASAP7_75t_SL g460 ( .A(n_396), .B(n_10), .Y(n_460) );
NAND2x1_ASAP7_75t_L g461 ( .A(n_395), .B(n_134), .Y(n_461) );
OAI21xp33_ASAP7_75t_SL g462 ( .A1(n_384), .A2(n_259), .B(n_255), .Y(n_462) );
OAI32xp33_ASAP7_75t_L g463 ( .A1(n_388), .A2(n_11), .A3(n_134), .B1(n_136), .B2(n_20), .Y(n_463) );
OAI22xp5_ASAP7_75t_L g464 ( .A1(n_431), .A2(n_134), .B1(n_136), .B2(n_256), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_427), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_380), .B(n_18), .Y(n_466) );
NOR3xp33_ASAP7_75t_L g467 ( .A(n_406), .B(n_253), .C(n_166), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_429), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_397), .Y(n_469) );
INVx1_ASAP7_75t_SL g470 ( .A(n_391), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_381), .Y(n_471) );
OAI211xp5_ASAP7_75t_SL g472 ( .A1(n_424), .A2(n_164), .B(n_162), .C(n_152), .Y(n_472) );
NAND3xp33_ASAP7_75t_L g473 ( .A(n_423), .B(n_157), .C(n_162), .Y(n_473) );
AOI21xp5_ASAP7_75t_L g474 ( .A1(n_419), .A2(n_253), .B(n_256), .Y(n_474) );
INVx1_ASAP7_75t_SL g475 ( .A(n_391), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_395), .Y(n_476) );
AOI22xp5_ASAP7_75t_L g477 ( .A1(n_407), .A2(n_157), .B1(n_152), .B2(n_202), .Y(n_477) );
INVx2_ASAP7_75t_L g478 ( .A(n_398), .Y(n_478) );
INVxp67_ASAP7_75t_L g479 ( .A(n_469), .Y(n_479) );
NOR3x1_ASAP7_75t_L g480 ( .A(n_454), .B(n_393), .C(n_419), .Y(n_480) );
INVxp67_ASAP7_75t_L g481 ( .A(n_448), .Y(n_481) );
INVx1_ASAP7_75t_SL g482 ( .A(n_444), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_441), .B(n_418), .Y(n_483) );
INVxp33_ASAP7_75t_L g484 ( .A(n_460), .Y(n_484) );
OAI21xp5_ASAP7_75t_L g485 ( .A1(n_440), .A2(n_431), .B(n_421), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_471), .B(n_443), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_435), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_449), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_450), .Y(n_489) );
OAI322xp33_ASAP7_75t_L g490 ( .A1(n_432), .A2(n_417), .A3(n_394), .B1(n_392), .B2(n_412), .C1(n_408), .C2(n_414), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_442), .B(n_399), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_456), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_457), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_434), .B(n_436), .Y(n_494) );
OAI221xp5_ASAP7_75t_SL g495 ( .A1(n_433), .A2(n_402), .B1(n_404), .B2(n_431), .C(n_398), .Y(n_495) );
OAI221xp5_ASAP7_75t_L g496 ( .A1(n_455), .A2(n_411), .B1(n_422), .B2(n_415), .C(n_421), .Y(n_496) );
NAND2xp5_ASAP7_75t_SL g497 ( .A(n_439), .B(n_411), .Y(n_497) );
NAND4xp25_ASAP7_75t_SL g498 ( .A(n_458), .B(n_422), .C(n_415), .D(n_411), .Y(n_498) );
NAND3xp33_ASAP7_75t_L g499 ( .A(n_458), .B(n_411), .C(n_416), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_478), .Y(n_500) );
NOR3x1_ASAP7_75t_L g501 ( .A(n_452), .B(n_416), .C(n_21), .Y(n_501) );
OAI22xp33_ASAP7_75t_L g502 ( .A1(n_470), .A2(n_416), .B1(n_157), .B2(n_256), .Y(n_502) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_445), .B(n_19), .Y(n_503) );
INVx2_ASAP7_75t_SL g504 ( .A(n_437), .Y(n_504) );
NOR2xp67_ASAP7_75t_L g505 ( .A(n_462), .B(n_25), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_446), .B(n_256), .Y(n_506) );
INVx2_ASAP7_75t_L g507 ( .A(n_476), .Y(n_507) );
CKINVDCx14_ASAP7_75t_R g508 ( .A(n_466), .Y(n_508) );
AOI221xp5_ASAP7_75t_L g509 ( .A1(n_447), .A2(n_451), .B1(n_465), .B2(n_468), .C(n_453), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_472), .A2(n_157), .B1(n_31), .B2(n_32), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_487), .Y(n_511) );
NOR2x1_ASAP7_75t_L g512 ( .A(n_498), .B(n_473), .Y(n_512) );
NAND4xp75_ASAP7_75t_L g513 ( .A(n_480), .B(n_453), .C(n_438), .D(n_477), .Y(n_513) );
AOI32xp33_ASAP7_75t_L g514 ( .A1(n_484), .A2(n_475), .A3(n_470), .B1(n_467), .B2(n_464), .Y(n_514) );
OAI22xp5_ASAP7_75t_L g515 ( .A1(n_508), .A2(n_475), .B1(n_464), .B2(n_446), .Y(n_515) );
AO21x1_ASAP7_75t_L g516 ( .A1(n_497), .A2(n_461), .B(n_474), .Y(n_516) );
XOR2x2_ASAP7_75t_L g517 ( .A(n_491), .B(n_459), .Y(n_517) );
INVx2_ASAP7_75t_L g518 ( .A(n_500), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_488), .Y(n_519) );
NOR2x1_ASAP7_75t_L g520 ( .A(n_497), .B(n_463), .Y(n_520) );
AOI22xp5_ASAP7_75t_L g521 ( .A1(n_508), .A2(n_157), .B1(n_256), .B2(n_45), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_484), .A2(n_157), .B(n_34), .Y(n_522) );
AOI22xp5_ASAP7_75t_L g523 ( .A1(n_483), .A2(n_28), .B1(n_46), .B2(n_49), .Y(n_523) );
A2O1A1Ixp33_ASAP7_75t_SL g524 ( .A1(n_503), .A2(n_50), .B(n_51), .C(n_52), .Y(n_524) );
INVx2_ASAP7_75t_SL g525 ( .A(n_482), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_489), .Y(n_526) );
INVx1_ASAP7_75t_SL g527 ( .A(n_504), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_492), .Y(n_528) );
O2A1O1Ixp33_ASAP7_75t_SL g529 ( .A1(n_485), .A2(n_53), .B(n_54), .C(n_56), .Y(n_529) );
NAND4xp25_ASAP7_75t_L g530 ( .A(n_501), .B(n_61), .C(n_62), .D(n_63), .Y(n_530) );
AOI221xp5_ASAP7_75t_L g531 ( .A1(n_515), .A2(n_490), .B1(n_495), .B2(n_479), .C(n_481), .Y(n_531) );
OAI221xp5_ASAP7_75t_L g532 ( .A1(n_514), .A2(n_509), .B1(n_499), .B2(n_496), .C(n_505), .Y(n_532) );
BUFx2_ASAP7_75t_L g533 ( .A(n_525), .Y(n_533) );
NAND3xp33_ASAP7_75t_SL g534 ( .A(n_516), .B(n_510), .C(n_503), .Y(n_534) );
AOI221xp5_ASAP7_75t_SL g535 ( .A1(n_527), .A2(n_486), .B1(n_494), .B2(n_493), .C(n_502), .Y(n_535) );
OAI221xp5_ASAP7_75t_SL g536 ( .A1(n_521), .A2(n_510), .B1(n_506), .B2(n_507), .C(n_500), .Y(n_536) );
AOI21xp33_ASAP7_75t_SL g537 ( .A1(n_521), .A2(n_513), .B(n_517), .Y(n_537) );
NAND4xp25_ASAP7_75t_SL g538 ( .A(n_512), .B(n_507), .C(n_68), .D(n_69), .Y(n_538) );
AOI221xp5_ASAP7_75t_L g539 ( .A1(n_511), .A2(n_67), .B1(n_70), .B2(n_71), .C(n_72), .Y(n_539) );
O2A1O1Ixp33_ASAP7_75t_L g540 ( .A1(n_520), .A2(n_74), .B(n_75), .C(n_78), .Y(n_540) );
OAI211xp5_ASAP7_75t_SL g541 ( .A1(n_523), .A2(n_151), .B(n_192), .C(n_529), .Y(n_541) );
HB1xp67_ASAP7_75t_L g542 ( .A(n_533), .Y(n_542) );
NAND3xp33_ASAP7_75t_SL g543 ( .A(n_537), .B(n_522), .C(n_524), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_531), .B(n_519), .Y(n_544) );
OR3x2_ASAP7_75t_L g545 ( .A(n_534), .B(n_530), .C(n_526), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_532), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_536), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_547), .A2(n_538), .B1(n_541), .B2(n_528), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_542), .Y(n_549) );
NOR2xp33_ASAP7_75t_SL g550 ( .A(n_543), .B(n_540), .Y(n_550) );
INVx3_ASAP7_75t_L g551 ( .A(n_549), .Y(n_551) );
NAND3xp33_ASAP7_75t_SL g552 ( .A(n_550), .B(n_546), .C(n_544), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_551), .Y(n_553) );
INVx2_ASAP7_75t_SL g554 ( .A(n_552), .Y(n_554) );
OAI22x1_ASAP7_75t_L g555 ( .A1(n_554), .A2(n_543), .B1(n_545), .B2(n_548), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_555), .A2(n_553), .B1(n_518), .B2(n_539), .Y(n_556) );
OAI21xp5_ASAP7_75t_L g557 ( .A1(n_556), .A2(n_535), .B(n_192), .Y(n_557) );
AOI22xp33_ASAP7_75t_SL g558 ( .A1(n_557), .A2(n_151), .B1(n_546), .B2(n_554), .Y(n_558) );
endmodule