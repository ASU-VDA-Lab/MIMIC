module fake_jpeg_776_n_113 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_113);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_113;

wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx11_ASAP7_75t_R g30 ( 
.A(n_20),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_21),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_22),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx16f_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_27),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_39),
.Y(n_40)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_39),
.Y(n_41)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_36),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_42),
.B(n_31),
.Y(n_51)
);

BUFx8_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_0),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_29),
.Y(n_52)
);

BUFx24_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx6_ASAP7_75t_SL g46 ( 
.A(n_45),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_43),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_32),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_52),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_45),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_62),
.Y(n_69)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_64),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_29),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_60),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_72),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_55),
.A2(n_32),
.B1(n_33),
.B2(n_37),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_70),
.A2(n_38),
.B1(n_50),
.B2(n_34),
.Y(n_77)
);

A2O1A1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_57),
.A2(n_37),
.B(n_33),
.C(n_35),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_71),
.B(n_50),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_61),
.A2(n_49),
.B(n_50),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_30),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_10),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_61),
.A2(n_38),
.B1(n_34),
.B2(n_35),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_75),
.A2(n_26),
.B1(n_24),
.B2(n_23),
.Y(n_85)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_78),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_73),
.B(n_0),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_79),
.B(n_80),
.Y(n_89)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_84),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_28),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_83),
.B(n_86),
.C(n_71),
.Y(n_88)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_85),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_SL g86 ( 
.A(n_69),
.B(n_18),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_88),
.B(n_91),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_82),
.A2(n_75),
.B1(n_70),
.B2(n_3),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_90),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_86),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_85),
.B(n_1),
.Y(n_95)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_95),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_79),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_96),
.A2(n_5),
.B(n_6),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_97),
.B(n_100),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_93),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_98),
.A2(n_102),
.B1(n_94),
.B2(n_90),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_SL g100 ( 
.A(n_93),
.B(n_4),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_103),
.B(n_104),
.C(n_100),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_99),
.B(n_87),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_106),
.A2(n_105),
.B1(n_101),
.B2(n_92),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_107),
.B(n_104),
.Y(n_108)
);

AOI31xp67_ASAP7_75t_SL g109 ( 
.A1(n_108),
.A2(n_88),
.A3(n_89),
.B(n_12),
.Y(n_109)
);

A2O1A1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_109),
.A2(n_13),
.B(n_17),
.C(n_8),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_6),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_111),
.B(n_7),
.C(n_8),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_112),
.B(n_7),
.Y(n_113)
);


endmodule