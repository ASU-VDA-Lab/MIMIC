module real_jpeg_5303_n_7 (n_5, n_4, n_0, n_1, n_2, n_6, n_28, n_29, n_3, n_7);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_6;
input n_28;
input n_29;
input n_3;

output n_7;

wire n_17;
wire n_8;
wire n_21;
wire n_10;
wire n_9;
wire n_12;
wire n_24;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_22;
wire n_18;
wire n_26;
wire n_20;
wire n_19;
wire n_16;
wire n_15;
wire n_13;

INVx5_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

AOI221xp5_ASAP7_75t_L g7 ( 
.A1(n_1),
.A2(n_8),
.B1(n_17),
.B2(n_19),
.C(n_23),
.Y(n_7)
);

OAI32xp33_ASAP7_75t_L g17 ( 
.A1(n_1),
.A2(n_2),
.A3(n_18),
.B1(n_19),
.B2(n_22),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_L g10 ( 
.A1(n_3),
.A2(n_11),
.B(n_14),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g12 ( 
.A(n_6),
.B(n_28),
.Y(n_12)
);

O2A1O1Ixp33_ASAP7_75t_L g23 ( 
.A1(n_8),
.A2(n_19),
.B(n_24),
.C(n_25),
.Y(n_23)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_9),
.Y(n_8)
);

MAJIxp5_ASAP7_75t_L g9 ( 
.A(n_10),
.B(n_15),
.C(n_16),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_SL g11 ( 
.A(n_12),
.B(n_13),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_12),
.B(n_13),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_18),
.B(n_22),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_18),
.B(n_22),
.Y(n_26)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_29),
.Y(n_13)
);


endmodule