module real_jpeg_28959_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_113;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_103;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_111;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_0),
.B(n_21),
.Y(n_40)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_0),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_1),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_1),
.A2(n_28),
.B1(n_50),
.B2(n_51),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_1),
.A2(n_21),
.B1(n_23),
.B2(n_28),
.Y(n_106)
);

BUFx8_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_3),
.A2(n_25),
.B1(n_26),
.B2(n_35),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

A2O1A1Ixp33_ASAP7_75t_L g56 ( 
.A1(n_3),
.A2(n_34),
.B(n_50),
.C(n_57),
.Y(n_56)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_3),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_4),
.A2(n_21),
.B1(n_23),
.B2(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_4),
.A2(n_25),
.B1(n_26),
.B2(n_38),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_5),
.A2(n_21),
.B1(n_23),
.B2(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

OAI32xp33_ASAP7_75t_L g89 ( 
.A1(n_6),
.A2(n_23),
.A3(n_25),
.B1(n_90),
.B2(n_91),
.Y(n_89)
);

BUFx24_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_8),
.A2(n_25),
.B1(n_26),
.B2(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_8),
.A2(n_21),
.B1(n_23),
.B2(n_30),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_9),
.A2(n_21),
.B1(n_23),
.B2(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_9),
.Y(n_76)
);

INVx11_ASAP7_75t_SL g22 ( 
.A(n_10),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_11),
.B(n_33),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_11),
.A2(n_50),
.B(n_53),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_11),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_11),
.A2(n_25),
.B(n_87),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_11),
.B(n_25),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_11),
.A2(n_39),
.B1(n_45),
.B2(n_106),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_81),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_79),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_46),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_15),
.B(n_46),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_31),
.C(n_36),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_16),
.A2(n_31),
.B1(n_32),
.B2(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_16),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_27),
.B2(n_29),
.Y(n_16)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_17),
.A2(n_18),
.B1(n_27),
.B2(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_24),
.Y(n_17)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_18),
.B(n_55),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_20),
.B1(n_21),
.B2(n_23),
.Y(n_18)
);

OAI22xp33_ASAP7_75t_L g24 ( 
.A1(n_19),
.A2(n_20),
.B1(n_25),
.B2(n_26),
.Y(n_24)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_20),
.B(n_21),
.Y(n_91)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_21),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_21),
.B(n_111),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_25),
.B(n_71),
.Y(n_70)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI32xp33_ASAP7_75t_L g69 ( 
.A1(n_26),
.A2(n_50),
.A3(n_54),
.B1(n_58),
.B2(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_29),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_34),
.A2(n_49),
.B1(n_56),
.B2(n_60),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_36),
.B(n_93),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_37),
.A2(n_39),
.B1(n_41),
.B2(n_43),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_37),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_39),
.A2(n_41),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_39),
.A2(n_73),
.B1(n_99),
.B2(n_106),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_40),
.A2(n_98),
.B1(n_100),
.B2(n_101),
.Y(n_97)
);

INVx5_ASAP7_75t_SL g43 ( 
.A(n_44),
.Y(n_43)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_47),
.A2(n_68),
.B1(n_77),
.B2(n_78),
.Y(n_46)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_61),
.B1(n_66),
.B2(n_67),
.Y(n_47)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_58),
.Y(n_57)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_51),
.B(n_55),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_55),
.B(n_112),
.Y(n_111)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_63),
.B1(n_64),
.B2(n_65),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_68),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_72),
.Y(n_68)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_73),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_82),
.A2(n_95),
.B(n_116),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_92),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_83),
.B(n_92),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_84),
.B(n_88),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_84),
.A2(n_85),
.B1(n_88),
.B2(n_89),
.Y(n_102)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_87),
.Y(n_90)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_103),
.B(n_115),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_102),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_97),
.B(n_102),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_104),
.A2(n_108),
.B(n_114),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_107),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_105),
.B(n_107),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_109),
.B(n_110),
.Y(n_108)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);


endmodule