module real_jpeg_1190_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_1),
.A2(n_58),
.B1(n_59),
.B2(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_1),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_1),
.A2(n_34),
.B1(n_36),
.B2(n_71),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_1),
.A2(n_28),
.B1(n_29),
.B2(n_71),
.Y(n_169)
);

OAI22xp33_ASAP7_75t_L g213 ( 
.A1(n_1),
.A2(n_45),
.B1(n_49),
.B2(n_71),
.Y(n_213)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_2),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_3),
.A2(n_58),
.B1(n_59),
.B2(n_177),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_3),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_3),
.A2(n_34),
.B1(n_36),
.B2(n_177),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_3),
.A2(n_28),
.B1(n_29),
.B2(n_177),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_3),
.A2(n_45),
.B1(n_49),
.B2(n_177),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_4),
.A2(n_34),
.B1(n_36),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_4),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_4),
.A2(n_38),
.B1(n_58),
.B2(n_59),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_4),
.A2(n_28),
.B1(n_29),
.B2(n_38),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_4),
.A2(n_38),
.B1(n_45),
.B2(n_49),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_6),
.A2(n_58),
.B1(n_59),
.B2(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_6),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_6),
.A2(n_34),
.B1(n_36),
.B2(n_151),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_6),
.A2(n_28),
.B1(n_29),
.B2(n_151),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_6),
.A2(n_45),
.B1(n_49),
.B2(n_151),
.Y(n_250)
);

BUFx8_ASAP7_75t_L g60 ( 
.A(n_7),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_8),
.A2(n_58),
.B1(n_59),
.B2(n_66),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_8),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_8),
.A2(n_34),
.B1(n_36),
.B2(n_66),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_8),
.A2(n_28),
.B1(n_29),
.B2(n_66),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_8),
.A2(n_45),
.B1(n_49),
.B2(n_66),
.Y(n_189)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_11),
.A2(n_58),
.B1(n_59),
.B2(n_196),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_11),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_11),
.A2(n_34),
.B1(n_36),
.B2(n_196),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_11),
.A2(n_28),
.B1(n_29),
.B2(n_196),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_11),
.A2(n_45),
.B1(n_49),
.B2(n_196),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_12),
.B(n_58),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_12),
.B(n_84),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_12),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_12),
.A2(n_58),
.B(n_186),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_12),
.B(n_27),
.Y(n_248)
);

AOI21xp33_ASAP7_75t_L g255 ( 
.A1(n_12),
.A2(n_36),
.B(n_256),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_12),
.B(n_45),
.C(n_48),
.Y(n_264)
);

OAI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_12),
.A2(n_28),
.B1(n_29),
.B2(n_222),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_12),
.B(n_102),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_12),
.B(n_43),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_13),
.A2(n_58),
.B1(n_59),
.B2(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_13),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_13),
.A2(n_34),
.B1(n_36),
.B2(n_68),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_13),
.A2(n_28),
.B1(n_29),
.B2(n_68),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_13),
.A2(n_45),
.B1(n_49),
.B2(n_68),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_14),
.A2(n_34),
.B1(n_36),
.B2(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_14),
.A2(n_28),
.B1(n_29),
.B2(n_41),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_14),
.A2(n_41),
.B1(n_45),
.B2(n_49),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_15),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_16),
.A2(n_58),
.B1(n_59),
.B2(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_16),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_16),
.A2(n_34),
.B1(n_36),
.B2(n_112),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_16),
.A2(n_28),
.B1(n_29),
.B2(n_112),
.Y(n_218)
);

OAI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_16),
.A2(n_45),
.B1(n_49),
.B2(n_112),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_90),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_88),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_77),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_21),
.B(n_77),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_69),
.C(n_72),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_22),
.A2(n_69),
.B1(n_120),
.B2(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_22),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_54),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_42),
.B2(n_53),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_25),
.B(n_42),
.C(n_54),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_37),
.B1(n_39),
.B2(n_40),
.Y(n_25)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_26),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_26),
.A2(n_39),
.B1(n_117),
.B2(n_146),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_26),
.A2(n_39),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_26),
.A2(n_39),
.B1(n_207),
.B2(n_208),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_26),
.A2(n_39),
.B1(n_192),
.B2(n_208),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_26),
.A2(n_39),
.B1(n_207),
.B2(n_255),
.Y(n_254)
);

OR2x2_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_33),
.Y(n_26)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_27),
.A2(n_74),
.B1(n_75),
.B2(n_76),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_27),
.A2(n_75),
.B(n_80),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_27),
.A2(n_74),
.B1(n_75),
.B2(n_116),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_27),
.A2(n_75),
.B1(n_147),
.B2(n_174),
.Y(n_173)
);

AO22x2_ASAP7_75t_SL g27 ( 
.A1(n_28),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_27)
);

OAI22xp33_ASAP7_75t_L g51 ( 
.A1(n_28),
.A2(n_29),
.B1(n_47),
.B2(n_48),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_28),
.B(n_32),
.Y(n_223)
);

INVx4_ASAP7_75t_SL g28 ( 
.A(n_29),
.Y(n_28)
);

OAI32xp33_ASAP7_75t_L g220 ( 
.A1(n_29),
.A2(n_31),
.A3(n_36),
.B1(n_221),
.B2(n_223),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_29),
.B(n_264),
.Y(n_263)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx3_ASAP7_75t_SL g32 ( 
.A(n_31),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g33 ( 
.A1(n_31),
.A2(n_32),
.B1(n_34),
.B2(n_36),
.Y(n_33)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

OA22x2_ASAP7_75t_L g64 ( 
.A1(n_34),
.A2(n_36),
.B1(n_61),
.B2(n_63),
.Y(n_64)
);

NAND2xp33_ASAP7_75t_SL g187 ( 
.A(n_34),
.B(n_61),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_34),
.B(n_222),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

AOI32xp33_ASAP7_75t_L g185 ( 
.A1(n_36),
.A2(n_59),
.A3(n_63),
.B1(n_186),
.B2(n_187),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_37),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_40),
.Y(n_80)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_42),
.B(n_69),
.C(n_73),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_42),
.A2(n_53),
.B1(n_73),
.B2(n_123),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_50),
.B(n_52),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_43),
.A2(n_50),
.B1(n_107),
.B2(n_108),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_43),
.A2(n_50),
.B1(n_52),
.B2(n_108),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_43),
.A2(n_50),
.B1(n_107),
.B2(n_143),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_43),
.A2(n_50),
.B1(n_216),
.B2(n_218),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_43),
.A2(n_50),
.B1(n_218),
.B2(n_238),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_43),
.A2(n_50),
.B1(n_246),
.B2(n_247),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_43),
.A2(n_50),
.B1(n_246),
.B2(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_51),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_44),
.A2(n_144),
.B1(n_169),
.B2(n_170),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_44),
.A2(n_170),
.B1(n_217),
.B2(n_258),
.Y(n_257)
);

OA22x2_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_44)
);

INVx4_ASAP7_75t_SL g49 ( 
.A(n_45),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_45),
.B(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_45),
.B(n_274),
.Y(n_273)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_50),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_64),
.B1(n_65),
.B2(n_67),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_55),
.A2(n_64),
.B1(n_65),
.B2(n_70),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_55),
.A2(n_64),
.B1(n_70),
.B2(n_111),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_55),
.A2(n_64),
.B1(n_111),
.B2(n_149),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_55),
.A2(n_64),
.B1(n_195),
.B2(n_197),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_55),
.A2(n_64),
.B1(n_195),
.B2(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_56),
.A2(n_82),
.B1(n_83),
.B2(n_84),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_56),
.A2(n_84),
.B1(n_150),
.B2(n_176),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_64),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_59),
.B1(n_61),
.B2(n_63),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_61),
.Y(n_63)
);

BUFx4f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_67),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_69),
.A2(n_120),
.B1(n_121),
.B2(n_122),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_69),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_72),
.B(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_73),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_87),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_81),
.B1(n_85),
.B2(n_86),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_79),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_81),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

AO21x1_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_157),
.B(n_314),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_152),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_94),
.B(n_126),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_94),
.B(n_126),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_113),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_95),
.B(n_119),
.C(n_124),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_109),
.B(n_110),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_96),
.A2(n_97),
.B1(n_129),
.B2(n_130),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_105),
.Y(n_97)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_98),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_98),
.A2(n_109),
.B1(n_110),
.B2(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_98),
.A2(n_105),
.B1(n_106),
.B2(n_109),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_101),
.B(n_103),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_99),
.A2(n_101),
.B1(n_140),
.B2(n_172),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_99),
.A2(n_101),
.B1(n_225),
.B2(n_227),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_99),
.A2(n_101),
.B1(n_284),
.B2(n_285),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_100),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_100),
.A2(n_102),
.B1(n_104),
.B2(n_139),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_100),
.A2(n_102),
.B1(n_189),
.B2(n_190),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_100),
.A2(n_102),
.B1(n_189),
.B2(n_213),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_100),
.A2(n_102),
.B1(n_226),
.B2(n_250),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_100),
.A2(n_102),
.B1(n_222),
.B2(n_276),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_100),
.A2(n_102),
.B1(n_276),
.B2(n_280),
.Y(n_279)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_110),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_119),
.B1(n_124),
.B2(n_125),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_114),
.Y(n_124)
);

OAI21xp33_ASAP7_75t_L g133 ( 
.A1(n_114),
.A2(n_115),
.B(n_118),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_118),
.Y(n_114)
);

INVxp33_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_119),
.Y(n_125)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_132),
.C(n_134),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_127),
.A2(n_128),
.B1(n_132),
.B2(n_133),
.Y(n_160)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_134),
.B(n_160),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_145),
.C(n_148),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_135),
.A2(n_136),
.B1(n_163),
.B2(n_164),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_141),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_137),
.A2(n_138),
.B1(n_141),
.B2(n_142),
.Y(n_198)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_145),
.B(n_148),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_152),
.A2(n_315),
.B(n_316),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_153),
.B(n_156),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_153),
.B(n_156),
.Y(n_316)
);

AO21x1_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_178),
.B(n_313),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_161),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_159),
.B(n_161),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_165),
.C(n_166),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_162),
.B(n_165),
.Y(n_200)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_163),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_166),
.B(n_200),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_173),
.C(n_175),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_167),
.B(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_168),
.B(n_171),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_168),
.B(n_171),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_169),
.Y(n_238)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_172),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_173),
.B(n_175),
.Y(n_182)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_174),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_176),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_201),
.B(n_312),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_199),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_180),
.B(n_199),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_183),
.C(n_198),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_181),
.B(n_198),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_183),
.B(n_299),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_191),
.C(n_194),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g301 ( 
.A(n_184),
.B(n_302),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_188),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_185),
.B(n_188),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_191),
.B(n_194),
.Y(n_302)
);

AOI31xp33_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_296),
.A3(n_305),
.B(n_309),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_241),
.B(n_295),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_228),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_204),
.B(n_228),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_215),
.C(n_219),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_205),
.B(n_292),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_209),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_206),
.B(n_210),
.C(n_214),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_211),
.B1(n_212),
.B2(n_214),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_212),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_213),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_215),
.B(n_219),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_224),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_220),
.B(n_224),
.Y(n_252)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_221),
.Y(n_256)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_232),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_230),
.B(n_231),
.C(n_232),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_235),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_233),
.B(n_236),
.C(n_240),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_237),
.B1(n_239),
.B2(n_240),
.Y(n_235)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_236),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_237),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_242),
.A2(n_290),
.B(n_294),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_259),
.B(n_289),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_251),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_244),
.B(n_251),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_248),
.C(n_249),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_245),
.B(n_248),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_247),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_249),
.B(n_269),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_250),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_252),
.B(n_254),
.C(n_257),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_257),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_260),
.A2(n_270),
.B(n_288),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_268),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_261),
.B(n_268),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_265),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_262),
.A2(n_263),
.B1(n_265),
.B2(n_266),
.Y(n_286)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_282),
.B(n_287),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_277),
.B(n_281),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_275),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_278),
.B(n_279),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_280),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_286),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_283),
.B(n_286),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_291),
.B(n_293),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_291),
.B(n_293),
.Y(n_294)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_297),
.A2(n_310),
.B(n_311),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_298),
.B(n_300),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_298),
.B(n_300),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_303),
.C(n_304),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_301),
.B(n_308),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_303),
.B(n_304),
.Y(n_308)
);

OR2x2_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_306),
.B(n_307),
.Y(n_310)
);


endmodule