module real_jpeg_14427_n_12 (n_5, n_4, n_8, n_0, n_280, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_280;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_78;
wire n_83;
wire n_249;
wire n_215;
wire n_176;
wire n_166;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_238;
wire n_178;
wire n_67;
wire n_79;
wire n_76;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_70;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_216;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_257;
wire n_25;
wire n_217;
wire n_210;
wire n_53;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;
wire n_16;

INVx4_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_2),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_3),
.A2(n_43),
.B1(n_45),
.B2(n_46),
.Y(n_42)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_3),
.A2(n_26),
.B1(n_27),
.B2(n_45),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_3),
.A2(n_45),
.B1(n_100),
.B2(n_101),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_3),
.A2(n_45),
.B1(n_149),
.B2(n_150),
.Y(n_183)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_5),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_6),
.A2(n_26),
.B1(n_27),
.B2(n_37),
.Y(n_36)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_6),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_6),
.A2(n_37),
.B1(n_43),
.B2(n_46),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_6),
.A2(n_37),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_6),
.A2(n_37),
.B1(n_149),
.B2(n_150),
.Y(n_162)
);

BUFx12_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_8),
.A2(n_26),
.B1(n_27),
.B2(n_30),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_8),
.B(n_55),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_8),
.B(n_27),
.C(n_48),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_8),
.A2(n_30),
.B1(n_43),
.B2(n_46),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_8),
.B(n_31),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_8),
.B(n_47),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_8),
.A2(n_30),
.B1(n_100),
.B2(n_101),
.Y(n_106)
);

O2A1O1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_8),
.A2(n_57),
.B(n_101),
.C(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_8),
.B(n_128),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_8),
.A2(n_30),
.B1(n_149),
.B2(n_150),
.Y(n_167)
);

BUFx2_ASAP7_75t_L g130 ( 
.A(n_9),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_10),
.A2(n_26),
.B1(n_27),
.B2(n_155),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_10),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_10),
.A2(n_43),
.B1(n_46),
.B2(n_155),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_10),
.A2(n_100),
.B1(n_101),
.B2(n_155),
.Y(n_254)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_257),
.Y(n_12)
);

AOI21xp5_ASAP7_75t_SL g13 ( 
.A1(n_14),
.A2(n_238),
.B(n_256),
.Y(n_13)
);

OAI21xp5_ASAP7_75t_SL g14 ( 
.A1(n_15),
.A2(n_217),
.B(n_237),
.Y(n_14)
);

AOI321xp33_ASAP7_75t_SL g15 ( 
.A1(n_16),
.A2(n_178),
.A3(n_210),
.B1(n_215),
.B2(n_216),
.C(n_280),
.Y(n_15)
);

OAI21xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_139),
.B(n_177),
.Y(n_16)
);

AOI21xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_116),
.B(n_138),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_93),
.B(n_115),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_71),
.B(n_92),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_62),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_21),
.B(n_62),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_38),
.B1(n_39),
.B2(n_61),
.Y(n_21)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_33),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_23),
.B(n_89),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_31),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_25),
.B(n_35),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_25),
.A2(n_32),
.B(n_35),
.Y(n_111)
);

AO22x1_ASAP7_75t_L g47 ( 
.A1(n_26),
.A2(n_27),
.B1(n_48),
.B2(n_49),
.Y(n_47)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_32),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_27),
.B(n_75),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI21xp33_ASAP7_75t_L g113 ( 
.A1(n_30),
.A2(n_46),
.B(n_58),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_30),
.B(n_101),
.C(n_129),
.Y(n_148)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_32),
.B(n_36),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_32),
.B(n_82),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_32),
.A2(n_89),
.B(n_154),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_34),
.B(n_81),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_36),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_35),
.B(n_82),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_35),
.A2(n_154),
.B(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_40),
.A2(n_54),
.B1(n_59),
.B2(n_60),
.Y(n_39)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_50),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_41),
.B(n_68),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_41),
.A2(n_175),
.B(n_204),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_42),
.B(n_47),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_42),
.B(n_51),
.Y(n_108)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_43),
.A2(n_46),
.B1(n_48),
.B2(n_49),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_43),
.A2(n_46),
.B1(n_57),
.B2(n_58),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_47),
.B(n_53),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_47),
.B(n_69),
.Y(n_120)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_47),
.Y(n_176)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_48),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_50),
.B(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_51),
.B(n_53),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_51),
.B(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_51),
.Y(n_175)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_54),
.B(n_59),
.C(n_61),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_55),
.B(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_55),
.B(n_106),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_55),
.A2(n_103),
.B(n_106),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_55),
.A2(n_171),
.B(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_56),
.B(n_105),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_56),
.B(n_133),
.Y(n_132)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_57),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_57),
.A2(n_58),
.B1(n_100),
.B2(n_101),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_66),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_63),
.A2(n_64),
.B1(n_66),
.B2(n_87),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_68),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_67),
.B(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_70),
.A2(n_175),
.B(n_176),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_85),
.B(n_91),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_79),
.B(n_84),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_76),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_78),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_78),
.B(n_81),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_80),
.B(n_83),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_80),
.B(n_83),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_81),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_88),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_86),
.B(n_88),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_90),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_95),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_95),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_109),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_107),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_97),
.B(n_107),
.C(n_109),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_102),
.Y(n_97)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_98),
.Y(n_172)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_99),
.Y(n_135)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_100),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_100),
.A2(n_101),
.B1(n_129),
.B2(n_130),
.Y(n_128)
);

INVxp33_ASAP7_75t_L g231 ( 
.A(n_102),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_103),
.B(n_106),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_104),
.B(n_135),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_104),
.B(n_133),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_104),
.A2(n_272),
.B(n_273),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_108),
.A2(n_176),
.B(n_204),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_108),
.B(n_120),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_111),
.B1(n_112),
.B2(n_114),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_110),
.A2(n_111),
.B1(n_234),
.B2(n_235),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_110),
.A2(n_111),
.B1(n_247),
.B2(n_248),
.Y(n_246)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_111),
.B(n_112),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_111),
.B(n_234),
.Y(n_245)
);

AOI21xp33_ASAP7_75t_L g262 ( 
.A1(n_111),
.A2(n_245),
.B(n_247),
.Y(n_262)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_112),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_117),
.B(n_137),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_117),
.B(n_137),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_124),
.B1(n_125),
.B2(n_136),
.Y(n_117)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_118),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_119),
.A2(n_121),
.B1(n_122),
.B2(n_123),
.Y(n_118)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_119),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_121),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_121),
.B(n_122),
.C(n_124),
.Y(n_140)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx24_ASAP7_75t_SL g278 ( 
.A(n_125),
.Y(n_278)
);

FAx1_ASAP7_75t_SL g125 ( 
.A(n_126),
.B(n_127),
.CI(n_131),
.CON(n_125),
.SN(n_125)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_126),
.B(n_127),
.C(n_131),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_128),
.B(n_162),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_128),
.B(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_128),
.B(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_128),
.B(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_128),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_129),
.A2(n_130),
.B1(n_149),
.B2(n_150),
.Y(n_166)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_134),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_132),
.B(n_231),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_132),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_134),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_141),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_140),
.B(n_141),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_142),
.A2(n_143),
.B1(n_157),
.B2(n_158),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_145),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_144),
.B(n_145),
.C(n_157),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_147),
.B1(n_153),
.B2(n_156),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_146),
.B(n_156),
.Y(n_188)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_148),
.B(n_149),
.Y(n_147)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx13_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx12f_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_153),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_168),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_159),
.B(n_170),
.C(n_173),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_163),
.Y(n_159)
);

INVxp33_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_161),
.B(n_197),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_162),
.B(n_165),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_163),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_164),
.B(n_167),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_164),
.A2(n_167),
.B(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_165),
.B(n_183),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_167),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_169),
.A2(n_170),
.B1(n_173),
.B2(n_174),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_173),
.A2(n_174),
.B1(n_271),
.B2(n_274),
.Y(n_270)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_179),
.B(n_205),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_179),
.B(n_205),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_189),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_180),
.B(n_190),
.C(n_201),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_185),
.C(n_188),
.Y(n_180)
);

FAx1_ASAP7_75t_SL g207 ( 
.A(n_181),
.B(n_185),
.CI(n_188),
.CON(n_207),
.SN(n_207)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_184),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_182),
.B(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_184),
.B(n_227),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_201),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_195),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_191),
.B(n_198),
.C(n_199),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_194),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_192),
.B(n_194),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_196),
.A2(n_198),
.B1(n_199),
.B2(n_200),
.Y(n_195)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_196),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_198),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_202),
.B(n_203),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_208),
.C(n_209),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_206),
.A2(n_207),
.B1(n_212),
.B2(n_213),
.Y(n_211)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

BUFx24_ASAP7_75t_SL g277 ( 
.A(n_207),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_208),
.B(n_209),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_211),
.B(n_214),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_211),
.B(n_214),
.Y(n_215)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_218),
.B(n_219),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_236),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_222),
.B1(n_232),
.B2(n_233),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_221),
.B(n_233),
.C(n_236),
.Y(n_239)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_223),
.B(n_225),
.C(n_230),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_225),
.A2(n_226),
.B1(n_229),
.B2(n_230),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_234),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_239),
.B(n_240),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_241),
.B(n_243),
.C(n_251),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_243),
.A2(n_244),
.B1(n_250),
.B2(n_251),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_252),
.A2(n_253),
.B(n_255),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_252),
.B(n_253),
.Y(n_255)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_254),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_255),
.A2(n_264),
.B1(n_265),
.B2(n_275),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_255),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_276),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_260),
.B(n_261),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_267),
.B1(n_269),
.B2(n_270),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_271),
.Y(n_274)
);


endmodule