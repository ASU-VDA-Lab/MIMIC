module real_aes_3013_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_453;
wire n_374;
wire n_379;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_330;
wire n_388;
wire n_395;
wire n_332;
wire n_292;
wire n_400;
wire n_116;
wire n_94;
wire n_462;
wire n_289;
wire n_280;
wire n_333;
wire n_213;
wire n_478;
wire n_356;
wire n_408;
wire n_184;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_174;
wire n_104;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_178;
wire n_409;
wire n_298;
wire n_439;
wire n_506;
wire n_297;
wire n_383;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_502;
wire n_434;
wire n_505;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_87;
wire n_171;
wire n_78;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_484;
wire n_326;
wire n_492;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_456;
wire n_359;
wire n_312;
wire n_266;
wire n_183;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_313;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_166;
wire n_103;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_0), .B(n_176), .Y(n_233) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_1), .A2(n_159), .B(n_209), .Y(n_208) );
AO22x2_ASAP7_75t_L g98 ( .A1(n_2), .A2(n_54), .B1(n_88), .B2(n_99), .Y(n_98) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_3), .B(n_166), .Y(n_222) );
INVx1_ASAP7_75t_L g142 ( .A(n_4), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_5), .B(n_166), .Y(n_186) );
AO22x2_ASAP7_75t_L g95 ( .A1(n_6), .A2(n_21), .B1(n_88), .B2(n_96), .Y(n_95) );
NAND2xp33_ASAP7_75t_L g203 ( .A(n_7), .B(n_170), .Y(n_203) );
INVx2_ASAP7_75t_L g156 ( .A(n_8), .Y(n_156) );
AOI221x1_ASAP7_75t_L g245 ( .A1(n_9), .A2(n_16), .B1(n_159), .B2(n_176), .C(n_246), .Y(n_245) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_10), .B(n_176), .Y(n_199) );
AO21x2_ASAP7_75t_L g196 ( .A1(n_11), .A2(n_197), .B(n_198), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_12), .B(n_189), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_13), .B(n_166), .Y(n_165) );
INVx1_ASAP7_75t_L g479 ( .A(n_13), .Y(n_479) );
AO21x1_ASAP7_75t_L g217 ( .A1(n_14), .A2(n_176), .B(n_218), .Y(n_217) );
AOI22xp5_ASAP7_75t_L g127 ( .A1(n_15), .A2(n_69), .B1(n_128), .B2(n_129), .Y(n_127) );
NAND2x1_ASAP7_75t_L g231 ( .A(n_17), .B(n_166), .Y(n_231) );
AO222x2_ASAP7_75t_L g83 ( .A1(n_18), .A2(n_23), .B1(n_55), .B2(n_84), .C1(n_100), .C2(n_103), .Y(n_83) );
NAND2x1_ASAP7_75t_L g185 ( .A(n_19), .B(n_170), .Y(n_185) );
AOI22xp33_ASAP7_75t_SL g132 ( .A1(n_20), .A2(n_59), .B1(n_133), .B2(n_134), .Y(n_132) );
OAI221xp5_ASAP7_75t_L g484 ( .A1(n_21), .A2(n_54), .B1(n_60), .B2(n_485), .C(n_487), .Y(n_484) );
AOI22xp33_ASAP7_75t_SL g114 ( .A1(n_22), .A2(n_48), .B1(n_115), .B2(n_118), .Y(n_114) );
OR2x2_ASAP7_75t_L g155 ( .A(n_24), .B(n_66), .Y(n_155) );
OA21x2_ASAP7_75t_L g194 ( .A1(n_24), .A2(n_66), .B(n_156), .Y(n_194) );
AOI22xp33_ASAP7_75t_L g108 ( .A1(n_25), .A2(n_26), .B1(n_109), .B2(n_112), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_27), .B(n_170), .Y(n_211) );
INVx3_ASAP7_75t_L g88 ( .A(n_28), .Y(n_88) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_29), .B(n_166), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_30), .B(n_170), .Y(n_221) );
AOI22xp5_ASAP7_75t_L g135 ( .A1(n_31), .A2(n_53), .B1(n_136), .B2(n_137), .Y(n_135) );
AOI21xp5_ASAP7_75t_L g263 ( .A1(n_32), .A2(n_159), .B(n_264), .Y(n_263) );
INVx1_ASAP7_75t_SL g89 ( .A(n_33), .Y(n_89) );
INVx1_ASAP7_75t_L g144 ( .A(n_34), .Y(n_144) );
AND2x2_ASAP7_75t_L g160 ( .A(n_34), .B(n_161), .Y(n_160) );
AND2x2_ASAP7_75t_L g174 ( .A(n_34), .B(n_142), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g267 ( .A(n_35), .B(n_176), .Y(n_267) );
INVx1_ASAP7_75t_L g508 ( .A(n_35), .Y(n_508) );
CKINVDCx20_ASAP7_75t_R g179 ( .A(n_36), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_37), .B(n_170), .Y(n_265) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_38), .A2(n_159), .B(n_184), .Y(n_183) );
AO22x2_ASAP7_75t_L g91 ( .A1(n_39), .A2(n_60), .B1(n_88), .B2(n_92), .Y(n_91) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_40), .B(n_170), .Y(n_232) );
INVx1_ASAP7_75t_L g163 ( .A(n_41), .Y(n_163) );
INVx1_ASAP7_75t_L g172 ( .A(n_41), .Y(n_172) );
AOI22xp33_ASAP7_75t_SL g123 ( .A1(n_42), .A2(n_44), .B1(n_124), .B2(n_125), .Y(n_123) );
INVx1_ASAP7_75t_L g90 ( .A(n_43), .Y(n_90) );
OAI22xp5_ASAP7_75t_L g469 ( .A1(n_45), .A2(n_470), .B1(n_471), .B2(n_472), .Y(n_469) );
INVx1_ASAP7_75t_L g471 ( .A(n_45), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_46), .B(n_166), .Y(n_248) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_47), .A2(n_159), .B(n_230), .Y(n_229) );
AOI22xp5_ASAP7_75t_L g476 ( .A1(n_49), .A2(n_62), .B1(n_477), .B2(n_478), .Y(n_476) );
INVx1_ASAP7_75t_L g478 ( .A(n_49), .Y(n_478) );
AO21x1_ASAP7_75t_L g219 ( .A1(n_50), .A2(n_159), .B(n_220), .Y(n_219) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_51), .B(n_176), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_52), .B(n_176), .Y(n_187) );
INVxp33_ASAP7_75t_L g489 ( .A(n_54), .Y(n_489) );
AND2x2_ASAP7_75t_L g268 ( .A(n_56), .B(n_190), .Y(n_268) );
INVx1_ASAP7_75t_L g161 ( .A(n_57), .Y(n_161) );
INVx1_ASAP7_75t_L g168 ( .A(n_57), .Y(n_168) );
AND2x2_ASAP7_75t_L g191 ( .A(n_58), .B(n_192), .Y(n_191) );
INVxp67_ASAP7_75t_L g488 ( .A(n_60), .Y(n_488) );
AOI22xp5_ASAP7_75t_L g79 ( .A1(n_61), .A2(n_80), .B1(n_81), .B2(n_138), .Y(n_79) );
CKINVDCx20_ASAP7_75t_R g138 ( .A(n_61), .Y(n_138) );
INVx1_ASAP7_75t_L g477 ( .A(n_62), .Y(n_477) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_63), .B(n_176), .Y(n_175) );
AND2x2_ASAP7_75t_L g205 ( .A(n_64), .B(n_192), .Y(n_205) );
AND2x2_ASAP7_75t_L g218 ( .A(n_65), .B(n_154), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_67), .B(n_170), .Y(n_169) );
AND2x2_ASAP7_75t_L g235 ( .A(n_68), .B(n_192), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_70), .B(n_166), .Y(n_266) );
AOI22xp5_ASAP7_75t_L g465 ( .A1(n_70), .A2(n_466), .B1(n_481), .B2(n_491), .Y(n_465) );
INVx1_ASAP7_75t_L g497 ( .A(n_70), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g158 ( .A1(n_71), .A2(n_159), .B(n_164), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_72), .B(n_170), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_73), .B(n_166), .Y(n_210) );
BUFx2_ASAP7_75t_L g470 ( .A(n_74), .Y(n_470) );
BUFx2_ASAP7_75t_SL g486 ( .A(n_75), .Y(n_486) );
AOI21xp5_ASAP7_75t_L g200 ( .A1(n_76), .A2(n_159), .B(n_201), .Y(n_200) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_139), .B1(n_145), .B2(n_462), .C(n_464), .Y(n_77) );
CKINVDCx20_ASAP7_75t_R g78 ( .A(n_79), .Y(n_78) );
OAI222xp33_ASAP7_75t_L g464 ( .A1(n_80), .A2(n_81), .B1(n_465), .B2(n_496), .C1(n_499), .C2(n_508), .Y(n_464) );
INVx1_ASAP7_75t_L g80 ( .A(n_81), .Y(n_80) );
NAND2x1_ASAP7_75t_L g81 ( .A(n_82), .B(n_121), .Y(n_81) );
NOR2x1_ASAP7_75t_L g82 ( .A(n_83), .B(n_107), .Y(n_82) );
AND2x4_ASAP7_75t_L g84 ( .A(n_85), .B(n_93), .Y(n_84) );
AND2x2_ASAP7_75t_L g112 ( .A(n_85), .B(n_113), .Y(n_112) );
AND2x2_ASAP7_75t_L g118 ( .A(n_85), .B(n_119), .Y(n_118) );
AND2x2_ASAP7_75t_L g85 ( .A(n_86), .B(n_91), .Y(n_85) );
HB1xp67_ASAP7_75t_L g101 ( .A(n_86), .Y(n_101) );
AND2x2_ASAP7_75t_L g105 ( .A(n_86), .B(n_106), .Y(n_105) );
INVx2_ASAP7_75t_L g111 ( .A(n_86), .Y(n_111) );
OAI22x1_ASAP7_75t_L g86 ( .A1(n_87), .A2(n_88), .B1(n_89), .B2(n_90), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
INVx1_ASAP7_75t_L g92 ( .A(n_88), .Y(n_92) );
INVx2_ASAP7_75t_L g96 ( .A(n_88), .Y(n_96) );
INVx1_ASAP7_75t_L g99 ( .A(n_88), .Y(n_99) );
INVx2_ASAP7_75t_L g106 ( .A(n_91), .Y(n_106) );
AND2x2_ASAP7_75t_L g110 ( .A(n_91), .B(n_111), .Y(n_110) );
BUFx2_ASAP7_75t_L g126 ( .A(n_91), .Y(n_126) );
AND2x6_ASAP7_75t_L g128 ( .A(n_93), .B(n_110), .Y(n_128) );
AND2x2_ASAP7_75t_L g133 ( .A(n_93), .B(n_105), .Y(n_133) );
AND2x2_ASAP7_75t_L g136 ( .A(n_93), .B(n_130), .Y(n_136) );
AND2x4_ASAP7_75t_L g93 ( .A(n_94), .B(n_97), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_95), .Y(n_94) );
AND2x2_ASAP7_75t_L g102 ( .A(n_95), .B(n_98), .Y(n_102) );
AND2x4_ASAP7_75t_L g104 ( .A(n_95), .B(n_97), .Y(n_104) );
INVx1_ASAP7_75t_L g117 ( .A(n_95), .Y(n_117) );
INVxp67_ASAP7_75t_L g113 ( .A(n_97), .Y(n_113) );
INVx2_ASAP7_75t_L g97 ( .A(n_98), .Y(n_97) );
AND2x2_ASAP7_75t_L g116 ( .A(n_98), .B(n_117), .Y(n_116) );
AND2x2_ASAP7_75t_SL g100 ( .A(n_101), .B(n_102), .Y(n_100) );
AND2x4_ASAP7_75t_L g125 ( .A(n_102), .B(n_126), .Y(n_125) );
AND2x4_ASAP7_75t_L g134 ( .A(n_102), .B(n_130), .Y(n_134) );
AND2x4_ASAP7_75t_L g103 ( .A(n_104), .B(n_105), .Y(n_103) );
AND2x2_ASAP7_75t_L g109 ( .A(n_104), .B(n_110), .Y(n_109) );
AND2x2_ASAP7_75t_L g137 ( .A(n_104), .B(n_130), .Y(n_137) );
AND2x4_ASAP7_75t_L g115 ( .A(n_105), .B(n_116), .Y(n_115) );
AND2x4_ASAP7_75t_L g130 ( .A(n_106), .B(n_111), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_108), .B(n_114), .Y(n_107) );
AND2x2_ASAP7_75t_SL g124 ( .A(n_110), .B(n_116), .Y(n_124) );
AND2x6_ASAP7_75t_L g129 ( .A(n_116), .B(n_130), .Y(n_129) );
HB1xp67_ASAP7_75t_L g120 ( .A(n_117), .Y(n_120) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
NOR2xp33_ASAP7_75t_L g121 ( .A(n_122), .B(n_131), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g122 ( .A(n_123), .B(n_127), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_132), .B(n_135), .Y(n_131) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
OR2x2_ASAP7_75t_SL g140 ( .A(n_141), .B(n_143), .Y(n_140) );
INVx1_ASAP7_75t_L g490 ( .A(n_141), .Y(n_490) );
HB1xp67_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
AND2x2_ASAP7_75t_L g162 ( .A(n_142), .B(n_163), .Y(n_162) );
AND3x1_ASAP7_75t_SL g483 ( .A(n_143), .B(n_484), .C(n_490), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_143), .B(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
NOR2x1p5_ASAP7_75t_L g503 ( .A(n_144), .B(n_504), .Y(n_503) );
HB1xp67_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
OR2x6_ASAP7_75t_L g146 ( .A(n_147), .B(n_360), .Y(n_146) );
NAND3xp33_ASAP7_75t_SL g147 ( .A(n_148), .B(n_272), .C(n_327), .Y(n_147) );
AOI221xp5_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_212), .B1(n_236), .B2(n_240), .C(n_250), .Y(n_148) );
AND2x2_ASAP7_75t_L g149 ( .A(n_150), .B(n_195), .Y(n_149) );
AND2x2_ASAP7_75t_SL g238 ( .A(n_150), .B(n_239), .Y(n_238) );
INVx2_ASAP7_75t_L g271 ( .A(n_150), .Y(n_271) );
AND2x2_ASAP7_75t_L g316 ( .A(n_150), .B(n_253), .Y(n_316) );
AND2x4_ASAP7_75t_L g150 ( .A(n_151), .B(n_180), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g304 ( .A(n_152), .Y(n_304) );
INVx1_ASAP7_75t_L g314 ( .A(n_152), .Y(n_314) );
AO21x2_ASAP7_75t_L g152 ( .A1(n_153), .A2(n_157), .B(n_178), .Y(n_152) );
NOR2xp33_ASAP7_75t_L g178 ( .A(n_153), .B(n_179), .Y(n_178) );
AO21x2_ASAP7_75t_L g278 ( .A1(n_153), .A2(n_157), .B(n_178), .Y(n_278) );
INVx1_ASAP7_75t_SL g153 ( .A(n_154), .Y(n_153) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_154), .A2(n_199), .B(n_200), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_154), .B(n_224), .Y(n_223) );
AND2x4_ASAP7_75t_L g154 ( .A(n_155), .B(n_156), .Y(n_154) );
AND2x2_ASAP7_75t_SL g190 ( .A(n_155), .B(n_156), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_158), .B(n_175), .Y(n_157) );
AND2x6_ASAP7_75t_L g159 ( .A(n_160), .B(n_162), .Y(n_159) );
AND2x6_ASAP7_75t_L g170 ( .A(n_161), .B(n_171), .Y(n_170) );
INVx2_ASAP7_75t_L g505 ( .A(n_161), .Y(n_505) );
AND2x4_ASAP7_75t_L g166 ( .A(n_163), .B(n_167), .Y(n_166) );
INVx2_ASAP7_75t_L g507 ( .A(n_163), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_169), .B(n_173), .Y(n_164) );
AND2x4_ASAP7_75t_L g177 ( .A(n_167), .B(n_171), .Y(n_177) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_173), .A2(n_185), .B(n_186), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_173), .A2(n_202), .B(n_203), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_173), .A2(n_210), .B(n_211), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_173), .A2(n_221), .B(n_222), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_173), .A2(n_231), .B(n_232), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_173), .A2(n_247), .B(n_248), .Y(n_246) );
AOI21xp5_ASAP7_75t_L g264 ( .A1(n_173), .A2(n_265), .B(n_266), .Y(n_264) );
INVx5_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
AND2x4_ASAP7_75t_L g176 ( .A(n_174), .B(n_177), .Y(n_176) );
HB1xp67_ASAP7_75t_L g463 ( .A(n_176), .Y(n_463) );
OR2x2_ASAP7_75t_L g293 ( .A(n_180), .B(n_196), .Y(n_293) );
NAND2x1p5_ASAP7_75t_L g324 ( .A(n_180), .B(n_239), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_180), .B(n_204), .Y(n_337) );
INVx2_ASAP7_75t_L g346 ( .A(n_180), .Y(n_346) );
AND2x2_ASAP7_75t_L g367 ( .A(n_180), .B(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g451 ( .A(n_180), .B(n_270), .Y(n_451) );
INVx4_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
AND2x2_ASAP7_75t_L g279 ( .A(n_181), .B(n_204), .Y(n_279) );
AND2x2_ASAP7_75t_L g412 ( .A(n_181), .B(n_239), .Y(n_412) );
HB1xp67_ASAP7_75t_L g438 ( .A(n_181), .Y(n_438) );
AO21x2_ASAP7_75t_L g181 ( .A1(n_182), .A2(n_188), .B(n_191), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_183), .B(n_187), .Y(n_182) );
CKINVDCx5p33_ASAP7_75t_R g188 ( .A(n_189), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_189), .A2(n_207), .B(n_208), .Y(n_206) );
OA21x2_ASAP7_75t_L g244 ( .A1(n_189), .A2(n_245), .B(n_249), .Y(n_244) );
OA21x2_ASAP7_75t_L g256 ( .A1(n_189), .A2(n_245), .B(n_249), .Y(n_256) );
BUFx6f_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVx3_ASAP7_75t_L g234 ( .A(n_192), .Y(n_234) );
INVx4_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
INVx3_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
BUFx4f_ASAP7_75t_L g197 ( .A(n_194), .Y(n_197) );
AND2x4_ASAP7_75t_L g366 ( .A(n_195), .B(n_367), .Y(n_366) );
AOI321xp33_ASAP7_75t_L g380 ( .A1(n_195), .A2(n_309), .A3(n_310), .B1(n_342), .B2(n_381), .C(n_384), .Y(n_380) );
AND2x2_ASAP7_75t_L g195 ( .A(n_196), .B(n_204), .Y(n_195) );
BUFx3_ASAP7_75t_L g237 ( .A(n_196), .Y(n_237) );
INVx2_ASAP7_75t_L g270 ( .A(n_196), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_196), .B(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g303 ( .A(n_196), .B(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g336 ( .A(n_196), .Y(n_336) );
INVx5_ASAP7_75t_L g239 ( .A(n_204), .Y(n_239) );
NOR2x1_ASAP7_75t_SL g288 ( .A(n_204), .B(n_278), .Y(n_288) );
BUFx2_ASAP7_75t_L g383 ( .A(n_204), .Y(n_383) );
OR2x6_ASAP7_75t_L g204 ( .A(n_205), .B(n_206), .Y(n_204) );
INVxp67_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_214), .B(n_225), .Y(n_213) );
NOR2xp33_ASAP7_75t_SL g281 ( .A(n_214), .B(n_282), .Y(n_281) );
NOR4xp25_ASAP7_75t_L g384 ( .A(n_214), .B(n_378), .C(n_382), .D(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g422 ( .A(n_214), .Y(n_422) );
AND2x2_ASAP7_75t_L g456 ( .A(n_214), .B(n_396), .Y(n_456) );
BUFx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
INVx2_ASAP7_75t_L g257 ( .A(n_215), .Y(n_257) );
INVx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
INVx2_ASAP7_75t_L g311 ( .A(n_216), .Y(n_311) );
OAI21x1_ASAP7_75t_SL g216 ( .A1(n_217), .A2(n_219), .B(n_223), .Y(n_216) );
INVx1_ASAP7_75t_L g224 ( .A(n_218), .Y(n_224) );
AOI33xp33_ASAP7_75t_L g452 ( .A1(n_225), .A2(n_254), .A3(n_285), .B1(n_301), .B2(n_407), .B3(n_453), .Y(n_452) );
INVx1_ASAP7_75t_SL g225 ( .A(n_226), .Y(n_225) );
AND2x2_ASAP7_75t_L g242 ( .A(n_226), .B(n_243), .Y(n_242) );
AND2x4_ASAP7_75t_L g252 ( .A(n_226), .B(n_253), .Y(n_252) );
BUFx3_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVx2_ASAP7_75t_L g259 ( .A(n_227), .Y(n_259) );
INVxp67_ASAP7_75t_L g340 ( .A(n_227), .Y(n_340) );
AND2x2_ASAP7_75t_L g396 ( .A(n_227), .B(n_261), .Y(n_396) );
AO21x2_ASAP7_75t_L g227 ( .A1(n_228), .A2(n_234), .B(n_235), .Y(n_227) );
AO21x2_ASAP7_75t_L g300 ( .A1(n_228), .A2(n_234), .B(n_235), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_229), .B(n_233), .Y(n_228) );
AO21x2_ASAP7_75t_L g261 ( .A1(n_234), .A2(n_262), .B(n_268), .Y(n_261) );
AO21x2_ASAP7_75t_L g297 ( .A1(n_234), .A2(n_262), .B(n_268), .Y(n_297) );
AOI21xp5_ASAP7_75t_L g417 ( .A1(n_236), .A2(n_418), .B(n_419), .Y(n_417) );
AND2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_238), .Y(n_236) );
AND2x2_ASAP7_75t_L g405 ( .A(n_237), .B(n_279), .Y(n_405) );
AND3x2_ASAP7_75t_L g407 ( .A(n_237), .B(n_291), .C(n_346), .Y(n_407) );
INVx3_ASAP7_75t_SL g359 ( .A(n_238), .Y(n_359) );
INVx4_ASAP7_75t_L g253 ( .A(n_239), .Y(n_253) );
AND2x2_ASAP7_75t_L g291 ( .A(n_239), .B(n_278), .Y(n_291) );
INVxp67_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
BUFx2_ASAP7_75t_L g285 ( .A(n_243), .Y(n_285) );
AND2x4_ASAP7_75t_L g310 ( .A(n_243), .B(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g373 ( .A(n_243), .B(n_261), .Y(n_373) );
INVx2_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
INVx2_ASAP7_75t_L g343 ( .A(n_244), .Y(n_343) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_244), .Y(n_365) );
O2A1O1Ixp33_ASAP7_75t_R g250 ( .A1(n_251), .A2(n_254), .B(n_258), .C(n_269), .Y(n_250) );
CKINVDCx16_ASAP7_75t_R g251 ( .A(n_252), .Y(n_251) );
AND2x2_ASAP7_75t_L g302 ( .A(n_253), .B(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_253), .B(n_314), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_253), .B(n_270), .Y(n_431) );
INVx1_ASAP7_75t_SL g254 ( .A(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g413 ( .A(n_255), .B(n_403), .Y(n_413) );
AND2x2_ASAP7_75t_SL g255 ( .A(n_256), .B(n_257), .Y(n_255) );
AND2x2_ASAP7_75t_L g260 ( .A(n_256), .B(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g282 ( .A(n_256), .B(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g298 ( .A(n_256), .B(n_299), .Y(n_298) );
AND2x4_ASAP7_75t_L g331 ( .A(n_256), .B(n_311), .Y(n_331) );
AND2x4_ASAP7_75t_L g296 ( .A(n_257), .B(n_297), .Y(n_296) );
OR2x2_ASAP7_75t_L g320 ( .A(n_257), .B(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g358 ( .A(n_257), .B(n_283), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_259), .B(n_260), .Y(n_258) );
AND2x2_ASAP7_75t_L g286 ( .A(n_259), .B(n_283), .Y(n_286) );
AND2x2_ASAP7_75t_L g301 ( .A(n_259), .B(n_261), .Y(n_301) );
BUFx2_ASAP7_75t_L g357 ( .A(n_259), .Y(n_357) );
AND2x2_ASAP7_75t_L g371 ( .A(n_259), .B(n_282), .Y(n_371) );
INVx2_ASAP7_75t_L g283 ( .A(n_261), .Y(n_283) );
NAND2xp5_ASAP7_75t_SL g262 ( .A(n_263), .B(n_267), .Y(n_262) );
OAI22xp33_ASAP7_75t_L g319 ( .A1(n_269), .A2(n_320), .B1(n_322), .B2(n_326), .Y(n_319) );
INVx2_ASAP7_75t_SL g350 ( .A(n_269), .Y(n_350) );
OR2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
AND2x2_ASAP7_75t_L g325 ( .A(n_270), .B(n_278), .Y(n_325) );
INVx1_ASAP7_75t_L g432 ( .A(n_271), .Y(n_432) );
NOR3xp33_ASAP7_75t_L g272 ( .A(n_273), .B(n_305), .C(n_319), .Y(n_272) );
OAI221xp5_ASAP7_75t_SL g273 ( .A1(n_274), .A2(n_280), .B1(n_284), .B2(n_287), .C(n_289), .Y(n_273) );
INVx1_ASAP7_75t_SL g274 ( .A(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g275 ( .A(n_276), .B(n_279), .Y(n_275) );
INVxp67_ASAP7_75t_SL g276 ( .A(n_277), .Y(n_276) );
INVx1_ASAP7_75t_L g333 ( .A(n_277), .Y(n_333) );
INVxp67_ASAP7_75t_SL g461 ( .A(n_277), .Y(n_461) );
INVx1_ASAP7_75t_L g424 ( .A(n_279), .Y(n_424) );
AND2x2_ASAP7_75t_SL g434 ( .A(n_279), .B(n_303), .Y(n_434) );
INVxp67_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_283), .B(n_311), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
OR2x2_ASAP7_75t_L g317 ( .A(n_285), .B(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g395 ( .A(n_285), .Y(n_395) );
AND2x2_ASAP7_75t_L g330 ( .A(n_286), .B(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g376 ( .A(n_288), .B(n_336), .Y(n_376) );
AND2x2_ASAP7_75t_L g453 ( .A(n_288), .B(n_451), .Y(n_453) );
AOI22xp5_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_294), .B1(n_301), .B2(n_302), .Y(n_289) );
AND2x4_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
INVx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
OR2x2_ASAP7_75t_L g312 ( .A(n_293), .B(n_313), .Y(n_312) );
INVx1_ASAP7_75t_SL g294 ( .A(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_296), .B(n_298), .Y(n_295) );
INVx2_ASAP7_75t_L g318 ( .A(n_296), .Y(n_318) );
AND2x4_ASAP7_75t_L g342 ( .A(n_296), .B(n_343), .Y(n_342) );
OAI21xp33_ASAP7_75t_SL g372 ( .A1(n_296), .A2(n_373), .B(n_374), .Y(n_372) );
AND2x2_ASAP7_75t_L g399 ( .A(n_296), .B(n_357), .Y(n_399) );
INVx2_ASAP7_75t_L g321 ( .A(n_297), .Y(n_321) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_297), .Y(n_354) );
INVx1_ASAP7_75t_SL g378 ( .A(n_298), .Y(n_378) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
BUFx2_ASAP7_75t_L g309 ( .A(n_300), .Y(n_309) );
AND2x4_ASAP7_75t_SL g403 ( .A(n_300), .B(n_321), .Y(n_403) );
AND2x2_ASAP7_75t_L g400 ( .A(n_303), .B(n_346), .Y(n_400) );
AND2x2_ASAP7_75t_L g426 ( .A(n_303), .B(n_412), .Y(n_426) );
HB1xp67_ASAP7_75t_L g348 ( .A(n_304), .Y(n_348) );
INVx1_ASAP7_75t_L g368 ( .A(n_304), .Y(n_368) );
OAI22xp33_ASAP7_75t_L g305 ( .A1(n_306), .A2(n_312), .B1(n_315), .B2(n_317), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g307 ( .A(n_308), .B(n_310), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_SL g326 ( .A(n_310), .B(n_321), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_310), .B(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g449 ( .A(n_310), .Y(n_449) );
INVx2_ASAP7_75t_SL g374 ( .A(n_312), .Y(n_374) );
AND2x2_ASAP7_75t_L g386 ( .A(n_314), .B(n_346), .Y(n_386) );
INVx2_ASAP7_75t_L g392 ( .A(n_314), .Y(n_392) );
INVxp33_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx2_ASAP7_75t_L g351 ( .A(n_317), .Y(n_351) );
NOR2xp33_ASAP7_75t_L g377 ( .A(n_320), .B(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g442 ( .A(n_320), .Y(n_442) );
INVx1_ASAP7_75t_L g370 ( .A(n_322), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_323), .B(n_325), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_323), .B(n_390), .Y(n_389) );
INVx2_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g381 ( .A(n_325), .B(n_382), .Y(n_381) );
AOI22xp5_ASAP7_75t_L g454 ( .A1(n_325), .A2(n_455), .B1(n_456), .B2(n_457), .Y(n_454) );
NOR3xp33_ASAP7_75t_L g327 ( .A(n_328), .B(n_349), .C(n_352), .Y(n_327) );
OAI221xp5_ASAP7_75t_L g328 ( .A1(n_329), .A2(n_332), .B1(n_334), .B2(n_338), .C(n_341), .Y(n_328) );
INVx1_ASAP7_75t_SL g329 ( .A(n_330), .Y(n_329) );
INVx1_ASAP7_75t_SL g447 ( .A(n_332), .Y(n_447) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g416 ( .A(n_333), .B(n_382), .Y(n_416) );
OR2x2_ASAP7_75t_L g334 ( .A(n_335), .B(n_337), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g347 ( .A(n_336), .B(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g418 ( .A(n_338), .Y(n_418) );
OR2x2_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
INVx1_ASAP7_75t_L g415 ( .A(n_339), .Y(n_415) );
INVx1_ASAP7_75t_L g421 ( .A(n_340), .Y(n_421) );
OR2x2_ASAP7_75t_L g444 ( .A(n_340), .B(n_445), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_342), .B(n_344), .Y(n_341) );
INVx1_ASAP7_75t_SL g353 ( .A(n_343), .Y(n_353) );
AND2x2_ASAP7_75t_L g423 ( .A(n_343), .B(n_403), .Y(n_423) );
AND2x2_ASAP7_75t_SL g455 ( .A(n_343), .B(n_356), .Y(n_455) );
INVx1_ASAP7_75t_SL g344 ( .A(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_346), .B(n_347), .Y(n_345) );
INVx1_ASAP7_75t_L g460 ( .A(n_346), .Y(n_460) );
INVx1_ASAP7_75t_L g410 ( .A(n_348), .Y(n_410) );
AND2x2_ASAP7_75t_L g349 ( .A(n_350), .B(n_351), .Y(n_349) );
O2A1O1Ixp33_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_354), .B(n_355), .C(n_359), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_353), .B(n_403), .Y(n_427) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_356), .B(n_407), .Y(n_406) );
AND2x2_ASAP7_75t_L g356 ( .A(n_357), .B(n_358), .Y(n_356) );
AND2x2_ASAP7_75t_L g364 ( .A(n_358), .B(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g445 ( .A(n_358), .Y(n_445) );
NAND4xp75_ASAP7_75t_L g360 ( .A(n_361), .B(n_417), .C(n_433), .D(n_454), .Y(n_360) );
NOR3x1_ASAP7_75t_L g361 ( .A(n_362), .B(n_379), .C(n_401), .Y(n_361) );
NAND4xp75_ASAP7_75t_L g362 ( .A(n_363), .B(n_369), .C(n_372), .D(n_375), .Y(n_362) );
NAND2xp5_ASAP7_75t_SL g363 ( .A(n_364), .B(n_366), .Y(n_363) );
AND2x2_ASAP7_75t_L g414 ( .A(n_365), .B(n_415), .Y(n_414) );
INVx1_ASAP7_75t_SL g439 ( .A(n_366), .Y(n_439) );
NAND2xp5_ASAP7_75t_SL g369 ( .A(n_370), .B(n_371), .Y(n_369) );
INVx1_ASAP7_75t_SL g428 ( .A(n_371), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_376), .B(n_377), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_380), .B(n_387), .Y(n_379) );
INVx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_383), .B(n_447), .Y(n_446) );
INVx1_ASAP7_75t_SL g385 ( .A(n_386), .Y(n_385) );
AOI21xp5_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_393), .B(n_397), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
OAI322xp33_ASAP7_75t_L g419 ( .A1(n_391), .A2(n_420), .A3(n_424), .B1(n_425), .B2(n_427), .C1(n_428), .C2(n_429), .Y(n_419) );
INVx2_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_392), .B(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_395), .B(n_396), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_395), .B(n_442), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_396), .B(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_399), .B(n_400), .Y(n_398) );
OAI211xp5_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_404), .B(n_406), .C(n_408), .Y(n_401) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
AOI22xp5_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_413), .B1(n_414), .B2(n_416), .Y(n_408) );
NOR2xp33_ASAP7_75t_SL g409 ( .A(n_410), .B(n_411), .Y(n_409) );
INVx2_ASAP7_75t_SL g411 ( .A(n_412), .Y(n_411) );
AOI21xp5_ASAP7_75t_L g420 ( .A1(n_421), .A2(n_422), .B(n_423), .Y(n_420) );
INVxp67_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
NOR2xp33_ASAP7_75t_L g458 ( .A(n_426), .B(n_459), .Y(n_458) );
NAND2xp5_ASAP7_75t_SL g429 ( .A(n_430), .B(n_432), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
OR2x2_ASAP7_75t_L g436 ( .A(n_431), .B(n_437), .Y(n_436) );
O2A1O1Ixp5_ASAP7_75t_L g433 ( .A1(n_434), .A2(n_435), .B(n_440), .C(n_443), .Y(n_433) );
NAND2xp5_ASAP7_75t_SL g435 ( .A(n_436), .B(n_439), .Y(n_435) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
OAI221xp5_ASAP7_75t_SL g443 ( .A1(n_444), .A2(n_446), .B1(n_448), .B2(n_450), .C(n_452), .Y(n_443) );
INVxp67_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
AND2x2_ASAP7_75t_L g459 ( .A(n_460), .B(n_461), .Y(n_459) );
HB1xp67_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
CKINVDCx20_ASAP7_75t_R g466 ( .A(n_467), .Y(n_466) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_467), .A2(n_483), .B1(n_497), .B2(n_498), .Y(n_496) );
AOI22xp5_ASAP7_75t_L g467 ( .A1(n_468), .A2(n_469), .B1(n_473), .B2(n_474), .Y(n_467) );
CKINVDCx20_ASAP7_75t_R g468 ( .A(n_469), .Y(n_468) );
CKINVDCx16_ASAP7_75t_R g472 ( .A(n_470), .Y(n_472) );
CKINVDCx20_ASAP7_75t_R g473 ( .A(n_474), .Y(n_473) );
OAI22xp5_ASAP7_75t_SL g474 ( .A1(n_475), .A2(n_476), .B1(n_479), .B2(n_480), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g480 ( .A(n_479), .Y(n_480) );
CKINVDCx20_ASAP7_75t_R g481 ( .A(n_482), .Y(n_481) );
CKINVDCx20_ASAP7_75t_R g482 ( .A(n_483), .Y(n_482) );
INVxp67_ASAP7_75t_L g495 ( .A(n_484), .Y(n_495) );
CKINVDCx8_ASAP7_75t_R g485 ( .A(n_486), .Y(n_485) );
NOR2xp33_ASAP7_75t_L g487 ( .A(n_488), .B(n_489), .Y(n_487) );
CKINVDCx16_ASAP7_75t_R g493 ( .A(n_490), .Y(n_493) );
AO21x1_ASAP7_75t_SL g501 ( .A1(n_490), .A2(n_502), .B(n_506), .Y(n_501) );
CKINVDCx20_ASAP7_75t_R g491 ( .A(n_492), .Y(n_491) );
CKINVDCx20_ASAP7_75t_R g498 ( .A(n_492), .Y(n_498) );
OR2x2_ASAP7_75t_L g492 ( .A(n_493), .B(n_494), .Y(n_492) );
CKINVDCx20_ASAP7_75t_R g499 ( .A(n_500), .Y(n_499) );
CKINVDCx20_ASAP7_75t_R g500 ( .A(n_501), .Y(n_500) );
HB1xp67_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx3_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
HB1xp67_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
endmodule