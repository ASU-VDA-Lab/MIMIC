module fake_jpeg_23320_n_342 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_342);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_342;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx4f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_3),
.B(n_14),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx11_ASAP7_75t_SL g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_36),
.A2(n_42),
.B1(n_48),
.B2(n_18),
.Y(n_50)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVxp67_ASAP7_75t_SL g60 ( 
.A(n_37),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_45),
.Y(n_53)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_24),
.B(n_0),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_44),
.B(n_22),
.Y(n_57)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx6_ASAP7_75t_SL g49 ( 
.A(n_40),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_49),
.B(n_51),
.Y(n_86)
);

INVxp67_ASAP7_75t_SL g94 ( 
.A(n_50),
.Y(n_94)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_36),
.A2(n_18),
.B1(n_23),
.B2(n_33),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_52),
.A2(n_64),
.B1(n_69),
.B2(n_73),
.Y(n_87)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_35),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_57),
.B(n_70),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_42),
.A2(n_23),
.B1(n_32),
.B2(n_21),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_58),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_113)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_42),
.A2(n_17),
.B1(n_34),
.B2(n_32),
.Y(n_64)
);

A2O1A1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_38),
.A2(n_26),
.B(n_28),
.C(n_34),
.Y(n_65)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

NAND2xp33_ASAP7_75t_SL g67 ( 
.A(n_40),
.B(n_26),
.Y(n_67)
);

AOI32xp33_ASAP7_75t_L g78 ( 
.A1(n_67),
.A2(n_43),
.A3(n_26),
.B1(n_35),
.B2(n_16),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_37),
.B(n_28),
.Y(n_68)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_68),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_48),
.A2(n_17),
.B1(n_34),
.B2(n_21),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_45),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_47),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_71),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_41),
.B(n_22),
.Y(n_72)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_72),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_48),
.A2(n_32),
.B1(n_21),
.B2(n_19),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_38),
.A2(n_32),
.B1(n_19),
.B2(n_16),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_74),
.A2(n_30),
.B1(n_35),
.B2(n_29),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_39),
.A2(n_32),
.B1(n_20),
.B2(n_31),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_75),
.A2(n_31),
.B1(n_30),
.B2(n_24),
.Y(n_82)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_76),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_43),
.B(n_20),
.Y(n_77)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_77),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_78),
.B(n_58),
.Y(n_119)
);

OA22x2_ASAP7_75t_L g79 ( 
.A1(n_60),
.A2(n_47),
.B1(n_26),
.B2(n_29),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_79),
.A2(n_83),
.B1(n_76),
.B2(n_63),
.Y(n_136)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_80),
.Y(n_117)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_81),
.B(n_84),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_82),
.A2(n_102),
.B(n_59),
.Y(n_132)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_51),
.A2(n_29),
.B1(n_27),
.B2(n_26),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_88),
.A2(n_113),
.B1(n_74),
.B2(n_76),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_57),
.B(n_0),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_89),
.B(n_96),
.Y(n_130)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_93),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_72),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_95),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_68),
.B(n_0),
.Y(n_96)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_70),
.Y(n_97)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_67),
.B(n_0),
.Y(n_99)
);

OAI21xp33_ASAP7_75t_L g116 ( 
.A1(n_99),
.A2(n_15),
.B(n_10),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_53),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_100),
.B(n_108),
.Y(n_134)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_55),
.Y(n_101)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_101),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_62),
.A2(n_9),
.B1(n_14),
.B2(n_13),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_55),
.Y(n_103)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_103),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_65),
.A2(n_9),
.B1(n_14),
.B2(n_13),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_104),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_49),
.Y(n_106)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_106),
.Y(n_121)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_77),
.Y(n_108)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_63),
.Y(n_109)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_109),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_L g110 ( 
.A1(n_65),
.A2(n_8),
.B1(n_13),
.B2(n_12),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_110),
.A2(n_59),
.B1(n_63),
.B2(n_61),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g112 ( 
.A(n_62),
.Y(n_112)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_112),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_62),
.A2(n_7),
.B1(n_11),
.B2(n_10),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_114),
.Y(n_126)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_53),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g120 ( 
.A(n_115),
.Y(n_120)
);

OR2x2_ASAP7_75t_SL g162 ( 
.A(n_116),
.B(n_108),
.Y(n_162)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_106),
.Y(n_118)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_118),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_119),
.B(n_87),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_80),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_127),
.B(n_129),
.Y(n_146)
);

OR2x2_ASAP7_75t_L g128 ( 
.A(n_86),
.B(n_73),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_128),
.B(n_133),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_132),
.A2(n_83),
.B(n_79),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_91),
.B(n_66),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_136),
.A2(n_81),
.B1(n_111),
.B2(n_109),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_113),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_137),
.B(n_142),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_91),
.B(n_56),
.C(n_61),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_139),
.B(n_90),
.C(n_105),
.Y(n_179)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_93),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_97),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_143),
.B(n_79),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_114),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_144),
.B(n_145),
.Y(n_163)
);

A2O1A1O1Ixp25_ASAP7_75t_L g147 ( 
.A1(n_119),
.A2(n_99),
.B(n_94),
.C(n_104),
.D(n_110),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_147),
.B(n_179),
.C(n_142),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_138),
.B(n_85),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_148),
.B(n_152),
.Y(n_186)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_118),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_149),
.B(n_158),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_150),
.A2(n_172),
.B1(n_174),
.B2(n_178),
.Y(n_184)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_135),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_133),
.A2(n_99),
.B(n_98),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_153),
.A2(n_141),
.B(n_140),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_139),
.B(n_96),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_154),
.A2(n_175),
.B(n_79),
.Y(n_207)
);

FAx1_ASAP7_75t_SL g156 ( 
.A(n_130),
.B(n_89),
.CI(n_98),
.CON(n_156),
.SN(n_156)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_156),
.B(n_160),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_157),
.B(n_130),
.Y(n_182)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_118),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_134),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_159),
.B(n_161),
.Y(n_189)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_135),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_134),
.Y(n_161)
);

OAI21xp33_ASAP7_75t_L g197 ( 
.A1(n_162),
.A2(n_105),
.B(n_123),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_132),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_164),
.B(n_168),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_121),
.B(n_92),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g188 ( 
.A(n_165),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_124),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_166),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_138),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_167),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_145),
.Y(n_168)
);

INVx4_ASAP7_75t_SL g169 ( 
.A(n_140),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_169),
.B(n_171),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_117),
.B(n_107),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_170),
.B(n_177),
.Y(n_183)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_121),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_137),
.A2(n_111),
.B1(n_101),
.B2(n_84),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_120),
.A2(n_59),
.B1(n_107),
.B2(n_90),
.Y(n_174)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_121),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_176),
.Y(n_190)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_136),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_125),
.A2(n_126),
.B1(n_117),
.B2(n_129),
.Y(n_178)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_180),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_182),
.B(n_207),
.Y(n_217)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_170),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_187),
.B(n_191),
.Y(n_227)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_155),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_151),
.B(n_128),
.Y(n_192)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_192),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_151),
.B(n_128),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_193),
.B(n_196),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_146),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_194),
.B(n_195),
.Y(n_229)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_150),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_178),
.B(n_179),
.Y(n_196)
);

OA22x2_ASAP7_75t_L g218 ( 
.A1(n_197),
.A2(n_206),
.B1(n_162),
.B2(n_154),
.Y(n_218)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_169),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_200),
.B(n_201),
.Y(n_226)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_163),
.Y(n_201)
);

INVx13_ASAP7_75t_L g202 ( 
.A(n_158),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_202),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_204),
.B(n_209),
.C(n_191),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_166),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_205),
.Y(n_233)
);

AND2x6_ASAP7_75t_L g206 ( 
.A(n_157),
.B(n_122),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_153),
.B(n_154),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_208),
.B(n_175),
.Y(n_221)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_152),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_210),
.B(n_159),
.Y(n_225)
);

BUFx2_ASAP7_75t_L g212 ( 
.A(n_149),
.Y(n_212)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_212),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_164),
.A2(n_122),
.B1(n_123),
.B2(n_143),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_213),
.A2(n_194),
.B1(n_201),
.B2(n_199),
.Y(n_234)
);

OAI32xp33_ASAP7_75t_L g238 ( 
.A1(n_214),
.A2(n_141),
.A3(n_131),
.B1(n_173),
.B2(n_124),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_211),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_215),
.B(n_205),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_188),
.B(n_161),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_216),
.B(n_223),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_218),
.A2(n_238),
.B(n_189),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_221),
.B(n_2),
.Y(n_266)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_203),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_185),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_224),
.B(n_200),
.Y(n_256)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_225),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_195),
.A2(n_168),
.B1(n_177),
.B2(n_147),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_228),
.A2(n_237),
.B1(n_240),
.B2(n_210),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_182),
.B(n_156),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_230),
.B(n_232),
.C(n_239),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_187),
.B(n_160),
.Y(n_231)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_231),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_208),
.B(n_156),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_234),
.A2(n_207),
.B(n_213),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_183),
.B(n_171),
.Y(n_235)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_235),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_184),
.A2(n_183),
.B1(n_192),
.B2(n_181),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_181),
.A2(n_131),
.B1(n_66),
.B2(n_54),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_204),
.B(n_66),
.C(n_54),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_241),
.B(n_212),
.C(n_54),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_193),
.B(n_214),
.Y(n_242)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_242),
.Y(n_261)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_243),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_233),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_244),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_246),
.B(n_252),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_247),
.A2(n_249),
.B1(n_258),
.B2(n_259),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_242),
.A2(n_220),
.B(n_222),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_248),
.B(n_254),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_234),
.A2(n_206),
.B1(n_196),
.B2(n_193),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_217),
.B(n_221),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_226),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_255),
.B(n_236),
.Y(n_270)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_256),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_220),
.A2(n_196),
.B1(n_190),
.B2(n_202),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_235),
.A2(n_190),
.B1(n_186),
.B2(n_198),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_260),
.B(n_224),
.C(n_240),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_237),
.A2(n_228),
.B1(n_229),
.B2(n_227),
.Y(n_262)
);

CKINVDCx14_ASAP7_75t_R g278 ( 
.A(n_262),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_222),
.A2(n_1),
.B(n_2),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_263),
.B(n_265),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_218),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_264)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_264),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_231),
.A2(n_8),
.B(n_10),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_266),
.B(n_241),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_250),
.B(n_217),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_269),
.B(n_275),
.Y(n_291)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_270),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_250),
.B(n_230),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_276),
.B(n_279),
.C(n_258),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_252),
.B(n_232),
.C(n_239),
.Y(n_279)
);

A2O1A1Ixp33_ASAP7_75t_L g280 ( 
.A1(n_249),
.A2(n_218),
.B(n_225),
.C(n_238),
.Y(n_280)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_280),
.Y(n_298)
);

XOR2x2_ASAP7_75t_L g282 ( 
.A(n_248),
.B(n_218),
.Y(n_282)
);

XNOR2x1_ASAP7_75t_L g302 ( 
.A(n_282),
.B(n_268),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_283),
.B(n_286),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_255),
.B(n_215),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_284),
.B(n_285),
.Y(n_301)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_256),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_266),
.B(n_219),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_287),
.B(n_293),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_279),
.C(n_283),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_288),
.B(n_289),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_275),
.B(n_246),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_276),
.B(n_251),
.C(n_257),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_290),
.B(n_292),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_267),
.B(n_251),
.C(n_257),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_267),
.B(n_261),
.C(n_245),
.Y(n_293)
);

NOR2x1_ASAP7_75t_SL g294 ( 
.A(n_282),
.B(n_259),
.Y(n_294)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_294),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_274),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_296),
.B(n_271),
.Y(n_304)
);

FAx1_ASAP7_75t_SL g297 ( 
.A(n_286),
.B(n_254),
.CI(n_264),
.CON(n_297),
.SN(n_297)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_297),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_278),
.A2(n_247),
.B1(n_263),
.B2(n_253),
.Y(n_299)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_299),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_302),
.A2(n_270),
.B(n_273),
.Y(n_311)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_304),
.Y(n_316)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_301),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_308),
.B(n_312),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_298),
.A2(n_280),
.B1(n_272),
.B2(n_281),
.Y(n_310)
);

O2A1O1Ixp33_ASAP7_75t_L g322 ( 
.A1(n_310),
.A2(n_314),
.B(n_300),
.C(n_291),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_311),
.B(n_5),
.Y(n_325)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_290),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_295),
.B(n_273),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_302),
.A2(n_260),
.B1(n_265),
.B2(n_269),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_315),
.B(n_287),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_318),
.A2(n_305),
.B1(n_306),
.B2(n_309),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_304),
.B(n_297),
.Y(n_319)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_319),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_303),
.A2(n_292),
.B1(n_293),
.B2(n_288),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_320),
.B(n_321),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_308),
.B(n_300),
.Y(n_321)
);

OAI21x1_ASAP7_75t_SL g330 ( 
.A1(n_322),
.A2(n_311),
.B(n_310),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_307),
.A2(n_291),
.B1(n_5),
.B2(n_4),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_323),
.B(n_324),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_313),
.B(n_15),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_325),
.B(n_5),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_316),
.B(n_309),
.C(n_314),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_327),
.A2(n_317),
.B(n_325),
.Y(n_334)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_328),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_330),
.A2(n_332),
.B(n_323),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_334),
.Y(n_338)
);

INVxp67_ASAP7_75t_SL g337 ( 
.A(n_335),
.Y(n_337)
);

AOI21xp33_ASAP7_75t_L g336 ( 
.A1(n_326),
.A2(n_320),
.B(n_322),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_338),
.A2(n_336),
.B(n_333),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_339),
.A2(n_337),
.B(n_327),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_329),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_341),
.A2(n_331),
.B(n_332),
.Y(n_342)
);


endmodule