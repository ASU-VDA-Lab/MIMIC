module real_aes_4213_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_357;
wire n_635;
wire n_287;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_580;
wire n_577;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_549;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_560;
wire n_260;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_453;
wire n_374;
wire n_379;
wire n_235;
wire n_399;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_570;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_547;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_250;
wire n_85;
wire n_605;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_171;
wire n_87;
wire n_78;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_557;
wire n_501;
wire n_488;
wire n_251;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_546;
wire n_151;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_601;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
INVx1_ASAP7_75t_L g245 ( .A(n_0), .Y(n_245) );
AOI22xp5_ASAP7_75t_L g221 ( .A1(n_1), .A2(n_12), .B1(n_84), .B2(n_198), .Y(n_221) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_2), .A2(n_60), .B1(n_585), .B2(n_586), .Y(n_584) );
INVx2_ASAP7_75t_L g178 ( .A(n_3), .Y(n_178) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_4), .A2(n_73), .B1(n_510), .B2(n_531), .Y(n_509) );
INVx1_ASAP7_75t_SL g118 ( .A(n_5), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_6), .B(n_236), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_7), .B(n_255), .Y(n_254) );
INVx1_ASAP7_75t_L g528 ( .A(n_8), .Y(n_528) );
INVxp67_ASAP7_75t_L g538 ( .A(n_8), .Y(n_538) );
NOR2xp33_ASAP7_75t_L g565 ( .A(n_8), .B(n_52), .Y(n_565) );
AOI22xp33_ASAP7_75t_L g249 ( .A1(n_9), .A2(n_38), .B1(n_250), .B2(n_251), .Y(n_249) );
OA21x2_ASAP7_75t_L g111 ( .A1(n_10), .A2(n_50), .B(n_112), .Y(n_111) );
OA21x2_ASAP7_75t_L g132 ( .A1(n_10), .A2(n_50), .B(n_112), .Y(n_132) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_11), .B(n_514), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_13), .B(n_156), .Y(n_209) );
HB1xp67_ASAP7_75t_L g625 ( .A(n_13), .Y(n_625) );
AOI22xp5_ASAP7_75t_L g170 ( .A1(n_14), .A2(n_57), .B1(n_171), .B2(n_172), .Y(n_170) );
INVx2_ASAP7_75t_L g202 ( .A(n_15), .Y(n_202) );
OAI22xp5_ASAP7_75t_L g620 ( .A1(n_16), .A2(n_506), .B1(n_507), .B2(n_621), .Y(n_620) );
CKINVDCx5p33_ASAP7_75t_R g621 ( .A(n_16), .Y(n_621) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_17), .A2(n_35), .B1(n_541), .B2(n_546), .Y(n_540) );
INVx1_ASAP7_75t_SL g601 ( .A(n_18), .Y(n_601) );
AOI22xp5_ASAP7_75t_L g222 ( .A1(n_19), .A2(n_23), .B1(n_116), .B2(n_153), .Y(n_222) );
BUFx3_ASAP7_75t_L g608 ( .A(n_20), .Y(n_608) );
O2A1O1Ixp5_ASAP7_75t_L g195 ( .A1(n_21), .A2(n_89), .B(n_196), .C(n_197), .Y(n_195) );
AOI22xp33_ASAP7_75t_L g174 ( .A1(n_22), .A2(n_45), .B1(n_175), .B2(n_176), .Y(n_174) );
CKINVDCx5p33_ASAP7_75t_R g597 ( .A(n_23), .Y(n_597) );
CKINVDCx5p33_ASAP7_75t_R g154 ( .A(n_24), .Y(n_154) );
BUFx6f_ASAP7_75t_L g514 ( .A(n_25), .Y(n_514) );
AOI22xp5_ASAP7_75t_L g257 ( .A1(n_26), .A2(n_59), .B1(n_258), .B2(n_260), .Y(n_257) );
INVx1_ASAP7_75t_L g191 ( .A(n_27), .Y(n_191) );
INVx1_ASAP7_75t_L g515 ( .A(n_28), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_28), .B(n_51), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_29), .B(n_187), .Y(n_240) );
INVx2_ASAP7_75t_L g199 ( .A(n_30), .Y(n_199) );
CKINVDCx5p33_ASAP7_75t_R g157 ( .A(n_31), .Y(n_157) );
INVx2_ASAP7_75t_L g208 ( .A(n_32), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_33), .B(n_238), .Y(n_237) );
INVx1_ASAP7_75t_SL g125 ( .A(n_34), .Y(n_125) );
INVx1_ASAP7_75t_L g149 ( .A(n_36), .Y(n_149) );
INVx1_ASAP7_75t_L g112 ( .A(n_37), .Y(n_112) );
AND2x4_ASAP7_75t_L g92 ( .A(n_39), .B(n_93), .Y(n_92) );
AND2x4_ASAP7_75t_L g143 ( .A(n_39), .B(n_93), .Y(n_143) );
HB1xp67_ASAP7_75t_L g618 ( .A(n_39), .Y(n_618) );
INVx1_ASAP7_75t_L g133 ( .A(n_40), .Y(n_133) );
BUFx6f_ASAP7_75t_L g90 ( .A(n_41), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g505 ( .A(n_42), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_43), .A2(n_46), .B1(n_580), .B2(n_583), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_44), .A2(n_68), .B1(n_571), .B2(n_577), .Y(n_570) );
NOR2xp33_ASAP7_75t_L g212 ( .A(n_47), .B(n_120), .Y(n_212) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_48), .A2(n_62), .B1(n_558), .B2(n_559), .Y(n_557) );
OA22x2_ASAP7_75t_L g519 ( .A1(n_49), .A2(n_52), .B1(n_514), .B2(n_518), .Y(n_519) );
INVx1_ASAP7_75t_L g551 ( .A(n_49), .Y(n_551) );
INVx1_ASAP7_75t_L g530 ( .A(n_51), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_51), .B(n_549), .Y(n_568) );
HB1xp67_ASAP7_75t_L g611 ( .A(n_51), .Y(n_611) );
OAI21xp33_ASAP7_75t_L g552 ( .A1(n_52), .A2(n_58), .B(n_539), .Y(n_552) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_53), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g189 ( .A(n_54), .Y(n_189) );
NAND2xp5_ASAP7_75t_SL g553 ( .A(n_55), .B(n_554), .Y(n_553) );
NOR2xp33_ASAP7_75t_L g128 ( .A(n_56), .B(n_117), .Y(n_128) );
INVx1_ASAP7_75t_L g517 ( .A(n_58), .Y(n_517) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_58), .B(n_74), .Y(n_566) );
BUFx6f_ASAP7_75t_L g85 ( .A(n_61), .Y(n_85) );
INVx1_ASAP7_75t_L g122 ( .A(n_61), .Y(n_122) );
BUFx5_ASAP7_75t_L g127 ( .A(n_61), .Y(n_127) );
HB1xp67_ASAP7_75t_L g593 ( .A(n_63), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_64), .A2(n_75), .B1(n_588), .B2(n_589), .Y(n_587) );
NOR2xp33_ASAP7_75t_L g119 ( .A(n_65), .B(n_120), .Y(n_119) );
INVx2_ASAP7_75t_L g211 ( .A(n_66), .Y(n_211) );
HB1xp67_ASAP7_75t_L g600 ( .A(n_67), .Y(n_600) );
INVx1_ASAP7_75t_L g215 ( .A(n_69), .Y(n_215) );
INVx2_ASAP7_75t_L g161 ( .A(n_70), .Y(n_161) );
INVx2_ASAP7_75t_SL g93 ( .A(n_71), .Y(n_93) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_72), .B(n_232), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_74), .B(n_523), .Y(n_522) );
AO32x2_ASAP7_75t_L g219 ( .A1(n_76), .A2(n_91), .A3(n_200), .B1(n_220), .B2(n_224), .Y(n_219) );
AO22x2_ASAP7_75t_L g313 ( .A1(n_76), .A2(n_220), .B1(n_314), .B2(n_316), .Y(n_313) );
AOI21xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_94), .B(n_501), .Y(n_77) );
BUFx4f_ASAP7_75t_SL g78 ( .A(n_79), .Y(n_78) );
AND2x2_ASAP7_75t_L g79 ( .A(n_80), .B(n_91), .Y(n_79) );
OA21x2_ASAP7_75t_L g628 ( .A1(n_80), .A2(n_629), .B(n_630), .Y(n_628) );
NOR2xp33_ASAP7_75t_L g80 ( .A(n_81), .B(n_86), .Y(n_80) );
CKINVDCx16_ASAP7_75t_R g81 ( .A(n_82), .Y(n_81) );
HB1xp67_ASAP7_75t_L g82 ( .A(n_83), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_84), .Y(n_83) );
INVx2_ASAP7_75t_L g193 ( .A(n_84), .Y(n_193) );
INVxp67_ASAP7_75t_SL g260 ( .A(n_84), .Y(n_260) );
INVx2_ASAP7_75t_L g84 ( .A(n_85), .Y(n_84) );
INVx3_ASAP7_75t_L g117 ( .A(n_85), .Y(n_117) );
INVx2_ASAP7_75t_L g147 ( .A(n_85), .Y(n_147) );
INVx6_ASAP7_75t_L g156 ( .A(n_85), .Y(n_156) );
CKINVDCx20_ASAP7_75t_R g86 ( .A(n_87), .Y(n_86) );
HB1xp67_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
NOR2xp33_ASAP7_75t_L g151 ( .A(n_88), .B(n_142), .Y(n_151) );
INVx4_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
OAI22xp5_ASAP7_75t_L g220 ( .A1(n_89), .A2(n_221), .B1(n_222), .B2(n_223), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_89), .A2(n_235), .B(n_237), .Y(n_234) );
BUFx6f_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
BUFx6f_ASAP7_75t_L g123 ( .A(n_90), .Y(n_123) );
INVx3_ASAP7_75t_L g129 ( .A(n_90), .Y(n_129) );
INVx4_ASAP7_75t_L g188 ( .A(n_90), .Y(n_188) );
INVx1_ASAP7_75t_L g262 ( .A(n_90), .Y(n_262) );
BUFx6f_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
INVx3_ASAP7_75t_L g113 ( .A(n_92), .Y(n_113) );
AND2x2_ASAP7_75t_L g167 ( .A(n_92), .B(n_168), .Y(n_167) );
AND2x2_ASAP7_75t_L g314 ( .A(n_92), .B(n_315), .Y(n_314) );
HB1xp67_ASAP7_75t_L g616 ( .A(n_93), .Y(n_616) );
INVx2_ASAP7_75t_L g94 ( .A(n_95), .Y(n_94) );
BUFx2_ASAP7_75t_L g95 ( .A(n_96), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_97), .Y(n_96) );
INVx2_ASAP7_75t_L g97 ( .A(n_98), .Y(n_97) );
INVx2_ASAP7_75t_SL g98 ( .A(n_99), .Y(n_98) );
NAND2x1p5_ASAP7_75t_L g99 ( .A(n_100), .B(n_386), .Y(n_99) );
AND3x1_ASAP7_75t_L g100 ( .A(n_101), .B(n_342), .C(n_370), .Y(n_100) );
NOR3xp33_ASAP7_75t_SL g101 ( .A(n_102), .B(n_279), .C(n_318), .Y(n_101) );
NAND2xp5_ASAP7_75t_L g102 ( .A(n_103), .B(n_263), .Y(n_102) );
A2O1A1Ixp33_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_163), .B(n_216), .C(n_228), .Y(n_103) );
HB1xp67_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
AND2x2_ASAP7_75t_L g306 ( .A(n_105), .B(n_307), .Y(n_306) );
AND2x4_ASAP7_75t_L g320 ( .A(n_105), .B(n_321), .Y(n_320) );
NAND2x1p5_ASAP7_75t_L g452 ( .A(n_105), .B(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g462 ( .A(n_105), .Y(n_462) );
AND2x2_ASAP7_75t_L g105 ( .A(n_106), .B(n_134), .Y(n_105) );
INVxp67_ASAP7_75t_SL g273 ( .A(n_106), .Y(n_273) );
OR2x2_ASAP7_75t_L g346 ( .A(n_106), .B(n_347), .Y(n_346) );
INVx2_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx2_ASAP7_75t_L g268 ( .A(n_107), .Y(n_268) );
AND2x2_ASAP7_75t_L g281 ( .A(n_107), .B(n_275), .Y(n_281) );
OR2x2_ASAP7_75t_L g289 ( .A(n_107), .B(n_134), .Y(n_289) );
HB1xp67_ASAP7_75t_L g293 ( .A(n_107), .Y(n_293) );
INVx1_ASAP7_75t_L g333 ( .A(n_107), .Y(n_333) );
INVx1_ASAP7_75t_L g403 ( .A(n_107), .Y(n_403) );
AO31x2_ASAP7_75t_L g107 ( .A1(n_108), .A2(n_114), .A3(n_124), .B(n_130), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g108 ( .A(n_109), .B(n_113), .Y(n_108) );
INVx2_ASAP7_75t_L g168 ( .A(n_109), .Y(n_168) );
INVx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
INVx4_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
BUFx3_ASAP7_75t_L g159 ( .A(n_111), .Y(n_159) );
INVx2_ASAP7_75t_L g179 ( .A(n_111), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_113), .B(n_132), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_113), .B(n_132), .Y(n_246) );
NOR2xp67_ASAP7_75t_L g253 ( .A(n_113), .B(n_132), .Y(n_253) );
A2O1A1Ixp33_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_118), .B(n_119), .C(n_123), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx2_ASAP7_75t_L g172 ( .A(n_117), .Y(n_172) );
INVx1_ASAP7_75t_L g236 ( .A(n_117), .Y(n_236) );
INVx1_ASAP7_75t_L g251 ( .A(n_117), .Y(n_251) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx2_ASAP7_75t_L g175 ( .A(n_121), .Y(n_175) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx2_ASAP7_75t_L g140 ( .A(n_122), .Y(n_140) );
INVx1_ASAP7_75t_L g173 ( .A(n_123), .Y(n_173) );
A2O1A1Ixp33_ASAP7_75t_L g210 ( .A1(n_123), .A2(n_139), .B(n_211), .C(n_212), .Y(n_210) );
INVx1_ASAP7_75t_L g223 ( .A(n_123), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g252 ( .A(n_123), .B(n_253), .Y(n_252) );
A2O1A1Ixp33_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_126), .B(n_128), .C(n_129), .Y(n_124) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx2_ASAP7_75t_L g153 ( .A(n_127), .Y(n_153) );
INVx2_ASAP7_75t_L g238 ( .A(n_127), .Y(n_238) );
INVx1_ASAP7_75t_L g242 ( .A(n_127), .Y(n_242) );
INVx2_ASAP7_75t_L g250 ( .A(n_127), .Y(n_250) );
INVx3_ASAP7_75t_L g144 ( .A(n_129), .Y(n_144) );
A2O1A1Ixp33_ASAP7_75t_L g206 ( .A1(n_129), .A2(n_207), .B(n_208), .C(n_209), .Y(n_206) );
NOR2xp33_ASAP7_75t_SL g130 ( .A(n_131), .B(n_133), .Y(n_130) );
NOR2xp33_ASAP7_75t_L g214 ( .A(n_131), .B(n_215), .Y(n_214) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx1_ASAP7_75t_L g162 ( .A(n_132), .Y(n_162) );
BUFx3_ASAP7_75t_L g255 ( .A(n_132), .Y(n_255) );
INVx1_ASAP7_75t_L g315 ( .A(n_132), .Y(n_315) );
INVx2_ASAP7_75t_L g266 ( .A(n_134), .Y(n_266) );
BUFx2_ASAP7_75t_L g448 ( .A(n_134), .Y(n_448) );
AO21x2_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_158), .B(n_160), .Y(n_134) );
AO21x2_ASAP7_75t_L g275 ( .A1(n_135), .A2(n_160), .B(n_276), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_136), .B(n_150), .Y(n_135) );
AOI22xp5_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_141), .B1(n_145), .B2(n_148), .Y(n_136) );
NOR2xp67_ASAP7_75t_L g137 ( .A(n_138), .B(n_139), .Y(n_137) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx2_ASAP7_75t_L g171 ( .A(n_140), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g141 ( .A(n_142), .B(n_144), .Y(n_141) );
NOR3xp33_ASAP7_75t_L g148 ( .A(n_142), .B(n_144), .C(n_149), .Y(n_148) );
AOI221x1_ASAP7_75t_L g182 ( .A1(n_142), .A2(n_183), .B1(n_186), .B2(n_190), .C(n_192), .Y(n_182) );
INVx4_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
OAI22xp5_ASAP7_75t_L g169 ( .A1(n_144), .A2(n_170), .B1(n_173), .B2(n_174), .Y(n_169) );
INVx1_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g259 ( .A(n_147), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_151), .B(n_152), .Y(n_150) );
OAI22xp33_ASAP7_75t_L g152 ( .A1(n_153), .A2(n_154), .B1(n_155), .B2(n_157), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_155), .B(n_244), .Y(n_243) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx1_ASAP7_75t_L g176 ( .A(n_156), .Y(n_176) );
INVx2_ASAP7_75t_L g185 ( .A(n_156), .Y(n_185) );
INVx2_ASAP7_75t_SL g198 ( .A(n_156), .Y(n_198) );
INVx3_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
NOR2xp33_ASAP7_75t_L g160 ( .A(n_161), .B(n_162), .Y(n_160) );
INVx1_ASAP7_75t_L g224 ( .A(n_162), .Y(n_224) );
AND2x2_ASAP7_75t_L g163 ( .A(n_164), .B(n_180), .Y(n_163) );
INVx2_ASAP7_75t_L g311 ( .A(n_164), .Y(n_311) );
NAND2xp5_ASAP7_75t_SL g327 ( .A(n_164), .B(n_180), .Y(n_327) );
INVx4_ASAP7_75t_L g355 ( .A(n_164), .Y(n_355) );
AND2x2_ASAP7_75t_L g495 ( .A(n_164), .B(n_340), .Y(n_495) );
BUFx3_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx1_ASAP7_75t_L g301 ( .A(n_165), .Y(n_301) );
INVx1_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx1_ASAP7_75t_L g227 ( .A(n_166), .Y(n_227) );
INVx1_ASAP7_75t_L g361 ( .A(n_166), .Y(n_361) );
AOI21x1_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_169), .B(n_177), .Y(n_166) );
INVx3_ASAP7_75t_L g196 ( .A(n_175), .Y(n_196) );
INVx1_ASAP7_75t_L g207 ( .A(n_176), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_178), .B(n_179), .Y(n_177) );
BUFx3_ASAP7_75t_L g200 ( .A(n_179), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g201 ( .A(n_179), .B(n_202), .Y(n_201) );
INVx3_ASAP7_75t_L g232 ( .A(n_179), .Y(n_232) );
AND2x2_ASAP7_75t_L g277 ( .A(n_180), .B(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g295 ( .A(n_180), .B(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g298 ( .A(n_180), .B(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g442 ( .A(n_180), .B(n_347), .Y(n_442) );
AND2x2_ASAP7_75t_L g180 ( .A(n_181), .B(n_203), .Y(n_180) );
INVx2_ASAP7_75t_L g226 ( .A(n_181), .Y(n_226) );
INVx1_ASAP7_75t_L g341 ( .A(n_181), .Y(n_341) );
AND2x2_ASAP7_75t_L g374 ( .A(n_181), .B(n_204), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_181), .B(n_361), .Y(n_422) );
OR2x2_ASAP7_75t_L g470 ( .A(n_181), .B(n_361), .Y(n_470) );
AO31x2_ASAP7_75t_L g181 ( .A1(n_182), .A2(n_194), .A3(n_200), .B(n_201), .Y(n_181) );
INVx1_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
AND2x2_ASAP7_75t_L g186 ( .A(n_187), .B(n_189), .Y(n_186) );
AND2x2_ASAP7_75t_L g190 ( .A(n_187), .B(n_191), .Y(n_190) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_188), .B(n_245), .Y(n_244) );
INVx1_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
INVx1_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_198), .B(n_199), .Y(n_197) );
INVx2_ASAP7_75t_L g316 ( .A(n_200), .Y(n_316) );
AND2x4_ASAP7_75t_L g351 ( .A(n_203), .B(n_313), .Y(n_351) );
AND2x2_ASAP7_75t_L g396 ( .A(n_203), .B(n_227), .Y(n_396) );
INVx2_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
AND2x4_ASAP7_75t_L g217 ( .A(n_204), .B(n_218), .Y(n_217) );
BUFx3_ASAP7_75t_L g317 ( .A(n_204), .Y(n_317) );
AND2x4_ASAP7_75t_L g340 ( .A(n_204), .B(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g367 ( .A(n_204), .Y(n_367) );
INVx3_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
AO31x2_ASAP7_75t_L g205 ( .A1(n_206), .A2(n_210), .A3(n_213), .B(n_214), .Y(n_205) );
AO22x1_ASAP7_75t_L g634 ( .A1(n_211), .A2(n_506), .B1(n_507), .B2(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_211), .Y(n_635) );
AND2x2_ASAP7_75t_L g216 ( .A(n_217), .B(n_225), .Y(n_216) );
INVx2_ASAP7_75t_L g385 ( .A(n_217), .Y(n_385) );
OAI21xp5_ASAP7_75t_L g404 ( .A1(n_217), .A2(n_405), .B(n_408), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_218), .B(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g356 ( .A(n_218), .B(n_357), .Y(n_356) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
BUFx8_ASAP7_75t_L g278 ( .A(n_219), .Y(n_278) );
AND2x2_ASAP7_75t_L g475 ( .A(n_219), .B(n_301), .Y(n_475) );
INVxp67_ASAP7_75t_L g276 ( .A(n_224), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_225), .B(n_351), .Y(n_437) );
AND2x2_ASAP7_75t_L g225 ( .A(n_226), .B(n_227), .Y(n_225) );
INVx2_ASAP7_75t_SL g357 ( .A(n_226), .Y(n_357) );
BUFx3_ASAP7_75t_L g395 ( .A(n_226), .Y(n_395) );
INVx1_ASAP7_75t_L g474 ( .A(n_226), .Y(n_474) );
HB1xp67_ASAP7_75t_L g321 ( .A(n_227), .Y(n_321) );
INVx2_ASAP7_75t_L g347 ( .A(n_227), .Y(n_347) );
INVx1_ASAP7_75t_L g358 ( .A(n_228), .Y(n_358) );
HB1xp67_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
AND2x2_ASAP7_75t_L g292 ( .A(n_229), .B(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g472 ( .A(n_229), .B(n_281), .Y(n_472) );
AND2x2_ASAP7_75t_L g229 ( .A(n_230), .B(n_247), .Y(n_229) );
INVx2_ASAP7_75t_L g270 ( .A(n_230), .Y(n_270) );
INVx1_ASAP7_75t_L g285 ( .A(n_230), .Y(n_285) );
HB1xp67_ASAP7_75t_L g291 ( .A(n_230), .Y(n_291) );
INVx1_ASAP7_75t_L g309 ( .A(n_230), .Y(n_309) );
AND2x2_ASAP7_75t_L g466 ( .A(n_230), .B(n_268), .Y(n_466) );
AND2x4_ASAP7_75t_L g230 ( .A(n_231), .B(n_233), .Y(n_230) );
OAI21xp5_ASAP7_75t_L g233 ( .A1(n_234), .A2(n_239), .B(n_246), .Y(n_233) );
OAI21xp5_ASAP7_75t_L g239 ( .A1(n_240), .A2(n_241), .B(n_243), .Y(n_239) );
INVx1_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
AND2x2_ASAP7_75t_L g269 ( .A(n_247), .B(n_270), .Y(n_269) );
INVx2_ASAP7_75t_L g304 ( .A(n_247), .Y(n_304) );
INVx1_ASAP7_75t_L g324 ( .A(n_247), .Y(n_324) );
INVx1_ASAP7_75t_L g380 ( .A(n_247), .Y(n_380) );
NAND2x1p5_ASAP7_75t_L g247 ( .A(n_248), .B(n_256), .Y(n_247) );
AND2x2_ASAP7_75t_SL g284 ( .A(n_248), .B(n_256), .Y(n_284) );
OA21x2_ASAP7_75t_L g248 ( .A1(n_249), .A2(n_252), .B(n_254), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_253), .B(n_262), .Y(n_261) );
OR2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_261), .Y(n_256) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
OAI21xp5_ASAP7_75t_L g263 ( .A1(n_264), .A2(n_271), .B(n_277), .Y(n_263) );
INVx2_ASAP7_75t_L g369 ( .A(n_264), .Y(n_369) );
AND2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_269), .Y(n_264) );
AND2x2_ASAP7_75t_L g302 ( .A(n_265), .B(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g400 ( .A(n_265), .B(n_401), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_265), .B(n_383), .Y(n_428) );
AND2x4_ASAP7_75t_L g436 ( .A(n_265), .B(n_308), .Y(n_436) );
AND2x4_ASAP7_75t_L g265 ( .A(n_266), .B(n_267), .Y(n_265) );
AND2x2_ASAP7_75t_L g493 ( .A(n_266), .B(n_304), .Y(n_493) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g426 ( .A(n_269), .B(n_281), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_269), .B(n_448), .Y(n_456) );
AND2x2_ASAP7_75t_L g477 ( .A(n_269), .B(n_478), .Y(n_477) );
OR2x2_ASAP7_75t_L g274 ( .A(n_270), .B(n_275), .Y(n_274) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
INVx2_ASAP7_75t_L g411 ( .A(n_272), .Y(n_411) );
OR2x6_ASAP7_75t_L g272 ( .A(n_273), .B(n_274), .Y(n_272) );
INVxp67_ASAP7_75t_SL g337 ( .A(n_274), .Y(n_337) );
INVxp67_ASAP7_75t_L g381 ( .A(n_274), .Y(n_381) );
AND2x2_ASAP7_75t_L g330 ( .A(n_275), .B(n_304), .Y(n_330) );
AND2x2_ASAP7_75t_L g350 ( .A(n_275), .B(n_309), .Y(n_350) );
AND2x2_ASAP7_75t_L g487 ( .A(n_275), .B(n_488), .Y(n_487) );
INVx2_ASAP7_75t_L g296 ( .A(n_278), .Y(n_296) );
INVx1_ASAP7_75t_L g326 ( .A(n_278), .Y(n_326) );
AND2x2_ASAP7_75t_SL g339 ( .A(n_278), .B(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g373 ( .A(n_278), .B(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g420 ( .A(n_278), .B(n_421), .Y(n_420) );
NAND4xp25_ASAP7_75t_L g431 ( .A(n_278), .B(n_349), .C(n_350), .D(n_395), .Y(n_431) );
BUFx3_ASAP7_75t_L g441 ( .A(n_278), .Y(n_441) );
OR2x2_ASAP7_75t_L g450 ( .A(n_278), .B(n_451), .Y(n_450) );
OAI211xp5_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_294), .B(n_297), .C(n_305), .Y(n_279) );
AOI221xp5_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_282), .B1(n_286), .B2(n_290), .C(n_292), .Y(n_280) );
OAI322xp33_ASAP7_75t_L g352 ( .A1(n_281), .A2(n_353), .A3(n_358), .B1(n_359), .B2(n_362), .C1(n_363), .C2(n_369), .Y(n_352) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
AND2x2_ASAP7_75t_L g401 ( .A(n_284), .B(n_285), .Y(n_401) );
INVx1_ASAP7_75t_L g453 ( .A(n_284), .Y(n_453) );
INVx2_ASAP7_75t_L g488 ( .A(n_284), .Y(n_488) );
INVx1_ASAP7_75t_L g384 ( .A(n_285), .Y(n_384) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g439 ( .A(n_288), .B(n_401), .Y(n_439) );
INVx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
OR2x2_ASAP7_75t_L g417 ( .A(n_289), .B(n_379), .Y(n_417) );
AND2x4_ASAP7_75t_L g492 ( .A(n_290), .B(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g331 ( .A(n_291), .B(n_332), .Y(n_331) );
INVx2_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_298), .B(n_302), .Y(n_297) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g407 ( .A(n_300), .Y(n_407) );
OR2x2_ASAP7_75t_L g414 ( .A(n_300), .B(n_415), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_303), .B(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g461 ( .A(n_303), .Y(n_461) );
BUFx2_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
HB1xp67_ASAP7_75t_L g336 ( .A(n_304), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_306), .B(n_310), .Y(n_305) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g489 ( .A(n_309), .B(n_403), .Y(n_489) );
AND2x2_ASAP7_75t_L g310 ( .A(n_311), .B(n_312), .Y(n_310) );
INVx2_ASAP7_75t_L g398 ( .A(n_312), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_312), .B(n_483), .Y(n_482) );
AND2x4_ASAP7_75t_L g312 ( .A(n_313), .B(n_317), .Y(n_312) );
AND2x2_ASAP7_75t_L g360 ( .A(n_313), .B(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g368 ( .A(n_313), .Y(n_368) );
INVx1_ASAP7_75t_L g392 ( .A(n_313), .Y(n_392) );
INVx2_ASAP7_75t_SL g491 ( .A(n_317), .Y(n_491) );
OAI322xp33_ASAP7_75t_L g318 ( .A1(n_319), .A2(n_322), .A3(n_325), .B1(n_327), .B2(n_328), .C1(n_334), .C2(n_338), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_320), .B(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
BUFx3_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g349 ( .A(n_324), .B(n_332), .Y(n_349) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
AND2x4_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
AOI21xp5_ASAP7_75t_L g370 ( .A1(n_330), .A2(n_371), .B(n_375), .Y(n_370) );
INVxp67_ASAP7_75t_L g478 ( .A(n_332), .Y(n_478) );
INVx2_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_335), .B(n_345), .Y(n_344) );
AND2x4_ASAP7_75t_L g335 ( .A(n_336), .B(n_337), .Y(n_335) );
INVx2_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_340), .B(n_360), .Y(n_359) );
INVx2_ASAP7_75t_L g451 ( .A(n_340), .Y(n_451) );
O2A1O1Ixp5_ASAP7_75t_L g342 ( .A1(n_343), .A2(n_348), .B(n_351), .C(n_352), .Y(n_342) );
INVxp33_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx2_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
OAI32xp33_ASAP7_75t_L g375 ( .A1(n_346), .A2(n_376), .A3(n_377), .B1(n_382), .B2(n_385), .Y(n_375) );
INVx1_ASAP7_75t_L g365 ( .A(n_347), .Y(n_365) );
BUFx3_ASAP7_75t_L g372 ( .A(n_347), .Y(n_372) );
AND2x2_ASAP7_75t_L g490 ( .A(n_347), .B(n_491), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_347), .B(n_357), .Y(n_497) );
AOI21xp33_ASAP7_75t_L g388 ( .A1(n_348), .A2(n_389), .B(n_397), .Y(n_388) );
AND2x4_ASAP7_75t_L g348 ( .A(n_349), .B(n_350), .Y(n_348) );
INVxp67_ASAP7_75t_R g362 ( .A(n_349), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_351), .B(n_355), .Y(n_444) );
AND2x4_ASAP7_75t_L g468 ( .A(n_351), .B(n_469), .Y(n_468) );
AND2x4_ASAP7_75t_L g479 ( .A(n_351), .B(n_395), .Y(n_479) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
AND2x4_ASAP7_75t_L g354 ( .A(n_355), .B(n_356), .Y(n_354) );
INVx1_ASAP7_75t_L g485 ( .A(n_357), .Y(n_485) );
AOI21xp33_ASAP7_75t_SL g443 ( .A1(n_359), .A2(n_444), .B(n_445), .Y(n_443) );
HB1xp67_ASAP7_75t_L g483 ( .A(n_361), .Y(n_483) );
OAI22xp5_ASAP7_75t_L g397 ( .A1(n_363), .A2(n_398), .B1(n_399), .B2(n_402), .Y(n_397) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_365), .B(n_366), .Y(n_364) );
AND2x4_ASAP7_75t_SL g366 ( .A(n_367), .B(n_368), .Y(n_366) );
AND2x2_ASAP7_75t_L g371 ( .A(n_372), .B(n_373), .Y(n_371) );
INVx1_ASAP7_75t_L g376 ( .A(n_373), .Y(n_376) );
INVxp67_ASAP7_75t_L g423 ( .A(n_373), .Y(n_423) );
AND2x2_ASAP7_75t_L g391 ( .A(n_374), .B(n_392), .Y(n_391) );
INVx2_ASAP7_75t_L g415 ( .A(n_374), .Y(n_415) );
INVx2_ASAP7_75t_L g455 ( .A(n_374), .Y(n_455) );
INVx1_ASAP7_75t_L g463 ( .A(n_376), .Y(n_463) );
INVx3_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
AOI22xp5_ASAP7_75t_L g438 ( .A1(n_378), .A2(n_439), .B1(n_440), .B2(n_442), .Y(n_438) );
AND2x4_ASAP7_75t_L g378 ( .A(n_379), .B(n_381), .Y(n_378) );
INVx1_ASAP7_75t_L g410 ( .A(n_379), .Y(n_410) );
INVx2_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AND2x2_ASAP7_75t_L g446 ( .A(n_383), .B(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
NOR3x1_ASAP7_75t_L g386 ( .A(n_387), .B(n_432), .C(n_480), .Y(n_386) );
NAND3xp33_ASAP7_75t_L g387 ( .A(n_388), .B(n_404), .C(n_412), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_390), .B(n_393), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
AND2x4_ASAP7_75t_L g430 ( .A(n_392), .B(n_421), .Y(n_430) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_395), .B(n_396), .Y(n_394) );
INVx2_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_407), .B(n_455), .Y(n_454) );
OAI21xp5_ASAP7_75t_SL g494 ( .A1(n_408), .A2(n_495), .B(n_496), .Y(n_494) );
AND2x4_ASAP7_75t_L g408 ( .A(n_409), .B(n_411), .Y(n_408) );
INVxp67_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
AOI221xp5_ASAP7_75t_L g412 ( .A1(n_413), .A2(n_416), .B1(n_418), .B2(n_424), .C(n_427), .Y(n_412) );
INVx1_ASAP7_75t_SL g413 ( .A(n_414), .Y(n_413) );
INVx2_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_419), .B(n_423), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
OA21x2_ASAP7_75t_L g481 ( .A1(n_425), .A2(n_482), .B(n_484), .Y(n_481) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
OAI21xp5_ASAP7_75t_L g427 ( .A1(n_428), .A2(n_429), .B(n_431), .Y(n_427) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
AOI22xp33_ASAP7_75t_L g476 ( .A1(n_430), .A2(n_472), .B1(n_477), .B2(n_479), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_433), .B(n_457), .Y(n_432) );
NOR3xp33_ASAP7_75t_L g433 ( .A(n_434), .B(n_443), .C(n_449), .Y(n_433) );
OAI21xp5_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_437), .B(n_438), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
AND2x2_ASAP7_75t_L g499 ( .A(n_439), .B(n_500), .Y(n_499) );
INVxp67_ASAP7_75t_SL g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
OAI22xp33_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_452), .B1(n_454), .B2(n_456), .Y(n_449) );
INVx1_ASAP7_75t_L g500 ( .A(n_455), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g457 ( .A1(n_458), .A2(n_463), .B(n_464), .Y(n_457) );
INVxp67_ASAP7_75t_SL g458 ( .A(n_459), .Y(n_458) );
INVxp67_ASAP7_75t_SL g459 ( .A(n_460), .Y(n_459) );
NOR2x1p5_ASAP7_75t_L g460 ( .A(n_461), .B(n_462), .Y(n_460) );
OAI211xp5_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_467), .B(n_471), .C(n_476), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_472), .B(n_473), .Y(n_471) );
AND2x4_ASAP7_75t_SL g473 ( .A(n_474), .B(n_475), .Y(n_473) );
NAND3xp33_ASAP7_75t_L g480 ( .A(n_481), .B(n_494), .C(n_498), .Y(n_480) );
AOI22xp5_ASAP7_75t_L g484 ( .A1(n_485), .A2(n_486), .B1(n_490), .B2(n_492), .Y(n_484) );
AND2x4_ASAP7_75t_L g486 ( .A(n_487), .B(n_489), .Y(n_486) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
OAI221xp5_ASAP7_75t_L g501 ( .A1(n_502), .A2(n_602), .B1(n_619), .B2(n_622), .C(n_624), .Y(n_501) );
XOR2xp5_ASAP7_75t_L g502 ( .A(n_503), .B(n_591), .Y(n_502) );
AOI22xp5_ASAP7_75t_L g503 ( .A1(n_504), .A2(n_506), .B1(n_507), .B2(n_590), .Y(n_503) );
CKINVDCx5p33_ASAP7_75t_R g590 ( .A(n_504), .Y(n_590) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
OR2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_569), .Y(n_507) );
NAND4xp25_ASAP7_75t_L g508 ( .A(n_509), .B(n_540), .C(n_553), .D(n_557), .Y(n_508) );
AND2x4_ASAP7_75t_L g510 ( .A(n_511), .B(n_520), .Y(n_510) );
AND2x2_ASAP7_75t_L g556 ( .A(n_511), .B(n_544), .Y(n_556) );
AND2x4_ASAP7_75t_L g580 ( .A(n_511), .B(n_581), .Y(n_580) );
AND2x4_ASAP7_75t_L g583 ( .A(n_511), .B(n_578), .Y(n_583) );
AND2x2_ASAP7_75t_L g511 ( .A(n_512), .B(n_519), .Y(n_511) );
INVx1_ASAP7_75t_L g543 ( .A(n_512), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_513), .B(n_516), .Y(n_512) );
NAND2xp33_ASAP7_75t_L g513 ( .A(n_514), .B(n_515), .Y(n_513) );
INVx2_ASAP7_75t_L g518 ( .A(n_514), .Y(n_518) );
INVx3_ASAP7_75t_L g523 ( .A(n_514), .Y(n_523) );
NAND2xp33_ASAP7_75t_L g529 ( .A(n_514), .B(n_530), .Y(n_529) );
HB1xp67_ASAP7_75t_L g534 ( .A(n_514), .Y(n_534) );
INVx1_ASAP7_75t_L g539 ( .A(n_514), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_515), .B(n_551), .Y(n_550) );
INVxp67_ASAP7_75t_L g612 ( .A(n_515), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_517), .B(n_518), .Y(n_516) );
OAI21xp5_ASAP7_75t_L g537 ( .A1(n_517), .A2(n_538), .B(n_539), .Y(n_537) );
AND2x2_ASAP7_75t_L g536 ( .A(n_519), .B(n_537), .Y(n_536) );
AND2x2_ASAP7_75t_L g542 ( .A(n_519), .B(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g573 ( .A(n_519), .Y(n_573) );
AND2x4_ASAP7_75t_L g558 ( .A(n_520), .B(n_542), .Y(n_558) );
AND2x4_ASAP7_75t_L g585 ( .A(n_520), .B(n_572), .Y(n_585) );
AND2x4_ASAP7_75t_L g520 ( .A(n_521), .B(n_525), .Y(n_520) );
AND2x2_ASAP7_75t_L g532 ( .A(n_521), .B(n_533), .Y(n_532) );
INVx2_ASAP7_75t_L g545 ( .A(n_521), .Y(n_545) );
OR2x2_ASAP7_75t_L g575 ( .A(n_521), .B(n_576), .Y(n_575) );
AND2x4_ASAP7_75t_L g581 ( .A(n_521), .B(n_582), .Y(n_581) );
AND2x4_ASAP7_75t_L g521 ( .A(n_522), .B(n_524), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_523), .B(n_528), .Y(n_527) );
INVxp67_ASAP7_75t_L g549 ( .A(n_523), .Y(n_549) );
NAND3xp33_ASAP7_75t_L g567 ( .A(n_524), .B(n_548), .C(n_568), .Y(n_567) );
AND2x4_ASAP7_75t_L g544 ( .A(n_525), .B(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g576 ( .A(n_526), .Y(n_576) );
AND2x2_ASAP7_75t_L g526 ( .A(n_527), .B(n_529), .Y(n_526) );
AND2x2_ASAP7_75t_L g531 ( .A(n_532), .B(n_536), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_534), .B(n_535), .Y(n_533) );
INVx1_ASAP7_75t_L g563 ( .A(n_534), .Y(n_563) );
HB1xp67_ASAP7_75t_L g609 ( .A(n_535), .Y(n_609) );
AND2x2_ASAP7_75t_L g541 ( .A(n_542), .B(n_544), .Y(n_541) );
AND2x4_ASAP7_75t_L g572 ( .A(n_543), .B(n_573), .Y(n_572) );
AND2x4_ASAP7_75t_L g546 ( .A(n_544), .B(n_547), .Y(n_546) );
AND2x4_ASAP7_75t_L g586 ( .A(n_544), .B(n_572), .Y(n_586) );
AND2x4_ASAP7_75t_L g577 ( .A(n_547), .B(n_578), .Y(n_577) );
AND2x4_ASAP7_75t_L g589 ( .A(n_547), .B(n_581), .Y(n_589) );
AND2x2_ASAP7_75t_L g547 ( .A(n_548), .B(n_552), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_549), .B(n_550), .Y(n_548) );
HB1xp67_ASAP7_75t_L g613 ( .A(n_551), .Y(n_613) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx4_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx3_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
AO21x2_ASAP7_75t_L g562 ( .A1(n_563), .A2(n_564), .B(n_567), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_565), .B(n_566), .Y(n_564) );
NAND4xp25_ASAP7_75t_L g569 ( .A(n_570), .B(n_579), .C(n_584), .D(n_587), .Y(n_569) );
AND2x4_ASAP7_75t_L g571 ( .A(n_572), .B(n_574), .Y(n_571) );
AND2x4_ASAP7_75t_L g588 ( .A(n_572), .B(n_581), .Y(n_588) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx2_ASAP7_75t_L g578 ( .A(n_575), .Y(n_578) );
INVx1_ASAP7_75t_L g582 ( .A(n_576), .Y(n_582) );
OAI22xp5_ASAP7_75t_L g591 ( .A1(n_592), .A2(n_593), .B1(n_594), .B2(n_595), .Y(n_591) );
CKINVDCx5p33_ASAP7_75t_R g592 ( .A(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
AOI22xp5_ASAP7_75t_L g595 ( .A1(n_596), .A2(n_597), .B1(n_598), .B2(n_599), .Y(n_595) );
CKINVDCx5p33_ASAP7_75t_R g596 ( .A(n_597), .Y(n_596) );
CKINVDCx20_ASAP7_75t_R g598 ( .A(n_599), .Y(n_598) );
XNOR2xp5_ASAP7_75t_L g599 ( .A(n_600), .B(n_601), .Y(n_599) );
INVx1_ASAP7_75t_SL g602 ( .A(n_603), .Y(n_602) );
BUFx2_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
CKINVDCx5p33_ASAP7_75t_R g604 ( .A(n_605), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_606), .B(n_614), .Y(n_605) );
INVxp67_ASAP7_75t_SL g606 ( .A(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g633 ( .A(n_607), .B(n_614), .Y(n_633) );
AOI211xp5_ASAP7_75t_L g607 ( .A1(n_608), .A2(n_609), .B(n_610), .C(n_613), .Y(n_607) );
NOR2xp33_ASAP7_75t_L g610 ( .A(n_611), .B(n_612), .Y(n_610) );
NOR2xp33_ASAP7_75t_L g614 ( .A(n_615), .B(n_617), .Y(n_614) );
OR2x2_ASAP7_75t_L g623 ( .A(n_615), .B(n_618), .Y(n_623) );
INVx1_ASAP7_75t_L g629 ( .A(n_615), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_615), .B(n_617), .Y(n_630) );
HB1xp67_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
BUFx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
AOI22xp5_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_626), .B1(n_631), .B2(n_634), .Y(n_624) );
CKINVDCx20_ASAP7_75t_R g626 ( .A(n_627), .Y(n_626) );
BUFx2_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
INVx1_ASAP7_75t_SL g632 ( .A(n_633), .Y(n_632) );
endmodule