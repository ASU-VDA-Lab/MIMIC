module fake_netlist_5_1973_n_5639 (n_924, n_1263, n_977, n_1378, n_611, n_1126, n_1423, n_1166, n_469, n_1508, n_82, n_785, n_549, n_532, n_1161, n_1150, n_226, n_1488, n_667, n_790, n_1055, n_1501, n_111, n_880, n_544, n_1007, n_155, n_552, n_1528, n_1370, n_1292, n_1198, n_1360, n_1099, n_956, n_564, n_423, n_21, n_105, n_1021, n_4, n_551, n_1323, n_1466, n_688, n_1353, n_800, n_1347, n_1535, n_671, n_819, n_1451, n_1022, n_915, n_1545, n_864, n_173, n_859, n_951, n_1264, n_447, n_247, n_1494, n_292, n_625, n_854, n_1462, n_1580, n_674, n_417, n_516, n_933, n_1152, n_497, n_1607, n_1563, n_606, n_275, n_26, n_877, n_2, n_755, n_1118, n_6, n_947, n_1285, n_373, n_307, n_1359, n_530, n_87, n_150, n_1107, n_556, n_1230, n_668, n_375, n_301, n_929, n_1124, n_902, n_1576, n_191, n_1104, n_1294, n_659, n_51, n_1257, n_171, n_1182, n_579, n_1261, n_938, n_1098, n_320, n_1154, n_1242, n_1135, n_24, n_406, n_519, n_1016, n_1243, n_546, n_101, n_1280, n_281, n_240, n_291, n_231, n_257, n_731, n_371, n_1483, n_1314, n_1512, n_709, n_1490, n_317, n_1236, n_569, n_227, n_920, n_1289, n_1517, n_94, n_335, n_370, n_976, n_343, n_1449, n_308, n_1566, n_297, n_156, n_1078, n_775, n_219, n_157, n_600, n_1484, n_1374, n_1328, n_223, n_264, n_1598, n_955, n_163, n_339, n_1146, n_882, n_183, n_243, n_1036, n_1097, n_347, n_59, n_550, n_696, n_897, n_215, n_350, n_196, n_798, n_646, n_1428, n_436, n_1394, n_1414, n_1216, n_290, n_580, n_1040, n_578, n_926, n_344, n_1218, n_422, n_475, n_777, n_1070, n_1547, n_1030, n_72, n_415, n_1071, n_485, n_1165, n_1267, n_1561, n_496, n_1391, n_958, n_1034, n_670, n_1513, n_1600, n_48, n_521, n_663, n_845, n_673, n_837, n_1239, n_528, n_680, n_1473, n_1587, n_395, n_164, n_553, n_901, n_813, n_1521, n_1284, n_1590, n_214, n_675, n_888, n_1167, n_1626, n_637, n_1384, n_1556, n_184, n_446, n_1064, n_144, n_858, n_114, n_96, n_923, n_691, n_1151, n_881, n_1405, n_468, n_213, n_129, n_342, n_464, n_363, n_1582, n_197, n_1069, n_1075, n_1450, n_1322, n_1471, n_1459, n_460, n_889, n_973, n_477, n_571, n_1585, n_461, n_1599, n_1211, n_1197, n_1523, n_907, n_1447, n_1377, n_190, n_989, n_1039, n_34, n_228, n_283, n_1403, n_488, n_736, n_892, n_1000, n_1202, n_1278, n_1002, n_1463, n_1581, n_49, n_310, n_54, n_593, n_12, n_748, n_586, n_1058, n_838, n_332, n_1053, n_1224, n_349, n_1248, n_230, n_1331, n_953, n_279, n_1014, n_1241, n_70, n_289, n_963, n_1052, n_954, n_627, n_1385, n_440, n_793, n_478, n_476, n_1527, n_534, n_884, n_345, n_944, n_1623, n_91, n_1565, n_182, n_143, n_647, n_237, n_407, n_1072, n_832, n_857, n_207, n_561, n_1319, n_1387, n_1532, n_18, n_1027, n_971, n_1156, n_117, n_326, n_794, n_404, n_686, n_847, n_1393, n_596, n_1368, n_558, n_702, n_1276, n_822, n_1412, n_728, n_266, n_1162, n_272, n_1538, n_1199, n_352, n_53, n_1038, n_520, n_1369, n_409, n_887, n_154, n_71, n_300, n_809, n_870, n_931, n_599, n_1481, n_434, n_1544, n_868, n_639, n_914, n_411, n_414, n_1293, n_965, n_935, n_121, n_1175, n_817, n_360, n_36, n_1479, n_64, n_759, n_28, n_806, n_1477, n_324, n_1571, n_187, n_1189, n_103, n_97, n_11, n_7, n_1259, n_706, n_746, n_747, n_52, n_784, n_110, n_1244, n_431, n_1194, n_615, n_851, n_843, n_523, n_913, n_1537, n_705, n_865, n_61, n_678, n_697, n_127, n_1222, n_75, n_776, n_1415, n_367, n_452, n_525, n_1260, n_1464, n_649, n_547, n_43, n_1444, n_1191, n_116, n_284, n_1128, n_139, n_744, n_590, n_629, n_1308, n_254, n_1233, n_23, n_1615, n_1529, n_526, n_293, n_372, n_677, n_244, n_47, n_1333, n_1121, n_314, n_368, n_433, n_604, n_8, n_949, n_100, n_1443, n_1008, n_946, n_1539, n_1001, n_1503, n_498, n_1468, n_1559, n_689, n_738, n_1624, n_640, n_1510, n_252, n_624, n_1380, n_1617, n_295, n_133, n_1010, n_1231, n_739, n_1279, n_1406, n_1195, n_610, n_936, n_568, n_1500, n_39, n_1090, n_757, n_633, n_439, n_106, n_259, n_448, n_758, n_999, n_93, n_1158, n_1509, n_563, n_1145, n_878, n_524, n_204, n_394, n_1049, n_1153, n_741, n_1306, n_1068, n_122, n_331, n_10, n_906, n_1163, n_1207, n_919, n_908, n_90, n_724, n_658, n_1362, n_1586, n_456, n_959, n_535, n_152, n_940, n_1445, n_9, n_1492, n_592, n_1169, n_45, n_1596, n_1017, n_123, n_978, n_1434, n_1054, n_1474, n_1269, n_1095, n_1614, n_267, n_514, n_457, n_1079, n_1045, n_1208, n_603, n_1431, n_484, n_1593, n_1033, n_442, n_131, n_636, n_660, n_1009, n_1148, n_109, n_742, n_750, n_995, n_454, n_1609, n_374, n_185, n_396, n_1383, n_1073, n_255, n_662, n_459, n_218, n_962, n_1215, n_1171, n_1578, n_723, n_1065, n_1592, n_1336, n_1574, n_473, n_1309, n_1426, n_1043, n_355, n_486, n_1548, n_614, n_337, n_1421, n_88, n_1286, n_1177, n_1355, n_168, n_974, n_727, n_1159, n_957, n_773, n_208, n_142, n_743, n_299, n_303, n_296, n_613, n_1119, n_1240, n_65, n_829, n_1612, n_1416, n_361, n_700, n_1237, n_573, n_69, n_1420, n_1132, n_388, n_1366, n_1300, n_1127, n_761, n_1568, n_1006, n_329, n_274, n_1270, n_1486, n_582, n_1332, n_1390, n_73, n_19, n_309, n_30, n_512, n_1591, n_84, n_130, n_322, n_1249, n_652, n_1111, n_1365, n_25, n_1349, n_1093, n_288, n_1031, n_263, n_609, n_1041, n_1265, n_44, n_224, n_1562, n_383, n_834, n_112, n_765, n_893, n_1015, n_1140, n_891, n_239, n_630, n_55, n_504, n_511, n_874, n_358, n_1101, n_77, n_102, n_1106, n_1456, n_1304, n_1324, n_987, n_261, n_174, n_1455, n_767, n_993, n_1407, n_1551, n_545, n_441, n_860, n_450, n_429, n_948, n_1217, n_628, n_365, n_729, n_1131, n_1084, n_970, n_911, n_1430, n_83, n_513, n_1094, n_1354, n_560, n_1534, n_340, n_1351, n_1044, n_1205, n_346, n_1209, n_1552, n_495, n_602, n_574, n_1435, n_879, n_16, n_58, n_623, n_405, n_824, n_359, n_490, n_1327, n_996, n_921, n_233, n_572, n_366, n_815, n_128, n_120, n_327, n_135, n_1381, n_1611, n_1037, n_1080, n_1274, n_1316, n_426, n_1438, n_1082, n_589, n_716, n_562, n_1436, n_62, n_952, n_1229, n_391, n_701, n_1437, n_1023, n_645, n_539, n_803, n_1092, n_238, n_531, n_890, n_764, n_1056, n_1424, n_162, n_960, n_222, n_1290, n_1123, n_1467, n_1047, n_634, n_199, n_32, n_1252, n_348, n_1382, n_1029, n_925, n_1206, n_424, n_1311, n_1519, n_256, n_950, n_1553, n_380, n_419, n_1346, n_444, n_1299, n_1060, n_1141, n_316, n_389, n_418, n_248, n_136, n_86, n_146, n_912, n_315, n_968, n_451, n_619, n_408, n_1386, n_376, n_967, n_1442, n_74, n_1139, n_515, n_57, n_351, n_885, n_397, n_1432, n_1357, n_483, n_683, n_1057, n_1051, n_1085, n_1066, n_721, n_1157, n_841, n_1050, n_22, n_802, n_46, n_1608, n_983, n_38, n_280, n_1305, n_873, n_378, n_1112, n_762, n_1283, n_17, n_690, n_33, n_583, n_302, n_1343, n_1203, n_821, n_321, n_1179, n_621, n_753, n_455, n_1048, n_1288, n_212, n_385, n_507, n_1560, n_1605, n_330, n_1228, n_972, n_692, n_820, n_1200, n_1301, n_1363, n_1185, n_991, n_828, n_779, n_576, n_1143, n_1579, n_1329, n_1312, n_1439, n_804, n_537, n_945, n_492, n_153, n_1504, n_943, n_341, n_250, n_992, n_543, n_260, n_842, n_650, n_984, n_694, n_286, n_883, n_470, n_325, n_449, n_1594, n_132, n_1214, n_1342, n_1400, n_900, n_856, n_918, n_942, n_189, n_1147, n_1557, n_1610, n_13, n_1077, n_1422, n_540, n_618, n_896, n_323, n_195, n_356, n_894, n_831, n_964, n_1373, n_1350, n_1511, n_1470, n_1096, n_234, n_1575, n_833, n_5, n_225, n_1307, n_988, n_814, n_192, n_1549, n_1201, n_1114, n_655, n_1616, n_1446, n_669, n_472, n_1458, n_1176, n_1472, n_387, n_1149, n_398, n_635, n_763, n_1020, n_1062, n_211, n_1219, n_3, n_1204, n_178, n_1035, n_287, n_555, n_783, n_1188, n_661, n_41, n_849, n_15, n_336, n_584, n_681, n_50, n_430, n_510, n_216, n_311, n_830, n_1296, n_1413, n_801, n_241, n_875, n_357, n_1110, n_445, n_749, n_1134, n_1358, n_717, n_165, n_939, n_482, n_1088, n_588, n_1173, n_789, n_1232, n_1603, n_734, n_638, n_866, n_107, n_969, n_1401, n_1019, n_1105, n_249, n_304, n_1338, n_577, n_1522, n_1419, n_338, n_149, n_693, n_1506, n_14, n_836, n_990, n_1389, n_975, n_1256, n_567, n_1465, n_778, n_1122, n_151, n_306, n_458, n_770, n_1375, n_1102, n_711, n_1499, n_85, n_1187, n_1441, n_1392, n_1597, n_1164, n_489, n_1174, n_1371, n_617, n_1303, n_1572, n_876, n_1516, n_1190, n_118, n_601, n_917, n_966, n_253, n_1116, n_1212, n_1541, n_172, n_206, n_217, n_726, n_982, n_1573, n_1453, n_818, n_861, n_1183, n_899, n_1253, n_210, n_774, n_1628, n_1335, n_1514, n_1059, n_1345, n_176, n_1133, n_557, n_1410, n_1005, n_607, n_1003, n_679, n_710, n_527, n_1168, n_707, n_937, n_1427, n_393, n_108, n_487, n_1584, n_665, n_66, n_1440, n_177, n_421, n_1356, n_910, n_768, n_1475, n_1302, n_205, n_1136, n_1313, n_1491, n_754, n_1496, n_179, n_1125, n_125, n_410, n_708, n_529, n_735, n_232, n_1109, n_126, n_895, n_1310, n_202, n_427, n_1399, n_1543, n_791, n_732, n_1533, n_193, n_808, n_797, n_1025, n_500, n_1067, n_148, n_435, n_159, n_766, n_1457, n_541, n_538, n_1117, n_799, n_687, n_715, n_1480, n_1482, n_1213, n_1266, n_536, n_872, n_594, n_200, n_1291, n_1297, n_1155, n_1418, n_89, n_1524, n_1485, n_115, n_1011, n_1184, n_985, n_869, n_810, n_416, n_827, n_401, n_1352, n_626, n_1144, n_1137, n_1570, n_1170, n_305, n_137, n_676, n_294, n_318, n_653, n_642, n_1602, n_194, n_855, n_1178, n_1461, n_850, n_684, n_124, n_268, n_664, n_503, n_235, n_1372, n_605, n_1273, n_353, n_620, n_643, n_916, n_1081, n_493, n_1235, n_703, n_698, n_980, n_1115, n_1282, n_1318, n_780, n_998, n_1454, n_467, n_1227, n_1531, n_840, n_1334, n_501, n_823, n_245, n_725, n_1388, n_1417, n_1295, n_672, n_581, n_382, n_554, n_1625, n_898, n_1013, n_1452, n_718, n_265, n_1120, n_719, n_443, n_198, n_714, n_909, n_1497, n_1530, n_997, n_932, n_612, n_1409, n_788, n_1326, n_119, n_1268, n_559, n_825, n_508, n_506, n_1320, n_737, n_986, n_509, n_1317, n_147, n_1518, n_1281, n_67, n_1192, n_1024, n_1063, n_209, n_1564, n_1613, n_733, n_1489, n_1376, n_941, n_981, n_1569, n_68, n_867, n_186, n_134, n_587, n_63, n_792, n_756, n_1429, n_399, n_1238, n_548, n_812, n_298, n_518, n_505, n_282, n_752, n_905, n_1476, n_1108, n_782, n_1100, n_1395, n_862, n_1425, n_760, n_1620, n_381, n_220, n_390, n_1330, n_31, n_481, n_1554, n_769, n_42, n_1046, n_271, n_934, n_1618, n_826, n_886, n_1221, n_654, n_1172, n_167, n_379, n_428, n_1341, n_570, n_1361, n_853, n_377, n_751, n_786, n_1083, n_1142, n_1129, n_392, n_158, n_704, n_787, n_138, n_961, n_771, n_276, n_95, n_1225, n_1520, n_169, n_522, n_1287, n_1262, n_400, n_930, n_181, n_1411, n_221, n_622, n_1577, n_1087, n_386, n_994, n_848, n_1550, n_1498, n_1223, n_1272, n_104, n_682, n_1567, n_56, n_141, n_1247, n_922, n_816, n_591, n_145, n_1536, n_1344, n_313, n_631, n_479, n_1246, n_1339, n_1478, n_432, n_839, n_1210, n_1364, n_328, n_140, n_1250, n_369, n_871, n_598, n_685, n_928, n_608, n_1367, n_78, n_1460, n_772, n_1555, n_499, n_1589, n_517, n_98, n_402, n_413, n_1086, n_796, n_1619, n_236, n_1502, n_1469, n_1012, n_1, n_1396, n_1348, n_903, n_1525, n_740, n_203, n_384, n_1404, n_80, n_35, n_1315, n_277, n_1061, n_92, n_333, n_1298, n_462, n_1193, n_1255, n_258, n_1113, n_29, n_79, n_1226, n_722, n_1277, n_188, n_844, n_201, n_471, n_852, n_1487, n_40, n_1028, n_1601, n_781, n_474, n_542, n_463, n_1546, n_595, n_502, n_466, n_420, n_1337, n_1495, n_632, n_699, n_979, n_1515, n_1627, n_1245, n_846, n_465, n_76, n_362, n_1321, n_170, n_27, n_161, n_273, n_585, n_270, n_616, n_81, n_745, n_1103, n_648, n_1379, n_312, n_1076, n_1091, n_1408, n_494, n_641, n_730, n_1325, n_1595, n_354, n_575, n_480, n_425, n_795, n_695, n_180, n_656, n_1606, n_1220, n_37, n_1540, n_229, n_437, n_60, n_403, n_453, n_1130, n_720, n_0, n_1526, n_863, n_805, n_1604, n_1275, n_113, n_712, n_246, n_1583, n_1042, n_1402, n_269, n_285, n_412, n_1493, n_657, n_644, n_1160, n_1397, n_491, n_1258, n_1074, n_1621, n_251, n_160, n_566, n_565, n_1448, n_1507, n_1398, n_597, n_1181, n_1505, n_1196, n_651, n_1340, n_334, n_811, n_1558, n_807, n_835, n_175, n_666, n_262, n_1433, n_99, n_1254, n_1026, n_1234, n_319, n_364, n_1138, n_927, n_20, n_1089, n_1004, n_1186, n_1032, n_242, n_1018, n_438, n_713, n_904, n_1588, n_1622, n_166, n_1180, n_1271, n_533, n_1542, n_1251, n_278, n_5639);

input n_924;
input n_1263;
input n_977;
input n_1378;
input n_611;
input n_1126;
input n_1423;
input n_1166;
input n_469;
input n_1508;
input n_82;
input n_785;
input n_549;
input n_532;
input n_1161;
input n_1150;
input n_226;
input n_1488;
input n_667;
input n_790;
input n_1055;
input n_1501;
input n_111;
input n_880;
input n_544;
input n_1007;
input n_155;
input n_552;
input n_1528;
input n_1370;
input n_1292;
input n_1198;
input n_1360;
input n_1099;
input n_956;
input n_564;
input n_423;
input n_21;
input n_105;
input n_1021;
input n_4;
input n_551;
input n_1323;
input n_1466;
input n_688;
input n_1353;
input n_800;
input n_1347;
input n_1535;
input n_671;
input n_819;
input n_1451;
input n_1022;
input n_915;
input n_1545;
input n_864;
input n_173;
input n_859;
input n_951;
input n_1264;
input n_447;
input n_247;
input n_1494;
input n_292;
input n_625;
input n_854;
input n_1462;
input n_1580;
input n_674;
input n_417;
input n_516;
input n_933;
input n_1152;
input n_497;
input n_1607;
input n_1563;
input n_606;
input n_275;
input n_26;
input n_877;
input n_2;
input n_755;
input n_1118;
input n_6;
input n_947;
input n_1285;
input n_373;
input n_307;
input n_1359;
input n_530;
input n_87;
input n_150;
input n_1107;
input n_556;
input n_1230;
input n_668;
input n_375;
input n_301;
input n_929;
input n_1124;
input n_902;
input n_1576;
input n_191;
input n_1104;
input n_1294;
input n_659;
input n_51;
input n_1257;
input n_171;
input n_1182;
input n_579;
input n_1261;
input n_938;
input n_1098;
input n_320;
input n_1154;
input n_1242;
input n_1135;
input n_24;
input n_406;
input n_519;
input n_1016;
input n_1243;
input n_546;
input n_101;
input n_1280;
input n_281;
input n_240;
input n_291;
input n_231;
input n_257;
input n_731;
input n_371;
input n_1483;
input n_1314;
input n_1512;
input n_709;
input n_1490;
input n_317;
input n_1236;
input n_569;
input n_227;
input n_920;
input n_1289;
input n_1517;
input n_94;
input n_335;
input n_370;
input n_976;
input n_343;
input n_1449;
input n_308;
input n_1566;
input n_297;
input n_156;
input n_1078;
input n_775;
input n_219;
input n_157;
input n_600;
input n_1484;
input n_1374;
input n_1328;
input n_223;
input n_264;
input n_1598;
input n_955;
input n_163;
input n_339;
input n_1146;
input n_882;
input n_183;
input n_243;
input n_1036;
input n_1097;
input n_347;
input n_59;
input n_550;
input n_696;
input n_897;
input n_215;
input n_350;
input n_196;
input n_798;
input n_646;
input n_1428;
input n_436;
input n_1394;
input n_1414;
input n_1216;
input n_290;
input n_580;
input n_1040;
input n_578;
input n_926;
input n_344;
input n_1218;
input n_422;
input n_475;
input n_777;
input n_1070;
input n_1547;
input n_1030;
input n_72;
input n_415;
input n_1071;
input n_485;
input n_1165;
input n_1267;
input n_1561;
input n_496;
input n_1391;
input n_958;
input n_1034;
input n_670;
input n_1513;
input n_1600;
input n_48;
input n_521;
input n_663;
input n_845;
input n_673;
input n_837;
input n_1239;
input n_528;
input n_680;
input n_1473;
input n_1587;
input n_395;
input n_164;
input n_553;
input n_901;
input n_813;
input n_1521;
input n_1284;
input n_1590;
input n_214;
input n_675;
input n_888;
input n_1167;
input n_1626;
input n_637;
input n_1384;
input n_1556;
input n_184;
input n_446;
input n_1064;
input n_144;
input n_858;
input n_114;
input n_96;
input n_923;
input n_691;
input n_1151;
input n_881;
input n_1405;
input n_468;
input n_213;
input n_129;
input n_342;
input n_464;
input n_363;
input n_1582;
input n_197;
input n_1069;
input n_1075;
input n_1450;
input n_1322;
input n_1471;
input n_1459;
input n_460;
input n_889;
input n_973;
input n_477;
input n_571;
input n_1585;
input n_461;
input n_1599;
input n_1211;
input n_1197;
input n_1523;
input n_907;
input n_1447;
input n_1377;
input n_190;
input n_989;
input n_1039;
input n_34;
input n_228;
input n_283;
input n_1403;
input n_488;
input n_736;
input n_892;
input n_1000;
input n_1202;
input n_1278;
input n_1002;
input n_1463;
input n_1581;
input n_49;
input n_310;
input n_54;
input n_593;
input n_12;
input n_748;
input n_586;
input n_1058;
input n_838;
input n_332;
input n_1053;
input n_1224;
input n_349;
input n_1248;
input n_230;
input n_1331;
input n_953;
input n_279;
input n_1014;
input n_1241;
input n_70;
input n_289;
input n_963;
input n_1052;
input n_954;
input n_627;
input n_1385;
input n_440;
input n_793;
input n_478;
input n_476;
input n_1527;
input n_534;
input n_884;
input n_345;
input n_944;
input n_1623;
input n_91;
input n_1565;
input n_182;
input n_143;
input n_647;
input n_237;
input n_407;
input n_1072;
input n_832;
input n_857;
input n_207;
input n_561;
input n_1319;
input n_1387;
input n_1532;
input n_18;
input n_1027;
input n_971;
input n_1156;
input n_117;
input n_326;
input n_794;
input n_404;
input n_686;
input n_847;
input n_1393;
input n_596;
input n_1368;
input n_558;
input n_702;
input n_1276;
input n_822;
input n_1412;
input n_728;
input n_266;
input n_1162;
input n_272;
input n_1538;
input n_1199;
input n_352;
input n_53;
input n_1038;
input n_520;
input n_1369;
input n_409;
input n_887;
input n_154;
input n_71;
input n_300;
input n_809;
input n_870;
input n_931;
input n_599;
input n_1481;
input n_434;
input n_1544;
input n_868;
input n_639;
input n_914;
input n_411;
input n_414;
input n_1293;
input n_965;
input n_935;
input n_121;
input n_1175;
input n_817;
input n_360;
input n_36;
input n_1479;
input n_64;
input n_759;
input n_28;
input n_806;
input n_1477;
input n_324;
input n_1571;
input n_187;
input n_1189;
input n_103;
input n_97;
input n_11;
input n_7;
input n_1259;
input n_706;
input n_746;
input n_747;
input n_52;
input n_784;
input n_110;
input n_1244;
input n_431;
input n_1194;
input n_615;
input n_851;
input n_843;
input n_523;
input n_913;
input n_1537;
input n_705;
input n_865;
input n_61;
input n_678;
input n_697;
input n_127;
input n_1222;
input n_75;
input n_776;
input n_1415;
input n_367;
input n_452;
input n_525;
input n_1260;
input n_1464;
input n_649;
input n_547;
input n_43;
input n_1444;
input n_1191;
input n_116;
input n_284;
input n_1128;
input n_139;
input n_744;
input n_590;
input n_629;
input n_1308;
input n_254;
input n_1233;
input n_23;
input n_1615;
input n_1529;
input n_526;
input n_293;
input n_372;
input n_677;
input n_244;
input n_47;
input n_1333;
input n_1121;
input n_314;
input n_368;
input n_433;
input n_604;
input n_8;
input n_949;
input n_100;
input n_1443;
input n_1008;
input n_946;
input n_1539;
input n_1001;
input n_1503;
input n_498;
input n_1468;
input n_1559;
input n_689;
input n_738;
input n_1624;
input n_640;
input n_1510;
input n_252;
input n_624;
input n_1380;
input n_1617;
input n_295;
input n_133;
input n_1010;
input n_1231;
input n_739;
input n_1279;
input n_1406;
input n_1195;
input n_610;
input n_936;
input n_568;
input n_1500;
input n_39;
input n_1090;
input n_757;
input n_633;
input n_439;
input n_106;
input n_259;
input n_448;
input n_758;
input n_999;
input n_93;
input n_1158;
input n_1509;
input n_563;
input n_1145;
input n_878;
input n_524;
input n_204;
input n_394;
input n_1049;
input n_1153;
input n_741;
input n_1306;
input n_1068;
input n_122;
input n_331;
input n_10;
input n_906;
input n_1163;
input n_1207;
input n_919;
input n_908;
input n_90;
input n_724;
input n_658;
input n_1362;
input n_1586;
input n_456;
input n_959;
input n_535;
input n_152;
input n_940;
input n_1445;
input n_9;
input n_1492;
input n_592;
input n_1169;
input n_45;
input n_1596;
input n_1017;
input n_123;
input n_978;
input n_1434;
input n_1054;
input n_1474;
input n_1269;
input n_1095;
input n_1614;
input n_267;
input n_514;
input n_457;
input n_1079;
input n_1045;
input n_1208;
input n_603;
input n_1431;
input n_484;
input n_1593;
input n_1033;
input n_442;
input n_131;
input n_636;
input n_660;
input n_1009;
input n_1148;
input n_109;
input n_742;
input n_750;
input n_995;
input n_454;
input n_1609;
input n_374;
input n_185;
input n_396;
input n_1383;
input n_1073;
input n_255;
input n_662;
input n_459;
input n_218;
input n_962;
input n_1215;
input n_1171;
input n_1578;
input n_723;
input n_1065;
input n_1592;
input n_1336;
input n_1574;
input n_473;
input n_1309;
input n_1426;
input n_1043;
input n_355;
input n_486;
input n_1548;
input n_614;
input n_337;
input n_1421;
input n_88;
input n_1286;
input n_1177;
input n_1355;
input n_168;
input n_974;
input n_727;
input n_1159;
input n_957;
input n_773;
input n_208;
input n_142;
input n_743;
input n_299;
input n_303;
input n_296;
input n_613;
input n_1119;
input n_1240;
input n_65;
input n_829;
input n_1612;
input n_1416;
input n_361;
input n_700;
input n_1237;
input n_573;
input n_69;
input n_1420;
input n_1132;
input n_388;
input n_1366;
input n_1300;
input n_1127;
input n_761;
input n_1568;
input n_1006;
input n_329;
input n_274;
input n_1270;
input n_1486;
input n_582;
input n_1332;
input n_1390;
input n_73;
input n_19;
input n_309;
input n_30;
input n_512;
input n_1591;
input n_84;
input n_130;
input n_322;
input n_1249;
input n_652;
input n_1111;
input n_1365;
input n_25;
input n_1349;
input n_1093;
input n_288;
input n_1031;
input n_263;
input n_609;
input n_1041;
input n_1265;
input n_44;
input n_224;
input n_1562;
input n_383;
input n_834;
input n_112;
input n_765;
input n_893;
input n_1015;
input n_1140;
input n_891;
input n_239;
input n_630;
input n_55;
input n_504;
input n_511;
input n_874;
input n_358;
input n_1101;
input n_77;
input n_102;
input n_1106;
input n_1456;
input n_1304;
input n_1324;
input n_987;
input n_261;
input n_174;
input n_1455;
input n_767;
input n_993;
input n_1407;
input n_1551;
input n_545;
input n_441;
input n_860;
input n_450;
input n_429;
input n_948;
input n_1217;
input n_628;
input n_365;
input n_729;
input n_1131;
input n_1084;
input n_970;
input n_911;
input n_1430;
input n_83;
input n_513;
input n_1094;
input n_1354;
input n_560;
input n_1534;
input n_340;
input n_1351;
input n_1044;
input n_1205;
input n_346;
input n_1209;
input n_1552;
input n_495;
input n_602;
input n_574;
input n_1435;
input n_879;
input n_16;
input n_58;
input n_623;
input n_405;
input n_824;
input n_359;
input n_490;
input n_1327;
input n_996;
input n_921;
input n_233;
input n_572;
input n_366;
input n_815;
input n_128;
input n_120;
input n_327;
input n_135;
input n_1381;
input n_1611;
input n_1037;
input n_1080;
input n_1274;
input n_1316;
input n_426;
input n_1438;
input n_1082;
input n_589;
input n_716;
input n_562;
input n_1436;
input n_62;
input n_952;
input n_1229;
input n_391;
input n_701;
input n_1437;
input n_1023;
input n_645;
input n_539;
input n_803;
input n_1092;
input n_238;
input n_531;
input n_890;
input n_764;
input n_1056;
input n_1424;
input n_162;
input n_960;
input n_222;
input n_1290;
input n_1123;
input n_1467;
input n_1047;
input n_634;
input n_199;
input n_32;
input n_1252;
input n_348;
input n_1382;
input n_1029;
input n_925;
input n_1206;
input n_424;
input n_1311;
input n_1519;
input n_256;
input n_950;
input n_1553;
input n_380;
input n_419;
input n_1346;
input n_444;
input n_1299;
input n_1060;
input n_1141;
input n_316;
input n_389;
input n_418;
input n_248;
input n_136;
input n_86;
input n_146;
input n_912;
input n_315;
input n_968;
input n_451;
input n_619;
input n_408;
input n_1386;
input n_376;
input n_967;
input n_1442;
input n_74;
input n_1139;
input n_515;
input n_57;
input n_351;
input n_885;
input n_397;
input n_1432;
input n_1357;
input n_483;
input n_683;
input n_1057;
input n_1051;
input n_1085;
input n_1066;
input n_721;
input n_1157;
input n_841;
input n_1050;
input n_22;
input n_802;
input n_46;
input n_1608;
input n_983;
input n_38;
input n_280;
input n_1305;
input n_873;
input n_378;
input n_1112;
input n_762;
input n_1283;
input n_17;
input n_690;
input n_33;
input n_583;
input n_302;
input n_1343;
input n_1203;
input n_821;
input n_321;
input n_1179;
input n_621;
input n_753;
input n_455;
input n_1048;
input n_1288;
input n_212;
input n_385;
input n_507;
input n_1560;
input n_1605;
input n_330;
input n_1228;
input n_972;
input n_692;
input n_820;
input n_1200;
input n_1301;
input n_1363;
input n_1185;
input n_991;
input n_828;
input n_779;
input n_576;
input n_1143;
input n_1579;
input n_1329;
input n_1312;
input n_1439;
input n_804;
input n_537;
input n_945;
input n_492;
input n_153;
input n_1504;
input n_943;
input n_341;
input n_250;
input n_992;
input n_543;
input n_260;
input n_842;
input n_650;
input n_984;
input n_694;
input n_286;
input n_883;
input n_470;
input n_325;
input n_449;
input n_1594;
input n_132;
input n_1214;
input n_1342;
input n_1400;
input n_900;
input n_856;
input n_918;
input n_942;
input n_189;
input n_1147;
input n_1557;
input n_1610;
input n_13;
input n_1077;
input n_1422;
input n_540;
input n_618;
input n_896;
input n_323;
input n_195;
input n_356;
input n_894;
input n_831;
input n_964;
input n_1373;
input n_1350;
input n_1511;
input n_1470;
input n_1096;
input n_234;
input n_1575;
input n_833;
input n_5;
input n_225;
input n_1307;
input n_988;
input n_814;
input n_192;
input n_1549;
input n_1201;
input n_1114;
input n_655;
input n_1616;
input n_1446;
input n_669;
input n_472;
input n_1458;
input n_1176;
input n_1472;
input n_387;
input n_1149;
input n_398;
input n_635;
input n_763;
input n_1020;
input n_1062;
input n_211;
input n_1219;
input n_3;
input n_1204;
input n_178;
input n_1035;
input n_287;
input n_555;
input n_783;
input n_1188;
input n_661;
input n_41;
input n_849;
input n_15;
input n_336;
input n_584;
input n_681;
input n_50;
input n_430;
input n_510;
input n_216;
input n_311;
input n_830;
input n_1296;
input n_1413;
input n_801;
input n_241;
input n_875;
input n_357;
input n_1110;
input n_445;
input n_749;
input n_1134;
input n_1358;
input n_717;
input n_165;
input n_939;
input n_482;
input n_1088;
input n_588;
input n_1173;
input n_789;
input n_1232;
input n_1603;
input n_734;
input n_638;
input n_866;
input n_107;
input n_969;
input n_1401;
input n_1019;
input n_1105;
input n_249;
input n_304;
input n_1338;
input n_577;
input n_1522;
input n_1419;
input n_338;
input n_149;
input n_693;
input n_1506;
input n_14;
input n_836;
input n_990;
input n_1389;
input n_975;
input n_1256;
input n_567;
input n_1465;
input n_778;
input n_1122;
input n_151;
input n_306;
input n_458;
input n_770;
input n_1375;
input n_1102;
input n_711;
input n_1499;
input n_85;
input n_1187;
input n_1441;
input n_1392;
input n_1597;
input n_1164;
input n_489;
input n_1174;
input n_1371;
input n_617;
input n_1303;
input n_1572;
input n_876;
input n_1516;
input n_1190;
input n_118;
input n_601;
input n_917;
input n_966;
input n_253;
input n_1116;
input n_1212;
input n_1541;
input n_172;
input n_206;
input n_217;
input n_726;
input n_982;
input n_1573;
input n_1453;
input n_818;
input n_861;
input n_1183;
input n_899;
input n_1253;
input n_210;
input n_774;
input n_1628;
input n_1335;
input n_1514;
input n_1059;
input n_1345;
input n_176;
input n_1133;
input n_557;
input n_1410;
input n_1005;
input n_607;
input n_1003;
input n_679;
input n_710;
input n_527;
input n_1168;
input n_707;
input n_937;
input n_1427;
input n_393;
input n_108;
input n_487;
input n_1584;
input n_665;
input n_66;
input n_1440;
input n_177;
input n_421;
input n_1356;
input n_910;
input n_768;
input n_1475;
input n_1302;
input n_205;
input n_1136;
input n_1313;
input n_1491;
input n_754;
input n_1496;
input n_179;
input n_1125;
input n_125;
input n_410;
input n_708;
input n_529;
input n_735;
input n_232;
input n_1109;
input n_126;
input n_895;
input n_1310;
input n_202;
input n_427;
input n_1399;
input n_1543;
input n_791;
input n_732;
input n_1533;
input n_193;
input n_808;
input n_797;
input n_1025;
input n_500;
input n_1067;
input n_148;
input n_435;
input n_159;
input n_766;
input n_1457;
input n_541;
input n_538;
input n_1117;
input n_799;
input n_687;
input n_715;
input n_1480;
input n_1482;
input n_1213;
input n_1266;
input n_536;
input n_872;
input n_594;
input n_200;
input n_1291;
input n_1297;
input n_1155;
input n_1418;
input n_89;
input n_1524;
input n_1485;
input n_115;
input n_1011;
input n_1184;
input n_985;
input n_869;
input n_810;
input n_416;
input n_827;
input n_401;
input n_1352;
input n_626;
input n_1144;
input n_1137;
input n_1570;
input n_1170;
input n_305;
input n_137;
input n_676;
input n_294;
input n_318;
input n_653;
input n_642;
input n_1602;
input n_194;
input n_855;
input n_1178;
input n_1461;
input n_850;
input n_684;
input n_124;
input n_268;
input n_664;
input n_503;
input n_235;
input n_1372;
input n_605;
input n_1273;
input n_353;
input n_620;
input n_643;
input n_916;
input n_1081;
input n_493;
input n_1235;
input n_703;
input n_698;
input n_980;
input n_1115;
input n_1282;
input n_1318;
input n_780;
input n_998;
input n_1454;
input n_467;
input n_1227;
input n_1531;
input n_840;
input n_1334;
input n_501;
input n_823;
input n_245;
input n_725;
input n_1388;
input n_1417;
input n_1295;
input n_672;
input n_581;
input n_382;
input n_554;
input n_1625;
input n_898;
input n_1013;
input n_1452;
input n_718;
input n_265;
input n_1120;
input n_719;
input n_443;
input n_198;
input n_714;
input n_909;
input n_1497;
input n_1530;
input n_997;
input n_932;
input n_612;
input n_1409;
input n_788;
input n_1326;
input n_119;
input n_1268;
input n_559;
input n_825;
input n_508;
input n_506;
input n_1320;
input n_737;
input n_986;
input n_509;
input n_1317;
input n_147;
input n_1518;
input n_1281;
input n_67;
input n_1192;
input n_1024;
input n_1063;
input n_209;
input n_1564;
input n_1613;
input n_733;
input n_1489;
input n_1376;
input n_941;
input n_981;
input n_1569;
input n_68;
input n_867;
input n_186;
input n_134;
input n_587;
input n_63;
input n_792;
input n_756;
input n_1429;
input n_399;
input n_1238;
input n_548;
input n_812;
input n_298;
input n_518;
input n_505;
input n_282;
input n_752;
input n_905;
input n_1476;
input n_1108;
input n_782;
input n_1100;
input n_1395;
input n_862;
input n_1425;
input n_760;
input n_1620;
input n_381;
input n_220;
input n_390;
input n_1330;
input n_31;
input n_481;
input n_1554;
input n_769;
input n_42;
input n_1046;
input n_271;
input n_934;
input n_1618;
input n_826;
input n_886;
input n_1221;
input n_654;
input n_1172;
input n_167;
input n_379;
input n_428;
input n_1341;
input n_570;
input n_1361;
input n_853;
input n_377;
input n_751;
input n_786;
input n_1083;
input n_1142;
input n_1129;
input n_392;
input n_158;
input n_704;
input n_787;
input n_138;
input n_961;
input n_771;
input n_276;
input n_95;
input n_1225;
input n_1520;
input n_169;
input n_522;
input n_1287;
input n_1262;
input n_400;
input n_930;
input n_181;
input n_1411;
input n_221;
input n_622;
input n_1577;
input n_1087;
input n_386;
input n_994;
input n_848;
input n_1550;
input n_1498;
input n_1223;
input n_1272;
input n_104;
input n_682;
input n_1567;
input n_56;
input n_141;
input n_1247;
input n_922;
input n_816;
input n_591;
input n_145;
input n_1536;
input n_1344;
input n_313;
input n_631;
input n_479;
input n_1246;
input n_1339;
input n_1478;
input n_432;
input n_839;
input n_1210;
input n_1364;
input n_328;
input n_140;
input n_1250;
input n_369;
input n_871;
input n_598;
input n_685;
input n_928;
input n_608;
input n_1367;
input n_78;
input n_1460;
input n_772;
input n_1555;
input n_499;
input n_1589;
input n_517;
input n_98;
input n_402;
input n_413;
input n_1086;
input n_796;
input n_1619;
input n_236;
input n_1502;
input n_1469;
input n_1012;
input n_1;
input n_1396;
input n_1348;
input n_903;
input n_1525;
input n_740;
input n_203;
input n_384;
input n_1404;
input n_80;
input n_35;
input n_1315;
input n_277;
input n_1061;
input n_92;
input n_333;
input n_1298;
input n_462;
input n_1193;
input n_1255;
input n_258;
input n_1113;
input n_29;
input n_79;
input n_1226;
input n_722;
input n_1277;
input n_188;
input n_844;
input n_201;
input n_471;
input n_852;
input n_1487;
input n_40;
input n_1028;
input n_1601;
input n_781;
input n_474;
input n_542;
input n_463;
input n_1546;
input n_595;
input n_502;
input n_466;
input n_420;
input n_1337;
input n_1495;
input n_632;
input n_699;
input n_979;
input n_1515;
input n_1627;
input n_1245;
input n_846;
input n_465;
input n_76;
input n_362;
input n_1321;
input n_170;
input n_27;
input n_161;
input n_273;
input n_585;
input n_270;
input n_616;
input n_81;
input n_745;
input n_1103;
input n_648;
input n_1379;
input n_312;
input n_1076;
input n_1091;
input n_1408;
input n_494;
input n_641;
input n_730;
input n_1325;
input n_1595;
input n_354;
input n_575;
input n_480;
input n_425;
input n_795;
input n_695;
input n_180;
input n_656;
input n_1606;
input n_1220;
input n_37;
input n_1540;
input n_229;
input n_437;
input n_60;
input n_403;
input n_453;
input n_1130;
input n_720;
input n_0;
input n_1526;
input n_863;
input n_805;
input n_1604;
input n_1275;
input n_113;
input n_712;
input n_246;
input n_1583;
input n_1042;
input n_1402;
input n_269;
input n_285;
input n_412;
input n_1493;
input n_657;
input n_644;
input n_1160;
input n_1397;
input n_491;
input n_1258;
input n_1074;
input n_1621;
input n_251;
input n_160;
input n_566;
input n_565;
input n_1448;
input n_1507;
input n_1398;
input n_597;
input n_1181;
input n_1505;
input n_1196;
input n_651;
input n_1340;
input n_334;
input n_811;
input n_1558;
input n_807;
input n_835;
input n_175;
input n_666;
input n_262;
input n_1433;
input n_99;
input n_1254;
input n_1026;
input n_1234;
input n_319;
input n_364;
input n_1138;
input n_927;
input n_20;
input n_1089;
input n_1004;
input n_1186;
input n_1032;
input n_242;
input n_1018;
input n_438;
input n_713;
input n_904;
input n_1588;
input n_1622;
input n_166;
input n_1180;
input n_1271;
input n_533;
input n_1542;
input n_1251;
input n_278;

output n_5639;

wire n_2253;
wire n_2417;
wire n_2756;
wire n_4706;
wire n_5567;
wire n_2380;
wire n_3241;
wire n_3006;
wire n_5287;
wire n_2327;
wire n_2899;
wire n_5484;
wire n_3619;
wire n_3541;
wire n_3622;
wire n_2395;
wire n_5161;
wire n_5512;
wire n_5207;
wire n_2347;
wire n_4963;
wire n_4240;
wire n_4508;
wire n_2021;
wire n_2391;
wire n_5035;
wire n_5282;
wire n_1960;
wire n_2843;
wire n_3615;
wire n_2059;
wire n_2487;
wire n_1695;
wire n_3202;
wire n_4977;
wire n_3813;
wire n_3341;
wire n_3587;
wire n_4128;
wire n_3445;
wire n_2001;
wire n_4145;
wire n_3785;
wire n_5033;
wire n_4211;
wire n_3448;
wire n_3019;
wire n_2096;
wire n_3776;
wire n_2530;
wire n_4517;
wire n_2483;
wire n_1696;
wire n_4425;
wire n_4950;
wire n_4988;
wire n_1860;
wire n_4615;
wire n_1728;
wire n_2076;
wire n_5480;
wire n_2147;
wire n_3010;
wire n_2770;
wire n_4131;
wire n_5402;
wire n_2584;
wire n_3188;
wire n_5509;
wire n_3403;
wire n_3624;
wire n_3461;
wire n_3082;
wire n_2189;
wire n_3796;
wire n_5154;
wire n_3283;
wire n_5469;
wire n_2323;
wire n_2597;
wire n_3340;
wire n_3277;
wire n_5453;
wire n_2052;
wire n_4499;
wire n_4927;
wire n_5202;
wire n_3214;
wire n_2091;
wire n_4311;
wire n_3631;
wire n_3806;
wire n_4691;
wire n_4678;
wire n_2032;
wire n_2587;
wire n_5406;
wire n_3947;
wire n_3490;
wire n_1948;
wire n_3868;
wire n_3183;
wire n_3437;
wire n_3353;
wire n_4203;
wire n_3687;
wire n_5241;
wire n_2384;
wire n_3156;
wire n_3376;
wire n_5037;
wire n_4468;
wire n_3653;
wire n_5562;
wire n_3702;
wire n_4976;
wire n_2202;
wire n_2648;
wire n_5008;
wire n_2159;
wire n_2976;
wire n_3876;
wire n_2353;
wire n_2439;
wire n_4811;
wire n_5398;
wire n_2276;
wire n_2089;
wire n_3420;
wire n_5144;
wire n_3361;
wire n_4758;
wire n_4255;
wire n_1796;
wire n_5577;
wire n_4484;
wire n_3668;
wire n_4237;
wire n_2934;
wire n_1672;
wire n_1880;
wire n_3550;
wire n_2079;
wire n_2238;
wire n_1706;
wire n_3418;
wire n_4901;
wire n_2859;
wire n_3395;
wire n_4917;
wire n_2863;
wire n_2072;
wire n_2738;
wire n_2968;
wire n_2684;
wire n_3593;
wire n_5343;
wire n_4421;
wire n_4836;
wire n_5062;
wire n_4020;
wire n_2730;
wire n_2251;
wire n_3915;
wire n_4469;
wire n_4414;
wire n_5184;
wire n_4532;
wire n_3339;
wire n_3349;
wire n_3735;
wire n_2248;
wire n_3007;
wire n_2622;
wire n_2062;
wire n_2668;
wire n_5463;
wire n_2100;
wire n_5236;
wire n_3310;
wire n_3487;
wire n_2258;
wire n_1667;
wire n_3983;
wire n_4405;
wire n_5433;
wire n_1926;
wire n_4195;
wire n_4969;
wire n_4504;
wire n_2776;
wire n_4408;
wire n_2140;
wire n_2385;
wire n_1819;
wire n_4531;
wire n_2987;
wire n_4567;
wire n_4164;
wire n_5315;
wire n_4234;
wire n_4130;
wire n_3611;
wire n_2862;
wire n_5348;
wire n_2175;
wire n_5055;
wire n_2324;
wire n_2606;
wire n_3187;
wire n_2828;
wire n_5397;
wire n_4471;
wire n_5031;
wire n_3392;
wire n_3975;
wire n_3430;
wire n_4444;
wire n_3208;
wire n_3331;
wire n_2379;
wire n_4983;
wire n_2911;
wire n_2154;
wire n_4916;
wire n_3649;
wire n_4302;
wire n_2514;
wire n_5189;
wire n_5381;
wire n_4786;
wire n_3257;
wire n_4160;
wire n_2293;
wire n_5516;
wire n_4051;
wire n_2028;
wire n_3009;
wire n_3981;
wire n_1841;
wire n_2581;
wire n_3224;
wire n_4647;
wire n_3752;
wire n_1711;
wire n_1891;
wire n_5254;
wire n_3526;
wire n_2546;
wire n_3790;
wire n_3491;
wire n_4613;
wire n_4649;
wire n_1888;
wire n_5615;
wire n_1963;
wire n_4795;
wire n_2226;
wire n_2891;
wire n_4028;
wire n_5479;
wire n_1690;
wire n_3819;
wire n_2449;
wire n_5083;
wire n_2297;
wire n_4186;
wire n_4731;
wire n_1759;
wire n_2177;
wire n_3747;
wire n_5592;
wire n_2227;
wire n_4618;
wire n_2190;
wire n_3346;
wire n_4742;
wire n_2876;
wire n_4099;
wire n_3484;
wire n_3620;
wire n_1746;
wire n_2479;
wire n_4295;
wire n_5303;
wire n_4694;
wire n_4533;
wire n_3038;
wire n_5081;
wire n_5124;
wire n_3068;
wire n_2871;
wire n_4244;
wire n_4603;
wire n_2943;
wire n_4254;
wire n_3143;
wire n_3168;
wire n_1680;
wire n_4697;
wire n_2607;
wire n_3994;
wire n_4190;
wire n_4810;
wire n_3317;
wire n_4391;
wire n_3263;
wire n_2582;
wire n_4157;
wire n_4283;
wire n_4681;
wire n_4638;
wire n_3455;
wire n_5047;
wire n_3452;
wire n_5346;
wire n_1994;
wire n_5517;
wire n_4707;
wire n_2577;
wire n_4527;
wire n_5109;
wire n_2796;
wire n_2342;
wire n_4156;
wire n_1851;
wire n_4848;
wire n_2937;
wire n_3095;
wire n_2805;
wire n_5624;
wire n_4918;
wire n_3856;
wire n_2914;
wire n_4898;
wire n_1964;
wire n_2869;
wire n_4002;
wire n_5010;
wire n_2406;
wire n_3623;
wire n_2846;
wire n_2925;
wire n_3773;
wire n_3918;
wire n_2398;
wire n_2857;
wire n_5358;
wire n_4528;
wire n_3932;
wire n_4619;
wire n_4673;
wire n_3516;
wire n_4822;
wire n_2155;
wire n_2516;
wire n_3797;
wire n_2947;
wire n_5580;
wire n_4299;
wire n_4801;
wire n_1665;
wire n_3515;
wire n_2886;
wire n_2093;
wire n_2473;
wire n_3287;
wire n_3378;
wire n_5435;
wire n_4279;
wire n_4769;
wire n_4632;
wire n_5373;
wire n_4294;
wire n_1732;
wire n_5279;
wire n_4125;
wire n_4232;
wire n_4949;
wire n_2941;
wire n_2457;
wire n_5493;
wire n_4790;
wire n_2536;
wire n_1758;
wire n_2952;
wire n_4847;
wire n_5321;
wire n_3058;
wire n_5096;
wire n_4365;
wire n_1878;
wire n_3505;
wire n_4610;
wire n_3730;
wire n_4489;
wire n_5210;
wire n_4967;
wire n_4992;
wire n_3001;
wire n_3945;
wire n_4542;
wire n_2729;
wire n_2261;
wire n_3597;
wire n_2897;
wire n_2077;
wire n_4198;
wire n_2909;
wire n_4534;
wire n_4500;
wire n_5014;
wire n_3185;
wire n_3523;
wire n_1785;
wire n_2829;
wire n_4597;
wire n_4329;
wire n_4087;
wire n_3811;
wire n_1664;
wire n_3200;
wire n_2231;
wire n_2017;
wire n_2604;
wire n_4257;
wire n_3453;
wire n_2390;
wire n_3213;
wire n_3077;
wire n_3474;
wire n_3984;
wire n_2151;
wire n_2106;
wire n_2716;
wire n_4665;
wire n_1913;
wire n_1823;
wire n_3679;
wire n_3422;
wire n_3888;
wire n_5638;
wire n_4189;
wire n_1875;
wire n_2803;
wire n_3707;
wire n_1846;
wire n_5584;
wire n_3429;
wire n_1903;
wire n_3849;
wire n_3946;
wire n_3229;
wire n_4463;
wire n_1805;
wire n_4687;
wire n_4670;
wire n_4084;
wire n_4703;
wire n_4037;
wire n_2922;
wire n_3275;
wire n_3499;
wire n_2645;
wire n_2727;
wire n_3421;
wire n_2240;
wire n_2436;
wire n_3618;
wire n_2593;
wire n_5262;
wire n_3683;
wire n_3642;
wire n_3286;
wire n_3808;
wire n_4763;
wire n_1684;
wire n_3590;
wire n_5310;
wire n_4594;
wire n_3424;
wire n_2301;
wire n_3583;
wire n_3560;
wire n_4076;
wire n_4714;
wire n_2419;
wire n_3215;
wire n_5146;
wire n_4776;
wire n_2122;
wire n_2512;
wire n_4102;
wire n_2786;
wire n_3171;
wire n_5213;
wire n_3020;
wire n_3677;
wire n_3462;
wire n_5441;
wire n_3468;
wire n_2910;
wire n_1893;
wire n_2163;
wire n_2254;
wire n_3546;
wire n_2647;
wire n_4443;
wire n_5461;
wire n_4507;
wire n_1811;
wire n_2443;
wire n_2624;
wire n_3012;
wire n_4575;
wire n_3244;
wire n_3130;
wire n_3822;
wire n_3569;
wire n_5629;
wire n_4452;
wire n_4348;
wire n_5634;
wire n_5430;
wire n_5362;
wire n_4355;
wire n_3494;
wire n_5050;
wire n_5063;
wire n_5229;
wire n_2125;
wire n_3771;
wire n_5199;
wire n_3110;
wire n_4572;
wire n_3073;
wire n_5527;
wire n_5609;
wire n_5416;
wire n_4026;
wire n_2265;
wire n_4104;
wire n_4512;
wire n_3554;
wire n_4377;
wire n_5266;
wire n_3178;
wire n_5355;
wire n_2334;
wire n_4521;
wire n_4488;
wire n_2289;
wire n_3051;
wire n_2783;
wire n_2263;
wire n_3750;
wire n_2341;
wire n_3632;
wire n_4588;
wire n_2733;
wire n_2785;
wire n_2415;
wire n_3299;
wire n_4519;
wire n_5551;
wire n_3715;
wire n_3040;
wire n_1938;
wire n_2499;
wire n_3568;
wire n_5475;
wire n_3737;
wire n_1967;
wire n_3255;
wire n_4856;
wire n_2997;
wire n_4400;
wire n_5168;
wire n_3326;
wire n_3734;
wire n_4778;
wire n_2429;
wire n_5322;
wire n_1793;
wire n_4352;
wire n_4441;
wire n_4761;
wire n_1804;
wire n_4347;
wire n_4095;
wire n_3196;
wire n_4593;
wire n_2533;
wire n_2364;
wire n_3492;
wire n_2780;
wire n_4727;
wire n_4568;
wire n_5371;
wire n_2291;
wire n_4043;
wire n_1636;
wire n_3601;
wire n_5418;
wire n_1865;
wire n_2973;
wire n_2094;
wire n_2393;
wire n_1697;
wire n_5316;
wire n_3831;
wire n_3801;
wire n_2043;
wire n_2751;
wire n_4893;
wire n_5032;
wire n_1934;
wire n_4948;
wire n_4000;
wire n_3240;
wire n_2025;
wire n_4406;
wire n_2758;
wire n_1807;
wire n_2618;
wire n_5112;
wire n_5386;
wire n_2559;
wire n_4748;
wire n_2295;
wire n_3931;
wire n_4010;
wire n_2840;
wire n_5017;
wire n_1814;
wire n_2822;
wire n_4710;
wire n_4607;
wire n_5123;
wire n_4117;
wire n_3636;
wire n_1722;
wire n_2441;
wire n_1802;
wire n_3083;
wire n_4487;
wire n_5001;
wire n_2795;
wire n_2981;
wire n_2282;
wire n_2800;
wire n_4817;
wire n_3380;
wire n_2098;
wire n_3460;
wire n_3409;
wire n_3538;
wire n_2068;
wire n_4849;
wire n_4867;
wire n_5424;
wire n_2641;
wire n_3198;
wire n_1895;
wire n_4728;
wire n_4247;
wire n_4933;
wire n_4018;
wire n_3900;
wire n_4902;
wire n_4518;
wire n_4409;
wire n_4411;
wire n_3872;
wire n_4336;
wire n_2270;
wire n_4777;
wire n_2653;
wire n_2496;
wire n_1908;
wire n_2259;
wire n_3877;
wire n_2995;
wire n_5496;
wire n_2494;
wire n_3547;
wire n_3977;
wire n_4052;
wire n_3459;
wire n_4398;
wire n_3155;
wire n_2633;
wire n_4954;
wire n_2435;
wire n_2097;
wire n_5460;
wire n_4304;
wire n_3911;
wire n_5333;
wire n_4431;
wire n_4192;
wire n_5570;
wire n_3736;
wire n_4805;
wire n_4885;
wire n_1661;
wire n_3565;
wire n_4701;
wire n_2575;
wire n_5040;
wire n_1658;
wire n_1904;
wire n_1899;
wire n_2067;
wire n_2219;
wire n_3533;
wire n_2877;
wire n_2148;
wire n_1726;
wire n_4631;
wire n_3035;
wire n_5194;
wire n_5464;
wire n_1657;
wire n_1725;
wire n_3639;
wire n_2501;
wire n_3079;
wire n_4965;
wire n_1915;
wire n_5610;
wire n_5239;
wire n_2605;
wire n_4747;
wire n_5197;
wire n_1979;
wire n_2924;
wire n_4111;
wire n_2484;
wire n_4587;
wire n_3731;
wire n_2946;
wire n_5305;
wire n_4538;
wire n_2754;
wire n_1742;
wire n_5376;
wire n_2489;
wire n_5204;
wire n_2012;
wire n_4094;
wire n_3503;
wire n_2866;
wire n_3561;
wire n_2917;
wire n_2425;
wire n_3536;
wire n_3661;
wire n_4150;
wire n_4878;
wire n_1703;
wire n_1650;
wire n_3934;
wire n_4985;
wire n_3922;
wire n_3846;
wire n_2103;
wire n_2160;
wire n_2498;
wire n_2697;
wire n_3074;
wire n_1999;
wire n_2372;
wire n_3673;
wire n_3768;
wire n_2861;
wire n_2630;
wire n_3943;
wire n_2430;
wire n_2433;
wire n_3293;
wire n_5508;
wire n_5582;
wire n_4022;
wire n_4852;
wire n_2528;
wire n_4869;
wire n_4700;
wire n_4035;
wire n_2316;
wire n_1898;
wire n_3294;
wire n_4426;
wire n_3415;
wire n_2284;
wire n_2817;
wire n_3139;
wire n_5292;
wire n_2598;
wire n_4601;
wire n_2687;
wire n_1890;
wire n_4220;
wire n_1944;
wire n_5630;
wire n_3431;
wire n_3169;
wire n_3151;
wire n_2078;
wire n_3284;
wire n_3070;
wire n_4066;
wire n_2884;
wire n_4515;
wire n_4351;
wire n_5264;
wire n_3126;
wire n_4403;
wire n_1981;
wire n_1663;
wire n_1718;
wire n_4509;
wire n_4858;
wire n_3700;
wire n_5504;
wire n_4223;
wire n_1889;
wire n_5025;
wire n_2966;
wire n_2326;
wire n_2188;
wire n_4644;
wire n_4456;
wire n_5060;
wire n_5334;
wire n_2448;
wire n_4346;
wire n_3170;
wire n_2748;
wire n_3311;
wire n_3272;
wire n_2898;
wire n_2717;
wire n_1861;
wire n_5581;
wire n_3691;
wire n_3628;
wire n_4235;
wire n_1867;
wire n_1945;
wire n_3018;
wire n_2573;
wire n_4435;
wire n_2939;
wire n_3807;
wire n_2447;
wire n_4764;
wire n_5394;
wire n_2774;
wire n_1707;
wire n_4655;
wire n_3161;
wire n_4581;
wire n_4827;
wire n_2488;
wire n_3477;
wire n_5421;
wire n_2476;
wire n_4399;
wire n_2781;
wire n_5309;
wire n_2778;
wire n_4782;
wire n_4363;
wire n_2887;
wire n_4864;
wire n_2691;
wire n_3054;
wire n_4335;
wire n_2526;
wire n_2703;
wire n_2167;
wire n_5428;
wire n_3391;
wire n_4259;
wire n_5541;
wire n_2709;
wire n_5543;
wire n_4865;
wire n_4056;
wire n_4564;
wire n_3840;
wire n_5085;
wire n_3518;
wire n_2956;
wire n_3733;
wire n_2173;
wire n_1842;
wire n_3738;
wire n_5116;
wire n_3464;
wire n_2018;
wire n_4526;
wire n_3245;
wire n_4417;
wire n_4899;
wire n_2119;
wire n_2552;
wire n_2157;
wire n_5411;
wire n_2453;
wire n_4798;
wire n_3509;
wire n_3352;
wire n_3076;
wire n_3535;
wire n_2182;
wire n_3251;
wire n_2931;
wire n_5185;
wire n_3118;
wire n_3511;
wire n_3443;
wire n_2146;
wire n_3644;
wire n_5076;
wire n_3336;
wire n_3935;
wire n_3521;
wire n_5379;
wire n_3562;
wire n_3948;
wire n_4750;
wire n_2918;
wire n_3232;
wire n_1673;
wire n_2112;
wire n_1739;
wire n_2958;
wire n_4981;
wire n_3114;
wire n_3125;
wire n_2394;
wire n_3612;
wire n_2954;
wire n_4835;
wire n_4430;
wire n_5565;
wire n_4081;
wire n_3132;
wire n_4407;
wire n_3951;
wire n_4894;
wire n_3238;
wire n_3210;
wire n_2036;
wire n_3267;
wire n_4995;
wire n_5524;
wire n_3964;
wire n_3772;
wire n_1956;
wire n_1642;
wire n_2279;
wire n_3373;
wire n_4446;
wire n_3884;
wire n_3726;
wire n_2525;
wire n_2892;
wire n_2907;
wire n_3577;
wire n_2820;
wire n_2049;
wire n_2273;
wire n_2719;
wire n_1741;
wire n_4057;
wire n_4332;
wire n_4314;
wire n_3347;
wire n_3216;
wire n_3809;
wire n_2113;
wire n_4288;
wire n_3567;
wire n_5066;
wire n_1634;
wire n_3939;
wire n_5401;
wire n_4241;
wire n_3321;
wire n_3212;
wire n_2256;
wire n_3152;
wire n_5106;
wire n_5468;
wire n_2920;
wire n_4265;
wire n_5319;
wire n_2247;
wire n_3705;
wire n_2802;
wire n_4705;
wire n_3159;
wire n_5455;
wire n_2268;
wire n_3778;
wire n_5337;
wire n_3304;
wire n_3912;
wire n_1729;
wire n_2739;
wire n_2771;
wire n_4604;
wire n_5223;
wire n_3795;
wire n_5020;
wire n_4419;
wire n_4477;
wire n_3179;
wire n_3256;
wire n_2386;
wire n_3086;
wire n_2369;
wire n_2927;
wire n_4217;
wire n_4395;
wire n_2821;
wire n_5074;
wire n_2568;
wire n_5364;
wire n_1738;
wire n_3728;
wire n_3064;
wire n_3088;
wire n_4639;
wire n_3713;
wire n_3663;
wire n_5046;
wire n_5166;
wire n_3246;
wire n_2495;
wire n_1789;
wire n_5088;
wire n_2302;
wire n_5457;
wire n_5532;
wire n_2069;
wire n_3434;
wire n_1806;
wire n_4227;
wire n_4033;
wire n_4289;
wire n_2024;
wire n_4780;
wire n_4243;
wire n_4982;
wire n_3695;
wire n_4330;
wire n_2482;
wire n_2677;
wire n_5544;
wire n_3832;
wire n_3987;
wire n_5352;
wire n_4991;
wire n_5538;
wire n_1698;
wire n_2329;
wire n_2142;
wire n_5410;
wire n_3332;
wire n_3048;
wire n_3937;
wire n_2203;
wire n_4525;
wire n_3782;
wire n_2978;
wire n_2058;
wire n_2458;
wire n_4208;
wire n_3786;
wire n_2888;
wire n_3638;
wire n_5503;
wire n_1633;
wire n_4177;
wire n_3763;
wire n_2669;
wire n_1778;
wire n_2306;
wire n_3022;
wire n_4264;
wire n_3087;
wire n_3489;
wire n_2566;
wire n_5129;
wire n_2149;
wire n_5500;
wire n_3060;
wire n_4276;
wire n_5219;
wire n_5605;
wire n_3013;
wire n_1984;
wire n_5170;
wire n_2408;
wire n_5320;
wire n_1877;
wire n_3049;
wire n_1723;
wire n_5107;
wire n_4485;
wire n_4626;
wire n_2659;
wire n_4975;
wire n_1852;
wire n_5602;
wire n_3089;
wire n_2470;
wire n_5405;
wire n_3985;
wire n_5253;
wire n_4760;
wire n_4652;
wire n_4624;
wire n_2551;
wire n_2682;
wire n_3440;
wire n_1748;
wire n_4569;
wire n_2699;
wire n_4897;
wire n_2769;
wire n_3542;
wire n_3436;
wire n_5491;
wire n_2615;
wire n_3940;
wire n_2985;
wire n_5636;
wire n_5065;
wire n_2753;
wire n_3637;
wire n_2842;
wire n_4523;
wire n_1836;
wire n_2868;
wire n_5492;
wire n_3141;
wire n_5084;
wire n_3164;
wire n_3570;
wire n_5260;
wire n_4919;
wire n_4025;
wire n_2712;
wire n_5328;
wire n_3936;
wire n_4503;
wire n_3507;
wire n_3821;
wire n_2700;
wire n_3367;
wire n_4464;
wire n_3096;
wire n_3496;
wire n_4114;
wire n_2544;
wire n_2356;
wire n_4556;
wire n_5454;
wire n_2620;
wire n_4089;
wire n_5621;
wire n_2919;
wire n_4327;
wire n_4218;
wire n_2150;
wire n_3146;
wire n_5165;
wire n_2241;
wire n_2757;
wire n_5573;
wire n_4353;
wire n_2042;
wire n_1754;
wire n_2921;
wire n_2720;
wire n_1854;
wire n_4990;
wire n_5529;
wire n_1856;
wire n_4959;
wire n_4161;
wire n_3992;
wire n_2616;
wire n_1906;
wire n_4103;
wire n_4466;
wire n_2262;
wire n_2462;
wire n_3625;
wire n_2798;
wire n_2945;
wire n_2331;
wire n_2837;
wire n_4844;
wire n_2979;
wire n_5257;
wire n_3655;
wire n_4688;
wire n_4765;
wire n_2548;
wire n_5180;
wire n_2108;
wire n_3640;
wire n_4388;
wire n_4206;
wire n_1779;
wire n_4738;
wire n_3909;
wire n_3207;
wire n_3944;
wire n_4434;
wire n_4837;
wire n_3042;
wire n_1942;
wire n_2510;
wire n_4219;
wire n_2804;
wire n_3659;
wire n_2120;
wire n_5012;
wire n_1876;
wire n_4620;
wire n_1810;
wire n_2813;
wire n_4438;
wire n_2009;
wire n_2222;
wire n_3510;
wire n_3218;
wire n_2667;
wire n_3150;
wire n_4325;
wire n_1733;
wire n_2413;
wire n_3775;
wire n_4133;
wire n_4184;
wire n_5203;
wire n_2518;
wire n_2629;
wire n_4481;
wire n_3416;
wire n_4379;
wire n_2181;
wire n_1829;
wire n_4030;
wire n_4490;
wire n_3138;
wire n_4397;
wire n_1710;
wire n_2928;
wire n_1734;
wire n_4820;
wire n_3770;
wire n_5094;
wire n_4938;
wire n_4179;
wire n_3469;
wire n_5336;
wire n_2723;
wire n_3220;
wire n_4641;
wire n_2539;
wire n_5548;
wire n_5601;
wire n_3855;
wire n_2054;
wire n_5339;
wire n_4931;
wire n_1765;
wire n_3158;
wire n_1744;
wire n_2623;
wire n_3113;
wire n_2718;
wire n_3760;
wire n_4078;
wire n_1760;
wire n_2856;
wire n_1832;
wire n_4146;
wire n_4360;
wire n_3666;
wire n_3828;
wire n_3288;
wire n_5514;
wire n_4404;
wire n_5091;
wire n_1874;
wire n_4787;
wire n_2060;
wire n_2613;
wire n_1987;
wire n_3667;
wire n_5486;
wire n_3703;
wire n_4903;
wire n_3558;
wire n_2545;
wire n_2787;
wire n_5599;
wire n_4356;
wire n_2061;
wire n_4432;
wire n_5251;
wire n_2378;
wire n_1740;
wire n_4291;
wire n_5403;
wire n_4386;
wire n_4149;
wire n_1692;
wire n_2982;
wire n_2481;
wire n_3545;
wire n_2507;
wire n_4019;
wire n_2900;
wire n_2339;
wire n_4637;
wire n_4935;
wire n_4785;
wire n_3426;
wire n_3454;
wire n_3820;
wire n_5608;
wire n_3741;
wire n_3410;
wire n_2029;
wire n_5298;
wire n_5596;
wire n_1887;
wire n_4413;
wire n_2346;
wire n_3990;
wire n_4493;
wire n_3475;
wire n_2882;
wire n_1721;
wire n_2338;
wire n_3672;
wire n_5290;
wire n_3197;
wire n_3109;
wire n_2721;
wire n_5095;
wire n_3002;
wire n_5324;
wire n_3897;
wire n_3845;
wire n_2081;
wire n_4570;
wire n_2156;
wire n_5101;
wire n_4296;
wire n_1820;
wire n_5019;
wire n_2418;
wire n_5589;
wire n_2179;
wire n_1724;
wire n_2521;
wire n_3458;
wire n_3330;
wire n_4606;
wire n_4774;
wire n_2477;
wire n_3887;
wire n_4093;
wire n_4672;
wire n_3519;
wire n_4174;
wire n_3374;
wire n_3045;
wire n_2367;
wire n_1870;
wire n_4766;
wire n_5633;
wire n_2896;
wire n_4074;
wire n_4600;
wire n_1927;
wire n_5583;
wire n_4460;
wire n_3645;
wire n_3223;
wire n_3929;
wire n_2255;
wire n_2272;
wire n_1965;
wire n_1902;
wire n_1941;
wire n_5501;
wire n_3938;
wire n_5377;
wire n_2878;
wire n_3498;
wire n_2015;
wire n_1982;
wire n_4110;
wire n_3189;
wire n_2066;
wire n_3154;
wire n_2905;
wire n_3965;
wire n_3566;
wire n_2220;
wire n_4349;
wire n_3788;
wire n_2410;
wire n_4313;
wire n_1935;
wire n_3366;
wire n_2696;
wire n_4863;
wire n_3242;
wire n_3525;
wire n_3486;
wire n_2405;
wire n_3995;
wire n_2953;
wire n_2088;
wire n_4036;
wire n_5100;
wire n_1795;
wire n_2578;
wire n_3483;
wire n_1821;
wire n_3894;
wire n_3478;
wire n_4015;
wire n_3890;
wire n_2740;
wire n_5367;
wire n_2656;
wire n_3524;
wire n_5616;
wire n_5034;
wire n_1708;
wire n_3549;
wire n_1691;
wire n_2092;
wire n_2075;
wire n_3658;
wire n_1776;
wire n_4807;
wire n_2281;
wire n_2131;
wire n_3026;
wire n_1757;
wire n_1919;
wire n_4230;
wire n_3419;
wire n_2053;
wire n_1958;
wire n_3784;
wire n_2969;
wire n_3941;
wire n_2864;
wire n_3195;
wire n_3190;
wire n_3678;
wire n_2664;
wire n_3456;
wire n_5628;
wire n_1808;
wire n_2266;
wire n_2650;
wire n_4428;
wire n_5003;
wire n_5252;
wire n_2731;
wire n_5614;
wire n_5134;
wire n_3953;
wire n_3166;
wire n_4122;
wire n_3976;
wire n_3979;
wire n_4582;
wire n_2998;
wire n_4684;
wire n_4840;
wire n_3162;
wire n_2760;
wire n_3377;
wire n_3749;
wire n_3962;
wire n_1826;
wire n_2304;
wire n_5325;
wire n_2637;
wire n_5375;
wire n_4384;
wire n_4423;
wire n_4096;
wire n_2881;
wire n_3282;
wire n_1763;
wire n_3231;
wire n_1966;
wire n_4996;
wire n_2475;
wire n_4598;
wire n_5064;
wire n_4478;
wire n_2646;
wire n_5536;
wire n_5173;
wire n_3920;
wire n_4890;
wire n_5027;
wire n_3203;
wire n_3866;
wire n_2903;
wire n_3921;
wire n_4106;
wire n_3717;
wire n_2743;
wire n_2675;
wire n_3052;
wire n_5215;
wire n_3743;
wire n_1932;
wire n_4721;
wire n_5597;
wire n_5635;
wire n_1983;
wire n_4029;
wire n_3870;
wire n_4496;
wire n_3529;
wire n_1977;
wire n_2153;
wire n_4338;
wire n_3094;
wire n_2310;
wire n_3952;
wire n_2287;
wire n_2860;
wire n_2056;
wire n_2318;
wire n_1735;
wire n_2502;
wire n_2504;
wire n_4495;
wire n_4762;
wire n_2974;
wire n_2901;
wire n_1940;
wire n_2793;
wire n_3442;
wire n_3998;
wire n_2285;
wire n_3147;
wire n_4141;
wire n_5121;
wire n_1824;
wire n_1917;
wire n_3386;
wire n_4107;
wire n_4667;
wire n_2325;
wire n_5555;
wire n_3488;
wire n_2446;
wire n_4547;
wire n_2893;
wire n_2588;
wire n_2962;
wire n_4004;
wire n_5576;
wire n_4668;
wire n_4953;
wire n_5466;
wire n_3898;
wire n_1786;
wire n_5284;
wire n_4997;
wire n_5308;
wire n_4274;
wire n_2627;
wire n_4759;
wire n_4467;
wire n_2080;
wire n_2377;
wire n_2340;
wire n_3552;
wire n_3684;
wire n_4735;
wire n_3137;
wire n_5578;
wire n_2361;
wire n_4113;
wire n_1998;
wire n_4686;
wire n_5530;
wire n_3759;
wire n_4321;
wire n_4342;
wire n_2034;
wire n_3933;
wire n_3206;
wire n_5506;
wire n_3966;
wire n_5243;
wire n_5449;
wire n_1702;
wire n_5221;
wire n_4183;
wire n_4068;
wire n_4872;
wire n_4233;
wire n_3192;
wire n_3764;
wire n_4709;
wire n_5038;
wire n_5311;
wire n_2649;
wire n_1929;
wire n_5575;
wire n_2807;
wire n_2542;
wire n_2313;
wire n_3324;
wire n_3914;
wire n_4625;
wire n_2558;
wire n_2063;
wire n_3803;
wire n_3742;
wire n_2252;
wire n_4819;
wire n_1685;
wire n_1714;
wire n_2576;
wire n_4900;
wire n_3390;
wire n_3746;
wire n_2373;
wire n_1713;
wire n_3817;
wire n_2745;
wire n_1737;
wire n_2493;
wire n_4930;
wire n_5276;
wire n_5078;
wire n_4537;
wire n_2885;
wire n_5011;
wire n_3318;
wire n_4070;
wire n_4282;
wire n_3485;
wire n_4180;
wire n_3839;
wire n_5205;
wire n_3333;
wire n_2845;
wire n_4143;
wire n_4659;
wire n_2602;
wire n_4579;
wire n_4616;
wire n_3014;
wire n_2547;
wire n_5023;
wire n_1812;
wire n_4105;
wire n_2532;
wire n_3791;
wire n_2665;
wire n_5351;
wire n_3905;
wire n_3368;
wire n_3530;
wire n_1930;
wire n_1955;
wire n_2765;
wire n_3329;
wire n_2994;
wire n_2401;
wire n_3135;
wire n_5476;
wire n_2003;
wire n_5446;
wire n_4895;
wire n_3573;
wire n_3148;
wire n_2264;
wire n_3534;
wire n_4275;
wire n_3970;
wire n_3438;
wire n_4098;
wire n_4789;
wire n_1972;
wire n_2806;
wire n_2184;
wire n_5312;
wire n_3217;
wire n_3404;
wire n_3425;
wire n_5111;
wire n_4055;
wire n_2926;
wire n_3540;
wire n_3670;
wire n_3973;
wire n_2023;
wire n_3249;
wire n_2351;
wire n_5113;
wire n_4442;
wire n_4698;
wire n_4779;
wire n_2286;
wire n_4966;
wire n_2065;
wire n_4017;
wire n_3397;
wire n_3740;
wire n_4418;
wire n_2549;
wire n_2705;
wire n_2332;
wire n_2977;
wire n_3723;
wire n_3600;
wire n_4134;
wire n_2836;
wire n_2130;
wire n_5167;
wire n_3239;
wire n_5117;
wire n_2773;
wire n_3365;
wire n_3476;
wire n_3686;
wire n_4913;
wire n_5612;
wire n_1791;
wire n_2850;
wire n_1747;
wire n_4251;
wire n_1817;
wire n_3982;
wire n_2654;
wire n_4621;
wire n_3176;
wire n_4559;
wire n_2186;
wire n_4368;
wire n_4740;
wire n_5301;
wire n_5007;
wire n_3581;
wire n_2562;
wire n_4077;
wire n_4642;
wire n_2221;
wire n_3576;
wire n_1792;
wire n_1868;
wire n_4049;
wire n_3862;
wire n_5214;
wire n_5487;
wire n_5563;
wire n_3495;
wire n_3879;
wire n_2348;
wire n_5497;
wire n_4724;
wire n_1772;
wire n_5526;
wire n_2818;
wire n_3646;
wire n_2129;
wire n_3345;
wire n_4546;
wire n_3584;
wire n_3756;
wire n_2889;
wire n_5593;
wire n_5021;
wire n_2772;
wire n_5444;
wire n_1675;
wire n_1924;
wire n_4382;
wire n_3999;
wire n_2844;
wire n_2138;
wire n_5211;
wire n_5230;
wire n_2260;
wire n_5389;
wire n_1813;
wire n_4833;
wire n_3056;
wire n_2345;
wire n_5110;
wire n_3295;
wire n_2382;
wire n_4719;
wire n_4178;
wire n_3062;
wire n_2317;
wire n_5425;
wire n_3289;
wire n_1973;
wire n_2579;
wire n_1770;
wire n_4228;
wire n_4401;
wire n_1756;
wire n_1716;
wire n_2788;
wire n_2984;
wire n_3364;
wire n_5560;
wire n_1873;
wire n_3201;
wire n_3472;
wire n_2874;
wire n_5179;
wire n_4605;
wire n_4877;
wire n_3235;
wire n_4968;
wire n_5030;
wire n_3949;
wire n_3543;
wire n_3050;
wire n_3903;
wire n_4834;
wire n_5272;
wire n_2742;
wire n_3314;
wire n_2183;
wire n_4158;
wire n_2360;
wire n_3254;
wire n_5361;
wire n_4171;
wire n_4045;
wire n_4562;
wire n_5068;
wire n_3634;
wire n_2834;
wire n_2531;
wire n_5015;
wire n_2702;
wire n_2030;
wire n_3115;
wire n_4749;
wire n_4390;
wire n_5302;
wire n_4979;
wire n_1794;
wire n_2234;
wire n_4804;
wire n_5545;
wire n_2209;
wire n_4270;
wire n_2797;
wire n_5152;
wire n_2321;
wire n_3680;
wire n_3497;
wire n_5409;
wire n_2940;
wire n_2612;
wire n_5128;
wire n_4566;
wire n_2841;
wire n_3322;
wire n_4576;
wire n_2505;
wire n_2427;
wire n_4061;
wire n_3250;
wire n_2070;
wire n_2594;
wire n_1914;
wire n_2335;
wire n_2904;
wire n_5307;
wire n_4767;
wire n_4328;
wire n_3004;
wire n_3112;
wire n_2349;
wire n_3874;
wire n_5415;
wire n_4676;
wire n_4544;
wire n_2170;
wire n_3175;
wire n_3522;
wire n_4429;
wire n_4591;
wire n_3266;
wire n_4646;
wire n_4563;
wire n_4725;
wire n_2210;
wire n_4169;
wire n_5331;
wire n_3247;
wire n_3091;
wire n_3066;
wire n_2426;
wire n_4320;
wire n_5341;
wire n_4881;
wire n_5271;
wire n_5089;
wire n_5263;
wire n_3613;
wire n_3444;
wire n_4012;
wire n_5518;
wire n_4636;
wire n_5637;
wire n_4584;
wire n_5622;
wire n_3910;
wire n_4711;
wire n_3319;
wire n_5240;
wire n_3335;
wire n_3413;
wire n_5495;
wire n_1969;
wire n_4680;
wire n_2044;
wire n_5546;
wire n_2689;
wire n_3259;
wire n_5482;
wire n_4191;
wire n_5224;
wire n_4293;
wire n_2010;
wire n_3688;
wire n_3016;
wire n_1693;
wire n_5393;
wire n_2599;
wire n_3338;
wire n_3414;
wire n_1827;
wire n_4671;
wire n_4209;
wire n_5041;
wire n_1751;
wire n_5431;
wire n_2200;
wire n_3261;
wire n_5026;
wire n_3863;
wire n_3027;
wire n_2746;
wire n_5059;
wire n_5505;
wire n_3127;
wire n_1780;
wire n_3732;
wire n_4250;
wire n_5329;
wire n_3596;
wire n_4699;
wire n_3906;
wire n_4127;
wire n_3297;
wire n_2683;
wire n_2388;
wire n_4292;
wire n_3641;
wire n_4577;
wire n_4854;
wire n_4202;
wire n_5212;
wire n_5000;
wire n_2853;
wire n_3766;
wire n_2880;
wire n_1666;
wire n_3350;
wire n_2389;
wire n_4165;
wire n_4866;
wire n_4038;
wire n_4109;
wire n_5297;
wire n_5420;
wire n_4412;
wire n_3407;
wire n_3599;
wire n_3621;
wire n_5234;
wire n_2244;
wire n_3815;
wire n_2257;
wire n_2538;
wire n_2105;
wire n_5259;
wire n_3163;
wire n_5440;
wire n_1686;
wire n_3710;
wire n_4155;
wire n_2031;
wire n_3891;
wire n_4144;
wire n_2165;
wire n_3379;
wire n_4374;
wire n_3532;
wire n_5131;
wire n_1818;
wire n_2127;
wire n_3531;
wire n_2963;
wire n_3834;
wire n_4548;
wire n_3258;
wire n_4989;
wire n_4622;
wire n_4315;
wire n_2959;
wire n_2047;
wire n_1845;
wire n_2193;
wire n_2478;
wire n_5140;
wire n_4816;
wire n_2983;
wire n_3810;
wire n_2715;
wire n_5598;
wire n_2085;
wire n_1669;
wire n_5306;
wire n_4483;
wire n_5342;
wire n_2782;
wire n_2672;
wire n_1670;
wire n_2651;
wire n_4358;
wire n_5147;
wire n_3656;
wire n_2071;
wire n_2643;
wire n_2561;
wire n_4793;
wire n_4168;
wire n_3446;
wire n_5511;
wire n_3028;
wire n_4806;
wire n_4350;
wire n_5533;
wire n_5280;
wire n_5235;
wire n_3836;
wire n_3963;
wire n_1872;
wire n_3389;
wire n_1931;
wire n_4187;
wire n_4166;
wire n_5206;
wire n_3222;
wire n_1801;
wire n_5419;
wire n_2970;
wire n_2235;
wire n_4937;
wire n_3980;
wire n_2791;
wire n_5103;
wire n_3755;
wire n_4258;
wire n_4498;
wire n_2174;
wire n_2714;
wire n_5285;
wire n_3563;
wire n_2506;
wire n_4064;
wire n_4936;
wire n_5387;
wire n_1863;
wire n_3841;
wire n_2118;
wire n_4770;
wire n_2944;
wire n_2407;
wire n_4907;
wire n_5058;
wire n_3262;
wire n_5018;
wire n_4006;
wire n_4861;
wire n_3690;
wire n_2358;
wire n_5192;
wire n_5141;
wire n_3716;
wire n_5133;
wire n_1700;
wire n_2833;
wire n_4712;
wire n_3191;
wire n_3837;
wire n_3193;
wire n_1971;
wire n_3252;
wire n_2275;
wire n_2855;
wire n_3273;
wire n_3544;
wire n_4310;
wire n_1950;
wire n_2370;
wire n_5159;
wire n_3954;
wire n_3025;
wire n_4674;
wire n_4908;
wire n_5097;
wire n_2750;
wire n_3899;
wire n_4159;
wire n_3714;
wire n_3071;
wire n_3739;
wire n_4069;
wire n_2784;
wire n_3718;
wire n_3092;
wire n_3470;
wire n_4862;
wire n_2557;
wire n_5300;
wire n_4850;
wire n_3781;
wire n_4813;
wire n_4912;
wire n_2590;
wire n_2330;
wire n_2942;
wire n_5525;
wire n_3106;
wire n_1882;
wire n_3328;
wire n_3889;
wire n_4256;
wire n_4224;
wire n_3508;
wire n_4024;
wire n_2267;
wire n_2218;
wire n_2636;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_5400;
wire n_2759;
wire n_4415;
wire n_5552;
wire n_4702;
wire n_4252;
wire n_4457;
wire n_5139;
wire n_2319;
wire n_3481;
wire n_5481;
wire n_2808;
wire n_2679;
wire n_1709;
wire n_2676;
wire n_4491;
wire n_2930;
wire n_1838;
wire n_3514;
wire n_2777;
wire n_2434;
wire n_4132;
wire n_2660;
wire n_2611;
wire n_4261;
wire n_1660;
wire n_4886;
wire n_4090;
wire n_2529;
wire n_2698;
wire n_5043;
wire n_1662;
wire n_4001;
wire n_3047;
wire n_2454;
wire n_4371;
wire n_5281;
wire n_4473;
wire n_3120;
wire n_4007;
wire n_1743;
wire n_4268;
wire n_5048;
wire n_5521;
wire n_5028;
wire n_4480;
wire n_2350;
wire n_3895;
wire n_4194;
wire n_5585;
wire n_4824;
wire n_1892;
wire n_4120;
wire n_4427;
wire n_3745;
wire n_2990;
wire n_1766;
wire n_3119;
wire n_4142;
wire n_4082;
wire n_5561;
wire n_3479;
wire n_4085;
wire n_4073;
wire n_4260;
wire n_1649;
wire n_4163;
wire n_4439;
wire n_2064;
wire n_3867;
wire n_4372;
wire n_3500;
wire n_3279;
wire n_2621;
wire n_5073;
wire n_5024;
wire n_4262;
wire n_2671;
wire n_1798;
wire n_1790;
wire n_4720;
wire n_1647;
wire n_4685;
wire n_2563;
wire n_2387;
wire n_4334;
wire n_1674;
wire n_1830;
wire n_2073;
wire n_4511;
wire n_5515;
wire n_4014;
wire n_5250;
wire n_3144;
wire n_4757;
wire n_2913;
wire n_2336;
wire n_5607;
wire n_4175;
wire n_2005;
wire n_1916;
wire n_4648;
wire n_5006;
wire n_4892;
wire n_3823;
wire n_1866;
wire n_4173;
wire n_4970;
wire n_3816;
wire n_5404;
wire n_4108;
wire n_4486;
wire n_2960;
wire n_5438;
wire n_4627;
wire n_2290;
wire n_2045;
wire n_3369;
wire n_3783;
wire n_2040;
wire n_3199;
wire n_3843;
wire n_2145;
wire n_1639;
wire n_3030;
wire n_2580;
wire n_3685;
wire n_4249;
wire n_5163;
wire n_2039;
wire n_4961;
wire n_3753;
wire n_2035;
wire n_4718;
wire n_3555;
wire n_3579;
wire n_5190;
wire n_2509;
wire n_3236;
wire n_4317;
wire n_4855;
wire n_3969;
wire n_2459;
wire n_4154;
wire n_3396;
wire n_4023;
wire n_4420;
wire n_1923;
wire n_5138;
wire n_5374;
wire n_2116;
wire n_1828;
wire n_2320;
wire n_5349;
wire n_2038;
wire n_2137;
wire n_4973;
wire n_4640;
wire n_2583;
wire n_4396;
wire n_5127;
wire n_4367;
wire n_2087;
wire n_5485;
wire n_5216;
wire n_1989;
wire n_3818;
wire n_2523;
wire n_4387;
wire n_4951;
wire n_4453;
wire n_4170;
wire n_3719;
wire n_1959;
wire n_3681;
wire n_2737;
wire n_2399;
wire n_4308;
wire n_2812;
wire n_2355;
wire n_2133;
wire n_3830;
wire n_2585;
wire n_2725;
wire n_5175;
wire n_3883;
wire n_2565;
wire n_4152;
wire n_4392;
wire n_4660;
wire n_3149;
wire n_5611;
wire n_3268;
wire n_4281;
wire n_4661;
wire n_4200;
wire n_3614;
wire n_2111;
wire n_3301;
wire n_3466;
wire n_4962;
wire n_2595;
wire n_3411;
wire n_4958;
wire n_4271;
wire n_5171;
wire n_3586;
wire n_5554;
wire n_4071;
wire n_4921;
wire n_1980;
wire n_5427;
wire n_3065;
wire n_4361;
wire n_5417;
wire n_4614;
wire n_2681;
wire n_3103;
wire n_4945;
wire n_2424;
wire n_4922;
wire n_4732;
wire n_1651;
wire n_2775;
wire n_4693;
wire n_5488;
wire n_4326;
wire n_3557;
wire n_2230;
wire n_5447;
wire n_5383;
wire n_4744;
wire n_2851;
wire n_4305;
wire n_2490;
wire n_4213;
wire n_2849;
wire n_3692;
wire n_2204;
wire n_4929;
wire n_1961;
wire n_4964;
wire n_4802;
wire n_4139;
wire n_3029;
wire n_2508;
wire n_4031;
wire n_2416;
wire n_5437;
wire n_3881;
wire n_2461;
wire n_2243;
wire n_4583;
wire n_4210;
wire n_5245;
wire n_4666;
wire n_2929;
wire n_3751;
wire n_2555;
wire n_2662;
wire n_2368;
wire n_2890;
wire n_2554;
wire n_3698;
wire n_3927;
wire n_1840;
wire n_4540;
wire n_3961;
wire n_1630;
wire n_4891;
wire n_5603;
wire n_3559;
wire n_2661;
wire n_2572;
wire n_3993;
wire n_4940;
wire n_5208;
wire n_3588;
wire n_2308;
wire n_4590;
wire n_5606;
wire n_4830;
wire n_5231;
wire n_5237;
wire n_4664;
wire n_3860;
wire n_5456;
wire n_3160;
wire n_2191;
wire n_5093;
wire n_2428;
wire n_3847;
wire n_4946;
wire n_4906;
wire n_2158;
wire n_3290;
wire n_4663;
wire n_5390;
wire n_5347;
wire n_2824;
wire n_3033;
wire n_3298;
wire n_2440;
wire n_4883;
wire n_2923;
wire n_4162;
wire n_3665;
wire n_5115;
wire n_3264;
wire n_2333;
wire n_2916;
wire n_4297;
wire n_1632;
wire n_3800;
wire n_2403;
wire n_5407;
wire n_4608;
wire n_5232;
wire n_2792;
wire n_2870;
wire n_3991;
wire n_3134;
wire n_4172;
wire n_4791;
wire n_4536;
wire n_5149;
wire n_2463;
wire n_5151;
wire n_4773;
wire n_5345;
wire n_5357;
wire n_4497;
wire n_2472;
wire n_4611;
wire n_4755;
wire n_1768;
wire n_2294;
wire n_4960;
wire n_2993;
wire n_1719;
wire n_3864;
wire n_4658;
wire n_5135;
wire n_2732;
wire n_2948;
wire n_2309;
wire n_5494;
wire n_4362;
wire n_4306;
wire n_2123;
wire n_3209;
wire n_3504;
wire n_2685;
wire n_2037;
wire n_1953;
wire n_4422;
wire n_2589;
wire n_3482;
wire n_2233;
wire n_4555;
wire n_2827;
wire n_5136;
wire n_5228;
wire n_3956;
wire n_5323;
wire n_3572;
wire n_4215;
wire n_4280;
wire n_3375;
wire n_4047;
wire n_5471;
wire n_5434;
wire n_2082;
wire n_1643;
wire n_3167;
wire n_5558;
wire n_5350;
wire n_3423;
wire n_2362;
wire n_2609;
wire n_5338;
wire n_1976;
wire n_2223;
wire n_3044;
wire n_3854;
wire n_2468;
wire n_3078;
wire n_3253;
wire n_4027;
wire n_2280;
wire n_4599;
wire n_3363;
wire n_4812;
wire n_3689;
wire n_2020;
wire n_4628;
wire n_1881;
wire n_2749;
wire n_3451;
wire n_4873;
wire n_5588;
wire n_4657;
wire n_2971;
wire n_2311;
wire n_3950;
wire n_4458;
wire n_4121;
wire n_5090;
wire n_4476;
wire n_5613;
wire n_2298;
wire n_4756;
wire n_3869;
wire n_4307;
wire n_5104;
wire n_5042;
wire n_4860;
wire n_4359;
wire n_2303;
wire n_2810;
wire n_2747;
wire n_1848;
wire n_5571;
wire n_2126;
wire n_4573;
wire n_5289;
wire n_4118;
wire n_5513;
wire n_4803;
wire n_4079;
wire n_4091;
wire n_1638;
wire n_2002;
wire n_5145;
wire n_3712;
wire n_2371;
wire n_2935;
wire n_5132;
wire n_5191;
wire n_3085;
wire n_1655;
wire n_5359;
wire n_2574;
wire n_5293;
wire n_4316;
wire n_3697;
wire n_2638;
wire n_4044;
wire n_4062;
wire n_4524;
wire n_4843;
wire n_3971;
wire n_5510;
wire n_2016;
wire n_2949;
wire n_2711;
wire n_5363;
wire n_5200;
wire n_1653;
wire n_5618;
wire n_2867;
wire n_1894;
wire n_2794;
wire n_3145;
wire n_3124;
wire n_4253;
wire n_5356;
wire n_5369;
wire n_2608;
wire n_5258;
wire n_2657;
wire n_5255;
wire n_2852;
wire n_2392;
wire n_3517;
wire n_3100;
wire n_2522;
wire n_1834;
wire n_3758;
wire n_3356;
wire n_2835;
wire n_1968;
wire n_3269;
wire n_5080;
wire n_3506;
wire n_1736;
wire n_3605;
wire n_2409;
wire n_3402;
wire n_5295;
wire n_4679;
wire n_4115;
wire n_4998;
wire n_2988;
wire n_1731;
wire n_1970;
wire n_2766;
wire n_5627;
wire n_2201;
wire n_2117;
wire n_4167;
wire n_1993;
wire n_5155;
wire n_3835;
wire n_2205;
wire n_1777;
wire n_1957;
wire n_3967;
wire n_5016;
wire n_1912;
wire n_3401;
wire n_3226;
wire n_3902;
wire n_4730;
wire n_2779;
wire n_3654;
wire n_2164;
wire n_2115;
wire n_2232;
wire n_5327;
wire n_1774;
wire n_4713;
wire n_5137;
wire n_2811;
wire n_3348;
wire n_3358;
wire n_2121;
wire n_1803;
wire n_4204;
wire n_5098;
wire n_1991;
wire n_2224;
wire n_4743;
wire n_3805;
wire n_3825;
wire n_3657;
wire n_4924;
wire n_3928;
wire n_4859;
wire n_2692;
wire n_2008;
wire n_4654;
wire n_5423;
wire n_4733;
wire n_3792;
wire n_4272;
wire n_3974;
wire n_3871;
wire n_1753;
wire n_2283;
wire n_3278;
wire n_1689;
wire n_4269;
wire n_4695;
wire n_1855;
wire n_3312;
wire n_2197;
wire n_2199;
wire n_5069;
wire n_3285;
wire n_3968;
wire n_5099;
wire n_2228;
wire n_4704;
wire n_4551;
wire n_5052;
wire n_2421;
wire n_2902;
wire n_4957;
wire n_2480;
wire n_2363;
wire n_4072;
wire n_5579;
wire n_4781;
wire n_3606;
wire n_5004;
wire n_2550;
wire n_4424;
wire n_3055;
wire n_3711;
wire n_3315;
wire n_3172;
wire n_3292;
wire n_4436;
wire n_3878;
wire n_4450;
wire n_3553;
wire n_4746;
wire n_1683;
wire n_3131;
wire n_5118;
wire n_5105;
wire n_3850;
wire n_4459;
wire n_2996;
wire n_5591;
wire n_4050;
wire n_2315;
wire n_3228;
wire n_2102;
wire n_5623;
wire n_4853;
wire n_2422;
wire n_2239;
wire n_5256;
wire n_2950;
wire n_5220;
wire n_3852;
wire n_5178;
wire n_4520;
wire n_2057;
wire n_4008;
wire n_5507;
wire n_5077;
wire n_3858;
wire n_1901;
wire n_4502;
wire n_3032;
wire n_4851;
wire n_3072;
wire n_3081;
wire n_3313;
wire n_2710;
wire n_1745;
wire n_3924;
wire n_4571;
wire n_2006;
wire n_5314;
wire n_2343;
wire n_3439;
wire n_5049;
wire n_2535;
wire n_4205;
wire n_2726;
wire n_5277;
wire n_4723;
wire n_5176;
wire n_2799;
wire n_4454;
wire n_4229;
wire n_4739;
wire n_2376;
wire n_5483;
wire n_3017;
wire n_2456;
wire n_3904;
wire n_5150;
wire n_2678;
wire n_4838;
wire n_2872;
wire n_2451;
wire n_5075;
wire n_4879;
wire n_5051;
wire n_3926;
wire n_1962;
wire n_3996;
wire n_4221;
wire n_2854;
wire n_1701;
wire n_4181;
wire n_2764;
wire n_4225;
wire n_2567;
wire n_5142;
wire n_3102;
wire n_1648;
wire n_4153;
wire n_5156;
wire n_3627;
wire n_4300;
wire n_3551;
wire n_1769;
wire n_4783;
wire n_2964;
wire n_3769;
wire n_2673;
wire n_4530;
wire n_4267;
wire n_2292;
wire n_3865;
wire n_3859;
wire n_3722;
wire n_2442;
wire n_1943;
wire n_3117;
wire n_3428;
wire n_2961;
wire n_3351;
wire n_3527;
wire n_2883;
wire n_1752;
wire n_4182;
wire n_2912;
wire n_4825;
wire n_4440;
wire n_4549;
wire n_1910;
wire n_3955;
wire n_5120;
wire n_5470;
wire n_4565;
wire n_4039;
wire n_3227;
wire n_3300;
wire n_4303;
wire n_4574;
wire n_4839;
wire n_5222;
wire n_4016;
wire n_3435;
wire n_3575;
wire n_4231;
wire n_3165;
wire n_4923;
wire n_3652;
wire n_4097;
wire n_4083;
wire n_1937;
wire n_4461;
wire n_3234;
wire n_5392;
wire n_2381;
wire n_3303;
wire n_1654;
wire n_3916;
wire n_2569;
wire n_3556;
wire n_4101;
wire n_2196;
wire n_3591;
wire n_4273;
wire n_3024;
wire n_5443;
wire n_3512;
wire n_5600;
wire n_4939;
wire n_5169;
wire n_4389;
wire n_3930;
wire n_4448;
wire n_2161;
wire n_2404;
wire n_2083;
wire n_2503;
wire n_1936;
wire n_5502;
wire n_2027;
wire n_5568;
wire n_2642;
wire n_2500;
wire n_1918;
wire n_4831;
wire n_2513;
wire n_2695;
wire n_3480;
wire n_3057;
wire n_3194;
wire n_2414;
wire n_3662;
wire n_4319;
wire n_5474;
wire n_2229;
wire n_4596;
wire n_5413;
wire n_2004;
wire n_5412;
wire n_3694;
wire n_2586;
wire n_4726;
wire n_1879;
wire n_4751;
wire n_4222;
wire n_2274;
wire n_2972;
wire n_3225;
wire n_4119;
wire n_3799;
wire n_4298;
wire n_5201;
wire n_4474;
wire n_5217;
wire n_2511;
wire n_1681;
wire n_3383;
wire n_3585;
wire n_2975;
wire n_5490;
wire n_5029;
wire n_2704;
wire n_4214;
wire n_5158;
wire n_4884;
wire n_4366;
wire n_4009;
wire n_4580;
wire n_4129;
wire n_4871;
wire n_2617;
wire n_4999;
wire n_1859;
wire n_1677;
wire n_5557;
wire n_5472;
wire n_2955;
wire n_4112;
wire n_4337;
wire n_4138;
wire n_5396;
wire n_5335;
wire n_2520;
wire n_2134;
wire n_4236;
wire n_2185;
wire n_3270;
wire n_2143;
wire n_5002;
wire n_3595;
wire n_5143;
wire n_4238;
wire n_2374;
wire n_1947;
wire n_2114;
wire n_3571;
wire n_2396;
wire n_1799;
wire n_4734;
wire n_1939;
wire n_2486;
wire n_4635;
wire n_3501;
wire n_1869;
wire n_4013;
wire n_3039;
wire n_2011;
wire n_4242;
wire n_4984;
wire n_3851;
wire n_2543;
wire n_3036;
wire n_1896;
wire n_3180;
wire n_5283;
wire n_5268;
wire n_1705;
wire n_4561;
wire n_2639;
wire n_3325;
wire n_3107;
wire n_4021;
wire n_3880;
wire n_5122;
wire n_3186;
wire n_4955;
wire n_5556;
wire n_5462;
wire n_4501;
wire n_3696;
wire n_3650;
wire n_2761;
wire n_3157;
wire n_2537;
wire n_2144;
wire n_2515;
wire n_2466;
wire n_2652;
wire n_2635;
wire n_5330;
wire n_4197;
wire n_4829;
wire n_1949;
wire n_2936;
wire n_1946;
wire n_4715;
wire n_5039;
wire n_2141;
wire n_4369;
wire n_5378;
wire n_4543;
wire n_2099;
wire n_4941;
wire n_5542;
wire n_1831;
wire n_4394;
wire n_1850;
wire n_5519;
wire n_1749;
wire n_3101;
wire n_3669;
wire n_5278;
wire n_2663;
wire n_5586;
wire n_2693;
wire n_3798;
wire n_4065;
wire n_5187;
wire n_4944;
wire n_2249;
wire n_2180;
wire n_4135;
wire n_2632;
wire n_1755;
wire n_2908;
wire n_3744;
wire n_4263;
wire n_1862;
wire n_2915;
wire n_2300;
wire n_3291;
wire n_4716;
wire n_4942;
wire n_2432;
wire n_3405;
wire n_4745;
wire n_2337;
wire n_3907;
wire n_5344;
wire n_4629;
wire n_2932;
wire n_2980;
wire n_5225;
wire n_3306;
wire n_1784;
wire n_4857;
wire n_3136;
wire n_4080;
wire n_4226;
wire n_4741;
wire n_2101;
wire n_1986;
wire n_4752;
wire n_5265;
wire n_1750;
wire n_3986;
wire n_4376;
wire n_4753;
wire n_4552;
wire n_3885;
wire n_2713;
wire n_5196;
wire n_5181;
wire n_2644;
wire n_2951;
wire n_3008;
wire n_3709;
wire n_5574;
wire n_5126;
wire n_2214;
wire n_2055;
wire n_3427;
wire n_4067;
wire n_5553;
wire n_4042;
wire n_4176;
wire n_4385;
wire n_3320;
wire n_5009;
wire n_2688;
wire n_5368;
wire n_5626;
wire n_3651;
wire n_4333;
wire n_3359;
wire n_2865;
wire n_2706;
wire n_5499;
wire n_3676;
wire n_4375;
wire n_4788;
wire n_4717;
wire n_4986;
wire n_5604;
wire n_3789;
wire n_2152;
wire n_3598;
wire n_4815;
wire n_4246;
wire n_3580;
wire n_2139;
wire n_4609;
wire n_5291;
wire n_5114;
wire n_2674;
wire n_4088;
wire n_3682;
wire n_4357;
wire n_3371;
wire n_1809;
wire n_4462;
wire n_4472;
wire n_3433;
wire n_5288;
wire n_2305;
wire n_5540;
wire n_2450;
wire n_3447;
wire n_3305;
wire n_4148;
wire n_4151;
wire n_1712;
wire n_3528;
wire n_4373;
wire n_4934;
wire n_5218;
wire n_2322;
wire n_2271;
wire n_2625;
wire n_4630;
wire n_5408;
wire n_4643;
wire n_4331;
wire n_3989;
wire n_4475;
wire n_4846;
wire n_3804;
wire n_4344;
wire n_1775;
wire n_3296;
wire n_2762;
wire n_4683;
wire n_5366;
wire n_1847;
wire n_2767;
wire n_2603;
wire n_3116;
wire n_1884;
wire n_3602;
wire n_2967;
wire n_1905;
wire n_2553;
wire n_3706;
wire n_2195;
wire n_5477;
wire n_5451;
wire n_3923;
wire n_4696;
wire n_2626;
wire n_3441;
wire n_1978;
wire n_5086;
wire n_1629;
wire n_2801;
wire n_4011;
wire n_4905;
wire n_2763;
wire n_2825;
wire n_3643;
wire n_4876;
wire n_1997;
wire n_3748;
wire n_3142;
wire n_4278;
wire n_1635;
wire n_4623;
wire n_4910;
wire n_2690;
wire n_4410;
wire n_3370;
wire n_2215;
wire n_5053;
wire n_4553;
wire n_3978;
wire n_4809;
wire n_5226;
wire n_1925;
wire n_3660;
wire n_1815;
wire n_1788;
wire n_2491;
wire n_5079;
wire n_5590;
wire n_3833;
wire n_5632;
wire n_1679;
wire n_4841;
wire n_2022;
wire n_3814;
wire n_2592;
wire n_2838;
wire n_4842;
wire n_4911;
wire n_4340;
wire n_3513;
wire n_3133;
wire n_4645;
wire n_2992;
wire n_3725;
wire n_1833;
wire n_4920;
wire n_4972;
wire n_2517;
wire n_3128;
wire n_5426;
wire n_2631;
wire n_2178;
wire n_1767;
wire n_2469;
wire n_5625;
wire n_3355;
wire n_2007;
wire n_3917;
wire n_3942;
wire n_2736;
wire n_3765;
wire n_5531;
wire n_3000;
wire n_5429;
wire n_3108;
wire n_3111;
wire n_1839;
wire n_1837;
wire n_4557;
wire n_5248;
wire n_4451;
wire n_2875;
wire n_3844;
wire n_3280;
wire n_4054;
wire n_5448;
wire n_3471;
wire n_5432;
wire n_3205;
wire n_2046;
wire n_2848;
wire n_5160;
wire n_2741;
wire n_3003;
wire n_3610;
wire n_1933;
wire n_1656;
wire n_3564;
wire n_3988;
wire n_3457;
wire n_1678;
wire n_4324;
wire n_4821;
wire n_1871;
wire n_5445;
wire n_3630;
wire n_3271;
wire n_4771;
wire n_4086;
wire n_2412;
wire n_4814;
wire n_1781;
wire n_2084;
wire n_3648;
wire n_3075;
wire n_3173;
wire n_5332;
wire n_5108;
wire n_4692;
wire n_3031;
wire n_3701;
wire n_1773;
wire n_3243;
wire n_2666;
wire n_3385;
wire n_2171;
wire n_4708;
wire n_2768;
wire n_2314;
wire n_4826;
wire n_2420;
wire n_3343;
wire n_5489;
wire n_3767;
wire n_2873;
wire n_2299;
wire n_2540;
wire n_4589;
wire n_5057;
wire n_4578;
wire n_1640;
wire n_2162;
wire n_2847;
wire n_2051;
wire n_3221;
wire n_5436;
wire n_2168;
wire n_2790;
wire n_5072;
wire n_3629;
wire n_3021;
wire n_2359;
wire n_3674;
wire n_5286;
wire n_3502;
wire n_3098;
wire n_5013;
wire n_2312;
wire n_3015;
wire n_1920;
wire n_5569;
wire n_5439;
wire n_5619;
wire n_4147;
wire n_2048;
wire n_3607;
wire n_4925;
wire n_1921;
wire n_4974;
wire n_1800;
wire n_4932;
wire n_4510;
wire n_2571;
wire n_3276;
wire n_3787;
wire n_5119;
wire n_2124;
wire n_3827;
wire n_2519;
wire n_3354;
wire n_2724;
wire n_4447;
wire n_4285;
wire n_4651;
wire n_4818;
wire n_4514;
wire n_4800;
wire n_3960;
wire n_3248;
wire n_2277;
wire n_2110;
wire n_4433;
wire n_2879;
wire n_2474;
wire n_2090;
wire n_3153;
wire n_2033;
wire n_4341;
wire n_1682;
wire n_4312;
wire n_2628;
wire n_3399;
wire n_2132;
wire n_2400;
wire n_4633;
wire n_3838;
wire n_1909;
wire n_4277;
wire n_4140;
wire n_3675;
wire n_5092;
wire n_3387;
wire n_5186;
wire n_4662;
wire n_3779;
wire n_2464;
wire n_2831;
wire n_4882;
wire n_4993;
wire n_2365;
wire n_4832;
wire n_4207;
wire n_4545;
wire n_3037;
wire n_4868;
wire n_1885;
wire n_2452;
wire n_3925;
wire n_2176;
wire n_1816;
wire n_5238;
wire n_4059;
wire n_2455;
wire n_4595;
wire n_1849;
wire n_5054;
wire n_5631;
wire n_2467;
wire n_2288;
wire n_4063;
wire n_5399;
wire n_3592;
wire n_4650;
wire n_4888;
wire n_5326;
wire n_3394;
wire n_4874;
wire n_3793;
wire n_4669;
wire n_4339;
wire n_1645;
wire n_4041;
wire n_5459;
wire n_2858;
wire n_4060;
wire n_2658;
wire n_1717;
wire n_2895;
wire n_2128;
wire n_5528;
wire n_3097;
wire n_5391;
wire n_4541;
wire n_3824;
wire n_5422;
wire n_3388;
wire n_5267;
wire n_4494;
wire n_3059;
wire n_5523;
wire n_3465;
wire n_4796;
wire n_3589;
wire n_2534;
wire n_4799;
wire n_5153;
wire n_3449;
wire n_2694;
wire n_2198;
wire n_2610;
wire n_2989;
wire n_2789;
wire n_4775;
wire n_2216;
wire n_5044;
wire n_1897;
wire n_5365;
wire n_2933;
wire n_5045;
wire n_4381;
wire n_4266;
wire n_3886;
wire n_5354;
wire n_4455;
wire n_2328;
wire n_4248;
wire n_5452;
wire n_4754;
wire n_4554;
wire n_5595;
wire n_4845;
wire n_3053;
wire n_3893;
wire n_2465;
wire n_3548;
wire n_4585;
wire n_1699;
wire n_3334;
wire n_2541;
wire n_4383;
wire n_5535;
wire n_3875;
wire n_5370;
wire n_4003;
wire n_5372;
wire n_5299;
wire n_2402;
wire n_5594;
wire n_4301;
wire n_4586;
wire n_1954;
wire n_4048;
wire n_1844;
wire n_3777;
wire n_4784;
wire n_2999;
wire n_1644;
wire n_5550;
wire n_5082;
wire n_4046;
wire n_1974;
wire n_2086;
wire n_3537;
wire n_5209;
wire n_3080;
wire n_4199;
wire n_2701;
wire n_3362;
wire n_1631;
wire n_5559;
wire n_3105;
wire n_5478;
wire n_4286;
wire n_5102;
wire n_2556;
wire n_2269;
wire n_3274;
wire n_3041;
wire n_4470;
wire n_2236;
wire n_2816;
wire n_1911;
wire n_3616;
wire n_2460;
wire n_4058;
wire n_3664;
wire n_4188;
wire n_1668;
wire n_3913;
wire n_3417;
wire n_4034;
wire n_1688;
wire n_3327;
wire n_5275;
wire n_4689;
wire n_5071;
wire n_3067;
wire n_2755;
wire n_3237;
wire n_1992;
wire n_4402;
wire n_4239;
wire n_3400;
wire n_4550;
wire n_3382;
wire n_3574;
wire n_5227;
wire n_2169;
wire n_4201;
wire n_3316;
wire n_5242;
wire n_3099;
wire n_3704;
wire n_2596;
wire n_1730;
wire n_3603;
wire n_4123;
wire n_2192;
wire n_5520;
wire n_3633;
wire n_4479;
wire n_2670;
wire n_1646;
wire n_4416;
wire n_3372;
wire n_4539;
wire n_2707;
wire n_2471;
wire n_1671;
wire n_3230;
wire n_3342;
wire n_4682;
wire n_5353;
wire n_3708;
wire n_5294;
wire n_3729;
wire n_4978;
wire n_4690;
wire n_4437;
wire n_5458;
wire n_3861;
wire n_5617;
wire n_4736;
wire n_3780;
wire n_1928;
wire n_5244;
wire n_5382;
wire n_3957;
wire n_5274;
wire n_3848;
wire n_4284;
wire n_2600;
wire n_3919;
wire n_5384;
wire n_3608;
wire n_4513;
wire n_3233;
wire n_3829;
wire n_3177;
wire n_4053;
wire n_2352;
wire n_5125;
wire n_4040;
wire n_2207;
wire n_5587;
wire n_2619;
wire n_2444;
wire n_3123;
wire n_5056;
wire n_5249;
wire n_3393;
wire n_5198;
wire n_5360;
wire n_5233;
wire n_4887;
wire n_4617;
wire n_5269;
wire n_3520;
wire n_2492;
wire n_4005;
wire n_1687;
wire n_1637;
wire n_4904;
wire n_4792;
wire n_3578;
wire n_3812;
wire n_1886;
wire n_4980;
wire n_4290;
wire n_5247;
wire n_3727;
wire n_5317;
wire n_3774;
wire n_3093;
wire n_1843;
wire n_3061;
wire n_1659;
wire n_2431;
wire n_4956;
wire n_5380;
wire n_2206;
wire n_3182;
wire n_2564;
wire n_4947;
wire n_4656;
wire n_3896;
wire n_3958;
wire n_3450;
wire n_4729;
wire n_4987;
wire n_5182;
wire n_4971;
wire n_2000;
wire n_2074;
wire n_3174;
wire n_2217;
wire n_3398;
wire n_2307;
wire n_3408;
wire n_2722;
wire n_5388;
wire n_2640;
wire n_4823;
wire n_4875;
wire n_3432;
wire n_1771;
wire n_3090;
wire n_2437;
wire n_3762;
wire n_5564;
wire n_2445;
wire n_1835;
wire n_1988;
wire n_1853;
wire n_1787;
wire n_4137;
wire n_2634;
wire n_4529;
wire n_4323;
wire n_3034;
wire n_2212;
wire n_3972;
wire n_5539;
wire n_3308;
wire n_5036;
wire n_5547;
wire n_4772;
wire n_3467;
wire n_4322;
wire n_1720;
wire n_2830;
wire n_4354;
wire n_4653;
wire n_2354;
wire n_2246;
wire n_5273;
wire n_4677;
wire n_3901;
wire n_5261;
wire n_3757;
wire n_3381;
wire n_5193;
wire n_1782;
wire n_2245;
wire n_4909;
wire n_2965;
wire n_3635;
wire n_5022;
wire n_5005;
wire n_2814;
wire n_3882;
wire n_3046;
wire n_2213;
wire n_3826;
wire n_3211;
wire n_2211;
wire n_2095;
wire n_3121;
wire n_4634;
wire n_3337;
wire n_2527;
wire n_5534;
wire n_3204;
wire n_2136;
wire n_5174;
wire n_1822;
wire n_4952;
wire n_5157;
wire n_3005;
wire n_4380;
wire n_3129;
wire n_4126;
wire n_1783;
wire n_2601;
wire n_5087;
wire n_3043;
wire n_3802;
wire n_2375;
wire n_4506;
wire n_4880;
wire n_1907;
wire n_2686;
wire n_2344;
wire n_3892;
wire n_4896;
wire n_5620;
wire n_5061;
wire n_5572;
wire n_1985;
wire n_2107;
wire n_3219;
wire n_2906;
wire n_4943;
wire n_2187;
wire n_1762;
wire n_3023;
wire n_4193;
wire n_4075;
wire n_3104;
wire n_4737;
wire n_3647;
wire n_2819;
wire n_5195;
wire n_3609;
wire n_4136;
wire n_1715;
wire n_1952;
wire n_4393;
wire n_3720;
wire n_4535;
wire n_1922;
wire n_2560;
wire n_4522;
wire n_4794;
wire n_3959;
wire n_3140;
wire n_5246;
wire n_3724;
wire n_2104;
wire n_3011;
wire n_5164;
wire n_4196;
wire n_4592;
wire n_4675;
wire n_5340;
wire n_3069;
wire n_5498;
wire n_4370;
wire n_1900;
wire n_5183;
wire n_3084;
wire n_1727;
wire n_2735;
wire n_2497;
wire n_3412;
wire n_1995;
wire n_5549;
wire n_2411;
wire n_3761;
wire n_4889;
wire n_2014;
wire n_2986;
wire n_5442;
wire n_1641;
wire n_3184;
wire n_4828;
wire n_5385;
wire n_4558;
wire n_2172;
wire n_4722;
wire n_3626;
wire n_4768;
wire n_4100;
wire n_2250;
wire n_4092;
wire n_3908;
wire n_2423;
wire n_3671;
wire n_3344;
wire n_2194;
wire n_4465;
wire n_3302;
wire n_5537;
wire n_5304;
wire n_2680;
wire n_5130;
wire n_3122;
wire n_5162;
wire n_4808;
wire n_3842;
wire n_3265;
wire n_1857;
wire n_4482;
wire n_2041;
wire n_1797;
wire n_2957;
wire n_2357;
wire n_3309;
wire n_3260;
wire n_4926;
wire n_3357;
wire n_4116;
wire n_2570;
wire n_1858;
wire n_2815;
wire n_5473;
wire n_3754;
wire n_4612;
wire n_2744;
wire n_4287;
wire n_2397;
wire n_2208;
wire n_3063;
wire n_5177;
wire n_3617;
wire n_1652;
wire n_4516;
wire n_3794;
wire n_2809;
wire n_2050;
wire n_4505;
wire n_1676;
wire n_2591;
wire n_3384;
wire n_4602;
wire n_5172;
wire n_4449;
wire n_1864;
wire n_5070;
wire n_4445;
wire n_5566;
wire n_5414;
wire n_4870;
wire n_2438;
wire n_2832;
wire n_1975;
wire n_2296;
wire n_3181;
wire n_2278;
wire n_4915;
wire n_5296;
wire n_2135;
wire n_5450;
wire n_3493;
wire n_5313;
wire n_3323;
wire n_2734;
wire n_4914;
wire n_2823;
wire n_1761;
wire n_5270;
wire n_4345;
wire n_5188;
wire n_3281;
wire n_3307;
wire n_1694;
wire n_4318;
wire n_2485;
wire n_2655;
wire n_4185;
wire n_4797;
wire n_2366;
wire n_3997;
wire n_5465;
wire n_4032;
wire n_1764;
wire n_3582;
wire n_2826;
wire n_3539;
wire n_4343;
wire n_4212;
wire n_4124;
wire n_5467;
wire n_5522;
wire n_4492;
wire n_2708;
wire n_5148;
wire n_4994;
wire n_4245;
wire n_4364;
wire n_4928;
wire n_2225;
wire n_4378;
wire n_2383;
wire n_1996;
wire n_3406;
wire n_3604;
wire n_3853;
wire n_4216;
wire n_2019;
wire n_2166;
wire n_2938;
wire n_4309;
wire n_3594;
wire n_1704;
wire n_3721;
wire n_2026;
wire n_2109;
wire n_2013;
wire n_1990;
wire n_2614;
wire n_2991;
wire n_2242;
wire n_2752;
wire n_2894;
wire n_3473;
wire n_4560;
wire n_5318;
wire n_2839;
wire n_5395;
wire n_2237;
wire n_3463;
wire n_3699;
wire n_5067;
wire n_3360;
wire n_2524;
wire n_3873;
wire n_3693;
wire n_2728;
wire n_3857;

CKINVDCx5p33_ASAP7_75t_R g1629 ( 
.A(n_1263),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1024),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_452),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_10),
.Y(n_1632)
);

CKINVDCx20_ASAP7_75t_R g1633 ( 
.A(n_1562),
.Y(n_1633)
);

CKINVDCx5p33_ASAP7_75t_R g1634 ( 
.A(n_409),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1190),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1044),
.Y(n_1636)
);

CKINVDCx5p33_ASAP7_75t_R g1637 ( 
.A(n_1529),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1004),
.Y(n_1638)
);

CKINVDCx5p33_ASAP7_75t_R g1639 ( 
.A(n_1012),
.Y(n_1639)
);

BUFx6f_ASAP7_75t_L g1640 ( 
.A(n_72),
.Y(n_1640)
);

CKINVDCx5p33_ASAP7_75t_R g1641 ( 
.A(n_440),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_913),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1402),
.Y(n_1643)
);

BUFx10_ASAP7_75t_L g1644 ( 
.A(n_932),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_405),
.Y(n_1645)
);

CKINVDCx5p33_ASAP7_75t_R g1646 ( 
.A(n_1505),
.Y(n_1646)
);

CKINVDCx5p33_ASAP7_75t_R g1647 ( 
.A(n_236),
.Y(n_1647)
);

CKINVDCx5p33_ASAP7_75t_R g1648 ( 
.A(n_1556),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_430),
.Y(n_1649)
);

CKINVDCx5p33_ASAP7_75t_R g1650 ( 
.A(n_327),
.Y(n_1650)
);

CKINVDCx5p33_ASAP7_75t_R g1651 ( 
.A(n_687),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_36),
.Y(n_1652)
);

CKINVDCx5p33_ASAP7_75t_R g1653 ( 
.A(n_500),
.Y(n_1653)
);

CKINVDCx5p33_ASAP7_75t_R g1654 ( 
.A(n_1539),
.Y(n_1654)
);

CKINVDCx5p33_ASAP7_75t_R g1655 ( 
.A(n_743),
.Y(n_1655)
);

CKINVDCx5p33_ASAP7_75t_R g1656 ( 
.A(n_153),
.Y(n_1656)
);

CKINVDCx5p33_ASAP7_75t_R g1657 ( 
.A(n_1355),
.Y(n_1657)
);

CKINVDCx5p33_ASAP7_75t_R g1658 ( 
.A(n_982),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1115),
.Y(n_1659)
);

CKINVDCx5p33_ASAP7_75t_R g1660 ( 
.A(n_491),
.Y(n_1660)
);

CKINVDCx5p33_ASAP7_75t_R g1661 ( 
.A(n_260),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_983),
.Y(n_1662)
);

CKINVDCx5p33_ASAP7_75t_R g1663 ( 
.A(n_911),
.Y(n_1663)
);

CKINVDCx5p33_ASAP7_75t_R g1664 ( 
.A(n_906),
.Y(n_1664)
);

CKINVDCx5p33_ASAP7_75t_R g1665 ( 
.A(n_149),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_260),
.Y(n_1666)
);

CKINVDCx5p33_ASAP7_75t_R g1667 ( 
.A(n_1482),
.Y(n_1667)
);

CKINVDCx5p33_ASAP7_75t_R g1668 ( 
.A(n_273),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_1046),
.Y(n_1669)
);

CKINVDCx5p33_ASAP7_75t_R g1670 ( 
.A(n_1491),
.Y(n_1670)
);

CKINVDCx20_ASAP7_75t_R g1671 ( 
.A(n_1351),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1421),
.Y(n_1672)
);

CKINVDCx5p33_ASAP7_75t_R g1673 ( 
.A(n_1105),
.Y(n_1673)
);

INVx1_ASAP7_75t_SL g1674 ( 
.A(n_1466),
.Y(n_1674)
);

CKINVDCx5p33_ASAP7_75t_R g1675 ( 
.A(n_770),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_1192),
.Y(n_1676)
);

CKINVDCx5p33_ASAP7_75t_R g1677 ( 
.A(n_957),
.Y(n_1677)
);

CKINVDCx5p33_ASAP7_75t_R g1678 ( 
.A(n_499),
.Y(n_1678)
);

CKINVDCx5p33_ASAP7_75t_R g1679 ( 
.A(n_948),
.Y(n_1679)
);

CKINVDCx5p33_ASAP7_75t_R g1680 ( 
.A(n_1509),
.Y(n_1680)
);

CKINVDCx16_ASAP7_75t_R g1681 ( 
.A(n_1005),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_734),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_193),
.Y(n_1683)
);

CKINVDCx5p33_ASAP7_75t_R g1684 ( 
.A(n_915),
.Y(n_1684)
);

CKINVDCx5p33_ASAP7_75t_R g1685 ( 
.A(n_1530),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1452),
.Y(n_1686)
);

BUFx2_ASAP7_75t_L g1687 ( 
.A(n_973),
.Y(n_1687)
);

CKINVDCx5p33_ASAP7_75t_R g1688 ( 
.A(n_1423),
.Y(n_1688)
);

CKINVDCx20_ASAP7_75t_R g1689 ( 
.A(n_255),
.Y(n_1689)
);

INVx2_ASAP7_75t_SL g1690 ( 
.A(n_101),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_958),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1202),
.Y(n_1692)
);

BUFx3_ASAP7_75t_L g1693 ( 
.A(n_972),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_570),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1476),
.Y(n_1695)
);

CKINVDCx5p33_ASAP7_75t_R g1696 ( 
.A(n_1492),
.Y(n_1696)
);

CKINVDCx5p33_ASAP7_75t_R g1697 ( 
.A(n_582),
.Y(n_1697)
);

CKINVDCx20_ASAP7_75t_R g1698 ( 
.A(n_1299),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1196),
.Y(n_1699)
);

CKINVDCx20_ASAP7_75t_R g1700 ( 
.A(n_1340),
.Y(n_1700)
);

BUFx6f_ASAP7_75t_L g1701 ( 
.A(n_1498),
.Y(n_1701)
);

CKINVDCx5p33_ASAP7_75t_R g1702 ( 
.A(n_1378),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_806),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_529),
.Y(n_1704)
);

INVx2_ASAP7_75t_SL g1705 ( 
.A(n_1537),
.Y(n_1705)
);

BUFx10_ASAP7_75t_L g1706 ( 
.A(n_744),
.Y(n_1706)
);

INVx1_ASAP7_75t_SL g1707 ( 
.A(n_737),
.Y(n_1707)
);

CKINVDCx5p33_ASAP7_75t_R g1708 ( 
.A(n_932),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_120),
.Y(n_1709)
);

CKINVDCx5p33_ASAP7_75t_R g1710 ( 
.A(n_99),
.Y(n_1710)
);

CKINVDCx5p33_ASAP7_75t_R g1711 ( 
.A(n_26),
.Y(n_1711)
);

CKINVDCx20_ASAP7_75t_R g1712 ( 
.A(n_1417),
.Y(n_1712)
);

CKINVDCx20_ASAP7_75t_R g1713 ( 
.A(n_1204),
.Y(n_1713)
);

CKINVDCx5p33_ASAP7_75t_R g1714 ( 
.A(n_410),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1495),
.Y(n_1715)
);

INVx1_ASAP7_75t_SL g1716 ( 
.A(n_61),
.Y(n_1716)
);

BUFx3_ASAP7_75t_L g1717 ( 
.A(n_1053),
.Y(n_1717)
);

CKINVDCx5p33_ASAP7_75t_R g1718 ( 
.A(n_310),
.Y(n_1718)
);

CKINVDCx5p33_ASAP7_75t_R g1719 ( 
.A(n_127),
.Y(n_1719)
);

CKINVDCx5p33_ASAP7_75t_R g1720 ( 
.A(n_324),
.Y(n_1720)
);

BUFx3_ASAP7_75t_L g1721 ( 
.A(n_1479),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1517),
.Y(n_1722)
);

CKINVDCx16_ASAP7_75t_R g1723 ( 
.A(n_1544),
.Y(n_1723)
);

CKINVDCx5p33_ASAP7_75t_R g1724 ( 
.A(n_252),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1561),
.Y(n_1725)
);

BUFx3_ASAP7_75t_L g1726 ( 
.A(n_1401),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1064),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_413),
.Y(n_1728)
);

CKINVDCx5p33_ASAP7_75t_R g1729 ( 
.A(n_544),
.Y(n_1729)
);

CKINVDCx5p33_ASAP7_75t_R g1730 ( 
.A(n_1259),
.Y(n_1730)
);

CKINVDCx5p33_ASAP7_75t_R g1731 ( 
.A(n_695),
.Y(n_1731)
);

CKINVDCx5p33_ASAP7_75t_R g1732 ( 
.A(n_842),
.Y(n_1732)
);

CKINVDCx5p33_ASAP7_75t_R g1733 ( 
.A(n_1561),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1205),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_534),
.Y(n_1735)
);

CKINVDCx5p33_ASAP7_75t_R g1736 ( 
.A(n_64),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_536),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1187),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1513),
.Y(n_1739)
);

CKINVDCx5p33_ASAP7_75t_R g1740 ( 
.A(n_823),
.Y(n_1740)
);

CKINVDCx5p33_ASAP7_75t_R g1741 ( 
.A(n_231),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1206),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_532),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_763),
.Y(n_1744)
);

CKINVDCx5p33_ASAP7_75t_R g1745 ( 
.A(n_116),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_671),
.Y(n_1746)
);

CKINVDCx5p33_ASAP7_75t_R g1747 ( 
.A(n_755),
.Y(n_1747)
);

CKINVDCx5p33_ASAP7_75t_R g1748 ( 
.A(n_1041),
.Y(n_1748)
);

BUFx6f_ASAP7_75t_L g1749 ( 
.A(n_460),
.Y(n_1749)
);

CKINVDCx5p33_ASAP7_75t_R g1750 ( 
.A(n_22),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_951),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1537),
.Y(n_1752)
);

CKINVDCx5p33_ASAP7_75t_R g1753 ( 
.A(n_291),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_944),
.Y(n_1754)
);

INVxp67_ASAP7_75t_L g1755 ( 
.A(n_1476),
.Y(n_1755)
);

CKINVDCx16_ASAP7_75t_R g1756 ( 
.A(n_1448),
.Y(n_1756)
);

INVx2_ASAP7_75t_L g1757 ( 
.A(n_983),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_108),
.Y(n_1758)
);

BUFx6f_ASAP7_75t_L g1759 ( 
.A(n_1532),
.Y(n_1759)
);

CKINVDCx5p33_ASAP7_75t_R g1760 ( 
.A(n_327),
.Y(n_1760)
);

CKINVDCx20_ASAP7_75t_R g1761 ( 
.A(n_1514),
.Y(n_1761)
);

CKINVDCx5p33_ASAP7_75t_R g1762 ( 
.A(n_380),
.Y(n_1762)
);

CKINVDCx5p33_ASAP7_75t_R g1763 ( 
.A(n_704),
.Y(n_1763)
);

CKINVDCx5p33_ASAP7_75t_R g1764 ( 
.A(n_1503),
.Y(n_1764)
);

INVx3_ASAP7_75t_L g1765 ( 
.A(n_1001),
.Y(n_1765)
);

BUFx2_ASAP7_75t_L g1766 ( 
.A(n_1121),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_741),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1018),
.Y(n_1768)
);

BUFx6f_ASAP7_75t_L g1769 ( 
.A(n_1534),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1462),
.Y(n_1770)
);

CKINVDCx5p33_ASAP7_75t_R g1771 ( 
.A(n_944),
.Y(n_1771)
);

BUFx3_ASAP7_75t_L g1772 ( 
.A(n_808),
.Y(n_1772)
);

CKINVDCx16_ASAP7_75t_R g1773 ( 
.A(n_1464),
.Y(n_1773)
);

CKINVDCx5p33_ASAP7_75t_R g1774 ( 
.A(n_1461),
.Y(n_1774)
);

CKINVDCx16_ASAP7_75t_R g1775 ( 
.A(n_351),
.Y(n_1775)
);

CKINVDCx5p33_ASAP7_75t_R g1776 ( 
.A(n_1189),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_11),
.Y(n_1777)
);

CKINVDCx5p33_ASAP7_75t_R g1778 ( 
.A(n_452),
.Y(n_1778)
);

CKINVDCx5p33_ASAP7_75t_R g1779 ( 
.A(n_1206),
.Y(n_1779)
);

INVx2_ASAP7_75t_L g1780 ( 
.A(n_840),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_660),
.Y(n_1781)
);

CKINVDCx5p33_ASAP7_75t_R g1782 ( 
.A(n_990),
.Y(n_1782)
);

BUFx10_ASAP7_75t_L g1783 ( 
.A(n_1283),
.Y(n_1783)
);

INVx2_ASAP7_75t_SL g1784 ( 
.A(n_334),
.Y(n_1784)
);

CKINVDCx5p33_ASAP7_75t_R g1785 ( 
.A(n_963),
.Y(n_1785)
);

CKINVDCx20_ASAP7_75t_R g1786 ( 
.A(n_749),
.Y(n_1786)
);

BUFx8_ASAP7_75t_SL g1787 ( 
.A(n_1243),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_270),
.Y(n_1788)
);

BUFx3_ASAP7_75t_L g1789 ( 
.A(n_1374),
.Y(n_1789)
);

CKINVDCx5p33_ASAP7_75t_R g1790 ( 
.A(n_214),
.Y(n_1790)
);

CKINVDCx5p33_ASAP7_75t_R g1791 ( 
.A(n_1105),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1040),
.Y(n_1792)
);

CKINVDCx5p33_ASAP7_75t_R g1793 ( 
.A(n_819),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_756),
.Y(n_1794)
);

CKINVDCx5p33_ASAP7_75t_R g1795 ( 
.A(n_1039),
.Y(n_1795)
);

CKINVDCx5p33_ASAP7_75t_R g1796 ( 
.A(n_1500),
.Y(n_1796)
);

CKINVDCx5p33_ASAP7_75t_R g1797 ( 
.A(n_382),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_652),
.Y(n_1798)
);

CKINVDCx5p33_ASAP7_75t_R g1799 ( 
.A(n_336),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_621),
.Y(n_1800)
);

INVx2_ASAP7_75t_L g1801 ( 
.A(n_1480),
.Y(n_1801)
);

CKINVDCx5p33_ASAP7_75t_R g1802 ( 
.A(n_1564),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_782),
.Y(n_1803)
);

CKINVDCx5p33_ASAP7_75t_R g1804 ( 
.A(n_547),
.Y(n_1804)
);

CKINVDCx20_ASAP7_75t_R g1805 ( 
.A(n_1250),
.Y(n_1805)
);

CKINVDCx20_ASAP7_75t_R g1806 ( 
.A(n_461),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1457),
.Y(n_1807)
);

CKINVDCx5p33_ASAP7_75t_R g1808 ( 
.A(n_1263),
.Y(n_1808)
);

CKINVDCx5p33_ASAP7_75t_R g1809 ( 
.A(n_207),
.Y(n_1809)
);

CKINVDCx5p33_ASAP7_75t_R g1810 ( 
.A(n_1502),
.Y(n_1810)
);

CKINVDCx5p33_ASAP7_75t_R g1811 ( 
.A(n_1481),
.Y(n_1811)
);

CKINVDCx14_ASAP7_75t_R g1812 ( 
.A(n_779),
.Y(n_1812)
);

INVx1_ASAP7_75t_SL g1813 ( 
.A(n_1499),
.Y(n_1813)
);

CKINVDCx5p33_ASAP7_75t_R g1814 ( 
.A(n_1036),
.Y(n_1814)
);

CKINVDCx5p33_ASAP7_75t_R g1815 ( 
.A(n_733),
.Y(n_1815)
);

INVx2_ASAP7_75t_SL g1816 ( 
.A(n_1540),
.Y(n_1816)
);

HB1xp67_ASAP7_75t_L g1817 ( 
.A(n_1048),
.Y(n_1817)
);

INVx1_ASAP7_75t_SL g1818 ( 
.A(n_1046),
.Y(n_1818)
);

BUFx6f_ASAP7_75t_L g1819 ( 
.A(n_927),
.Y(n_1819)
);

CKINVDCx5p33_ASAP7_75t_R g1820 ( 
.A(n_19),
.Y(n_1820)
);

INVx1_ASAP7_75t_SL g1821 ( 
.A(n_1542),
.Y(n_1821)
);

CKINVDCx5p33_ASAP7_75t_R g1822 ( 
.A(n_258),
.Y(n_1822)
);

CKINVDCx5p33_ASAP7_75t_R g1823 ( 
.A(n_123),
.Y(n_1823)
);

BUFx10_ASAP7_75t_L g1824 ( 
.A(n_322),
.Y(n_1824)
);

CKINVDCx5p33_ASAP7_75t_R g1825 ( 
.A(n_204),
.Y(n_1825)
);

BUFx2_ASAP7_75t_L g1826 ( 
.A(n_224),
.Y(n_1826)
);

INVx2_ASAP7_75t_SL g1827 ( 
.A(n_1122),
.Y(n_1827)
);

CKINVDCx5p33_ASAP7_75t_R g1828 ( 
.A(n_1208),
.Y(n_1828)
);

BUFx6f_ASAP7_75t_L g1829 ( 
.A(n_939),
.Y(n_1829)
);

CKINVDCx5p33_ASAP7_75t_R g1830 ( 
.A(n_800),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_137),
.Y(n_1831)
);

CKINVDCx5p33_ASAP7_75t_R g1832 ( 
.A(n_1622),
.Y(n_1832)
);

CKINVDCx5p33_ASAP7_75t_R g1833 ( 
.A(n_1342),
.Y(n_1833)
);

CKINVDCx5p33_ASAP7_75t_R g1834 ( 
.A(n_1573),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1457),
.Y(n_1835)
);

CKINVDCx16_ASAP7_75t_R g1836 ( 
.A(n_1022),
.Y(n_1836)
);

CKINVDCx5p33_ASAP7_75t_R g1837 ( 
.A(n_1360),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_968),
.Y(n_1838)
);

CKINVDCx20_ASAP7_75t_R g1839 ( 
.A(n_1023),
.Y(n_1839)
);

CKINVDCx5p33_ASAP7_75t_R g1840 ( 
.A(n_693),
.Y(n_1840)
);

CKINVDCx5p33_ASAP7_75t_R g1841 ( 
.A(n_424),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1471),
.Y(n_1842)
);

CKINVDCx5p33_ASAP7_75t_R g1843 ( 
.A(n_986),
.Y(n_1843)
);

CKINVDCx5p33_ASAP7_75t_R g1844 ( 
.A(n_1539),
.Y(n_1844)
);

BUFx6f_ASAP7_75t_L g1845 ( 
.A(n_1574),
.Y(n_1845)
);

CKINVDCx5p33_ASAP7_75t_R g1846 ( 
.A(n_72),
.Y(n_1846)
);

INVx2_ASAP7_75t_SL g1847 ( 
.A(n_1089),
.Y(n_1847)
);

INVx2_ASAP7_75t_SL g1848 ( 
.A(n_53),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1161),
.Y(n_1849)
);

CKINVDCx16_ASAP7_75t_R g1850 ( 
.A(n_143),
.Y(n_1850)
);

CKINVDCx20_ASAP7_75t_R g1851 ( 
.A(n_924),
.Y(n_1851)
);

CKINVDCx5p33_ASAP7_75t_R g1852 ( 
.A(n_993),
.Y(n_1852)
);

CKINVDCx5p33_ASAP7_75t_R g1853 ( 
.A(n_690),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1510),
.Y(n_1854)
);

INVx1_ASAP7_75t_SL g1855 ( 
.A(n_176),
.Y(n_1855)
);

CKINVDCx5p33_ASAP7_75t_R g1856 ( 
.A(n_229),
.Y(n_1856)
);

CKINVDCx5p33_ASAP7_75t_R g1857 ( 
.A(n_136),
.Y(n_1857)
);

BUFx2_ASAP7_75t_L g1858 ( 
.A(n_545),
.Y(n_1858)
);

CKINVDCx5p33_ASAP7_75t_R g1859 ( 
.A(n_449),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1484),
.Y(n_1860)
);

INVxp67_ASAP7_75t_L g1861 ( 
.A(n_722),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_768),
.Y(n_1862)
);

CKINVDCx5p33_ASAP7_75t_R g1863 ( 
.A(n_1343),
.Y(n_1863)
);

INVx2_ASAP7_75t_L g1864 ( 
.A(n_1020),
.Y(n_1864)
);

BUFx10_ASAP7_75t_L g1865 ( 
.A(n_531),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1545),
.Y(n_1866)
);

CKINVDCx5p33_ASAP7_75t_R g1867 ( 
.A(n_1447),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1341),
.Y(n_1868)
);

CKINVDCx5p33_ASAP7_75t_R g1869 ( 
.A(n_290),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1535),
.Y(n_1870)
);

CKINVDCx5p33_ASAP7_75t_R g1871 ( 
.A(n_109),
.Y(n_1871)
);

CKINVDCx5p33_ASAP7_75t_R g1872 ( 
.A(n_1515),
.Y(n_1872)
);

CKINVDCx5p33_ASAP7_75t_R g1873 ( 
.A(n_1538),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1373),
.Y(n_1874)
);

CKINVDCx5p33_ASAP7_75t_R g1875 ( 
.A(n_114),
.Y(n_1875)
);

CKINVDCx5p33_ASAP7_75t_R g1876 ( 
.A(n_544),
.Y(n_1876)
);

CKINVDCx5p33_ASAP7_75t_R g1877 ( 
.A(n_992),
.Y(n_1877)
);

CKINVDCx5p33_ASAP7_75t_R g1878 ( 
.A(n_134),
.Y(n_1878)
);

CKINVDCx5p33_ASAP7_75t_R g1879 ( 
.A(n_601),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1000),
.Y(n_1880)
);

CKINVDCx5p33_ASAP7_75t_R g1881 ( 
.A(n_580),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1558),
.Y(n_1882)
);

CKINVDCx5p33_ASAP7_75t_R g1883 ( 
.A(n_718),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_927),
.Y(n_1884)
);

CKINVDCx5p33_ASAP7_75t_R g1885 ( 
.A(n_1527),
.Y(n_1885)
);

CKINVDCx5p33_ASAP7_75t_R g1886 ( 
.A(n_610),
.Y(n_1886)
);

CKINVDCx5p33_ASAP7_75t_R g1887 ( 
.A(n_1447),
.Y(n_1887)
);

CKINVDCx5p33_ASAP7_75t_R g1888 ( 
.A(n_1528),
.Y(n_1888)
);

CKINVDCx5p33_ASAP7_75t_R g1889 ( 
.A(n_605),
.Y(n_1889)
);

CKINVDCx5p33_ASAP7_75t_R g1890 ( 
.A(n_1200),
.Y(n_1890)
);

CKINVDCx5p33_ASAP7_75t_R g1891 ( 
.A(n_368),
.Y(n_1891)
);

BUFx2_ASAP7_75t_L g1892 ( 
.A(n_1254),
.Y(n_1892)
);

CKINVDCx5p33_ASAP7_75t_R g1893 ( 
.A(n_798),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_915),
.Y(n_1894)
);

CKINVDCx5p33_ASAP7_75t_R g1895 ( 
.A(n_1446),
.Y(n_1895)
);

CKINVDCx5p33_ASAP7_75t_R g1896 ( 
.A(n_283),
.Y(n_1896)
);

CKINVDCx5p33_ASAP7_75t_R g1897 ( 
.A(n_332),
.Y(n_1897)
);

CKINVDCx5p33_ASAP7_75t_R g1898 ( 
.A(n_541),
.Y(n_1898)
);

CKINVDCx5p33_ASAP7_75t_R g1899 ( 
.A(n_123),
.Y(n_1899)
);

CKINVDCx5p33_ASAP7_75t_R g1900 ( 
.A(n_127),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_512),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_4),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_282),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1536),
.Y(n_1904)
);

CKINVDCx5p33_ASAP7_75t_R g1905 ( 
.A(n_1061),
.Y(n_1905)
);

CKINVDCx5p33_ASAP7_75t_R g1906 ( 
.A(n_441),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_332),
.Y(n_1907)
);

CKINVDCx5p33_ASAP7_75t_R g1908 ( 
.A(n_1309),
.Y(n_1908)
);

CKINVDCx5p33_ASAP7_75t_R g1909 ( 
.A(n_1348),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_636),
.Y(n_1910)
);

CKINVDCx20_ASAP7_75t_R g1911 ( 
.A(n_46),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_333),
.Y(n_1912)
);

CKINVDCx20_ASAP7_75t_R g1913 ( 
.A(n_931),
.Y(n_1913)
);

CKINVDCx5p33_ASAP7_75t_R g1914 ( 
.A(n_1019),
.Y(n_1914)
);

CKINVDCx20_ASAP7_75t_R g1915 ( 
.A(n_890),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1617),
.Y(n_1916)
);

CKINVDCx5p33_ASAP7_75t_R g1917 ( 
.A(n_1536),
.Y(n_1917)
);

CKINVDCx5p33_ASAP7_75t_R g1918 ( 
.A(n_347),
.Y(n_1918)
);

CKINVDCx5p33_ASAP7_75t_R g1919 ( 
.A(n_528),
.Y(n_1919)
);

CKINVDCx5p33_ASAP7_75t_R g1920 ( 
.A(n_723),
.Y(n_1920)
);

CKINVDCx20_ASAP7_75t_R g1921 ( 
.A(n_1201),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1572),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1048),
.Y(n_1923)
);

CKINVDCx5p33_ASAP7_75t_R g1924 ( 
.A(n_896),
.Y(n_1924)
);

BUFx8_ASAP7_75t_SL g1925 ( 
.A(n_1288),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_986),
.Y(n_1926)
);

CKINVDCx5p33_ASAP7_75t_R g1927 ( 
.A(n_1128),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_648),
.Y(n_1928)
);

INVx1_ASAP7_75t_SL g1929 ( 
.A(n_202),
.Y(n_1929)
);

BUFx6f_ASAP7_75t_L g1930 ( 
.A(n_471),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_831),
.Y(n_1931)
);

CKINVDCx5p33_ASAP7_75t_R g1932 ( 
.A(n_247),
.Y(n_1932)
);

CKINVDCx5p33_ASAP7_75t_R g1933 ( 
.A(n_1454),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_420),
.Y(n_1934)
);

CKINVDCx20_ASAP7_75t_R g1935 ( 
.A(n_734),
.Y(n_1935)
);

CKINVDCx16_ASAP7_75t_R g1936 ( 
.A(n_378),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_792),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_848),
.Y(n_1938)
);

BUFx6f_ASAP7_75t_L g1939 ( 
.A(n_1425),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_418),
.Y(n_1940)
);

INVx2_ASAP7_75t_L g1941 ( 
.A(n_604),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_473),
.Y(n_1942)
);

CKINVDCx5p33_ASAP7_75t_R g1943 ( 
.A(n_291),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1245),
.Y(n_1944)
);

CKINVDCx16_ASAP7_75t_R g1945 ( 
.A(n_1256),
.Y(n_1945)
);

CKINVDCx5p33_ASAP7_75t_R g1946 ( 
.A(n_1112),
.Y(n_1946)
);

CKINVDCx5p33_ASAP7_75t_R g1947 ( 
.A(n_325),
.Y(n_1947)
);

CKINVDCx5p33_ASAP7_75t_R g1948 ( 
.A(n_1602),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_348),
.Y(n_1949)
);

CKINVDCx20_ASAP7_75t_R g1950 ( 
.A(n_714),
.Y(n_1950)
);

CKINVDCx20_ASAP7_75t_R g1951 ( 
.A(n_1469),
.Y(n_1951)
);

CKINVDCx20_ASAP7_75t_R g1952 ( 
.A(n_77),
.Y(n_1952)
);

CKINVDCx5p33_ASAP7_75t_R g1953 ( 
.A(n_443),
.Y(n_1953)
);

BUFx2_ASAP7_75t_L g1954 ( 
.A(n_709),
.Y(n_1954)
);

INVx1_ASAP7_75t_SL g1955 ( 
.A(n_368),
.Y(n_1955)
);

CKINVDCx5p33_ASAP7_75t_R g1956 ( 
.A(n_596),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_733),
.Y(n_1957)
);

BUFx6f_ASAP7_75t_L g1958 ( 
.A(n_1535),
.Y(n_1958)
);

CKINVDCx5p33_ASAP7_75t_R g1959 ( 
.A(n_768),
.Y(n_1959)
);

CKINVDCx5p33_ASAP7_75t_R g1960 ( 
.A(n_831),
.Y(n_1960)
);

CKINVDCx20_ASAP7_75t_R g1961 ( 
.A(n_79),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_954),
.Y(n_1962)
);

CKINVDCx5p33_ASAP7_75t_R g1963 ( 
.A(n_1252),
.Y(n_1963)
);

CKINVDCx5p33_ASAP7_75t_R g1964 ( 
.A(n_1540),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1488),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_22),
.Y(n_1966)
);

CKINVDCx5p33_ASAP7_75t_R g1967 ( 
.A(n_1213),
.Y(n_1967)
);

BUFx6f_ASAP7_75t_L g1968 ( 
.A(n_400),
.Y(n_1968)
);

BUFx6f_ASAP7_75t_L g1969 ( 
.A(n_871),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1516),
.Y(n_1970)
);

CKINVDCx5p33_ASAP7_75t_R g1971 ( 
.A(n_1154),
.Y(n_1971)
);

CKINVDCx5p33_ASAP7_75t_R g1972 ( 
.A(n_1346),
.Y(n_1972)
);

CKINVDCx5p33_ASAP7_75t_R g1973 ( 
.A(n_1135),
.Y(n_1973)
);

CKINVDCx5p33_ASAP7_75t_R g1974 ( 
.A(n_1467),
.Y(n_1974)
);

CKINVDCx5p33_ASAP7_75t_R g1975 ( 
.A(n_66),
.Y(n_1975)
);

CKINVDCx16_ASAP7_75t_R g1976 ( 
.A(n_515),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1551),
.Y(n_1977)
);

CKINVDCx5p33_ASAP7_75t_R g1978 ( 
.A(n_610),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1483),
.Y(n_1979)
);

CKINVDCx5p33_ASAP7_75t_R g1980 ( 
.A(n_1576),
.Y(n_1980)
);

CKINVDCx5p33_ASAP7_75t_R g1981 ( 
.A(n_318),
.Y(n_1981)
);

CKINVDCx5p33_ASAP7_75t_R g1982 ( 
.A(n_221),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1512),
.Y(n_1983)
);

CKINVDCx5p33_ASAP7_75t_R g1984 ( 
.A(n_1349),
.Y(n_1984)
);

CKINVDCx5p33_ASAP7_75t_R g1985 ( 
.A(n_1280),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_350),
.Y(n_1986)
);

HB1xp67_ASAP7_75t_L g1987 ( 
.A(n_1248),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_421),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_514),
.Y(n_1989)
);

CKINVDCx20_ASAP7_75t_R g1990 ( 
.A(n_1284),
.Y(n_1990)
);

CKINVDCx5p33_ASAP7_75t_R g1991 ( 
.A(n_342),
.Y(n_1991)
);

CKINVDCx5p33_ASAP7_75t_R g1992 ( 
.A(n_1211),
.Y(n_1992)
);

CKINVDCx5p33_ASAP7_75t_R g1993 ( 
.A(n_516),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1578),
.Y(n_1994)
);

CKINVDCx20_ASAP7_75t_R g1995 ( 
.A(n_1113),
.Y(n_1995)
);

CKINVDCx5p33_ASAP7_75t_R g1996 ( 
.A(n_1496),
.Y(n_1996)
);

CKINVDCx5p33_ASAP7_75t_R g1997 ( 
.A(n_808),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1378),
.Y(n_1998)
);

CKINVDCx5p33_ASAP7_75t_R g1999 ( 
.A(n_913),
.Y(n_1999)
);

CKINVDCx5p33_ASAP7_75t_R g2000 ( 
.A(n_1028),
.Y(n_2000)
);

INVx2_ASAP7_75t_L g2001 ( 
.A(n_1616),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1397),
.Y(n_2002)
);

CKINVDCx5p33_ASAP7_75t_R g2003 ( 
.A(n_454),
.Y(n_2003)
);

CKINVDCx5p33_ASAP7_75t_R g2004 ( 
.A(n_1056),
.Y(n_2004)
);

CKINVDCx5p33_ASAP7_75t_R g2005 ( 
.A(n_1361),
.Y(n_2005)
);

CKINVDCx5p33_ASAP7_75t_R g2006 ( 
.A(n_1260),
.Y(n_2006)
);

CKINVDCx5p33_ASAP7_75t_R g2007 ( 
.A(n_1052),
.Y(n_2007)
);

BUFx5_ASAP7_75t_L g2008 ( 
.A(n_222),
.Y(n_2008)
);

CKINVDCx5p33_ASAP7_75t_R g2009 ( 
.A(n_1483),
.Y(n_2009)
);

CKINVDCx5p33_ASAP7_75t_R g2010 ( 
.A(n_1501),
.Y(n_2010)
);

CKINVDCx20_ASAP7_75t_R g2011 ( 
.A(n_985),
.Y(n_2011)
);

CKINVDCx5p33_ASAP7_75t_R g2012 ( 
.A(n_175),
.Y(n_2012)
);

CKINVDCx5p33_ASAP7_75t_R g2013 ( 
.A(n_32),
.Y(n_2013)
);

CKINVDCx5p33_ASAP7_75t_R g2014 ( 
.A(n_1313),
.Y(n_2014)
);

BUFx3_ASAP7_75t_L g2015 ( 
.A(n_263),
.Y(n_2015)
);

BUFx10_ASAP7_75t_L g2016 ( 
.A(n_298),
.Y(n_2016)
);

BUFx2_ASAP7_75t_L g2017 ( 
.A(n_894),
.Y(n_2017)
);

CKINVDCx5p33_ASAP7_75t_R g2018 ( 
.A(n_1524),
.Y(n_2018)
);

INVx2_ASAP7_75t_SL g2019 ( 
.A(n_702),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1485),
.Y(n_2020)
);

CKINVDCx5p33_ASAP7_75t_R g2021 ( 
.A(n_636),
.Y(n_2021)
);

INVx1_ASAP7_75t_SL g2022 ( 
.A(n_99),
.Y(n_2022)
);

CKINVDCx5p33_ASAP7_75t_R g2023 ( 
.A(n_1014),
.Y(n_2023)
);

CKINVDCx5p33_ASAP7_75t_R g2024 ( 
.A(n_859),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1554),
.Y(n_2025)
);

CKINVDCx5p33_ASAP7_75t_R g2026 ( 
.A(n_218),
.Y(n_2026)
);

CKINVDCx5p33_ASAP7_75t_R g2027 ( 
.A(n_796),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1489),
.Y(n_2028)
);

CKINVDCx5p33_ASAP7_75t_R g2029 ( 
.A(n_1555),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1456),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1318),
.Y(n_2031)
);

CKINVDCx5p33_ASAP7_75t_R g2032 ( 
.A(n_1559),
.Y(n_2032)
);

INVx2_ASAP7_75t_L g2033 ( 
.A(n_991),
.Y(n_2033)
);

CKINVDCx5p33_ASAP7_75t_R g2034 ( 
.A(n_1586),
.Y(n_2034)
);

CKINVDCx5p33_ASAP7_75t_R g2035 ( 
.A(n_130),
.Y(n_2035)
);

INVx2_ASAP7_75t_SL g2036 ( 
.A(n_912),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_897),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1428),
.Y(n_2038)
);

CKINVDCx5p33_ASAP7_75t_R g2039 ( 
.A(n_548),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_820),
.Y(n_2040)
);

CKINVDCx5p33_ASAP7_75t_R g2041 ( 
.A(n_664),
.Y(n_2041)
);

CKINVDCx5p33_ASAP7_75t_R g2042 ( 
.A(n_1142),
.Y(n_2042)
);

BUFx6f_ASAP7_75t_L g2043 ( 
.A(n_1572),
.Y(n_2043)
);

CKINVDCx20_ASAP7_75t_R g2044 ( 
.A(n_440),
.Y(n_2044)
);

INVx2_ASAP7_75t_L g2045 ( 
.A(n_1197),
.Y(n_2045)
);

INVxp33_ASAP7_75t_L g2046 ( 
.A(n_1399),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1459),
.Y(n_2047)
);

CKINVDCx5p33_ASAP7_75t_R g2048 ( 
.A(n_1237),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1273),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_865),
.Y(n_2050)
);

CKINVDCx5p33_ASAP7_75t_R g2051 ( 
.A(n_231),
.Y(n_2051)
);

BUFx10_ASAP7_75t_L g2052 ( 
.A(n_723),
.Y(n_2052)
);

BUFx3_ASAP7_75t_L g2053 ( 
.A(n_447),
.Y(n_2053)
);

INVx2_ASAP7_75t_SL g2054 ( 
.A(n_540),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_1487),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_310),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_651),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_788),
.Y(n_2058)
);

BUFx6f_ASAP7_75t_L g2059 ( 
.A(n_1559),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1603),
.Y(n_2060)
);

CKINVDCx20_ASAP7_75t_R g2061 ( 
.A(n_147),
.Y(n_2061)
);

INVx2_ASAP7_75t_L g2062 ( 
.A(n_1478),
.Y(n_2062)
);

CKINVDCx5p33_ASAP7_75t_R g2063 ( 
.A(n_895),
.Y(n_2063)
);

CKINVDCx5p33_ASAP7_75t_R g2064 ( 
.A(n_274),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_950),
.Y(n_2065)
);

CKINVDCx5p33_ASAP7_75t_R g2066 ( 
.A(n_58),
.Y(n_2066)
);

CKINVDCx20_ASAP7_75t_R g2067 ( 
.A(n_427),
.Y(n_2067)
);

CKINVDCx5p33_ASAP7_75t_R g2068 ( 
.A(n_160),
.Y(n_2068)
);

BUFx3_ASAP7_75t_L g2069 ( 
.A(n_97),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_1240),
.Y(n_2070)
);

CKINVDCx16_ASAP7_75t_R g2071 ( 
.A(n_227),
.Y(n_2071)
);

BUFx6f_ASAP7_75t_L g2072 ( 
.A(n_909),
.Y(n_2072)
);

INVx1_ASAP7_75t_SL g2073 ( 
.A(n_277),
.Y(n_2073)
);

CKINVDCx5p33_ASAP7_75t_R g2074 ( 
.A(n_1225),
.Y(n_2074)
);

BUFx2_ASAP7_75t_L g2075 ( 
.A(n_950),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_867),
.Y(n_2076)
);

CKINVDCx5p33_ASAP7_75t_R g2077 ( 
.A(n_740),
.Y(n_2077)
);

CKINVDCx5p33_ASAP7_75t_R g2078 ( 
.A(n_662),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_299),
.Y(n_2079)
);

CKINVDCx16_ASAP7_75t_R g2080 ( 
.A(n_727),
.Y(n_2080)
);

CKINVDCx20_ASAP7_75t_R g2081 ( 
.A(n_1506),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_574),
.Y(n_2082)
);

INVx2_ASAP7_75t_L g2083 ( 
.A(n_607),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_1352),
.Y(n_2084)
);

CKINVDCx5p33_ASAP7_75t_R g2085 ( 
.A(n_101),
.Y(n_2085)
);

CKINVDCx14_ASAP7_75t_R g2086 ( 
.A(n_451),
.Y(n_2086)
);

CKINVDCx5p33_ASAP7_75t_R g2087 ( 
.A(n_470),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_683),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_1577),
.Y(n_2089)
);

CKINVDCx5p33_ASAP7_75t_R g2090 ( 
.A(n_476),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_946),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_775),
.Y(n_2092)
);

CKINVDCx5p33_ASAP7_75t_R g2093 ( 
.A(n_262),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_1562),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_1057),
.Y(n_2095)
);

BUFx3_ASAP7_75t_L g2096 ( 
.A(n_86),
.Y(n_2096)
);

CKINVDCx5p33_ASAP7_75t_R g2097 ( 
.A(n_283),
.Y(n_2097)
);

CKINVDCx20_ASAP7_75t_R g2098 ( 
.A(n_46),
.Y(n_2098)
);

CKINVDCx5p33_ASAP7_75t_R g2099 ( 
.A(n_1621),
.Y(n_2099)
);

INVx2_ASAP7_75t_L g2100 ( 
.A(n_1616),
.Y(n_2100)
);

CKINVDCx20_ASAP7_75t_R g2101 ( 
.A(n_179),
.Y(n_2101)
);

CKINVDCx5p33_ASAP7_75t_R g2102 ( 
.A(n_997),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_117),
.Y(n_2103)
);

CKINVDCx5p33_ASAP7_75t_R g2104 ( 
.A(n_1197),
.Y(n_2104)
);

INVxp67_ASAP7_75t_L g2105 ( 
.A(n_1156),
.Y(n_2105)
);

CKINVDCx5p33_ASAP7_75t_R g2106 ( 
.A(n_1427),
.Y(n_2106)
);

CKINVDCx5p33_ASAP7_75t_R g2107 ( 
.A(n_1123),
.Y(n_2107)
);

CKINVDCx5p33_ASAP7_75t_R g2108 ( 
.A(n_947),
.Y(n_2108)
);

CKINVDCx16_ASAP7_75t_R g2109 ( 
.A(n_235),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_113),
.Y(n_2110)
);

CKINVDCx5p33_ASAP7_75t_R g2111 ( 
.A(n_108),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_152),
.Y(n_2112)
);

INVx2_ASAP7_75t_SL g2113 ( 
.A(n_739),
.Y(n_2113)
);

CKINVDCx5p33_ASAP7_75t_R g2114 ( 
.A(n_1393),
.Y(n_2114)
);

CKINVDCx5p33_ASAP7_75t_R g2115 ( 
.A(n_209),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_91),
.Y(n_2116)
);

CKINVDCx20_ASAP7_75t_R g2117 ( 
.A(n_1494),
.Y(n_2117)
);

CKINVDCx5p33_ASAP7_75t_R g2118 ( 
.A(n_1445),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_253),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_769),
.Y(n_2120)
);

CKINVDCx5p33_ASAP7_75t_R g2121 ( 
.A(n_1465),
.Y(n_2121)
);

CKINVDCx5p33_ASAP7_75t_R g2122 ( 
.A(n_423),
.Y(n_2122)
);

CKINVDCx5p33_ASAP7_75t_R g2123 ( 
.A(n_284),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_968),
.Y(n_2124)
);

CKINVDCx5p33_ASAP7_75t_R g2125 ( 
.A(n_1125),
.Y(n_2125)
);

INVxp67_ASAP7_75t_L g2126 ( 
.A(n_1531),
.Y(n_2126)
);

CKINVDCx5p33_ASAP7_75t_R g2127 ( 
.A(n_740),
.Y(n_2127)
);

CKINVDCx5p33_ASAP7_75t_R g2128 ( 
.A(n_1511),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_1497),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_1070),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_1579),
.Y(n_2131)
);

CKINVDCx20_ASAP7_75t_R g2132 ( 
.A(n_815),
.Y(n_2132)
);

CKINVDCx20_ASAP7_75t_R g2133 ( 
.A(n_37),
.Y(n_2133)
);

CKINVDCx5p33_ASAP7_75t_R g2134 ( 
.A(n_413),
.Y(n_2134)
);

CKINVDCx5p33_ASAP7_75t_R g2135 ( 
.A(n_1493),
.Y(n_2135)
);

CKINVDCx5p33_ASAP7_75t_R g2136 ( 
.A(n_520),
.Y(n_2136)
);

CKINVDCx5p33_ASAP7_75t_R g2137 ( 
.A(n_313),
.Y(n_2137)
);

CKINVDCx5p33_ASAP7_75t_R g2138 ( 
.A(n_700),
.Y(n_2138)
);

CKINVDCx5p33_ASAP7_75t_R g2139 ( 
.A(n_1445),
.Y(n_2139)
);

CKINVDCx20_ASAP7_75t_R g2140 ( 
.A(n_896),
.Y(n_2140)
);

BUFx2_ASAP7_75t_L g2141 ( 
.A(n_1133),
.Y(n_2141)
);

CKINVDCx5p33_ASAP7_75t_R g2142 ( 
.A(n_546),
.Y(n_2142)
);

CKINVDCx5p33_ASAP7_75t_R g2143 ( 
.A(n_307),
.Y(n_2143)
);

CKINVDCx5p33_ASAP7_75t_R g2144 ( 
.A(n_94),
.Y(n_2144)
);

BUFx6f_ASAP7_75t_L g2145 ( 
.A(n_346),
.Y(n_2145)
);

CKINVDCx5p33_ASAP7_75t_R g2146 ( 
.A(n_680),
.Y(n_2146)
);

CKINVDCx5p33_ASAP7_75t_R g2147 ( 
.A(n_191),
.Y(n_2147)
);

CKINVDCx5p33_ASAP7_75t_R g2148 ( 
.A(n_431),
.Y(n_2148)
);

CKINVDCx5p33_ASAP7_75t_R g2149 ( 
.A(n_573),
.Y(n_2149)
);

CKINVDCx5p33_ASAP7_75t_R g2150 ( 
.A(n_282),
.Y(n_2150)
);

CKINVDCx5p33_ASAP7_75t_R g2151 ( 
.A(n_802),
.Y(n_2151)
);

CKINVDCx20_ASAP7_75t_R g2152 ( 
.A(n_848),
.Y(n_2152)
);

CKINVDCx5p33_ASAP7_75t_R g2153 ( 
.A(n_842),
.Y(n_2153)
);

BUFx10_ASAP7_75t_L g2154 ( 
.A(n_1255),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_169),
.Y(n_2155)
);

INVxp67_ASAP7_75t_L g2156 ( 
.A(n_1214),
.Y(n_2156)
);

CKINVDCx5p33_ASAP7_75t_R g2157 ( 
.A(n_926),
.Y(n_2157)
);

CKINVDCx5p33_ASAP7_75t_R g2158 ( 
.A(n_1490),
.Y(n_2158)
);

CKINVDCx5p33_ASAP7_75t_R g2159 ( 
.A(n_234),
.Y(n_2159)
);

CKINVDCx5p33_ASAP7_75t_R g2160 ( 
.A(n_517),
.Y(n_2160)
);

CKINVDCx5p33_ASAP7_75t_R g2161 ( 
.A(n_1449),
.Y(n_2161)
);

CKINVDCx5p33_ASAP7_75t_R g2162 ( 
.A(n_326),
.Y(n_2162)
);

CKINVDCx5p33_ASAP7_75t_R g2163 ( 
.A(n_583),
.Y(n_2163)
);

INVx2_ASAP7_75t_SL g2164 ( 
.A(n_1472),
.Y(n_2164)
);

CKINVDCx5p33_ASAP7_75t_R g2165 ( 
.A(n_270),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_258),
.Y(n_2166)
);

CKINVDCx5p33_ASAP7_75t_R g2167 ( 
.A(n_1095),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_1204),
.Y(n_2168)
);

BUFx10_ASAP7_75t_L g2169 ( 
.A(n_1453),
.Y(n_2169)
);

CKINVDCx5p33_ASAP7_75t_R g2170 ( 
.A(n_846),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_76),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_1328),
.Y(n_2172)
);

CKINVDCx5p33_ASAP7_75t_R g2173 ( 
.A(n_1569),
.Y(n_2173)
);

CKINVDCx5p33_ASAP7_75t_R g2174 ( 
.A(n_1518),
.Y(n_2174)
);

CKINVDCx5p33_ASAP7_75t_R g2175 ( 
.A(n_1155),
.Y(n_2175)
);

CKINVDCx5p33_ASAP7_75t_R g2176 ( 
.A(n_770),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_1133),
.Y(n_2177)
);

BUFx3_ASAP7_75t_L g2178 ( 
.A(n_1508),
.Y(n_2178)
);

CKINVDCx5p33_ASAP7_75t_R g2179 ( 
.A(n_781),
.Y(n_2179)
);

CKINVDCx5p33_ASAP7_75t_R g2180 ( 
.A(n_663),
.Y(n_2180)
);

CKINVDCx5p33_ASAP7_75t_R g2181 ( 
.A(n_51),
.Y(n_2181)
);

CKINVDCx5p33_ASAP7_75t_R g2182 ( 
.A(n_1078),
.Y(n_2182)
);

CKINVDCx5p33_ASAP7_75t_R g2183 ( 
.A(n_1411),
.Y(n_2183)
);

CKINVDCx5p33_ASAP7_75t_R g2184 ( 
.A(n_1367),
.Y(n_2184)
);

CKINVDCx5p33_ASAP7_75t_R g2185 ( 
.A(n_940),
.Y(n_2185)
);

CKINVDCx5p33_ASAP7_75t_R g2186 ( 
.A(n_1232),
.Y(n_2186)
);

INVxp67_ASAP7_75t_SL g2187 ( 
.A(n_1112),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_581),
.Y(n_2188)
);

CKINVDCx5p33_ASAP7_75t_R g2189 ( 
.A(n_83),
.Y(n_2189)
);

CKINVDCx5p33_ASAP7_75t_R g2190 ( 
.A(n_25),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_451),
.Y(n_2191)
);

CKINVDCx5p33_ASAP7_75t_R g2192 ( 
.A(n_769),
.Y(n_2192)
);

CKINVDCx5p33_ASAP7_75t_R g2193 ( 
.A(n_496),
.Y(n_2193)
);

CKINVDCx5p33_ASAP7_75t_R g2194 ( 
.A(n_1290),
.Y(n_2194)
);

CKINVDCx5p33_ASAP7_75t_R g2195 ( 
.A(n_611),
.Y(n_2195)
);

CKINVDCx5p33_ASAP7_75t_R g2196 ( 
.A(n_881),
.Y(n_2196)
);

CKINVDCx5p33_ASAP7_75t_R g2197 ( 
.A(n_1302),
.Y(n_2197)
);

CKINVDCx5p33_ASAP7_75t_R g2198 ( 
.A(n_1051),
.Y(n_2198)
);

CKINVDCx5p33_ASAP7_75t_R g2199 ( 
.A(n_1237),
.Y(n_2199)
);

BUFx3_ASAP7_75t_L g2200 ( 
.A(n_34),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_260),
.Y(n_2201)
);

CKINVDCx5p33_ASAP7_75t_R g2202 ( 
.A(n_1625),
.Y(n_2202)
);

CKINVDCx5p33_ASAP7_75t_R g2203 ( 
.A(n_278),
.Y(n_2203)
);

CKINVDCx5p33_ASAP7_75t_R g2204 ( 
.A(n_1275),
.Y(n_2204)
);

CKINVDCx5p33_ASAP7_75t_R g2205 ( 
.A(n_1458),
.Y(n_2205)
);

CKINVDCx14_ASAP7_75t_R g2206 ( 
.A(n_429),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_1242),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_105),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_1088),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_909),
.Y(n_2210)
);

CKINVDCx5p33_ASAP7_75t_R g2211 ( 
.A(n_1553),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_494),
.Y(n_2212)
);

CKINVDCx5p33_ASAP7_75t_R g2213 ( 
.A(n_1623),
.Y(n_2213)
);

INVx2_ASAP7_75t_SL g2214 ( 
.A(n_1104),
.Y(n_2214)
);

CKINVDCx5p33_ASAP7_75t_R g2215 ( 
.A(n_1522),
.Y(n_2215)
);

CKINVDCx5p33_ASAP7_75t_R g2216 ( 
.A(n_1568),
.Y(n_2216)
);

CKINVDCx5p33_ASAP7_75t_R g2217 ( 
.A(n_1380),
.Y(n_2217)
);

CKINVDCx5p33_ASAP7_75t_R g2218 ( 
.A(n_1575),
.Y(n_2218)
);

CKINVDCx5p33_ASAP7_75t_R g2219 ( 
.A(n_499),
.Y(n_2219)
);

CKINVDCx5p33_ASAP7_75t_R g2220 ( 
.A(n_490),
.Y(n_2220)
);

BUFx6f_ASAP7_75t_L g2221 ( 
.A(n_361),
.Y(n_2221)
);

CKINVDCx20_ASAP7_75t_R g2222 ( 
.A(n_1376),
.Y(n_2222)
);

CKINVDCx20_ASAP7_75t_R g2223 ( 
.A(n_1571),
.Y(n_2223)
);

CKINVDCx5p33_ASAP7_75t_R g2224 ( 
.A(n_1107),
.Y(n_2224)
);

CKINVDCx5p33_ASAP7_75t_R g2225 ( 
.A(n_1180),
.Y(n_2225)
);

CKINVDCx20_ASAP7_75t_R g2226 ( 
.A(n_1552),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_50),
.Y(n_2227)
);

BUFx3_ASAP7_75t_L g2228 ( 
.A(n_22),
.Y(n_2228)
);

CKINVDCx5p33_ASAP7_75t_R g2229 ( 
.A(n_1019),
.Y(n_2229)
);

CKINVDCx5p33_ASAP7_75t_R g2230 ( 
.A(n_1092),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_691),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_976),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_1395),
.Y(n_2233)
);

CKINVDCx5p33_ASAP7_75t_R g2234 ( 
.A(n_553),
.Y(n_2234)
);

CKINVDCx5p33_ASAP7_75t_R g2235 ( 
.A(n_626),
.Y(n_2235)
);

CKINVDCx5p33_ASAP7_75t_R g2236 ( 
.A(n_99),
.Y(n_2236)
);

CKINVDCx5p33_ASAP7_75t_R g2237 ( 
.A(n_1605),
.Y(n_2237)
);

CKINVDCx5p33_ASAP7_75t_R g2238 ( 
.A(n_384),
.Y(n_2238)
);

INVx1_ASAP7_75t_SL g2239 ( 
.A(n_1100),
.Y(n_2239)
);

CKINVDCx5p33_ASAP7_75t_R g2240 ( 
.A(n_38),
.Y(n_2240)
);

CKINVDCx20_ASAP7_75t_R g2241 ( 
.A(n_1519),
.Y(n_2241)
);

CKINVDCx20_ASAP7_75t_R g2242 ( 
.A(n_214),
.Y(n_2242)
);

CKINVDCx5p33_ASAP7_75t_R g2243 ( 
.A(n_869),
.Y(n_2243)
);

CKINVDCx5p33_ASAP7_75t_R g2244 ( 
.A(n_1601),
.Y(n_2244)
);

CKINVDCx5p33_ASAP7_75t_R g2245 ( 
.A(n_1521),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_275),
.Y(n_2246)
);

CKINVDCx5p33_ASAP7_75t_R g2247 ( 
.A(n_1151),
.Y(n_2247)
);

CKINVDCx5p33_ASAP7_75t_R g2248 ( 
.A(n_952),
.Y(n_2248)
);

CKINVDCx5p33_ASAP7_75t_R g2249 ( 
.A(n_17),
.Y(n_2249)
);

CKINVDCx5p33_ASAP7_75t_R g2250 ( 
.A(n_1533),
.Y(n_2250)
);

CKINVDCx5p33_ASAP7_75t_R g2251 ( 
.A(n_137),
.Y(n_2251)
);

CKINVDCx5p33_ASAP7_75t_R g2252 ( 
.A(n_1242),
.Y(n_2252)
);

CKINVDCx5p33_ASAP7_75t_R g2253 ( 
.A(n_1219),
.Y(n_2253)
);

CKINVDCx5p33_ASAP7_75t_R g2254 ( 
.A(n_1560),
.Y(n_2254)
);

CKINVDCx20_ASAP7_75t_R g2255 ( 
.A(n_669),
.Y(n_2255)
);

CKINVDCx20_ASAP7_75t_R g2256 ( 
.A(n_631),
.Y(n_2256)
);

CKINVDCx5p33_ASAP7_75t_R g2257 ( 
.A(n_1437),
.Y(n_2257)
);

CKINVDCx5p33_ASAP7_75t_R g2258 ( 
.A(n_1451),
.Y(n_2258)
);

CKINVDCx5p33_ASAP7_75t_R g2259 ( 
.A(n_1468),
.Y(n_2259)
);

CKINVDCx5p33_ASAP7_75t_R g2260 ( 
.A(n_1178),
.Y(n_2260)
);

CKINVDCx5p33_ASAP7_75t_R g2261 ( 
.A(n_1486),
.Y(n_2261)
);

CKINVDCx5p33_ASAP7_75t_R g2262 ( 
.A(n_649),
.Y(n_2262)
);

CKINVDCx5p33_ASAP7_75t_R g2263 ( 
.A(n_539),
.Y(n_2263)
);

CKINVDCx5p33_ASAP7_75t_R g2264 ( 
.A(n_687),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_443),
.Y(n_2265)
);

INVx1_ASAP7_75t_SL g2266 ( 
.A(n_1523),
.Y(n_2266)
);

CKINVDCx16_ASAP7_75t_R g2267 ( 
.A(n_1249),
.Y(n_2267)
);

CKINVDCx5p33_ASAP7_75t_R g2268 ( 
.A(n_773),
.Y(n_2268)
);

CKINVDCx20_ASAP7_75t_R g2269 ( 
.A(n_466),
.Y(n_2269)
);

CKINVDCx5p33_ASAP7_75t_R g2270 ( 
.A(n_402),
.Y(n_2270)
);

CKINVDCx5p33_ASAP7_75t_R g2271 ( 
.A(n_1199),
.Y(n_2271)
);

CKINVDCx20_ASAP7_75t_R g2272 ( 
.A(n_940),
.Y(n_2272)
);

INVx1_ASAP7_75t_SL g2273 ( 
.A(n_1191),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_1424),
.Y(n_2274)
);

INVx1_ASAP7_75t_L g2275 ( 
.A(n_1525),
.Y(n_2275)
);

CKINVDCx5p33_ASAP7_75t_R g2276 ( 
.A(n_1220),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_241),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_255),
.Y(n_2278)
);

BUFx10_ASAP7_75t_L g2279 ( 
.A(n_1016),
.Y(n_2279)
);

INVx1_ASAP7_75t_SL g2280 ( 
.A(n_1475),
.Y(n_2280)
);

INVx1_ASAP7_75t_SL g2281 ( 
.A(n_673),
.Y(n_2281)
);

CKINVDCx5p33_ASAP7_75t_R g2282 ( 
.A(n_27),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_960),
.Y(n_2283)
);

CKINVDCx20_ASAP7_75t_R g2284 ( 
.A(n_58),
.Y(n_2284)
);

CKINVDCx5p33_ASAP7_75t_R g2285 ( 
.A(n_1414),
.Y(n_2285)
);

CKINVDCx5p33_ASAP7_75t_R g2286 ( 
.A(n_696),
.Y(n_2286)
);

CKINVDCx5p33_ASAP7_75t_R g2287 ( 
.A(n_127),
.Y(n_2287)
);

INVx2_ASAP7_75t_SL g2288 ( 
.A(n_787),
.Y(n_2288)
);

CKINVDCx5p33_ASAP7_75t_R g2289 ( 
.A(n_328),
.Y(n_2289)
);

CKINVDCx5p33_ASAP7_75t_R g2290 ( 
.A(n_864),
.Y(n_2290)
);

CKINVDCx5p33_ASAP7_75t_R g2291 ( 
.A(n_1607),
.Y(n_2291)
);

INVx2_ASAP7_75t_SL g2292 ( 
.A(n_1184),
.Y(n_2292)
);

CKINVDCx20_ASAP7_75t_R g2293 ( 
.A(n_184),
.Y(n_2293)
);

CKINVDCx14_ASAP7_75t_R g2294 ( 
.A(n_1010),
.Y(n_2294)
);

CKINVDCx5p33_ASAP7_75t_R g2295 ( 
.A(n_318),
.Y(n_2295)
);

CKINVDCx5p33_ASAP7_75t_R g2296 ( 
.A(n_533),
.Y(n_2296)
);

INVx2_ASAP7_75t_SL g2297 ( 
.A(n_340),
.Y(n_2297)
);

CKINVDCx5p33_ASAP7_75t_R g2298 ( 
.A(n_1496),
.Y(n_2298)
);

CKINVDCx5p33_ASAP7_75t_R g2299 ( 
.A(n_1143),
.Y(n_2299)
);

CKINVDCx5p33_ASAP7_75t_R g2300 ( 
.A(n_1226),
.Y(n_2300)
);

CKINVDCx5p33_ASAP7_75t_R g2301 ( 
.A(n_898),
.Y(n_2301)
);

BUFx6f_ASAP7_75t_L g2302 ( 
.A(n_796),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_8),
.Y(n_2303)
);

CKINVDCx5p33_ASAP7_75t_R g2304 ( 
.A(n_1463),
.Y(n_2304)
);

CKINVDCx5p33_ASAP7_75t_R g2305 ( 
.A(n_1092),
.Y(n_2305)
);

CKINVDCx5p33_ASAP7_75t_R g2306 ( 
.A(n_703),
.Y(n_2306)
);

INVx1_ASAP7_75t_L g2307 ( 
.A(n_1565),
.Y(n_2307)
);

CKINVDCx20_ASAP7_75t_R g2308 ( 
.A(n_1458),
.Y(n_2308)
);

CKINVDCx20_ASAP7_75t_R g2309 ( 
.A(n_1543),
.Y(n_2309)
);

CKINVDCx5p33_ASAP7_75t_R g2310 ( 
.A(n_1319),
.Y(n_2310)
);

CKINVDCx5p33_ASAP7_75t_R g2311 ( 
.A(n_1085),
.Y(n_2311)
);

CKINVDCx5p33_ASAP7_75t_R g2312 ( 
.A(n_1566),
.Y(n_2312)
);

CKINVDCx5p33_ASAP7_75t_R g2313 ( 
.A(n_1082),
.Y(n_2313)
);

CKINVDCx5p33_ASAP7_75t_R g2314 ( 
.A(n_639),
.Y(n_2314)
);

CKINVDCx5p33_ASAP7_75t_R g2315 ( 
.A(n_739),
.Y(n_2315)
);

CKINVDCx5p33_ASAP7_75t_R g2316 ( 
.A(n_1523),
.Y(n_2316)
);

INVx1_ASAP7_75t_L g2317 ( 
.A(n_1106),
.Y(n_2317)
);

INVx2_ASAP7_75t_L g2318 ( 
.A(n_525),
.Y(n_2318)
);

CKINVDCx20_ASAP7_75t_R g2319 ( 
.A(n_194),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_144),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_1472),
.Y(n_2321)
);

INVx1_ASAP7_75t_L g2322 ( 
.A(n_685),
.Y(n_2322)
);

INVx2_ASAP7_75t_SL g2323 ( 
.A(n_1438),
.Y(n_2323)
);

BUFx3_ASAP7_75t_L g2324 ( 
.A(n_876),
.Y(n_2324)
);

CKINVDCx5p33_ASAP7_75t_R g2325 ( 
.A(n_181),
.Y(n_2325)
);

INVx1_ASAP7_75t_L g2326 ( 
.A(n_257),
.Y(n_2326)
);

BUFx3_ASAP7_75t_L g2327 ( 
.A(n_28),
.Y(n_2327)
);

BUFx2_ASAP7_75t_L g2328 ( 
.A(n_8),
.Y(n_2328)
);

INVx2_ASAP7_75t_L g2329 ( 
.A(n_577),
.Y(n_2329)
);

HB1xp67_ASAP7_75t_L g2330 ( 
.A(n_1058),
.Y(n_2330)
);

INVx1_ASAP7_75t_SL g2331 ( 
.A(n_573),
.Y(n_2331)
);

CKINVDCx5p33_ASAP7_75t_R g2332 ( 
.A(n_498),
.Y(n_2332)
);

CKINVDCx5p33_ASAP7_75t_R g2333 ( 
.A(n_921),
.Y(n_2333)
);

CKINVDCx20_ASAP7_75t_R g2334 ( 
.A(n_552),
.Y(n_2334)
);

INVx2_ASAP7_75t_L g2335 ( 
.A(n_1611),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_1580),
.Y(n_2336)
);

INVx1_ASAP7_75t_L g2337 ( 
.A(n_898),
.Y(n_2337)
);

INVx1_ASAP7_75t_L g2338 ( 
.A(n_1247),
.Y(n_2338)
);

CKINVDCx14_ASAP7_75t_R g2339 ( 
.A(n_553),
.Y(n_2339)
);

BUFx3_ASAP7_75t_L g2340 ( 
.A(n_892),
.Y(n_2340)
);

CKINVDCx5p33_ASAP7_75t_R g2341 ( 
.A(n_160),
.Y(n_2341)
);

BUFx3_ASAP7_75t_L g2342 ( 
.A(n_171),
.Y(n_2342)
);

HB1xp67_ASAP7_75t_L g2343 ( 
.A(n_719),
.Y(n_2343)
);

INVx1_ASAP7_75t_L g2344 ( 
.A(n_14),
.Y(n_2344)
);

CKINVDCx5p33_ASAP7_75t_R g2345 ( 
.A(n_1128),
.Y(n_2345)
);

INVxp33_ASAP7_75t_SL g2346 ( 
.A(n_6),
.Y(n_2346)
);

CKINVDCx5p33_ASAP7_75t_R g2347 ( 
.A(n_1557),
.Y(n_2347)
);

CKINVDCx5p33_ASAP7_75t_R g2348 ( 
.A(n_881),
.Y(n_2348)
);

CKINVDCx5p33_ASAP7_75t_R g2349 ( 
.A(n_1076),
.Y(n_2349)
);

CKINVDCx5p33_ASAP7_75t_R g2350 ( 
.A(n_1273),
.Y(n_2350)
);

CKINVDCx5p33_ASAP7_75t_R g2351 ( 
.A(n_1338),
.Y(n_2351)
);

INVx1_ASAP7_75t_L g2352 ( 
.A(n_1061),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_486),
.Y(n_2353)
);

BUFx10_ASAP7_75t_L g2354 ( 
.A(n_299),
.Y(n_2354)
);

CKINVDCx5p33_ASAP7_75t_R g2355 ( 
.A(n_134),
.Y(n_2355)
);

CKINVDCx5p33_ASAP7_75t_R g2356 ( 
.A(n_1549),
.Y(n_2356)
);

INVx1_ASAP7_75t_SL g2357 ( 
.A(n_628),
.Y(n_2357)
);

CKINVDCx20_ASAP7_75t_R g2358 ( 
.A(n_282),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_802),
.Y(n_2359)
);

CKINVDCx20_ASAP7_75t_R g2360 ( 
.A(n_1154),
.Y(n_2360)
);

CKINVDCx5p33_ASAP7_75t_R g2361 ( 
.A(n_1012),
.Y(n_2361)
);

CKINVDCx12_ASAP7_75t_R g2362 ( 
.A(n_447),
.Y(n_2362)
);

CKINVDCx5p33_ASAP7_75t_R g2363 ( 
.A(n_86),
.Y(n_2363)
);

INVx1_ASAP7_75t_L g2364 ( 
.A(n_1548),
.Y(n_2364)
);

CKINVDCx5p33_ASAP7_75t_R g2365 ( 
.A(n_88),
.Y(n_2365)
);

CKINVDCx5p33_ASAP7_75t_R g2366 ( 
.A(n_790),
.Y(n_2366)
);

CKINVDCx20_ASAP7_75t_R g2367 ( 
.A(n_754),
.Y(n_2367)
);

INVx1_ASAP7_75t_L g2368 ( 
.A(n_1221),
.Y(n_2368)
);

CKINVDCx20_ASAP7_75t_R g2369 ( 
.A(n_568),
.Y(n_2369)
);

CKINVDCx5p33_ASAP7_75t_R g2370 ( 
.A(n_1064),
.Y(n_2370)
);

INVxp67_ASAP7_75t_L g2371 ( 
.A(n_1014),
.Y(n_2371)
);

INVx1_ASAP7_75t_L g2372 ( 
.A(n_830),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_1470),
.Y(n_2373)
);

INVx1_ASAP7_75t_SL g2374 ( 
.A(n_54),
.Y(n_2374)
);

CKINVDCx5p33_ASAP7_75t_R g2375 ( 
.A(n_220),
.Y(n_2375)
);

CKINVDCx5p33_ASAP7_75t_R g2376 ( 
.A(n_1455),
.Y(n_2376)
);

CKINVDCx5p33_ASAP7_75t_R g2377 ( 
.A(n_852),
.Y(n_2377)
);

INVx1_ASAP7_75t_L g2378 ( 
.A(n_409),
.Y(n_2378)
);

CKINVDCx5p33_ASAP7_75t_R g2379 ( 
.A(n_1460),
.Y(n_2379)
);

INVx1_ASAP7_75t_L g2380 ( 
.A(n_236),
.Y(n_2380)
);

INVx1_ASAP7_75t_L g2381 ( 
.A(n_1526),
.Y(n_2381)
);

BUFx8_ASAP7_75t_SL g2382 ( 
.A(n_238),
.Y(n_2382)
);

CKINVDCx20_ASAP7_75t_R g2383 ( 
.A(n_77),
.Y(n_2383)
);

CKINVDCx5p33_ASAP7_75t_R g2384 ( 
.A(n_403),
.Y(n_2384)
);

CKINVDCx5p33_ASAP7_75t_R g2385 ( 
.A(n_2),
.Y(n_2385)
);

CKINVDCx20_ASAP7_75t_R g2386 ( 
.A(n_854),
.Y(n_2386)
);

CKINVDCx5p33_ASAP7_75t_R g2387 ( 
.A(n_519),
.Y(n_2387)
);

CKINVDCx5p33_ASAP7_75t_R g2388 ( 
.A(n_1541),
.Y(n_2388)
);

CKINVDCx5p33_ASAP7_75t_R g2389 ( 
.A(n_1547),
.Y(n_2389)
);

CKINVDCx5p33_ASAP7_75t_R g2390 ( 
.A(n_1388),
.Y(n_2390)
);

CKINVDCx5p33_ASAP7_75t_R g2391 ( 
.A(n_959),
.Y(n_2391)
);

CKINVDCx5p33_ASAP7_75t_R g2392 ( 
.A(n_584),
.Y(n_2392)
);

BUFx3_ASAP7_75t_L g2393 ( 
.A(n_1450),
.Y(n_2393)
);

BUFx3_ASAP7_75t_L g2394 ( 
.A(n_53),
.Y(n_2394)
);

CKINVDCx5p33_ASAP7_75t_R g2395 ( 
.A(n_925),
.Y(n_2395)
);

CKINVDCx20_ASAP7_75t_R g2396 ( 
.A(n_368),
.Y(n_2396)
);

INVx1_ASAP7_75t_L g2397 ( 
.A(n_1368),
.Y(n_2397)
);

CKINVDCx20_ASAP7_75t_R g2398 ( 
.A(n_1346),
.Y(n_2398)
);

INVx1_ASAP7_75t_L g2399 ( 
.A(n_1135),
.Y(n_2399)
);

CKINVDCx20_ASAP7_75t_R g2400 ( 
.A(n_1444),
.Y(n_2400)
);

INVx2_ASAP7_75t_L g2401 ( 
.A(n_513),
.Y(n_2401)
);

INVx2_ASAP7_75t_L g2402 ( 
.A(n_1473),
.Y(n_2402)
);

INVx1_ASAP7_75t_L g2403 ( 
.A(n_1164),
.Y(n_2403)
);

INVx2_ASAP7_75t_L g2404 ( 
.A(n_1413),
.Y(n_2404)
);

CKINVDCx5p33_ASAP7_75t_R g2405 ( 
.A(n_1205),
.Y(n_2405)
);

CKINVDCx16_ASAP7_75t_R g2406 ( 
.A(n_729),
.Y(n_2406)
);

CKINVDCx5p33_ASAP7_75t_R g2407 ( 
.A(n_1575),
.Y(n_2407)
);

CKINVDCx5p33_ASAP7_75t_R g2408 ( 
.A(n_61),
.Y(n_2408)
);

INVx1_ASAP7_75t_SL g2409 ( 
.A(n_571),
.Y(n_2409)
);

INVx1_ASAP7_75t_L g2410 ( 
.A(n_118),
.Y(n_2410)
);

CKINVDCx5p33_ASAP7_75t_R g2411 ( 
.A(n_1491),
.Y(n_2411)
);

INVx1_ASAP7_75t_L g2412 ( 
.A(n_304),
.Y(n_2412)
);

BUFx10_ASAP7_75t_L g2413 ( 
.A(n_50),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_378),
.Y(n_2414)
);

CKINVDCx5p33_ASAP7_75t_R g2415 ( 
.A(n_1570),
.Y(n_2415)
);

BUFx2_ASAP7_75t_L g2416 ( 
.A(n_1000),
.Y(n_2416)
);

INVx1_ASAP7_75t_SL g2417 ( 
.A(n_1532),
.Y(n_2417)
);

INVx1_ASAP7_75t_L g2418 ( 
.A(n_1504),
.Y(n_2418)
);

INVxp67_ASAP7_75t_L g2419 ( 
.A(n_1591),
.Y(n_2419)
);

INVx2_ASAP7_75t_L g2420 ( 
.A(n_399),
.Y(n_2420)
);

INVx1_ASAP7_75t_L g2421 ( 
.A(n_1617),
.Y(n_2421)
);

INVx1_ASAP7_75t_L g2422 ( 
.A(n_1270),
.Y(n_2422)
);

INVx1_ASAP7_75t_L g2423 ( 
.A(n_805),
.Y(n_2423)
);

INVx1_ASAP7_75t_L g2424 ( 
.A(n_1104),
.Y(n_2424)
);

CKINVDCx5p33_ASAP7_75t_R g2425 ( 
.A(n_1474),
.Y(n_2425)
);

CKINVDCx5p33_ASAP7_75t_R g2426 ( 
.A(n_1563),
.Y(n_2426)
);

INVx1_ASAP7_75t_SL g2427 ( 
.A(n_1390),
.Y(n_2427)
);

INVx2_ASAP7_75t_L g2428 ( 
.A(n_1408),
.Y(n_2428)
);

INVx2_ASAP7_75t_L g2429 ( 
.A(n_428),
.Y(n_2429)
);

CKINVDCx5p33_ASAP7_75t_R g2430 ( 
.A(n_1507),
.Y(n_2430)
);

CKINVDCx5p33_ASAP7_75t_R g2431 ( 
.A(n_444),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_175),
.Y(n_2432)
);

CKINVDCx5p33_ASAP7_75t_R g2433 ( 
.A(n_872),
.Y(n_2433)
);

INVx1_ASAP7_75t_SL g2434 ( 
.A(n_1233),
.Y(n_2434)
);

CKINVDCx16_ASAP7_75t_R g2435 ( 
.A(n_123),
.Y(n_2435)
);

CKINVDCx20_ASAP7_75t_R g2436 ( 
.A(n_1109),
.Y(n_2436)
);

INVx1_ASAP7_75t_L g2437 ( 
.A(n_1520),
.Y(n_2437)
);

INVx1_ASAP7_75t_L g2438 ( 
.A(n_1469),
.Y(n_2438)
);

BUFx10_ASAP7_75t_L g2439 ( 
.A(n_1567),
.Y(n_2439)
);

CKINVDCx5p33_ASAP7_75t_R g2440 ( 
.A(n_358),
.Y(n_2440)
);

CKINVDCx5p33_ASAP7_75t_R g2441 ( 
.A(n_1244),
.Y(n_2441)
);

CKINVDCx20_ASAP7_75t_R g2442 ( 
.A(n_1160),
.Y(n_2442)
);

CKINVDCx5p33_ASAP7_75t_R g2443 ( 
.A(n_580),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_1497),
.Y(n_2444)
);

CKINVDCx5p33_ASAP7_75t_R g2445 ( 
.A(n_1117),
.Y(n_2445)
);

CKINVDCx5p33_ASAP7_75t_R g2446 ( 
.A(n_1358),
.Y(n_2446)
);

CKINVDCx5p33_ASAP7_75t_R g2447 ( 
.A(n_1550),
.Y(n_2447)
);

INVx1_ASAP7_75t_L g2448 ( 
.A(n_3),
.Y(n_2448)
);

INVx2_ASAP7_75t_L g2449 ( 
.A(n_935),
.Y(n_2449)
);

INVx1_ASAP7_75t_SL g2450 ( 
.A(n_1436),
.Y(n_2450)
);

CKINVDCx5p33_ASAP7_75t_R g2451 ( 
.A(n_1477),
.Y(n_2451)
);

INVxp67_ASAP7_75t_L g2452 ( 
.A(n_1509),
.Y(n_2452)
);

INVx1_ASAP7_75t_L g2453 ( 
.A(n_286),
.Y(n_2453)
);

HB1xp67_ASAP7_75t_L g2454 ( 
.A(n_1317),
.Y(n_2454)
);

BUFx10_ASAP7_75t_L g2455 ( 
.A(n_817),
.Y(n_2455)
);

BUFx5_ASAP7_75t_L g2456 ( 
.A(n_179),
.Y(n_2456)
);

CKINVDCx5p33_ASAP7_75t_R g2457 ( 
.A(n_1546),
.Y(n_2457)
);

CKINVDCx5p33_ASAP7_75t_R g2458 ( 
.A(n_223),
.Y(n_2458)
);

CKINVDCx5p33_ASAP7_75t_R g2459 ( 
.A(n_810),
.Y(n_2459)
);

CKINVDCx5p33_ASAP7_75t_R g2460 ( 
.A(n_1471),
.Y(n_2460)
);

INVx1_ASAP7_75t_L g2461 ( 
.A(n_377),
.Y(n_2461)
);

INVx1_ASAP7_75t_L g2462 ( 
.A(n_1230),
.Y(n_2462)
);

BUFx6f_ASAP7_75t_L g2463 ( 
.A(n_1044),
.Y(n_2463)
);

INVx2_ASAP7_75t_L g2464 ( 
.A(n_999),
.Y(n_2464)
);

INVx1_ASAP7_75t_L g2465 ( 
.A(n_183),
.Y(n_2465)
);

CKINVDCx5p33_ASAP7_75t_R g2466 ( 
.A(n_824),
.Y(n_2466)
);

BUFx10_ASAP7_75t_L g2467 ( 
.A(n_113),
.Y(n_2467)
);

CKINVDCx5p33_ASAP7_75t_R g2468 ( 
.A(n_727),
.Y(n_2468)
);

INVxp67_ASAP7_75t_SL g2469 ( 
.A(n_1765),
.Y(n_2469)
);

INVx1_ASAP7_75t_L g2470 ( 
.A(n_2008),
.Y(n_2470)
);

INVx1_ASAP7_75t_L g2471 ( 
.A(n_2008),
.Y(n_2471)
);

CKINVDCx5p33_ASAP7_75t_R g2472 ( 
.A(n_2382),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_2008),
.Y(n_2473)
);

HB1xp67_ASAP7_75t_L g2474 ( 
.A(n_2362),
.Y(n_2474)
);

INVx1_ASAP7_75t_L g2475 ( 
.A(n_2008),
.Y(n_2475)
);

INVx1_ASAP7_75t_L g2476 ( 
.A(n_2008),
.Y(n_2476)
);

CKINVDCx20_ASAP7_75t_R g2477 ( 
.A(n_1812),
.Y(n_2477)
);

CKINVDCx20_ASAP7_75t_R g2478 ( 
.A(n_2086),
.Y(n_2478)
);

CKINVDCx20_ASAP7_75t_R g2479 ( 
.A(n_2206),
.Y(n_2479)
);

INVx2_ASAP7_75t_L g2480 ( 
.A(n_2456),
.Y(n_2480)
);

CKINVDCx16_ASAP7_75t_R g2481 ( 
.A(n_1775),
.Y(n_2481)
);

INVx1_ASAP7_75t_L g2482 ( 
.A(n_2456),
.Y(n_2482)
);

INVx1_ASAP7_75t_L g2483 ( 
.A(n_2456),
.Y(n_2483)
);

CKINVDCx5p33_ASAP7_75t_R g2484 ( 
.A(n_1787),
.Y(n_2484)
);

INVxp33_ASAP7_75t_L g2485 ( 
.A(n_1826),
.Y(n_2485)
);

CKINVDCx5p33_ASAP7_75t_R g2486 ( 
.A(n_1925),
.Y(n_2486)
);

INVx2_ASAP7_75t_L g2487 ( 
.A(n_2456),
.Y(n_2487)
);

BUFx3_ASAP7_75t_L g2488 ( 
.A(n_2015),
.Y(n_2488)
);

CKINVDCx20_ASAP7_75t_R g2489 ( 
.A(n_2294),
.Y(n_2489)
);

CKINVDCx5p33_ASAP7_75t_R g2490 ( 
.A(n_1850),
.Y(n_2490)
);

INVx1_ASAP7_75t_L g2491 ( 
.A(n_2465),
.Y(n_2491)
);

INVx1_ASAP7_75t_L g2492 ( 
.A(n_1632),
.Y(n_2492)
);

INVx1_ASAP7_75t_L g2493 ( 
.A(n_1652),
.Y(n_2493)
);

INVxp67_ASAP7_75t_L g2494 ( 
.A(n_2328),
.Y(n_2494)
);

CKINVDCx20_ASAP7_75t_R g2495 ( 
.A(n_2339),
.Y(n_2495)
);

INVxp67_ASAP7_75t_SL g2496 ( 
.A(n_1640),
.Y(n_2496)
);

INVx2_ASAP7_75t_L g2497 ( 
.A(n_1666),
.Y(n_2497)
);

INVx1_ASAP7_75t_L g2498 ( 
.A(n_1683),
.Y(n_2498)
);

NAND2xp33_ASAP7_75t_R g2499 ( 
.A(n_2346),
.B(n_0),
.Y(n_2499)
);

INVx1_ASAP7_75t_L g2500 ( 
.A(n_1709),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_2461),
.Y(n_2501)
);

CKINVDCx20_ASAP7_75t_R g2502 ( 
.A(n_1681),
.Y(n_2502)
);

CKINVDCx5p33_ASAP7_75t_R g2503 ( 
.A(n_2071),
.Y(n_2503)
);

INVx2_ASAP7_75t_L g2504 ( 
.A(n_1758),
.Y(n_2504)
);

CKINVDCx5p33_ASAP7_75t_R g2505 ( 
.A(n_2109),
.Y(n_2505)
);

INVx2_ASAP7_75t_L g2506 ( 
.A(n_1777),
.Y(n_2506)
);

INVx1_ASAP7_75t_L g2507 ( 
.A(n_1788),
.Y(n_2507)
);

INVxp67_ASAP7_75t_SL g2508 ( 
.A(n_1640),
.Y(n_2508)
);

CKINVDCx5p33_ASAP7_75t_R g2509 ( 
.A(n_2435),
.Y(n_2509)
);

CKINVDCx5p33_ASAP7_75t_R g2510 ( 
.A(n_1723),
.Y(n_2510)
);

INVx1_ASAP7_75t_L g2511 ( 
.A(n_1831),
.Y(n_2511)
);

CKINVDCx20_ASAP7_75t_R g2512 ( 
.A(n_1756),
.Y(n_2512)
);

CKINVDCx5p33_ASAP7_75t_R g2513 ( 
.A(n_1773),
.Y(n_2513)
);

CKINVDCx14_ASAP7_75t_R g2514 ( 
.A(n_1687),
.Y(n_2514)
);

INVxp67_ASAP7_75t_SL g2515 ( 
.A(n_2145),
.Y(n_2515)
);

INVxp67_ASAP7_75t_SL g2516 ( 
.A(n_2145),
.Y(n_2516)
);

CKINVDCx20_ASAP7_75t_R g2517 ( 
.A(n_1836),
.Y(n_2517)
);

CKINVDCx20_ASAP7_75t_R g2518 ( 
.A(n_1936),
.Y(n_2518)
);

CKINVDCx20_ASAP7_75t_R g2519 ( 
.A(n_1945),
.Y(n_2519)
);

INVxp67_ASAP7_75t_SL g2520 ( 
.A(n_2145),
.Y(n_2520)
);

INVxp67_ASAP7_75t_L g2521 ( 
.A(n_1766),
.Y(n_2521)
);

CKINVDCx5p33_ASAP7_75t_R g2522 ( 
.A(n_1976),
.Y(n_2522)
);

CKINVDCx20_ASAP7_75t_R g2523 ( 
.A(n_2080),
.Y(n_2523)
);

INVx1_ASAP7_75t_L g2524 ( 
.A(n_1902),
.Y(n_2524)
);

BUFx3_ASAP7_75t_L g2525 ( 
.A(n_2069),
.Y(n_2525)
);

INVx2_ASAP7_75t_L g2526 ( 
.A(n_1903),
.Y(n_2526)
);

INVxp33_ASAP7_75t_L g2527 ( 
.A(n_1817),
.Y(n_2527)
);

CKINVDCx5p33_ASAP7_75t_R g2528 ( 
.A(n_2267),
.Y(n_2528)
);

INVx1_ASAP7_75t_L g2529 ( 
.A(n_1907),
.Y(n_2529)
);

INVx1_ASAP7_75t_L g2530 ( 
.A(n_1912),
.Y(n_2530)
);

INVxp67_ASAP7_75t_SL g2531 ( 
.A(n_2221),
.Y(n_2531)
);

INVxp67_ASAP7_75t_L g2532 ( 
.A(n_1858),
.Y(n_2532)
);

INVx1_ASAP7_75t_L g2533 ( 
.A(n_1949),
.Y(n_2533)
);

INVxp33_ASAP7_75t_SL g2534 ( 
.A(n_1987),
.Y(n_2534)
);

INVxp67_ASAP7_75t_SL g2535 ( 
.A(n_2221),
.Y(n_2535)
);

INVx1_ASAP7_75t_L g2536 ( 
.A(n_1966),
.Y(n_2536)
);

INVx1_ASAP7_75t_L g2537 ( 
.A(n_1986),
.Y(n_2537)
);

CKINVDCx5p33_ASAP7_75t_R g2538 ( 
.A(n_2406),
.Y(n_2538)
);

CKINVDCx5p33_ASAP7_75t_R g2539 ( 
.A(n_1647),
.Y(n_2539)
);

INVx1_ASAP7_75t_L g2540 ( 
.A(n_2056),
.Y(n_2540)
);

INVxp67_ASAP7_75t_SL g2541 ( 
.A(n_2221),
.Y(n_2541)
);

CKINVDCx5p33_ASAP7_75t_R g2542 ( 
.A(n_1650),
.Y(n_2542)
);

INVx1_ASAP7_75t_L g2543 ( 
.A(n_2079),
.Y(n_2543)
);

INVx1_ASAP7_75t_L g2544 ( 
.A(n_2103),
.Y(n_2544)
);

INVx1_ASAP7_75t_L g2545 ( 
.A(n_2110),
.Y(n_2545)
);

INVx1_ASAP7_75t_L g2546 ( 
.A(n_2112),
.Y(n_2546)
);

INVx1_ASAP7_75t_L g2547 ( 
.A(n_2116),
.Y(n_2547)
);

INVx2_ASAP7_75t_L g2548 ( 
.A(n_2119),
.Y(n_2548)
);

INVx2_ASAP7_75t_SL g2549 ( 
.A(n_1824),
.Y(n_2549)
);

INVx1_ASAP7_75t_L g2550 ( 
.A(n_2155),
.Y(n_2550)
);

INVx1_ASAP7_75t_L g2551 ( 
.A(n_2166),
.Y(n_2551)
);

INVx1_ASAP7_75t_L g2552 ( 
.A(n_2171),
.Y(n_2552)
);

INVx1_ASAP7_75t_L g2553 ( 
.A(n_2201),
.Y(n_2553)
);

CKINVDCx5p33_ASAP7_75t_R g2554 ( 
.A(n_1656),
.Y(n_2554)
);

HB1xp67_ASAP7_75t_L g2555 ( 
.A(n_2330),
.Y(n_2555)
);

INVxp67_ASAP7_75t_SL g2556 ( 
.A(n_2343),
.Y(n_2556)
);

INVx1_ASAP7_75t_L g2557 ( 
.A(n_2208),
.Y(n_2557)
);

CKINVDCx5p33_ASAP7_75t_R g2558 ( 
.A(n_1661),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_2227),
.Y(n_2559)
);

BUFx6f_ASAP7_75t_L g2560 ( 
.A(n_1701),
.Y(n_2560)
);

INVx1_ASAP7_75t_L g2561 ( 
.A(n_2246),
.Y(n_2561)
);

INVx1_ASAP7_75t_L g2562 ( 
.A(n_2277),
.Y(n_2562)
);

BUFx2_ASAP7_75t_L g2563 ( 
.A(n_1892),
.Y(n_2563)
);

HB1xp67_ASAP7_75t_L g2564 ( 
.A(n_2454),
.Y(n_2564)
);

INVx1_ASAP7_75t_L g2565 ( 
.A(n_2278),
.Y(n_2565)
);

INVx2_ASAP7_75t_L g2566 ( 
.A(n_2303),
.Y(n_2566)
);

CKINVDCx20_ASAP7_75t_R g2567 ( 
.A(n_1633),
.Y(n_2567)
);

CKINVDCx20_ASAP7_75t_R g2568 ( 
.A(n_1671),
.Y(n_2568)
);

INVxp33_ASAP7_75t_SL g2569 ( 
.A(n_1665),
.Y(n_2569)
);

CKINVDCx5p33_ASAP7_75t_R g2570 ( 
.A(n_1668),
.Y(n_2570)
);

INVx1_ASAP7_75t_L g2571 ( 
.A(n_2320),
.Y(n_2571)
);

CKINVDCx5p33_ASAP7_75t_R g2572 ( 
.A(n_1710),
.Y(n_2572)
);

INVx1_ASAP7_75t_L g2573 ( 
.A(n_2326),
.Y(n_2573)
);

CKINVDCx5p33_ASAP7_75t_R g2574 ( 
.A(n_1711),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_2344),
.Y(n_2575)
);

INVx1_ASAP7_75t_L g2576 ( 
.A(n_2380),
.Y(n_2576)
);

INVxp33_ASAP7_75t_L g2577 ( 
.A(n_1954),
.Y(n_2577)
);

INVx1_ASAP7_75t_L g2578 ( 
.A(n_2453),
.Y(n_2578)
);

INVx1_ASAP7_75t_L g2579 ( 
.A(n_2410),
.Y(n_2579)
);

INVx1_ASAP7_75t_L g2580 ( 
.A(n_2412),
.Y(n_2580)
);

INVx1_ASAP7_75t_L g2581 ( 
.A(n_2432),
.Y(n_2581)
);

CKINVDCx5p33_ASAP7_75t_R g2582 ( 
.A(n_1718),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_2448),
.Y(n_2583)
);

CKINVDCx5p33_ASAP7_75t_R g2584 ( 
.A(n_1719),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_2096),
.Y(n_2585)
);

CKINVDCx5p33_ASAP7_75t_R g2586 ( 
.A(n_1720),
.Y(n_2586)
);

INVx1_ASAP7_75t_L g2587 ( 
.A(n_2200),
.Y(n_2587)
);

CKINVDCx20_ASAP7_75t_R g2588 ( 
.A(n_1698),
.Y(n_2588)
);

CKINVDCx14_ASAP7_75t_R g2589 ( 
.A(n_2017),
.Y(n_2589)
);

CKINVDCx20_ASAP7_75t_R g2590 ( 
.A(n_1700),
.Y(n_2590)
);

BUFx3_ASAP7_75t_L g2591 ( 
.A(n_2228),
.Y(n_2591)
);

INVx1_ASAP7_75t_L g2592 ( 
.A(n_2327),
.Y(n_2592)
);

CKINVDCx20_ASAP7_75t_R g2593 ( 
.A(n_1712),
.Y(n_2593)
);

INVx1_ASAP7_75t_L g2594 ( 
.A(n_2342),
.Y(n_2594)
);

INVx1_ASAP7_75t_L g2595 ( 
.A(n_2394),
.Y(n_2595)
);

INVxp67_ASAP7_75t_SL g2596 ( 
.A(n_1701),
.Y(n_2596)
);

CKINVDCx5p33_ASAP7_75t_R g2597 ( 
.A(n_1724),
.Y(n_2597)
);

CKINVDCx20_ASAP7_75t_R g2598 ( 
.A(n_1713),
.Y(n_2598)
);

INVx1_ASAP7_75t_L g2599 ( 
.A(n_1701),
.Y(n_2599)
);

CKINVDCx5p33_ASAP7_75t_R g2600 ( 
.A(n_1736),
.Y(n_2600)
);

INVx1_ASAP7_75t_L g2601 ( 
.A(n_1749),
.Y(n_2601)
);

INVxp67_ASAP7_75t_L g2602 ( 
.A(n_2075),
.Y(n_2602)
);

INVx1_ASAP7_75t_L g2603 ( 
.A(n_1749),
.Y(n_2603)
);

INVxp67_ASAP7_75t_SL g2604 ( 
.A(n_1759),
.Y(n_2604)
);

CKINVDCx5p33_ASAP7_75t_R g2605 ( 
.A(n_1741),
.Y(n_2605)
);

INVx1_ASAP7_75t_L g2606 ( 
.A(n_1759),
.Y(n_2606)
);

INVx2_ASAP7_75t_L g2607 ( 
.A(n_1759),
.Y(n_2607)
);

INVx1_ASAP7_75t_L g2608 ( 
.A(n_1769),
.Y(n_2608)
);

BUFx3_ASAP7_75t_L g2609 ( 
.A(n_1693),
.Y(n_2609)
);

INVxp67_ASAP7_75t_L g2610 ( 
.A(n_2141),
.Y(n_2610)
);

INVx1_ASAP7_75t_L g2611 ( 
.A(n_1769),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_1769),
.Y(n_2612)
);

INVx1_ASAP7_75t_L g2613 ( 
.A(n_1819),
.Y(n_2613)
);

INVx2_ASAP7_75t_L g2614 ( 
.A(n_2463),
.Y(n_2614)
);

INVxp33_ASAP7_75t_L g2615 ( 
.A(n_2416),
.Y(n_2615)
);

INVx1_ASAP7_75t_SL g2616 ( 
.A(n_2319),
.Y(n_2616)
);

INVx1_ASAP7_75t_L g2617 ( 
.A(n_1829),
.Y(n_2617)
);

INVx1_ASAP7_75t_L g2618 ( 
.A(n_1829),
.Y(n_2618)
);

INVx1_ASAP7_75t_L g2619 ( 
.A(n_1845),
.Y(n_2619)
);

INVx1_ASAP7_75t_L g2620 ( 
.A(n_1845),
.Y(n_2620)
);

CKINVDCx20_ASAP7_75t_R g2621 ( 
.A(n_1761),
.Y(n_2621)
);

HB1xp67_ASAP7_75t_L g2622 ( 
.A(n_1745),
.Y(n_2622)
);

INVxp67_ASAP7_75t_SL g2623 ( 
.A(n_1845),
.Y(n_2623)
);

INVxp67_ASAP7_75t_L g2624 ( 
.A(n_2413),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_1930),
.Y(n_2625)
);

INVx1_ASAP7_75t_L g2626 ( 
.A(n_1930),
.Y(n_2626)
);

INVx1_ASAP7_75t_L g2627 ( 
.A(n_1930),
.Y(n_2627)
);

HB1xp67_ASAP7_75t_L g2628 ( 
.A(n_1750),
.Y(n_2628)
);

INVx1_ASAP7_75t_L g2629 ( 
.A(n_1939),
.Y(n_2629)
);

INVx1_ASAP7_75t_L g2630 ( 
.A(n_1939),
.Y(n_2630)
);

INVx1_ASAP7_75t_L g2631 ( 
.A(n_1939),
.Y(n_2631)
);

INVx1_ASAP7_75t_SL g2632 ( 
.A(n_1689),
.Y(n_2632)
);

INVx1_ASAP7_75t_L g2633 ( 
.A(n_1958),
.Y(n_2633)
);

INVx1_ASAP7_75t_L g2634 ( 
.A(n_1958),
.Y(n_2634)
);

INVx1_ASAP7_75t_L g2635 ( 
.A(n_1958),
.Y(n_2635)
);

INVx1_ASAP7_75t_L g2636 ( 
.A(n_1968),
.Y(n_2636)
);

CKINVDCx5p33_ASAP7_75t_R g2637 ( 
.A(n_1753),
.Y(n_2637)
);

INVxp33_ASAP7_75t_L g2638 ( 
.A(n_2046),
.Y(n_2638)
);

HB1xp67_ASAP7_75t_L g2639 ( 
.A(n_2458),
.Y(n_2639)
);

INVx1_ASAP7_75t_L g2640 ( 
.A(n_1968),
.Y(n_2640)
);

HB1xp67_ASAP7_75t_L g2641 ( 
.A(n_1760),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_1969),
.Y(n_2642)
);

BUFx3_ASAP7_75t_L g2643 ( 
.A(n_1717),
.Y(n_2643)
);

CKINVDCx5p33_ASAP7_75t_R g2644 ( 
.A(n_1790),
.Y(n_2644)
);

INVx1_ASAP7_75t_L g2645 ( 
.A(n_1969),
.Y(n_2645)
);

INVxp33_ASAP7_75t_SL g2646 ( 
.A(n_1799),
.Y(n_2646)
);

BUFx6f_ASAP7_75t_L g2647 ( 
.A(n_2463),
.Y(n_2647)
);

INVxp33_ASAP7_75t_SL g2648 ( 
.A(n_1809),
.Y(n_2648)
);

INVx1_ASAP7_75t_L g2649 ( 
.A(n_1969),
.Y(n_2649)
);

INVxp67_ASAP7_75t_SL g2650 ( 
.A(n_2043),
.Y(n_2650)
);

INVx1_ASAP7_75t_L g2651 ( 
.A(n_2043),
.Y(n_2651)
);

INVx1_ASAP7_75t_L g2652 ( 
.A(n_2059),
.Y(n_2652)
);

CKINVDCx20_ASAP7_75t_R g2653 ( 
.A(n_1786),
.Y(n_2653)
);

CKINVDCx5p33_ASAP7_75t_R g2654 ( 
.A(n_1820),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_2072),
.Y(n_2655)
);

BUFx2_ASAP7_75t_L g2656 ( 
.A(n_1822),
.Y(n_2656)
);

INVx1_ASAP7_75t_L g2657 ( 
.A(n_2072),
.Y(n_2657)
);

INVx1_ASAP7_75t_L g2658 ( 
.A(n_2072),
.Y(n_2658)
);

INVx1_ASAP7_75t_L g2659 ( 
.A(n_2302),
.Y(n_2659)
);

INVx1_ASAP7_75t_L g2660 ( 
.A(n_2302),
.Y(n_2660)
);

INVx1_ASAP7_75t_L g2661 ( 
.A(n_2302),
.Y(n_2661)
);

INVx1_ASAP7_75t_L g2662 ( 
.A(n_1721),
.Y(n_2662)
);

CKINVDCx20_ASAP7_75t_R g2663 ( 
.A(n_1805),
.Y(n_2663)
);

BUFx2_ASAP7_75t_SL g2664 ( 
.A(n_2016),
.Y(n_2664)
);

CKINVDCx20_ASAP7_75t_R g2665 ( 
.A(n_1806),
.Y(n_2665)
);

INVxp33_ASAP7_75t_SL g2666 ( 
.A(n_1823),
.Y(n_2666)
);

INVx1_ASAP7_75t_L g2667 ( 
.A(n_1726),
.Y(n_2667)
);

CKINVDCx5p33_ASAP7_75t_R g2668 ( 
.A(n_1825),
.Y(n_2668)
);

HB1xp67_ASAP7_75t_L g2669 ( 
.A(n_1846),
.Y(n_2669)
);

INVx3_ASAP7_75t_L g2670 ( 
.A(n_1772),
.Y(n_2670)
);

INVx2_ASAP7_75t_L g2671 ( 
.A(n_1789),
.Y(n_2671)
);

INVx1_ASAP7_75t_L g2672 ( 
.A(n_2053),
.Y(n_2672)
);

INVx1_ASAP7_75t_L g2673 ( 
.A(n_2178),
.Y(n_2673)
);

INVx1_ASAP7_75t_L g2674 ( 
.A(n_2324),
.Y(n_2674)
);

INVxp67_ASAP7_75t_L g2675 ( 
.A(n_2016),
.Y(n_2675)
);

INVx1_ASAP7_75t_L g2676 ( 
.A(n_2340),
.Y(n_2676)
);

INVx1_ASAP7_75t_L g2677 ( 
.A(n_2393),
.Y(n_2677)
);

INVxp67_ASAP7_75t_SL g2678 ( 
.A(n_1755),
.Y(n_2678)
);

CKINVDCx16_ASAP7_75t_R g2679 ( 
.A(n_2354),
.Y(n_2679)
);

INVx1_ASAP7_75t_L g2680 ( 
.A(n_2462),
.Y(n_2680)
);

OAI22xp5_ASAP7_75t_L g2681 ( 
.A1(n_2534),
.A2(n_1857),
.B1(n_1869),
.B2(n_1856),
.Y(n_2681)
);

AND2x4_ASAP7_75t_L g2682 ( 
.A(n_2556),
.B(n_1690),
.Y(n_2682)
);

INVx2_ASAP7_75t_L g2683 ( 
.A(n_2607),
.Y(n_2683)
);

INVx6_ASAP7_75t_L g2684 ( 
.A(n_2488),
.Y(n_2684)
);

INVx2_ASAP7_75t_L g2685 ( 
.A(n_2614),
.Y(n_2685)
);

INVx1_ASAP7_75t_L g2686 ( 
.A(n_2596),
.Y(n_2686)
);

BUFx6f_ASAP7_75t_L g2687 ( 
.A(n_2560),
.Y(n_2687)
);

AND2x4_ASAP7_75t_L g2688 ( 
.A(n_2494),
.B(n_1784),
.Y(n_2688)
);

NOR2xp33_ASAP7_75t_L g2689 ( 
.A(n_2569),
.B(n_1848),
.Y(n_2689)
);

BUFx2_ASAP7_75t_L g2690 ( 
.A(n_2502),
.Y(n_2690)
);

BUFx6f_ASAP7_75t_L g2691 ( 
.A(n_2560),
.Y(n_2691)
);

NOR2x1_ASAP7_75t_L g2692 ( 
.A(n_2470),
.B(n_1631),
.Y(n_2692)
);

BUFx2_ASAP7_75t_L g2693 ( 
.A(n_2512),
.Y(n_2693)
);

NAND2xp5_ASAP7_75t_L g2694 ( 
.A(n_2469),
.B(n_2297),
.Y(n_2694)
);

INVx3_ASAP7_75t_L g2695 ( 
.A(n_2647),
.Y(n_2695)
);

INVx4_ASAP7_75t_L g2696 ( 
.A(n_2539),
.Y(n_2696)
);

CKINVDCx5p33_ASAP7_75t_R g2697 ( 
.A(n_2484),
.Y(n_2697)
);

HB1xp67_ASAP7_75t_L g2698 ( 
.A(n_2510),
.Y(n_2698)
);

AOI22xp5_ASAP7_75t_L g2699 ( 
.A1(n_2513),
.A2(n_1875),
.B1(n_1878),
.B2(n_1871),
.Y(n_2699)
);

BUFx2_ASAP7_75t_L g2700 ( 
.A(n_2517),
.Y(n_2700)
);

INVx1_ASAP7_75t_L g2701 ( 
.A(n_2604),
.Y(n_2701)
);

INVx1_ASAP7_75t_L g2702 ( 
.A(n_2623),
.Y(n_2702)
);

INVxp33_ASAP7_75t_SL g2703 ( 
.A(n_2472),
.Y(n_2703)
);

BUFx2_ASAP7_75t_L g2704 ( 
.A(n_2518),
.Y(n_2704)
);

AND2x2_ASAP7_75t_L g2705 ( 
.A(n_2638),
.B(n_2354),
.Y(n_2705)
);

INVx5_ASAP7_75t_L g2706 ( 
.A(n_2549),
.Y(n_2706)
);

INVx2_ASAP7_75t_L g2707 ( 
.A(n_2647),
.Y(n_2707)
);

INVx2_ASAP7_75t_L g2708 ( 
.A(n_2480),
.Y(n_2708)
);

INVx1_ASAP7_75t_L g2709 ( 
.A(n_2650),
.Y(n_2709)
);

INVx2_ASAP7_75t_L g2710 ( 
.A(n_2487),
.Y(n_2710)
);

AOI22xp5_ASAP7_75t_L g2711 ( 
.A1(n_2522),
.A2(n_1896),
.B1(n_1897),
.B2(n_1891),
.Y(n_2711)
);

INVx3_ASAP7_75t_L g2712 ( 
.A(n_2525),
.Y(n_2712)
);

INVx1_ASAP7_75t_L g2713 ( 
.A(n_2496),
.Y(n_2713)
);

INVx3_ASAP7_75t_L g2714 ( 
.A(n_2591),
.Y(n_2714)
);

INVx2_ASAP7_75t_L g2715 ( 
.A(n_2471),
.Y(n_2715)
);

INVx2_ASAP7_75t_L g2716 ( 
.A(n_2473),
.Y(n_2716)
);

NAND2xp5_ASAP7_75t_L g2717 ( 
.A(n_2508),
.B(n_1705),
.Y(n_2717)
);

BUFx6f_ASAP7_75t_L g2718 ( 
.A(n_2497),
.Y(n_2718)
);

OAI22xp5_ASAP7_75t_SL g2719 ( 
.A1(n_2519),
.A2(n_1952),
.B1(n_1961),
.B2(n_1911),
.Y(n_2719)
);

CKINVDCx6p67_ASAP7_75t_R g2720 ( 
.A(n_2477),
.Y(n_2720)
);

NOR2xp33_ASAP7_75t_L g2721 ( 
.A(n_2646),
.B(n_2648),
.Y(n_2721)
);

AND2x4_ASAP7_75t_L g2722 ( 
.A(n_2521),
.B(n_1816),
.Y(n_2722)
);

BUFx6f_ASAP7_75t_L g2723 ( 
.A(n_2504),
.Y(n_2723)
);

INVx1_ASAP7_75t_L g2724 ( 
.A(n_2515),
.Y(n_2724)
);

HB1xp67_ASAP7_75t_L g2725 ( 
.A(n_2528),
.Y(n_2725)
);

HB1xp67_ASAP7_75t_L g2726 ( 
.A(n_2538),
.Y(n_2726)
);

AOI22xp5_ASAP7_75t_L g2727 ( 
.A1(n_2490),
.A2(n_1900),
.B1(n_1918),
.B2(n_1899),
.Y(n_2727)
);

OAI21x1_ASAP7_75t_L g2728 ( 
.A1(n_2475),
.A2(n_1669),
.B(n_1635),
.Y(n_2728)
);

BUFx8_ASAP7_75t_SL g2729 ( 
.A(n_2486),
.Y(n_2729)
);

INVx1_ASAP7_75t_L g2730 ( 
.A(n_2516),
.Y(n_2730)
);

INVx2_ASAP7_75t_L g2731 ( 
.A(n_2476),
.Y(n_2731)
);

INVx6_ASAP7_75t_L g2732 ( 
.A(n_2609),
.Y(n_2732)
);

INVx1_ASAP7_75t_L g2733 ( 
.A(n_2520),
.Y(n_2733)
);

OA21x2_ASAP7_75t_L g2734 ( 
.A1(n_2482),
.A2(n_1704),
.B(n_1676),
.Y(n_2734)
);

INVx3_ASAP7_75t_L g2735 ( 
.A(n_2643),
.Y(n_2735)
);

BUFx8_ASAP7_75t_L g2736 ( 
.A(n_2563),
.Y(n_2736)
);

INVx1_ASAP7_75t_L g2737 ( 
.A(n_2531),
.Y(n_2737)
);

INVx2_ASAP7_75t_L g2738 ( 
.A(n_2483),
.Y(n_2738)
);

BUFx6f_ASAP7_75t_L g2739 ( 
.A(n_2506),
.Y(n_2739)
);

INVx2_ASAP7_75t_L g2740 ( 
.A(n_2599),
.Y(n_2740)
);

AND2x4_ASAP7_75t_L g2741 ( 
.A(n_2532),
.B(n_1827),
.Y(n_2741)
);

INVx2_ASAP7_75t_L g2742 ( 
.A(n_2601),
.Y(n_2742)
);

NAND2xp5_ASAP7_75t_L g2743 ( 
.A(n_2535),
.B(n_1847),
.Y(n_2743)
);

INVx1_ASAP7_75t_L g2744 ( 
.A(n_2541),
.Y(n_2744)
);

AND2x4_ASAP7_75t_L g2745 ( 
.A(n_2602),
.B(n_2019),
.Y(n_2745)
);

CKINVDCx5p33_ASAP7_75t_R g2746 ( 
.A(n_2542),
.Y(n_2746)
);

CKINVDCx5p33_ASAP7_75t_R g2747 ( 
.A(n_2554),
.Y(n_2747)
);

CKINVDCx5p33_ASAP7_75t_R g2748 ( 
.A(n_2558),
.Y(n_2748)
);

OAI22xp5_ASAP7_75t_L g2749 ( 
.A1(n_2514),
.A2(n_1932),
.B1(n_1947),
.B2(n_1943),
.Y(n_2749)
);

AND2x2_ASAP7_75t_L g2750 ( 
.A(n_2656),
.B(n_2413),
.Y(n_2750)
);

INVx2_ASAP7_75t_SL g2751 ( 
.A(n_2570),
.Y(n_2751)
);

INVx3_ASAP7_75t_L g2752 ( 
.A(n_2670),
.Y(n_2752)
);

INVx2_ASAP7_75t_L g2753 ( 
.A(n_2603),
.Y(n_2753)
);

INVx1_ASAP7_75t_L g2754 ( 
.A(n_2606),
.Y(n_2754)
);

INVx2_ASAP7_75t_L g2755 ( 
.A(n_2608),
.Y(n_2755)
);

NOR2xp33_ASAP7_75t_L g2756 ( 
.A(n_2666),
.B(n_1975),
.Y(n_2756)
);

INVx2_ASAP7_75t_L g2757 ( 
.A(n_2611),
.Y(n_2757)
);

NAND2xp5_ASAP7_75t_L g2758 ( 
.A(n_2678),
.B(n_2036),
.Y(n_2758)
);

INVx1_ASAP7_75t_L g2759 ( 
.A(n_2612),
.Y(n_2759)
);

AND2x4_ASAP7_75t_L g2760 ( 
.A(n_2610),
.B(n_2474),
.Y(n_2760)
);

BUFx6f_ASAP7_75t_L g2761 ( 
.A(n_2526),
.Y(n_2761)
);

INVx1_ASAP7_75t_L g2762 ( 
.A(n_2613),
.Y(n_2762)
);

INVx2_ASAP7_75t_L g2763 ( 
.A(n_2617),
.Y(n_2763)
);

OAI21x1_ASAP7_75t_L g2764 ( 
.A1(n_2618),
.A2(n_1737),
.B(n_1734),
.Y(n_2764)
);

BUFx6f_ASAP7_75t_L g2765 ( 
.A(n_2548),
.Y(n_2765)
);

INVx2_ASAP7_75t_SL g2766 ( 
.A(n_2572),
.Y(n_2766)
);

NOR2xp33_ASAP7_75t_SL g2767 ( 
.A(n_2478),
.B(n_1644),
.Y(n_2767)
);

INVx3_ASAP7_75t_L g2768 ( 
.A(n_2670),
.Y(n_2768)
);

INVx1_ASAP7_75t_L g2769 ( 
.A(n_2619),
.Y(n_2769)
);

NOR2x1_ASAP7_75t_L g2770 ( 
.A(n_2620),
.B(n_2625),
.Y(n_2770)
);

INVx2_ASAP7_75t_L g2771 ( 
.A(n_2626),
.Y(n_2771)
);

INVx2_ASAP7_75t_L g2772 ( 
.A(n_2627),
.Y(n_2772)
);

AOI22xp5_ASAP7_75t_L g2773 ( 
.A1(n_2503),
.A2(n_1982),
.B1(n_1991),
.B2(n_1981),
.Y(n_2773)
);

BUFx12f_ASAP7_75t_L g2774 ( 
.A(n_2505),
.Y(n_2774)
);

INVx3_ASAP7_75t_L g2775 ( 
.A(n_2671),
.Y(n_2775)
);

AND2x6_ASAP7_75t_L g2776 ( 
.A(n_2585),
.B(n_1716),
.Y(n_2776)
);

INVx1_ASAP7_75t_L g2777 ( 
.A(n_2629),
.Y(n_2777)
);

INVx1_ASAP7_75t_L g2778 ( 
.A(n_2630),
.Y(n_2778)
);

AND2x6_ASAP7_75t_L g2779 ( 
.A(n_2587),
.B(n_1855),
.Y(n_2779)
);

OA21x2_ASAP7_75t_L g2780 ( 
.A1(n_2631),
.A2(n_1780),
.B(n_1757),
.Y(n_2780)
);

BUFx6f_ASAP7_75t_L g2781 ( 
.A(n_2566),
.Y(n_2781)
);

CKINVDCx11_ASAP7_75t_R g2782 ( 
.A(n_2567),
.Y(n_2782)
);

INVx2_ASAP7_75t_L g2783 ( 
.A(n_2633),
.Y(n_2783)
);

INVx1_ASAP7_75t_L g2784 ( 
.A(n_2634),
.Y(n_2784)
);

INVx4_ASAP7_75t_L g2785 ( 
.A(n_2574),
.Y(n_2785)
);

BUFx6f_ASAP7_75t_L g2786 ( 
.A(n_2635),
.Y(n_2786)
);

INVx2_ASAP7_75t_L g2787 ( 
.A(n_2636),
.Y(n_2787)
);

BUFx3_ASAP7_75t_L g2788 ( 
.A(n_2662),
.Y(n_2788)
);

OAI22x1_ASAP7_75t_SL g2789 ( 
.A1(n_2568),
.A2(n_2098),
.B1(n_2101),
.B2(n_2061),
.Y(n_2789)
);

AOI22x1_ASAP7_75t_SL g2790 ( 
.A1(n_2523),
.A2(n_2242),
.B1(n_2284),
.B2(n_2133),
.Y(n_2790)
);

BUFx6f_ASAP7_75t_L g2791 ( 
.A(n_2640),
.Y(n_2791)
);

INVx1_ASAP7_75t_L g2792 ( 
.A(n_2642),
.Y(n_2792)
);

OAI21x1_ASAP7_75t_L g2793 ( 
.A1(n_2645),
.A2(n_1798),
.B(n_1794),
.Y(n_2793)
);

INVx1_ASAP7_75t_L g2794 ( 
.A(n_2649),
.Y(n_2794)
);

HB1xp67_ASAP7_75t_L g2795 ( 
.A(n_2509),
.Y(n_2795)
);

INVx1_ASAP7_75t_L g2796 ( 
.A(n_2651),
.Y(n_2796)
);

AND2x4_ASAP7_75t_L g2797 ( 
.A(n_2622),
.B(n_2054),
.Y(n_2797)
);

INVx1_ASAP7_75t_L g2798 ( 
.A(n_2652),
.Y(n_2798)
);

AND2x2_ASAP7_75t_L g2799 ( 
.A(n_2628),
.B(n_2467),
.Y(n_2799)
);

AND2x4_ASAP7_75t_L g2800 ( 
.A(n_2639),
.B(n_2113),
.Y(n_2800)
);

BUFx6f_ASAP7_75t_L g2801 ( 
.A(n_2655),
.Y(n_2801)
);

AND2x2_ASAP7_75t_L g2802 ( 
.A(n_2641),
.B(n_2467),
.Y(n_2802)
);

AND2x4_ASAP7_75t_L g2803 ( 
.A(n_2669),
.B(n_2555),
.Y(n_2803)
);

OAI21x1_ASAP7_75t_L g2804 ( 
.A1(n_2657),
.A2(n_1864),
.B(n_1801),
.Y(n_2804)
);

INVx6_ASAP7_75t_L g2805 ( 
.A(n_2679),
.Y(n_2805)
);

INVx3_ASAP7_75t_L g2806 ( 
.A(n_2658),
.Y(n_2806)
);

AND2x4_ASAP7_75t_L g2807 ( 
.A(n_2564),
.B(n_2624),
.Y(n_2807)
);

AND2x4_ASAP7_75t_L g2808 ( 
.A(n_2675),
.B(n_2164),
.Y(n_2808)
);

BUFx6f_ASAP7_75t_L g2809 ( 
.A(n_2659),
.Y(n_2809)
);

CKINVDCx5p33_ASAP7_75t_R g2810 ( 
.A(n_2582),
.Y(n_2810)
);

INVx1_ASAP7_75t_L g2811 ( 
.A(n_2660),
.Y(n_2811)
);

BUFx6f_ASAP7_75t_L g2812 ( 
.A(n_2661),
.Y(n_2812)
);

OAI22x1_ASAP7_75t_SL g2813 ( 
.A1(n_2588),
.A2(n_2358),
.B1(n_2383),
.B2(n_2293),
.Y(n_2813)
);

INVx2_ASAP7_75t_L g2814 ( 
.A(n_2491),
.Y(n_2814)
);

INVx2_ASAP7_75t_L g2815 ( 
.A(n_2492),
.Y(n_2815)
);

INVx2_ASAP7_75t_L g2816 ( 
.A(n_2493),
.Y(n_2816)
);

INVx1_ASAP7_75t_L g2817 ( 
.A(n_2680),
.Y(n_2817)
);

NAND2xp5_ASAP7_75t_L g2818 ( 
.A(n_2584),
.B(n_2214),
.Y(n_2818)
);

BUFx2_ASAP7_75t_L g2819 ( 
.A(n_2479),
.Y(n_2819)
);

OAI22xp5_ASAP7_75t_L g2820 ( 
.A1(n_2589),
.A2(n_2012),
.B1(n_2026),
.B2(n_2013),
.Y(n_2820)
);

INVx2_ASAP7_75t_L g2821 ( 
.A(n_2498),
.Y(n_2821)
);

INVx2_ASAP7_75t_L g2822 ( 
.A(n_2500),
.Y(n_2822)
);

INVx2_ASAP7_75t_L g2823 ( 
.A(n_2501),
.Y(n_2823)
);

NAND2xp5_ASAP7_75t_L g2824 ( 
.A(n_2586),
.B(n_2288),
.Y(n_2824)
);

INVx4_ASAP7_75t_L g2825 ( 
.A(n_2597),
.Y(n_2825)
);

BUFx6f_ASAP7_75t_L g2826 ( 
.A(n_2507),
.Y(n_2826)
);

NAND2xp5_ASAP7_75t_L g2827 ( 
.A(n_2600),
.B(n_2292),
.Y(n_2827)
);

AOI22xp5_ASAP7_75t_L g2828 ( 
.A1(n_2481),
.A2(n_2051),
.B1(n_2064),
.B2(n_2035),
.Y(n_2828)
);

BUFx6f_ASAP7_75t_L g2829 ( 
.A(n_2511),
.Y(n_2829)
);

OAI22xp5_ASAP7_75t_SL g2830 ( 
.A1(n_2489),
.A2(n_2396),
.B1(n_1839),
.B2(n_1851),
.Y(n_2830)
);

INVx3_ASAP7_75t_L g2831 ( 
.A(n_2592),
.Y(n_2831)
);

INVx1_ASAP7_75t_L g2832 ( 
.A(n_2524),
.Y(n_2832)
);

AOI22xp5_ASAP7_75t_L g2833 ( 
.A1(n_2495),
.A2(n_2068),
.B1(n_2085),
.B2(n_2066),
.Y(n_2833)
);

INVx3_ASAP7_75t_L g2834 ( 
.A(n_2594),
.Y(n_2834)
);

INVx2_ASAP7_75t_L g2835 ( 
.A(n_2529),
.Y(n_2835)
);

INVx2_ASAP7_75t_L g2836 ( 
.A(n_2530),
.Y(n_2836)
);

AND2x4_ASAP7_75t_L g2837 ( 
.A(n_2595),
.B(n_2323),
.Y(n_2837)
);

BUFx3_ASAP7_75t_L g2838 ( 
.A(n_2667),
.Y(n_2838)
);

NAND2xp5_ASAP7_75t_L g2839 ( 
.A(n_2605),
.B(n_2093),
.Y(n_2839)
);

BUFx2_ASAP7_75t_L g2840 ( 
.A(n_2637),
.Y(n_2840)
);

NAND2xp5_ASAP7_75t_L g2841 ( 
.A(n_2644),
.B(n_2097),
.Y(n_2841)
);

INVx2_ASAP7_75t_L g2842 ( 
.A(n_2533),
.Y(n_2842)
);

BUFx3_ASAP7_75t_L g2843 ( 
.A(n_2672),
.Y(n_2843)
);

INVx1_ASAP7_75t_L g2844 ( 
.A(n_2536),
.Y(n_2844)
);

INVx2_ASAP7_75t_L g2845 ( 
.A(n_2537),
.Y(n_2845)
);

AOI22xp5_ASAP7_75t_L g2846 ( 
.A1(n_2654),
.A2(n_2115),
.B1(n_2123),
.B2(n_2111),
.Y(n_2846)
);

OAI22xp5_ASAP7_75t_L g2847 ( 
.A1(n_2577),
.A2(n_2143),
.B1(n_2144),
.B2(n_2137),
.Y(n_2847)
);

NAND2xp5_ASAP7_75t_L g2848 ( 
.A(n_2668),
.B(n_2147),
.Y(n_2848)
);

INVx1_ASAP7_75t_L g2849 ( 
.A(n_2540),
.Y(n_2849)
);

INVx4_ASAP7_75t_L g2850 ( 
.A(n_2673),
.Y(n_2850)
);

INVx1_ASAP7_75t_L g2851 ( 
.A(n_2543),
.Y(n_2851)
);

INVx3_ASAP7_75t_L g2852 ( 
.A(n_2674),
.Y(n_2852)
);

INVx1_ASAP7_75t_L g2853 ( 
.A(n_2544),
.Y(n_2853)
);

INVx2_ASAP7_75t_L g2854 ( 
.A(n_2545),
.Y(n_2854)
);

NOR2xp33_ASAP7_75t_R g2855 ( 
.A(n_2697),
.B(n_2746),
.Y(n_2855)
);

INVx1_ASAP7_75t_L g2856 ( 
.A(n_2817),
.Y(n_2856)
);

BUFx6f_ASAP7_75t_L g2857 ( 
.A(n_2687),
.Y(n_2857)
);

CKINVDCx5p33_ASAP7_75t_R g2858 ( 
.A(n_2747),
.Y(n_2858)
);

CKINVDCx5p33_ASAP7_75t_R g2859 ( 
.A(n_2748),
.Y(n_2859)
);

CKINVDCx5p33_ASAP7_75t_R g2860 ( 
.A(n_2810),
.Y(n_2860)
);

BUFx3_ASAP7_75t_L g2861 ( 
.A(n_2684),
.Y(n_2861)
);

INVx2_ASAP7_75t_SL g2862 ( 
.A(n_2705),
.Y(n_2862)
);

CKINVDCx5p33_ASAP7_75t_R g2863 ( 
.A(n_2782),
.Y(n_2863)
);

CKINVDCx5p33_ASAP7_75t_R g2864 ( 
.A(n_2729),
.Y(n_2864)
);

CKINVDCx5p33_ASAP7_75t_R g2865 ( 
.A(n_2703),
.Y(n_2865)
);

CKINVDCx20_ASAP7_75t_R g2866 ( 
.A(n_2720),
.Y(n_2866)
);

INVx2_ASAP7_75t_L g2867 ( 
.A(n_2707),
.Y(n_2867)
);

CKINVDCx20_ASAP7_75t_R g2868 ( 
.A(n_2690),
.Y(n_2868)
);

INVx2_ASAP7_75t_L g2869 ( 
.A(n_2683),
.Y(n_2869)
);

CKINVDCx5p33_ASAP7_75t_R g2870 ( 
.A(n_2774),
.Y(n_2870)
);

CKINVDCx5p33_ASAP7_75t_R g2871 ( 
.A(n_2840),
.Y(n_2871)
);

CKINVDCx20_ASAP7_75t_R g2872 ( 
.A(n_2693),
.Y(n_2872)
);

CKINVDCx5p33_ASAP7_75t_R g2873 ( 
.A(n_2696),
.Y(n_2873)
);

INVx1_ASAP7_75t_L g2874 ( 
.A(n_2832),
.Y(n_2874)
);

CKINVDCx5p33_ASAP7_75t_R g2875 ( 
.A(n_2785),
.Y(n_2875)
);

CKINVDCx5p33_ASAP7_75t_R g2876 ( 
.A(n_2825),
.Y(n_2876)
);

NOR2xp33_ASAP7_75t_R g2877 ( 
.A(n_2751),
.B(n_2590),
.Y(n_2877)
);

INVxp67_ASAP7_75t_L g2878 ( 
.A(n_2756),
.Y(n_2878)
);

INVx2_ASAP7_75t_L g2879 ( 
.A(n_2685),
.Y(n_2879)
);

CKINVDCx5p33_ASAP7_75t_R g2880 ( 
.A(n_2766),
.Y(n_2880)
);

NAND2xp5_ASAP7_75t_SL g2881 ( 
.A(n_2706),
.B(n_2721),
.Y(n_2881)
);

BUFx10_ASAP7_75t_L g2882 ( 
.A(n_2805),
.Y(n_2882)
);

CKINVDCx5p33_ASAP7_75t_R g2883 ( 
.A(n_2700),
.Y(n_2883)
);

CKINVDCx5p33_ASAP7_75t_R g2884 ( 
.A(n_2704),
.Y(n_2884)
);

BUFx3_ASAP7_75t_L g2885 ( 
.A(n_2732),
.Y(n_2885)
);

BUFx3_ASAP7_75t_L g2886 ( 
.A(n_2712),
.Y(n_2886)
);

INVx1_ASAP7_75t_L g2887 ( 
.A(n_2844),
.Y(n_2887)
);

INVx1_ASAP7_75t_L g2888 ( 
.A(n_2849),
.Y(n_2888)
);

CKINVDCx5p33_ASAP7_75t_R g2889 ( 
.A(n_2819),
.Y(n_2889)
);

CKINVDCx20_ASAP7_75t_R g2890 ( 
.A(n_2795),
.Y(n_2890)
);

INVx3_ASAP7_75t_L g2891 ( 
.A(n_2715),
.Y(n_2891)
);

INVx3_ASAP7_75t_L g2892 ( 
.A(n_2716),
.Y(n_2892)
);

AOI21x1_ASAP7_75t_L g2893 ( 
.A1(n_2708),
.A2(n_2710),
.B(n_2731),
.Y(n_2893)
);

AND2x2_ASAP7_75t_L g2894 ( 
.A(n_2799),
.B(n_2802),
.Y(n_2894)
);

NOR2xp33_ASAP7_75t_R g2895 ( 
.A(n_2713),
.B(n_2593),
.Y(n_2895)
);

NAND2xp5_ASAP7_75t_L g2896 ( 
.A(n_2686),
.B(n_2676),
.Y(n_2896)
);

CKINVDCx5p33_ASAP7_75t_R g2897 ( 
.A(n_2698),
.Y(n_2897)
);

CKINVDCx5p33_ASAP7_75t_R g2898 ( 
.A(n_2725),
.Y(n_2898)
);

CKINVDCx5p33_ASAP7_75t_R g2899 ( 
.A(n_2726),
.Y(n_2899)
);

CKINVDCx5p33_ASAP7_75t_R g2900 ( 
.A(n_2839),
.Y(n_2900)
);

INVx1_ASAP7_75t_L g2901 ( 
.A(n_2851),
.Y(n_2901)
);

INVx1_ASAP7_75t_L g2902 ( 
.A(n_2853),
.Y(n_2902)
);

INVx1_ASAP7_75t_L g2903 ( 
.A(n_2826),
.Y(n_2903)
);

CKINVDCx5p33_ASAP7_75t_R g2904 ( 
.A(n_2841),
.Y(n_2904)
);

BUFx6f_ASAP7_75t_L g2905 ( 
.A(n_2691),
.Y(n_2905)
);

CKINVDCx5p33_ASAP7_75t_R g2906 ( 
.A(n_2848),
.Y(n_2906)
);

CKINVDCx5p33_ASAP7_75t_R g2907 ( 
.A(n_2830),
.Y(n_2907)
);

INVx1_ASAP7_75t_L g2908 ( 
.A(n_2829),
.Y(n_2908)
);

CKINVDCx5p33_ASAP7_75t_R g2909 ( 
.A(n_2736),
.Y(n_2909)
);

CKINVDCx5p33_ASAP7_75t_R g2910 ( 
.A(n_2735),
.Y(n_2910)
);

CKINVDCx20_ASAP7_75t_R g2911 ( 
.A(n_2719),
.Y(n_2911)
);

CKINVDCx5p33_ASAP7_75t_R g2912 ( 
.A(n_2714),
.Y(n_2912)
);

INVx1_ASAP7_75t_L g2913 ( 
.A(n_2738),
.Y(n_2913)
);

BUFx2_ASAP7_75t_L g2914 ( 
.A(n_2776),
.Y(n_2914)
);

CKINVDCx16_ASAP7_75t_R g2915 ( 
.A(n_2767),
.Y(n_2915)
);

CKINVDCx5p33_ASAP7_75t_R g2916 ( 
.A(n_2749),
.Y(n_2916)
);

BUFx2_ASAP7_75t_L g2917 ( 
.A(n_2776),
.Y(n_2917)
);

NAND2xp5_ASAP7_75t_SL g2918 ( 
.A(n_2689),
.B(n_2615),
.Y(n_2918)
);

AND2x6_ASAP7_75t_L g2919 ( 
.A(n_2750),
.B(n_2692),
.Y(n_2919)
);

CKINVDCx5p33_ASAP7_75t_R g2920 ( 
.A(n_2820),
.Y(n_2920)
);

AND3x2_ASAP7_75t_L g2921 ( 
.A(n_2807),
.B(n_2105),
.C(n_1861),
.Y(n_2921)
);

CKINVDCx5p33_ASAP7_75t_R g2922 ( 
.A(n_2846),
.Y(n_2922)
);

BUFx3_ASAP7_75t_L g2923 ( 
.A(n_2788),
.Y(n_2923)
);

AND2x6_ASAP7_75t_L g2924 ( 
.A(n_2682),
.B(n_1630),
.Y(n_2924)
);

CKINVDCx20_ASAP7_75t_R g2925 ( 
.A(n_2833),
.Y(n_2925)
);

NAND2xp5_ASAP7_75t_L g2926 ( 
.A(n_2701),
.B(n_2677),
.Y(n_2926)
);

CKINVDCx5p33_ASAP7_75t_R g2927 ( 
.A(n_2818),
.Y(n_2927)
);

CKINVDCx5p33_ASAP7_75t_R g2928 ( 
.A(n_2824),
.Y(n_2928)
);

CKINVDCx5p33_ASAP7_75t_R g2929 ( 
.A(n_2827),
.Y(n_2929)
);

INVx1_ASAP7_75t_L g2930 ( 
.A(n_2838),
.Y(n_2930)
);

CKINVDCx5p33_ASAP7_75t_R g2931 ( 
.A(n_2789),
.Y(n_2931)
);

CKINVDCx5p33_ASAP7_75t_R g2932 ( 
.A(n_2813),
.Y(n_2932)
);

INVxp67_ASAP7_75t_SL g2933 ( 
.A(n_2752),
.Y(n_2933)
);

NAND2xp33_ASAP7_75t_R g2934 ( 
.A(n_2803),
.B(n_2760),
.Y(n_2934)
);

CKINVDCx20_ASAP7_75t_R g2935 ( 
.A(n_2828),
.Y(n_2935)
);

CKINVDCx20_ASAP7_75t_R g2936 ( 
.A(n_2790),
.Y(n_2936)
);

INVx1_ASAP7_75t_L g2937 ( 
.A(n_2843),
.Y(n_2937)
);

CKINVDCx20_ASAP7_75t_R g2938 ( 
.A(n_2699),
.Y(n_2938)
);

BUFx6f_ASAP7_75t_L g2939 ( 
.A(n_2728),
.Y(n_2939)
);

CKINVDCx5p33_ASAP7_75t_R g2940 ( 
.A(n_2711),
.Y(n_2940)
);

INVx2_ASAP7_75t_L g2941 ( 
.A(n_2718),
.Y(n_2941)
);

CKINVDCx5p33_ASAP7_75t_R g2942 ( 
.A(n_2727),
.Y(n_2942)
);

INVxp33_ASAP7_75t_L g2943 ( 
.A(n_2847),
.Y(n_2943)
);

BUFx6f_ASAP7_75t_L g2944 ( 
.A(n_2764),
.Y(n_2944)
);

CKINVDCx5p33_ASAP7_75t_R g2945 ( 
.A(n_2773),
.Y(n_2945)
);

INVx1_ASAP7_75t_L g2946 ( 
.A(n_2723),
.Y(n_2946)
);

CKINVDCx5p33_ASAP7_75t_R g2947 ( 
.A(n_2681),
.Y(n_2947)
);

CKINVDCx5p33_ASAP7_75t_R g2948 ( 
.A(n_2724),
.Y(n_2948)
);

CKINVDCx5p33_ASAP7_75t_R g2949 ( 
.A(n_2730),
.Y(n_2949)
);

CKINVDCx16_ASAP7_75t_R g2950 ( 
.A(n_2797),
.Y(n_2950)
);

XOR2xp5_ASAP7_75t_L g2951 ( 
.A(n_2800),
.B(n_2598),
.Y(n_2951)
);

CKINVDCx5p33_ASAP7_75t_R g2952 ( 
.A(n_2733),
.Y(n_2952)
);

INVx1_ASAP7_75t_L g2953 ( 
.A(n_2739),
.Y(n_2953)
);

INVx1_ASAP7_75t_L g2954 ( 
.A(n_2761),
.Y(n_2954)
);

AND2x2_ASAP7_75t_L g2955 ( 
.A(n_2768),
.B(n_2664),
.Y(n_2955)
);

INVx1_ASAP7_75t_L g2956 ( 
.A(n_2765),
.Y(n_2956)
);

BUFx3_ASAP7_75t_L g2957 ( 
.A(n_2734),
.Y(n_2957)
);

CKINVDCx5p33_ASAP7_75t_R g2958 ( 
.A(n_2737),
.Y(n_2958)
);

CKINVDCx5p33_ASAP7_75t_R g2959 ( 
.A(n_2744),
.Y(n_2959)
);

CKINVDCx5p33_ASAP7_75t_R g2960 ( 
.A(n_2702),
.Y(n_2960)
);

INVx1_ASAP7_75t_L g2961 ( 
.A(n_2781),
.Y(n_2961)
);

CKINVDCx5p33_ASAP7_75t_R g2962 ( 
.A(n_2709),
.Y(n_2962)
);

INVx2_ASAP7_75t_L g2963 ( 
.A(n_2740),
.Y(n_2963)
);

CKINVDCx20_ASAP7_75t_R g2964 ( 
.A(n_2694),
.Y(n_2964)
);

NOR2xp67_ASAP7_75t_L g2965 ( 
.A(n_2775),
.B(n_2546),
.Y(n_2965)
);

HB1xp67_ASAP7_75t_L g2966 ( 
.A(n_2695),
.Y(n_2966)
);

AND3x2_ASAP7_75t_L g2967 ( 
.A(n_2808),
.B(n_2156),
.C(n_2126),
.Y(n_2967)
);

INVx1_ASAP7_75t_L g2968 ( 
.A(n_2780),
.Y(n_2968)
);

CKINVDCx5p33_ASAP7_75t_R g2969 ( 
.A(n_2779),
.Y(n_2969)
);

CKINVDCx5p33_ASAP7_75t_R g2970 ( 
.A(n_2779),
.Y(n_2970)
);

CKINVDCx5p33_ASAP7_75t_R g2971 ( 
.A(n_2758),
.Y(n_2971)
);

CKINVDCx5p33_ASAP7_75t_R g2972 ( 
.A(n_2722),
.Y(n_2972)
);

CKINVDCx20_ASAP7_75t_R g2973 ( 
.A(n_2717),
.Y(n_2973)
);

CKINVDCx5p33_ASAP7_75t_R g2974 ( 
.A(n_2741),
.Y(n_2974)
);

CKINVDCx16_ASAP7_75t_R g2975 ( 
.A(n_2688),
.Y(n_2975)
);

INVx2_ASAP7_75t_L g2976 ( 
.A(n_2742),
.Y(n_2976)
);

NOR2xp67_ASAP7_75t_L g2977 ( 
.A(n_2850),
.B(n_2547),
.Y(n_2977)
);

CKINVDCx5p33_ASAP7_75t_R g2978 ( 
.A(n_2745),
.Y(n_2978)
);

CKINVDCx20_ASAP7_75t_R g2979 ( 
.A(n_2743),
.Y(n_2979)
);

BUFx10_ASAP7_75t_L g2980 ( 
.A(n_2837),
.Y(n_2980)
);

CKINVDCx5p33_ASAP7_75t_R g2981 ( 
.A(n_2786),
.Y(n_2981)
);

INVx1_ASAP7_75t_L g2982 ( 
.A(n_2814),
.Y(n_2982)
);

NOR2xp33_ASAP7_75t_R g2983 ( 
.A(n_2831),
.B(n_2621),
.Y(n_2983)
);

BUFx2_ASAP7_75t_L g2984 ( 
.A(n_2834),
.Y(n_2984)
);

BUFx2_ASAP7_75t_L g2985 ( 
.A(n_2852),
.Y(n_2985)
);

NAND2xp5_ASAP7_75t_L g2986 ( 
.A(n_2754),
.B(n_2550),
.Y(n_2986)
);

CKINVDCx5p33_ASAP7_75t_R g2987 ( 
.A(n_2791),
.Y(n_2987)
);

INVx1_ASAP7_75t_L g2988 ( 
.A(n_2815),
.Y(n_2988)
);

CKINVDCx16_ASAP7_75t_R g2989 ( 
.A(n_2770),
.Y(n_2989)
);

INVx1_ASAP7_75t_L g2990 ( 
.A(n_2816),
.Y(n_2990)
);

BUFx16f_ASAP7_75t_R g2991 ( 
.A(n_2821),
.Y(n_2991)
);

NAND2xp5_ASAP7_75t_L g2992 ( 
.A(n_2759),
.B(n_2551),
.Y(n_2992)
);

CKINVDCx5p33_ASAP7_75t_R g2993 ( 
.A(n_2801),
.Y(n_2993)
);

INVx2_ASAP7_75t_SL g2994 ( 
.A(n_2809),
.Y(n_2994)
);

CKINVDCx5p33_ASAP7_75t_R g2995 ( 
.A(n_2812),
.Y(n_2995)
);

INVx1_ASAP7_75t_L g2996 ( 
.A(n_2822),
.Y(n_2996)
);

NAND2xp33_ASAP7_75t_R g2997 ( 
.A(n_2823),
.B(n_2150),
.Y(n_2997)
);

INVx1_ASAP7_75t_L g2998 ( 
.A(n_2835),
.Y(n_2998)
);

INVx2_ASAP7_75t_SL g2999 ( 
.A(n_2836),
.Y(n_2999)
);

CKINVDCx20_ASAP7_75t_R g3000 ( 
.A(n_2842),
.Y(n_3000)
);

CKINVDCx5p33_ASAP7_75t_R g3001 ( 
.A(n_2845),
.Y(n_3001)
);

BUFx6f_ASAP7_75t_L g3002 ( 
.A(n_2793),
.Y(n_3002)
);

CKINVDCx20_ASAP7_75t_R g3003 ( 
.A(n_2854),
.Y(n_3003)
);

INVx2_ASAP7_75t_L g3004 ( 
.A(n_2753),
.Y(n_3004)
);

HB1xp67_ASAP7_75t_L g3005 ( 
.A(n_2806),
.Y(n_3005)
);

CKINVDCx5p33_ASAP7_75t_R g3006 ( 
.A(n_2755),
.Y(n_3006)
);

AND2x4_ASAP7_75t_L g3007 ( 
.A(n_2762),
.B(n_2552),
.Y(n_3007)
);

CKINVDCx5p33_ASAP7_75t_R g3008 ( 
.A(n_2757),
.Y(n_3008)
);

CKINVDCx5p33_ASAP7_75t_R g3009 ( 
.A(n_2763),
.Y(n_3009)
);

CKINVDCx5p33_ASAP7_75t_R g3010 ( 
.A(n_2771),
.Y(n_3010)
);

CKINVDCx5p33_ASAP7_75t_R g3011 ( 
.A(n_2772),
.Y(n_3011)
);

CKINVDCx5p33_ASAP7_75t_R g3012 ( 
.A(n_2783),
.Y(n_3012)
);

CKINVDCx5p33_ASAP7_75t_R g3013 ( 
.A(n_2787),
.Y(n_3013)
);

CKINVDCx5p33_ASAP7_75t_R g3014 ( 
.A(n_2769),
.Y(n_3014)
);

AND3x1_ASAP7_75t_L g3015 ( 
.A(n_2777),
.B(n_1638),
.C(n_1636),
.Y(n_3015)
);

AND2x4_ASAP7_75t_L g3016 ( 
.A(n_2778),
.B(n_2553),
.Y(n_3016)
);

CKINVDCx5p33_ASAP7_75t_R g3017 ( 
.A(n_2784),
.Y(n_3017)
);

CKINVDCx5p33_ASAP7_75t_R g3018 ( 
.A(n_2792),
.Y(n_3018)
);

CKINVDCx5p33_ASAP7_75t_R g3019 ( 
.A(n_2794),
.Y(n_3019)
);

INVx1_ASAP7_75t_L g3020 ( 
.A(n_2796),
.Y(n_3020)
);

CKINVDCx5p33_ASAP7_75t_R g3021 ( 
.A(n_2798),
.Y(n_3021)
);

INVx1_ASAP7_75t_L g3022 ( 
.A(n_2811),
.Y(n_3022)
);

CKINVDCx5p33_ASAP7_75t_R g3023 ( 
.A(n_2804),
.Y(n_3023)
);

CKINVDCx20_ASAP7_75t_R g3024 ( 
.A(n_2782),
.Y(n_3024)
);

CKINVDCx5p33_ASAP7_75t_R g3025 ( 
.A(n_2746),
.Y(n_3025)
);

NAND2xp5_ASAP7_75t_L g3026 ( 
.A(n_2708),
.B(n_2557),
.Y(n_3026)
);

CKINVDCx5p33_ASAP7_75t_R g3027 ( 
.A(n_2746),
.Y(n_3027)
);

CKINVDCx20_ASAP7_75t_R g3028 ( 
.A(n_2782),
.Y(n_3028)
);

CKINVDCx5p33_ASAP7_75t_R g3029 ( 
.A(n_2746),
.Y(n_3029)
);

INVx2_ASAP7_75t_L g3030 ( 
.A(n_2707),
.Y(n_3030)
);

CKINVDCx20_ASAP7_75t_R g3031 ( 
.A(n_2782),
.Y(n_3031)
);

CKINVDCx5p33_ASAP7_75t_R g3032 ( 
.A(n_2746),
.Y(n_3032)
);

AND2x2_ASAP7_75t_L g3033 ( 
.A(n_2705),
.B(n_2485),
.Y(n_3033)
);

BUFx3_ASAP7_75t_L g3034 ( 
.A(n_2684),
.Y(n_3034)
);

CKINVDCx5p33_ASAP7_75t_R g3035 ( 
.A(n_2746),
.Y(n_3035)
);

CKINVDCx20_ASAP7_75t_R g3036 ( 
.A(n_2782),
.Y(n_3036)
);

INVxp67_ASAP7_75t_SL g3037 ( 
.A(n_2712),
.Y(n_3037)
);

NAND2xp33_ASAP7_75t_R g3038 ( 
.A(n_2690),
.B(n_2159),
.Y(n_3038)
);

NAND2xp33_ASAP7_75t_R g3039 ( 
.A(n_2690),
.B(n_2162),
.Y(n_3039)
);

INVx2_ASAP7_75t_L g3040 ( 
.A(n_2893),
.Y(n_3040)
);

HB1xp67_ASAP7_75t_SL g3041 ( 
.A(n_2864),
.Y(n_3041)
);

INVx2_ASAP7_75t_L g3042 ( 
.A(n_2869),
.Y(n_3042)
);

NAND2xp5_ASAP7_75t_L g3043 ( 
.A(n_2900),
.B(n_2904),
.Y(n_3043)
);

CKINVDCx20_ASAP7_75t_R g3044 ( 
.A(n_3024),
.Y(n_3044)
);

AND2x2_ASAP7_75t_L g3045 ( 
.A(n_2894),
.B(n_2616),
.Y(n_3045)
);

INVx2_ASAP7_75t_L g3046 ( 
.A(n_2879),
.Y(n_3046)
);

NAND2xp5_ASAP7_75t_L g3047 ( 
.A(n_2906),
.B(n_2187),
.Y(n_3047)
);

INVx1_ASAP7_75t_L g3048 ( 
.A(n_2856),
.Y(n_3048)
);

BUFx6f_ASAP7_75t_L g3049 ( 
.A(n_2857),
.Y(n_3049)
);

INVx1_ASAP7_75t_L g3050 ( 
.A(n_2874),
.Y(n_3050)
);

BUFx2_ASAP7_75t_L g3051 ( 
.A(n_2983),
.Y(n_3051)
);

OR2x6_ASAP7_75t_SL g3052 ( 
.A(n_2907),
.B(n_2165),
.Y(n_3052)
);

NAND2xp5_ASAP7_75t_SL g3053 ( 
.A(n_2971),
.B(n_2632),
.Y(n_3053)
);

INVx1_ASAP7_75t_L g3054 ( 
.A(n_2887),
.Y(n_3054)
);

OR2x2_ASAP7_75t_L g3055 ( 
.A(n_2918),
.B(n_2527),
.Y(n_3055)
);

INVx1_ASAP7_75t_L g3056 ( 
.A(n_2888),
.Y(n_3056)
);

INVx2_ASAP7_75t_L g3057 ( 
.A(n_2891),
.Y(n_3057)
);

INVx2_ASAP7_75t_L g3058 ( 
.A(n_2891),
.Y(n_3058)
);

AND2x2_ASAP7_75t_SL g3059 ( 
.A(n_2915),
.B(n_1941),
.Y(n_3059)
);

INVx5_ASAP7_75t_L g3060 ( 
.A(n_2882),
.Y(n_3060)
);

AND2x2_ASAP7_75t_L g3061 ( 
.A(n_2955),
.B(n_2653),
.Y(n_3061)
);

NAND2xp5_ASAP7_75t_SL g3062 ( 
.A(n_2927),
.B(n_1629),
.Y(n_3062)
);

BUFx6f_ASAP7_75t_L g3063 ( 
.A(n_2857),
.Y(n_3063)
);

AND2x4_ASAP7_75t_L g3064 ( 
.A(n_2885),
.B(n_2559),
.Y(n_3064)
);

CKINVDCx16_ASAP7_75t_R g3065 ( 
.A(n_2877),
.Y(n_3065)
);

INVx1_ASAP7_75t_L g3066 ( 
.A(n_2901),
.Y(n_3066)
);

INVx4_ASAP7_75t_L g3067 ( 
.A(n_2981),
.Y(n_3067)
);

INVx1_ASAP7_75t_L g3068 ( 
.A(n_2902),
.Y(n_3068)
);

NOR2xp33_ASAP7_75t_L g3069 ( 
.A(n_2878),
.B(n_2663),
.Y(n_3069)
);

INVx5_ASAP7_75t_L g3070 ( 
.A(n_2882),
.Y(n_3070)
);

NAND3x1_ASAP7_75t_L g3071 ( 
.A(n_2931),
.B(n_1643),
.C(n_1642),
.Y(n_3071)
);

INVxp67_ASAP7_75t_SL g3072 ( 
.A(n_2957),
.Y(n_3072)
);

NOR2xp33_ASAP7_75t_L g3073 ( 
.A(n_2928),
.B(n_2665),
.Y(n_3073)
);

HB1xp67_ASAP7_75t_L g3074 ( 
.A(n_2862),
.Y(n_3074)
);

AND2x4_ASAP7_75t_L g3075 ( 
.A(n_3034),
.B(n_2561),
.Y(n_3075)
);

BUFx10_ASAP7_75t_L g3076 ( 
.A(n_2909),
.Y(n_3076)
);

NAND3xp33_ASAP7_75t_L g3077 ( 
.A(n_2948),
.B(n_2952),
.C(n_2949),
.Y(n_3077)
);

AND2x6_ASAP7_75t_L g3078 ( 
.A(n_2930),
.B(n_1929),
.Y(n_3078)
);

BUFx3_ASAP7_75t_L g3079 ( 
.A(n_2886),
.Y(n_3079)
);

INVx2_ASAP7_75t_L g3080 ( 
.A(n_2892),
.Y(n_3080)
);

AOI22xp33_ASAP7_75t_L g3081 ( 
.A1(n_2943),
.A2(n_2033),
.B1(n_2045),
.B2(n_2001),
.Y(n_3081)
);

AND2x6_ASAP7_75t_L g3082 ( 
.A(n_2937),
.B(n_2923),
.Y(n_3082)
);

NOR2xp33_ASAP7_75t_L g3083 ( 
.A(n_2929),
.B(n_1674),
.Y(n_3083)
);

BUFx3_ASAP7_75t_L g3084 ( 
.A(n_2987),
.Y(n_3084)
);

NAND2xp5_ASAP7_75t_L g3085 ( 
.A(n_2968),
.B(n_2562),
.Y(n_3085)
);

AND2x2_ASAP7_75t_L g3086 ( 
.A(n_2984),
.B(n_2565),
.Y(n_3086)
);

INVx3_ASAP7_75t_L g3087 ( 
.A(n_2905),
.Y(n_3087)
);

INVx3_ASAP7_75t_L g3088 ( 
.A(n_2905),
.Y(n_3088)
);

INVx2_ASAP7_75t_L g3089 ( 
.A(n_2963),
.Y(n_3089)
);

NOR2xp33_ASAP7_75t_L g3090 ( 
.A(n_2958),
.B(n_1707),
.Y(n_3090)
);

AND2x2_ASAP7_75t_L g3091 ( 
.A(n_2985),
.B(n_2571),
.Y(n_3091)
);

NAND2xp5_ASAP7_75t_L g3092 ( 
.A(n_2913),
.B(n_2573),
.Y(n_3092)
);

INVx2_ASAP7_75t_L g3093 ( 
.A(n_2976),
.Y(n_3093)
);

INVx2_ASAP7_75t_L g3094 ( 
.A(n_3004),
.Y(n_3094)
);

INVx1_ASAP7_75t_L g3095 ( 
.A(n_3020),
.Y(n_3095)
);

INVx2_ASAP7_75t_L g3096 ( 
.A(n_2982),
.Y(n_3096)
);

INVx1_ASAP7_75t_L g3097 ( 
.A(n_3022),
.Y(n_3097)
);

NAND2xp5_ASAP7_75t_L g3098 ( 
.A(n_2933),
.B(n_2575),
.Y(n_3098)
);

AOI22xp33_ASAP7_75t_L g3099 ( 
.A1(n_3023),
.A2(n_2083),
.B1(n_2100),
.B2(n_2062),
.Y(n_3099)
);

NAND2xp5_ASAP7_75t_L g3100 ( 
.A(n_2959),
.B(n_2576),
.Y(n_3100)
);

AND2x6_ASAP7_75t_L g3101 ( 
.A(n_2941),
.B(n_1955),
.Y(n_3101)
);

INVx2_ASAP7_75t_L g3102 ( 
.A(n_2988),
.Y(n_3102)
);

NOR2xp33_ASAP7_75t_L g3103 ( 
.A(n_2960),
.B(n_1813),
.Y(n_3103)
);

NOR2xp33_ASAP7_75t_L g3104 ( 
.A(n_2962),
.B(n_1818),
.Y(n_3104)
);

INVx1_ASAP7_75t_L g3105 ( 
.A(n_2990),
.Y(n_3105)
);

AND2x4_ASAP7_75t_L g3106 ( 
.A(n_2994),
.B(n_2578),
.Y(n_3106)
);

INVx2_ASAP7_75t_L g3107 ( 
.A(n_2996),
.Y(n_3107)
);

BUFx6f_ASAP7_75t_L g3108 ( 
.A(n_2905),
.Y(n_3108)
);

AND2x4_ASAP7_75t_L g3109 ( 
.A(n_2946),
.B(n_2579),
.Y(n_3109)
);

NOR2xp33_ASAP7_75t_L g3110 ( 
.A(n_2964),
.B(n_1821),
.Y(n_3110)
);

INVx1_ASAP7_75t_L g3111 ( 
.A(n_2998),
.Y(n_3111)
);

INVx1_ASAP7_75t_L g3112 ( 
.A(n_3007),
.Y(n_3112)
);

INVx2_ASAP7_75t_L g3113 ( 
.A(n_2867),
.Y(n_3113)
);

INVx3_ASAP7_75t_L g3114 ( 
.A(n_3007),
.Y(n_3114)
);

AND2x2_ASAP7_75t_L g3115 ( 
.A(n_2880),
.B(n_2580),
.Y(n_3115)
);

BUFx10_ASAP7_75t_L g3116 ( 
.A(n_2865),
.Y(n_3116)
);

INVx1_ASAP7_75t_L g3117 ( 
.A(n_3016),
.Y(n_3117)
);

BUFx6f_ASAP7_75t_L g3118 ( 
.A(n_3016),
.Y(n_3118)
);

INVx1_ASAP7_75t_L g3119 ( 
.A(n_2999),
.Y(n_3119)
);

INVx3_ASAP7_75t_L g3120 ( 
.A(n_2993),
.Y(n_3120)
);

AND2x2_ASAP7_75t_L g3121 ( 
.A(n_2950),
.B(n_2581),
.Y(n_3121)
);

NAND2xp5_ASAP7_75t_SL g3122 ( 
.A(n_2873),
.B(n_1634),
.Y(n_3122)
);

AND2x2_ASAP7_75t_L g3123 ( 
.A(n_2914),
.B(n_2583),
.Y(n_3123)
);

INVx5_ASAP7_75t_L g3124 ( 
.A(n_2980),
.Y(n_3124)
);

OR2x2_ASAP7_75t_L g3125 ( 
.A(n_2975),
.B(n_2022),
.Y(n_3125)
);

BUFx10_ASAP7_75t_L g3126 ( 
.A(n_2870),
.Y(n_3126)
);

OR2x2_ASAP7_75t_L g3127 ( 
.A(n_2917),
.B(n_2972),
.Y(n_3127)
);

BUFx3_ASAP7_75t_L g3128 ( 
.A(n_2995),
.Y(n_3128)
);

NAND2xp5_ASAP7_75t_L g3129 ( 
.A(n_2924),
.B(n_1637),
.Y(n_3129)
);

INVx3_ASAP7_75t_L g3130 ( 
.A(n_2953),
.Y(n_3130)
);

INVx3_ASAP7_75t_L g3131 ( 
.A(n_2954),
.Y(n_3131)
);

INVx2_ASAP7_75t_L g3132 ( 
.A(n_3030),
.Y(n_3132)
);

AND2x6_ASAP7_75t_L g3133 ( 
.A(n_2956),
.B(n_2073),
.Y(n_3133)
);

INVx2_ASAP7_75t_L g3134 ( 
.A(n_3026),
.Y(n_3134)
);

INVx1_ASAP7_75t_L g3135 ( 
.A(n_2966),
.Y(n_3135)
);

NAND2xp33_ASAP7_75t_L g3136 ( 
.A(n_2919),
.B(n_2181),
.Y(n_3136)
);

NAND2xp5_ASAP7_75t_SL g3137 ( 
.A(n_2875),
.B(n_2876),
.Y(n_3137)
);

AND2x6_ASAP7_75t_L g3138 ( 
.A(n_2961),
.B(n_2374),
.Y(n_3138)
);

AND2x6_ASAP7_75t_L g3139 ( 
.A(n_2903),
.B(n_1645),
.Y(n_3139)
);

NAND2xp5_ASAP7_75t_L g3140 ( 
.A(n_2924),
.B(n_1639),
.Y(n_3140)
);

BUFx6f_ASAP7_75t_L g3141 ( 
.A(n_2980),
.Y(n_3141)
);

INVx1_ASAP7_75t_L g3142 ( 
.A(n_2986),
.Y(n_3142)
);

INVx1_ASAP7_75t_L g3143 ( 
.A(n_2992),
.Y(n_3143)
);

BUFx2_ASAP7_75t_L g3144 ( 
.A(n_2895),
.Y(n_3144)
);

INVx1_ASAP7_75t_L g3145 ( 
.A(n_3005),
.Y(n_3145)
);

BUFx10_ASAP7_75t_L g3146 ( 
.A(n_2863),
.Y(n_3146)
);

NAND2xp5_ASAP7_75t_L g3147 ( 
.A(n_2924),
.B(n_1641),
.Y(n_3147)
);

BUFx6f_ASAP7_75t_L g3148 ( 
.A(n_2944),
.Y(n_3148)
);

NAND2xp5_ASAP7_75t_SL g3149 ( 
.A(n_3001),
.B(n_1646),
.Y(n_3149)
);

AND2x2_ASAP7_75t_L g3150 ( 
.A(n_2910),
.B(n_1644),
.Y(n_3150)
);

NAND2xp5_ASAP7_75t_L g3151 ( 
.A(n_2919),
.B(n_1648),
.Y(n_3151)
);

INVx1_ASAP7_75t_L g3152 ( 
.A(n_2965),
.Y(n_3152)
);

INVx1_ASAP7_75t_L g3153 ( 
.A(n_2896),
.Y(n_3153)
);

BUFx3_ASAP7_75t_L g3154 ( 
.A(n_3000),
.Y(n_3154)
);

INVx6_ASAP7_75t_L g3155 ( 
.A(n_2989),
.Y(n_3155)
);

OR2x2_ASAP7_75t_L g3156 ( 
.A(n_2974),
.B(n_2239),
.Y(n_3156)
);

NAND2xp5_ASAP7_75t_L g3157 ( 
.A(n_2919),
.B(n_1651),
.Y(n_3157)
);

BUFx10_ASAP7_75t_L g3158 ( 
.A(n_2858),
.Y(n_3158)
);

NAND2xp5_ASAP7_75t_L g3159 ( 
.A(n_3037),
.B(n_1653),
.Y(n_3159)
);

BUFx6f_ASAP7_75t_L g3160 ( 
.A(n_2944),
.Y(n_3160)
);

AND2x4_ASAP7_75t_L g3161 ( 
.A(n_2908),
.B(n_1649),
.Y(n_3161)
);

NAND2xp5_ASAP7_75t_L g3162 ( 
.A(n_2926),
.B(n_1654),
.Y(n_3162)
);

BUFx6f_ASAP7_75t_L g3163 ( 
.A(n_2944),
.Y(n_3163)
);

INVx2_ASAP7_75t_SL g3164 ( 
.A(n_3006),
.Y(n_3164)
);

AND2x2_ASAP7_75t_L g3165 ( 
.A(n_2912),
.B(n_1706),
.Y(n_3165)
);

INVx2_ASAP7_75t_SL g3166 ( 
.A(n_3008),
.Y(n_3166)
);

INVx2_ASAP7_75t_L g3167 ( 
.A(n_2939),
.Y(n_3167)
);

AOI22x1_ASAP7_75t_L g3168 ( 
.A1(n_2939),
.A2(n_2190),
.B1(n_2203),
.B2(n_2189),
.Y(n_3168)
);

INVx4_ASAP7_75t_L g3169 ( 
.A(n_3009),
.Y(n_3169)
);

BUFx6f_ASAP7_75t_L g3170 ( 
.A(n_3002),
.Y(n_3170)
);

NAND2xp5_ASAP7_75t_SL g3171 ( 
.A(n_3014),
.B(n_1655),
.Y(n_3171)
);

NOR2xp33_ASAP7_75t_L g3172 ( 
.A(n_2973),
.B(n_2266),
.Y(n_3172)
);

INVx4_ASAP7_75t_L g3173 ( 
.A(n_3010),
.Y(n_3173)
);

BUFx2_ASAP7_75t_L g3174 ( 
.A(n_2868),
.Y(n_3174)
);

NAND2xp5_ASAP7_75t_L g3175 ( 
.A(n_3011),
.B(n_1657),
.Y(n_3175)
);

AND2x2_ASAP7_75t_L g3176 ( 
.A(n_2871),
.B(n_1706),
.Y(n_3176)
);

INVx3_ASAP7_75t_L g3177 ( 
.A(n_3012),
.Y(n_3177)
);

INVx2_ASAP7_75t_L g3178 ( 
.A(n_3002),
.Y(n_3178)
);

INVx1_ASAP7_75t_L g3179 ( 
.A(n_3013),
.Y(n_3179)
);

INVx2_ASAP7_75t_L g3180 ( 
.A(n_3002),
.Y(n_3180)
);

INVx1_ASAP7_75t_L g3181 ( 
.A(n_3017),
.Y(n_3181)
);

INVx1_ASAP7_75t_L g3182 ( 
.A(n_3018),
.Y(n_3182)
);

NOR2x1p5_ASAP7_75t_L g3183 ( 
.A(n_2969),
.B(n_2970),
.Y(n_3183)
);

NAND2xp5_ASAP7_75t_SL g3184 ( 
.A(n_3019),
.B(n_1658),
.Y(n_3184)
);

OAI22xp5_ASAP7_75t_L g3185 ( 
.A1(n_2922),
.A2(n_2419),
.B1(n_2452),
.B2(n_2371),
.Y(n_3185)
);

INVx2_ASAP7_75t_L g3186 ( 
.A(n_3021),
.Y(n_3186)
);

NOR2xp33_ASAP7_75t_L g3187 ( 
.A(n_2979),
.B(n_2273),
.Y(n_3187)
);

INVx1_ASAP7_75t_L g3188 ( 
.A(n_3003),
.Y(n_3188)
);

OAI22xp5_ASAP7_75t_L g3189 ( 
.A1(n_2947),
.A2(n_2281),
.B1(n_2331),
.B2(n_2280),
.Y(n_3189)
);

INVx1_ASAP7_75t_L g3190 ( 
.A(n_2977),
.Y(n_3190)
);

INVx2_ASAP7_75t_L g3191 ( 
.A(n_3015),
.Y(n_3191)
);

NAND2xp5_ASAP7_75t_L g3192 ( 
.A(n_2978),
.B(n_1660),
.Y(n_3192)
);

NOR2xp33_ASAP7_75t_L g3193 ( 
.A(n_2940),
.B(n_2357),
.Y(n_3193)
);

NOR2xp33_ASAP7_75t_L g3194 ( 
.A(n_2942),
.B(n_2409),
.Y(n_3194)
);

NAND2xp5_ASAP7_75t_SL g3195 ( 
.A(n_2945),
.B(n_1663),
.Y(n_3195)
);

OR2x2_ASAP7_75t_L g3196 ( 
.A(n_2951),
.B(n_2883),
.Y(n_3196)
);

NAND2xp5_ASAP7_75t_SL g3197 ( 
.A(n_2916),
.B(n_1664),
.Y(n_3197)
);

HB1xp67_ASAP7_75t_L g3198 ( 
.A(n_2934),
.Y(n_3198)
);

AOI22xp33_ASAP7_75t_L g3199 ( 
.A1(n_2920),
.A2(n_2329),
.B1(n_2335),
.B2(n_2318),
.Y(n_3199)
);

INVx1_ASAP7_75t_L g3200 ( 
.A(n_2967),
.Y(n_3200)
);

NOR2xp33_ASAP7_75t_L g3201 ( 
.A(n_2881),
.B(n_2417),
.Y(n_3201)
);

INVx2_ASAP7_75t_L g3202 ( 
.A(n_2921),
.Y(n_3202)
);

NOR2xp33_ASAP7_75t_L g3203 ( 
.A(n_2859),
.B(n_2427),
.Y(n_3203)
);

CKINVDCx5p33_ASAP7_75t_R g3204 ( 
.A(n_2855),
.Y(n_3204)
);

AND3x2_ASAP7_75t_L g3205 ( 
.A(n_2991),
.B(n_2402),
.C(n_2401),
.Y(n_3205)
);

NOR2x1p5_ASAP7_75t_L g3206 ( 
.A(n_2860),
.B(n_3025),
.Y(n_3206)
);

INVx3_ASAP7_75t_L g3207 ( 
.A(n_2884),
.Y(n_3207)
);

INVx1_ASAP7_75t_L g3208 ( 
.A(n_2897),
.Y(n_3208)
);

INVx1_ASAP7_75t_L g3209 ( 
.A(n_2898),
.Y(n_3209)
);

INVx1_ASAP7_75t_SL g3210 ( 
.A(n_2872),
.Y(n_3210)
);

NOR3xp33_ASAP7_75t_L g3211 ( 
.A(n_2899),
.B(n_2450),
.C(n_2434),
.Y(n_3211)
);

OAI21xp33_ASAP7_75t_SL g3212 ( 
.A1(n_2997),
.A2(n_1662),
.B(n_1659),
.Y(n_3212)
);

INVx2_ASAP7_75t_L g3213 ( 
.A(n_2938),
.Y(n_3213)
);

AND2x2_ASAP7_75t_L g3214 ( 
.A(n_3027),
.B(n_3029),
.Y(n_3214)
);

INVx2_ASAP7_75t_L g3215 ( 
.A(n_2935),
.Y(n_3215)
);

NAND2xp5_ASAP7_75t_L g3216 ( 
.A(n_3032),
.B(n_1667),
.Y(n_3216)
);

INVx3_ASAP7_75t_L g3217 ( 
.A(n_2889),
.Y(n_3217)
);

AND2x4_ASAP7_75t_L g3218 ( 
.A(n_2890),
.B(n_1672),
.Y(n_3218)
);

INVx2_ASAP7_75t_L g3219 ( 
.A(n_2925),
.Y(n_3219)
);

AND2x6_ASAP7_75t_L g3220 ( 
.A(n_3038),
.B(n_1682),
.Y(n_3220)
);

INVx3_ASAP7_75t_L g3221 ( 
.A(n_3035),
.Y(n_3221)
);

AND2x2_ASAP7_75t_L g3222 ( 
.A(n_2911),
.B(n_1783),
.Y(n_3222)
);

AND2x6_ASAP7_75t_L g3223 ( 
.A(n_3039),
.B(n_1686),
.Y(n_3223)
);

AND2x2_ASAP7_75t_L g3224 ( 
.A(n_2866),
.B(n_1783),
.Y(n_3224)
);

INVx1_ASAP7_75t_L g3225 ( 
.A(n_2932),
.Y(n_3225)
);

BUFx3_ASAP7_75t_L g3226 ( 
.A(n_3028),
.Y(n_3226)
);

AOI22xp33_ASAP7_75t_L g3227 ( 
.A1(n_2936),
.A2(n_2420),
.B1(n_2428),
.B2(n_2404),
.Y(n_3227)
);

AOI22xp5_ASAP7_75t_L g3228 ( 
.A1(n_3036),
.A2(n_2499),
.B1(n_1915),
.B2(n_1921),
.Y(n_3228)
);

INVx1_ASAP7_75t_L g3229 ( 
.A(n_3031),
.Y(n_3229)
);

INVx1_ASAP7_75t_L g3230 ( 
.A(n_2856),
.Y(n_3230)
);

INVx2_ASAP7_75t_L g3231 ( 
.A(n_2893),
.Y(n_3231)
);

INVx2_ASAP7_75t_L g3232 ( 
.A(n_2893),
.Y(n_3232)
);

AND2x6_ASAP7_75t_L g3233 ( 
.A(n_2894),
.B(n_1691),
.Y(n_3233)
);

CKINVDCx20_ASAP7_75t_R g3234 ( 
.A(n_3024),
.Y(n_3234)
);

NAND2xp5_ASAP7_75t_L g3235 ( 
.A(n_2900),
.B(n_1670),
.Y(n_3235)
);

INVx1_ASAP7_75t_L g3236 ( 
.A(n_2856),
.Y(n_3236)
);

NAND2xp5_ASAP7_75t_L g3237 ( 
.A(n_2900),
.B(n_1673),
.Y(n_3237)
);

BUFx3_ASAP7_75t_L g3238 ( 
.A(n_2861),
.Y(n_3238)
);

BUFx3_ASAP7_75t_L g3239 ( 
.A(n_2861),
.Y(n_3239)
);

AND2x4_ASAP7_75t_L g3240 ( 
.A(n_2861),
.B(n_1692),
.Y(n_3240)
);

AND2x6_ASAP7_75t_L g3241 ( 
.A(n_2894),
.B(n_1694),
.Y(n_3241)
);

INVx1_ASAP7_75t_SL g3242 ( 
.A(n_3033),
.Y(n_3242)
);

OR2x2_ASAP7_75t_L g3243 ( 
.A(n_3033),
.B(n_2236),
.Y(n_3243)
);

NAND2xp5_ASAP7_75t_L g3244 ( 
.A(n_2900),
.B(n_1675),
.Y(n_3244)
);

INVx1_ASAP7_75t_L g3245 ( 
.A(n_2856),
.Y(n_3245)
);

NAND2xp5_ASAP7_75t_L g3246 ( 
.A(n_2900),
.B(n_1677),
.Y(n_3246)
);

NAND2xp5_ASAP7_75t_L g3247 ( 
.A(n_2900),
.B(n_1678),
.Y(n_3247)
);

OAI22xp33_ASAP7_75t_L g3248 ( 
.A1(n_2943),
.A2(n_2249),
.B1(n_2251),
.B2(n_2240),
.Y(n_3248)
);

NOR2xp33_ASAP7_75t_L g3249 ( 
.A(n_2878),
.B(n_2282),
.Y(n_3249)
);

INVx1_ASAP7_75t_L g3250 ( 
.A(n_2856),
.Y(n_3250)
);

NOR2xp33_ASAP7_75t_L g3251 ( 
.A(n_2878),
.B(n_2287),
.Y(n_3251)
);

AND2x4_ASAP7_75t_L g3252 ( 
.A(n_2861),
.B(n_1695),
.Y(n_3252)
);

AND2x4_ASAP7_75t_L g3253 ( 
.A(n_2861),
.B(n_1699),
.Y(n_3253)
);

NAND2xp5_ASAP7_75t_L g3254 ( 
.A(n_2900),
.B(n_1679),
.Y(n_3254)
);

NOR2xp33_ASAP7_75t_L g3255 ( 
.A(n_2878),
.B(n_2289),
.Y(n_3255)
);

INVx1_ASAP7_75t_L g3256 ( 
.A(n_2856),
.Y(n_3256)
);

BUFx3_ASAP7_75t_L g3257 ( 
.A(n_2861),
.Y(n_3257)
);

INVx1_ASAP7_75t_L g3258 ( 
.A(n_2856),
.Y(n_3258)
);

AND2x4_ASAP7_75t_L g3259 ( 
.A(n_2861),
.B(n_1703),
.Y(n_3259)
);

OR2x2_ASAP7_75t_L g3260 ( 
.A(n_3033),
.B(n_2295),
.Y(n_3260)
);

NAND2xp5_ASAP7_75t_SL g3261 ( 
.A(n_2971),
.B(n_1680),
.Y(n_3261)
);

INVx3_ASAP7_75t_L g3262 ( 
.A(n_2857),
.Y(n_3262)
);

NAND2xp33_ASAP7_75t_SL g3263 ( 
.A(n_2914),
.B(n_1913),
.Y(n_3263)
);

INVx1_ASAP7_75t_L g3264 ( 
.A(n_2856),
.Y(n_3264)
);

INVx1_ASAP7_75t_L g3265 ( 
.A(n_2856),
.Y(n_3265)
);

OR2x6_ASAP7_75t_L g3266 ( 
.A(n_2861),
.B(n_2429),
.Y(n_3266)
);

INVx2_ASAP7_75t_L g3267 ( 
.A(n_2893),
.Y(n_3267)
);

INVx4_ASAP7_75t_L g3268 ( 
.A(n_2981),
.Y(n_3268)
);

AND2x6_ASAP7_75t_L g3269 ( 
.A(n_2894),
.B(n_1715),
.Y(n_3269)
);

BUFx6f_ASAP7_75t_L g3270 ( 
.A(n_2857),
.Y(n_3270)
);

INVx1_ASAP7_75t_L g3271 ( 
.A(n_2856),
.Y(n_3271)
);

INVxp33_ASAP7_75t_L g3272 ( 
.A(n_3033),
.Y(n_3272)
);

INVx1_ASAP7_75t_L g3273 ( 
.A(n_2856),
.Y(n_3273)
);

OR2x6_ASAP7_75t_L g3274 ( 
.A(n_2861),
.B(n_2449),
.Y(n_3274)
);

BUFx3_ASAP7_75t_L g3275 ( 
.A(n_2861),
.Y(n_3275)
);

AND2x4_ASAP7_75t_L g3276 ( 
.A(n_2861),
.B(n_1722),
.Y(n_3276)
);

BUFx3_ASAP7_75t_L g3277 ( 
.A(n_2861),
.Y(n_3277)
);

AND2x2_ASAP7_75t_L g3278 ( 
.A(n_2894),
.B(n_1865),
.Y(n_3278)
);

INVx3_ASAP7_75t_L g3279 ( 
.A(n_3049),
.Y(n_3279)
);

NAND2xp5_ASAP7_75t_SL g3280 ( 
.A(n_3077),
.B(n_1935),
.Y(n_3280)
);

INVx1_ASAP7_75t_L g3281 ( 
.A(n_3048),
.Y(n_3281)
);

NOR3xp33_ASAP7_75t_L g3282 ( 
.A(n_3193),
.B(n_1685),
.C(n_1684),
.Y(n_3282)
);

NOR2xp33_ASAP7_75t_L g3283 ( 
.A(n_3043),
.B(n_1950),
.Y(n_3283)
);

NAND2xp5_ASAP7_75t_L g3284 ( 
.A(n_3153),
.B(n_1688),
.Y(n_3284)
);

NOR2xp67_ASAP7_75t_L g3285 ( 
.A(n_3060),
.B(n_2325),
.Y(n_3285)
);

NAND3xp33_ASAP7_75t_L g3286 ( 
.A(n_3083),
.B(n_1697),
.C(n_1696),
.Y(n_3286)
);

AND2x2_ASAP7_75t_L g3287 ( 
.A(n_3045),
.B(n_1865),
.Y(n_3287)
);

NAND2xp33_ASAP7_75t_L g3288 ( 
.A(n_3148),
.B(n_2341),
.Y(n_3288)
);

NOR2xp33_ASAP7_75t_L g3289 ( 
.A(n_3194),
.B(n_1951),
.Y(n_3289)
);

NAND2xp5_ASAP7_75t_L g3290 ( 
.A(n_3143),
.B(n_1702),
.Y(n_3290)
);

NAND2xp5_ASAP7_75t_SL g3291 ( 
.A(n_3186),
.B(n_1990),
.Y(n_3291)
);

INVx2_ASAP7_75t_L g3292 ( 
.A(n_3231),
.Y(n_3292)
);

NAND2xp5_ASAP7_75t_SL g3293 ( 
.A(n_3177),
.B(n_1995),
.Y(n_3293)
);

AOI22xp33_ASAP7_75t_L g3294 ( 
.A1(n_3134),
.A2(n_2044),
.B1(n_2067),
.B2(n_2011),
.Y(n_3294)
);

NAND2xp5_ASAP7_75t_L g3295 ( 
.A(n_3090),
.B(n_1708),
.Y(n_3295)
);

AND2x2_ASAP7_75t_L g3296 ( 
.A(n_3103),
.B(n_2052),
.Y(n_3296)
);

NAND2xp5_ASAP7_75t_L g3297 ( 
.A(n_3104),
.B(n_1714),
.Y(n_3297)
);

INVx2_ASAP7_75t_L g3298 ( 
.A(n_3232),
.Y(n_3298)
);

NAND2xp5_ASAP7_75t_L g3299 ( 
.A(n_3249),
.B(n_3251),
.Y(n_3299)
);

O2A1O1Ixp5_ASAP7_75t_L g3300 ( 
.A1(n_3085),
.A2(n_2464),
.B(n_1727),
.C(n_1728),
.Y(n_3300)
);

A2O1A1Ixp33_ASAP7_75t_L g3301 ( 
.A1(n_3255),
.A2(n_1735),
.B(n_1738),
.C(n_1725),
.Y(n_3301)
);

INVx2_ASAP7_75t_L g3302 ( 
.A(n_3267),
.Y(n_3302)
);

INVx2_ASAP7_75t_SL g3303 ( 
.A(n_3121),
.Y(n_3303)
);

INVx8_ASAP7_75t_L g3304 ( 
.A(n_3060),
.Y(n_3304)
);

INVx1_ASAP7_75t_L g3305 ( 
.A(n_3050),
.Y(n_3305)
);

CKINVDCx5p33_ASAP7_75t_R g3306 ( 
.A(n_3204),
.Y(n_3306)
);

BUFx3_ASAP7_75t_L g3307 ( 
.A(n_3128),
.Y(n_3307)
);

AOI22xp33_ASAP7_75t_L g3308 ( 
.A1(n_3191),
.A2(n_2117),
.B1(n_2132),
.B2(n_2081),
.Y(n_3308)
);

INVx2_ASAP7_75t_SL g3309 ( 
.A(n_3064),
.Y(n_3309)
);

NAND2xp5_ASAP7_75t_SL g3310 ( 
.A(n_3164),
.B(n_2140),
.Y(n_3310)
);

NOR2xp33_ASAP7_75t_L g3311 ( 
.A(n_3203),
.B(n_2152),
.Y(n_3311)
);

OAI22xp5_ASAP7_75t_L g3312 ( 
.A1(n_3167),
.A2(n_2223),
.B1(n_2226),
.B2(n_2222),
.Y(n_3312)
);

NOR2xp33_ASAP7_75t_L g3313 ( 
.A(n_3272),
.B(n_2241),
.Y(n_3313)
);

INVx2_ASAP7_75t_L g3314 ( 
.A(n_3042),
.Y(n_3314)
);

NOR2xp33_ASAP7_75t_R g3315 ( 
.A(n_3044),
.B(n_2255),
.Y(n_3315)
);

INVx2_ASAP7_75t_L g3316 ( 
.A(n_3046),
.Y(n_3316)
);

NOR2xp33_ASAP7_75t_L g3317 ( 
.A(n_3053),
.B(n_2256),
.Y(n_3317)
);

NAND2xp5_ASAP7_75t_SL g3318 ( 
.A(n_3166),
.B(n_2269),
.Y(n_3318)
);

OR2x6_ASAP7_75t_L g3319 ( 
.A(n_3067),
.B(n_1739),
.Y(n_3319)
);

NAND2xp5_ASAP7_75t_L g3320 ( 
.A(n_3047),
.B(n_1729),
.Y(n_3320)
);

NAND2xp5_ASAP7_75t_L g3321 ( 
.A(n_3054),
.B(n_1730),
.Y(n_3321)
);

NAND2xp5_ASAP7_75t_L g3322 ( 
.A(n_3056),
.B(n_1731),
.Y(n_3322)
);

OAI22xp33_ASAP7_75t_SL g3323 ( 
.A1(n_3151),
.A2(n_2363),
.B1(n_2365),
.B2(n_2355),
.Y(n_3323)
);

NAND2xp5_ASAP7_75t_SL g3324 ( 
.A(n_3118),
.B(n_2272),
.Y(n_3324)
);

NAND2xp5_ASAP7_75t_SL g3325 ( 
.A(n_3235),
.B(n_3237),
.Y(n_3325)
);

INVx1_ASAP7_75t_L g3326 ( 
.A(n_3066),
.Y(n_3326)
);

NAND2xp5_ASAP7_75t_L g3327 ( 
.A(n_3068),
.B(n_1732),
.Y(n_3327)
);

NAND2x1_ASAP7_75t_L g3328 ( 
.A(n_3148),
.B(n_3160),
.Y(n_3328)
);

INVxp33_ASAP7_75t_SL g3329 ( 
.A(n_3214),
.Y(n_3329)
);

O2A1O1Ixp33_ASAP7_75t_L g3330 ( 
.A1(n_3212),
.A2(n_1743),
.B(n_1744),
.C(n_1742),
.Y(n_3330)
);

INVx1_ASAP7_75t_L g3331 ( 
.A(n_3095),
.Y(n_3331)
);

NAND2xp5_ASAP7_75t_SL g3332 ( 
.A(n_3244),
.B(n_2308),
.Y(n_3332)
);

BUFx6f_ASAP7_75t_L g3333 ( 
.A(n_3049),
.Y(n_3333)
);

A2O1A1Ixp33_ASAP7_75t_L g3334 ( 
.A1(n_3201),
.A2(n_1751),
.B(n_1752),
.C(n_1746),
.Y(n_3334)
);

NAND2xp5_ASAP7_75t_L g3335 ( 
.A(n_3097),
.B(n_1733),
.Y(n_3335)
);

NAND2xp5_ASAP7_75t_SL g3336 ( 
.A(n_3246),
.B(n_2309),
.Y(n_3336)
);

NAND2xp5_ASAP7_75t_SL g3337 ( 
.A(n_3247),
.B(n_2334),
.Y(n_3337)
);

NAND2xp5_ASAP7_75t_L g3338 ( 
.A(n_3230),
.B(n_1740),
.Y(n_3338)
);

INVx2_ASAP7_75t_SL g3339 ( 
.A(n_3075),
.Y(n_3339)
);

BUFx2_ASAP7_75t_L g3340 ( 
.A(n_3154),
.Y(n_3340)
);

NOR2xp33_ASAP7_75t_SL g3341 ( 
.A(n_3065),
.B(n_3158),
.Y(n_3341)
);

NAND2xp5_ASAP7_75t_L g3342 ( 
.A(n_3236),
.B(n_1747),
.Y(n_3342)
);

NAND2xp5_ASAP7_75t_L g3343 ( 
.A(n_3245),
.B(n_1748),
.Y(n_3343)
);

OR2x2_ASAP7_75t_L g3344 ( 
.A(n_3242),
.B(n_3055),
.Y(n_3344)
);

NOR2xp33_ASAP7_75t_L g3345 ( 
.A(n_3254),
.B(n_2360),
.Y(n_3345)
);

INVx1_ASAP7_75t_L g3346 ( 
.A(n_3250),
.Y(n_3346)
);

NOR2xp33_ASAP7_75t_L g3347 ( 
.A(n_3069),
.B(n_3181),
.Y(n_3347)
);

AND2x2_ASAP7_75t_L g3348 ( 
.A(n_3115),
.B(n_2052),
.Y(n_3348)
);

NOR2xp33_ASAP7_75t_SL g3349 ( 
.A(n_3116),
.B(n_2367),
.Y(n_3349)
);

NOR2xp33_ASAP7_75t_L g3350 ( 
.A(n_3182),
.B(n_2369),
.Y(n_3350)
);

INVx2_ASAP7_75t_L g3351 ( 
.A(n_3089),
.Y(n_3351)
);

NAND2xp5_ASAP7_75t_SL g3352 ( 
.A(n_3059),
.B(n_2386),
.Y(n_3352)
);

NAND2xp5_ASAP7_75t_L g3353 ( 
.A(n_3256),
.B(n_3258),
.Y(n_3353)
);

NAND2xp5_ASAP7_75t_SL g3354 ( 
.A(n_3179),
.B(n_2398),
.Y(n_3354)
);

NAND2xp5_ASAP7_75t_SL g3355 ( 
.A(n_3114),
.B(n_2400),
.Y(n_3355)
);

INVx3_ASAP7_75t_L g3356 ( 
.A(n_3063),
.Y(n_3356)
);

OAI21xp5_ASAP7_75t_L g3357 ( 
.A1(n_3178),
.A2(n_1767),
.B(n_1754),
.Y(n_3357)
);

AND2x2_ASAP7_75t_L g3358 ( 
.A(n_3086),
.B(n_2154),
.Y(n_3358)
);

INVx2_ASAP7_75t_L g3359 ( 
.A(n_3093),
.Y(n_3359)
);

OR2x2_ASAP7_75t_L g3360 ( 
.A(n_3125),
.B(n_2375),
.Y(n_3360)
);

BUFx8_ASAP7_75t_L g3361 ( 
.A(n_3174),
.Y(n_3361)
);

NAND2xp5_ASAP7_75t_SL g3362 ( 
.A(n_3169),
.B(n_2436),
.Y(n_3362)
);

AND2x2_ASAP7_75t_L g3363 ( 
.A(n_3091),
.B(n_2154),
.Y(n_3363)
);

AND2x4_ASAP7_75t_L g3364 ( 
.A(n_3070),
.B(n_3238),
.Y(n_3364)
);

NAND2xp5_ASAP7_75t_L g3365 ( 
.A(n_3264),
.B(n_1762),
.Y(n_3365)
);

NAND2xp5_ASAP7_75t_L g3366 ( 
.A(n_3265),
.B(n_1763),
.Y(n_3366)
);

AOI21xp5_ASAP7_75t_L g3367 ( 
.A1(n_3160),
.A2(n_1770),
.B(n_1768),
.Y(n_3367)
);

NAND2xp5_ASAP7_75t_SL g3368 ( 
.A(n_3173),
.B(n_3100),
.Y(n_3368)
);

NOR2xp33_ASAP7_75t_L g3369 ( 
.A(n_3110),
.B(n_2442),
.Y(n_3369)
);

INVx1_ASAP7_75t_L g3370 ( 
.A(n_3271),
.Y(n_3370)
);

O2A1O1Ixp5_ASAP7_75t_L g3371 ( 
.A1(n_3273),
.A2(n_1792),
.B(n_1800),
.C(n_1781),
.Y(n_3371)
);

OAI22xp5_ASAP7_75t_L g3372 ( 
.A1(n_3180),
.A2(n_1771),
.B1(n_1774),
.B2(n_1764),
.Y(n_3372)
);

INVx2_ASAP7_75t_SL g3373 ( 
.A(n_3123),
.Y(n_3373)
);

AOI22xp5_ASAP7_75t_L g3374 ( 
.A1(n_3136),
.A2(n_1778),
.B1(n_1779),
.B2(n_1776),
.Y(n_3374)
);

INVx1_ASAP7_75t_L g3375 ( 
.A(n_3105),
.Y(n_3375)
);

INVx2_ASAP7_75t_L g3376 ( 
.A(n_3094),
.Y(n_3376)
);

NOR2xp33_ASAP7_75t_L g3377 ( 
.A(n_3172),
.B(n_1782),
.Y(n_3377)
);

NOR2xp33_ASAP7_75t_L g3378 ( 
.A(n_3187),
.B(n_1785),
.Y(n_3378)
);

INVx2_ASAP7_75t_L g3379 ( 
.A(n_3113),
.Y(n_3379)
);

AOI22xp33_ASAP7_75t_L g3380 ( 
.A1(n_3220),
.A2(n_3223),
.B1(n_3241),
.B2(n_3233),
.Y(n_3380)
);

NAND2xp5_ASAP7_75t_SL g3381 ( 
.A(n_3190),
.B(n_1791),
.Y(n_3381)
);

NAND2xp5_ASAP7_75t_L g3382 ( 
.A(n_3163),
.B(n_1793),
.Y(n_3382)
);

AND2x4_ASAP7_75t_L g3383 ( 
.A(n_3070),
.B(n_1803),
.Y(n_3383)
);

INVx2_ASAP7_75t_L g3384 ( 
.A(n_3132),
.Y(n_3384)
);

INVx1_ASAP7_75t_L g3385 ( 
.A(n_3111),
.Y(n_3385)
);

AND2x6_ASAP7_75t_SL g3386 ( 
.A(n_3073),
.B(n_1807),
.Y(n_3386)
);

OAI22xp5_ASAP7_75t_L g3387 ( 
.A1(n_3163),
.A2(n_1796),
.B1(n_1797),
.B2(n_1795),
.Y(n_3387)
);

NOR2xp33_ASAP7_75t_L g3388 ( 
.A(n_3198),
.B(n_1802),
.Y(n_3388)
);

NOR2xp33_ASAP7_75t_L g3389 ( 
.A(n_3216),
.B(n_1804),
.Y(n_3389)
);

NOR2xp33_ASAP7_75t_L g3390 ( 
.A(n_3156),
.B(n_3197),
.Y(n_3390)
);

INVx2_ASAP7_75t_L g3391 ( 
.A(n_3096),
.Y(n_3391)
);

BUFx6f_ASAP7_75t_L g3392 ( 
.A(n_3063),
.Y(n_3392)
);

INVx2_ASAP7_75t_L g3393 ( 
.A(n_3102),
.Y(n_3393)
);

INVx2_ASAP7_75t_L g3394 ( 
.A(n_3107),
.Y(n_3394)
);

NAND2xp5_ASAP7_75t_L g3395 ( 
.A(n_3170),
.B(n_1808),
.Y(n_3395)
);

NAND2xp5_ASAP7_75t_SL g3396 ( 
.A(n_3144),
.B(n_1810),
.Y(n_3396)
);

NAND2xp5_ASAP7_75t_L g3397 ( 
.A(n_3162),
.B(n_1811),
.Y(n_3397)
);

INVx2_ASAP7_75t_L g3398 ( 
.A(n_3057),
.Y(n_3398)
);

INVx2_ASAP7_75t_L g3399 ( 
.A(n_3058),
.Y(n_3399)
);

NAND2xp5_ASAP7_75t_L g3400 ( 
.A(n_3098),
.B(n_1814),
.Y(n_3400)
);

NAND2xp5_ASAP7_75t_L g3401 ( 
.A(n_3099),
.B(n_3159),
.Y(n_3401)
);

CKINVDCx5p33_ASAP7_75t_R g3402 ( 
.A(n_3041),
.Y(n_3402)
);

NAND2xp5_ASAP7_75t_L g3403 ( 
.A(n_3278),
.B(n_1815),
.Y(n_3403)
);

AOI22xp5_ASAP7_75t_L g3404 ( 
.A1(n_3157),
.A2(n_3061),
.B1(n_3117),
.B2(n_3112),
.Y(n_3404)
);

AND2x6_ASAP7_75t_SL g3405 ( 
.A(n_3225),
.B(n_3222),
.Y(n_3405)
);

INVx1_ASAP7_75t_L g3406 ( 
.A(n_3092),
.Y(n_3406)
);

A2O1A1Ixp33_ASAP7_75t_L g3407 ( 
.A1(n_3129),
.A2(n_1838),
.B(n_1842),
.C(n_1835),
.Y(n_3407)
);

NAND2xp5_ASAP7_75t_SL g3408 ( 
.A(n_3175),
.B(n_3120),
.Y(n_3408)
);

OR2x6_ASAP7_75t_L g3409 ( 
.A(n_3268),
.B(n_1849),
.Y(n_3409)
);

OR2x6_ASAP7_75t_L g3410 ( 
.A(n_3155),
.B(n_1854),
.Y(n_3410)
);

INVx2_ASAP7_75t_L g3411 ( 
.A(n_3080),
.Y(n_3411)
);

INVx3_ASAP7_75t_L g3412 ( 
.A(n_3108),
.Y(n_3412)
);

INVx3_ASAP7_75t_L g3413 ( 
.A(n_3270),
.Y(n_3413)
);

NAND3xp33_ASAP7_75t_L g3414 ( 
.A(n_3189),
.B(n_1830),
.C(n_1828),
.Y(n_3414)
);

NOR2xp33_ASAP7_75t_L g3415 ( 
.A(n_3261),
.B(n_1832),
.Y(n_3415)
);

OR2x6_ASAP7_75t_L g3416 ( 
.A(n_3141),
.B(n_1860),
.Y(n_3416)
);

O2A1O1Ixp33_ASAP7_75t_L g3417 ( 
.A1(n_3185),
.A2(n_1866),
.B(n_1868),
.C(n_1862),
.Y(n_3417)
);

INVx1_ASAP7_75t_L g3418 ( 
.A(n_3109),
.Y(n_3418)
);

AOI21x1_ASAP7_75t_L g3419 ( 
.A1(n_3152),
.A2(n_1874),
.B(n_1870),
.Y(n_3419)
);

INVx2_ASAP7_75t_L g3420 ( 
.A(n_3119),
.Y(n_3420)
);

AOI22xp5_ASAP7_75t_L g3421 ( 
.A1(n_3233),
.A2(n_3269),
.B1(n_3241),
.B2(n_3140),
.Y(n_3421)
);

AOI22xp5_ASAP7_75t_L g3422 ( 
.A1(n_3269),
.A2(n_1834),
.B1(n_1837),
.B2(n_1833),
.Y(n_3422)
);

INVx4_ASAP7_75t_L g3423 ( 
.A(n_3141),
.Y(n_3423)
);

NAND2xp5_ASAP7_75t_L g3424 ( 
.A(n_3220),
.B(n_1840),
.Y(n_3424)
);

NAND2xp5_ASAP7_75t_L g3425 ( 
.A(n_3223),
.B(n_1841),
.Y(n_3425)
);

NAND2xp5_ASAP7_75t_L g3426 ( 
.A(n_3243),
.B(n_1843),
.Y(n_3426)
);

INVxp67_ASAP7_75t_L g3427 ( 
.A(n_3150),
.Y(n_3427)
);

INVx1_ASAP7_75t_L g3428 ( 
.A(n_3161),
.Y(n_3428)
);

NAND2xp5_ASAP7_75t_L g3429 ( 
.A(n_3260),
.B(n_1844),
.Y(n_3429)
);

INVx1_ASAP7_75t_L g3430 ( 
.A(n_3145),
.Y(n_3430)
);

NAND2xp5_ASAP7_75t_SL g3431 ( 
.A(n_3124),
.B(n_1852),
.Y(n_3431)
);

OR2x2_ASAP7_75t_L g3432 ( 
.A(n_3210),
.B(n_2385),
.Y(n_3432)
);

CKINVDCx5p33_ASAP7_75t_R g3433 ( 
.A(n_3234),
.Y(n_3433)
);

NAND2xp5_ASAP7_75t_L g3434 ( 
.A(n_3074),
.B(n_1853),
.Y(n_3434)
);

NAND2xp5_ASAP7_75t_L g3435 ( 
.A(n_3147),
.B(n_1859),
.Y(n_3435)
);

NOR2xp33_ASAP7_75t_SL g3436 ( 
.A(n_3126),
.B(n_2169),
.Y(n_3436)
);

NOR2xp33_ASAP7_75t_L g3437 ( 
.A(n_3062),
.B(n_1863),
.Y(n_3437)
);

AND2x2_ASAP7_75t_L g3438 ( 
.A(n_3165),
.B(n_3176),
.Y(n_3438)
);

INVx1_ASAP7_75t_L g3439 ( 
.A(n_3135),
.Y(n_3439)
);

NAND2xp5_ASAP7_75t_L g3440 ( 
.A(n_3081),
.B(n_1867),
.Y(n_3440)
);

INVx1_ASAP7_75t_L g3441 ( 
.A(n_3130),
.Y(n_3441)
);

NAND2xp5_ASAP7_75t_SL g3442 ( 
.A(n_3124),
.B(n_1872),
.Y(n_3442)
);

INVx2_ASAP7_75t_L g3443 ( 
.A(n_3131),
.Y(n_3443)
);

NOR2xp33_ASAP7_75t_L g3444 ( 
.A(n_3195),
.B(n_1873),
.Y(n_3444)
);

AOI22xp33_ASAP7_75t_L g3445 ( 
.A1(n_3168),
.A2(n_3248),
.B1(n_3199),
.B2(n_3211),
.Y(n_3445)
);

NOR2xp33_ASAP7_75t_L g3446 ( 
.A(n_3137),
.B(n_1876),
.Y(n_3446)
);

OR2x6_ASAP7_75t_L g3447 ( 
.A(n_3221),
.B(n_1880),
.Y(n_3447)
);

BUFx3_ASAP7_75t_L g3448 ( 
.A(n_3239),
.Y(n_3448)
);

INVx1_ASAP7_75t_L g3449 ( 
.A(n_3106),
.Y(n_3449)
);

INVx4_ASAP7_75t_L g3450 ( 
.A(n_3270),
.Y(n_3450)
);

INVx3_ASAP7_75t_L g3451 ( 
.A(n_3257),
.Y(n_3451)
);

NAND2xp5_ASAP7_75t_SL g3452 ( 
.A(n_3207),
.B(n_1877),
.Y(n_3452)
);

AOI22xp33_ASAP7_75t_L g3453 ( 
.A1(n_3227),
.A2(n_1884),
.B1(n_1894),
.B2(n_1882),
.Y(n_3453)
);

OAI221xp5_ASAP7_75t_L g3454 ( 
.A1(n_3263),
.A2(n_3192),
.B1(n_3184),
.B2(n_3171),
.C(n_3149),
.Y(n_3454)
);

NOR2xp33_ASAP7_75t_L g3455 ( 
.A(n_3208),
.B(n_1879),
.Y(n_3455)
);

INVx1_ASAP7_75t_L g3456 ( 
.A(n_3087),
.Y(n_3456)
);

INVx1_ASAP7_75t_L g3457 ( 
.A(n_3088),
.Y(n_3457)
);

INVx1_ASAP7_75t_L g3458 ( 
.A(n_3262),
.Y(n_3458)
);

INVxp33_ASAP7_75t_L g3459 ( 
.A(n_3218),
.Y(n_3459)
);

O2A1O1Ixp33_ASAP7_75t_L g3460 ( 
.A1(n_3122),
.A2(n_1904),
.B(n_1910),
.C(n_1901),
.Y(n_3460)
);

INVx2_ASAP7_75t_L g3461 ( 
.A(n_3079),
.Y(n_3461)
);

NOR3xp33_ASAP7_75t_L g3462 ( 
.A(n_3209),
.B(n_1883),
.C(n_1881),
.Y(n_3462)
);

INVx2_ASAP7_75t_L g3463 ( 
.A(n_3240),
.Y(n_3463)
);

INVx1_ASAP7_75t_L g3464 ( 
.A(n_3252),
.Y(n_3464)
);

NOR2xp33_ASAP7_75t_L g3465 ( 
.A(n_3051),
.B(n_3228),
.Y(n_3465)
);

INVx1_ASAP7_75t_L g3466 ( 
.A(n_3253),
.Y(n_3466)
);

INVx2_ASAP7_75t_SL g3467 ( 
.A(n_3259),
.Y(n_3467)
);

AND2x2_ASAP7_75t_L g3468 ( 
.A(n_3217),
.B(n_2279),
.Y(n_3468)
);

AND2x2_ASAP7_75t_L g3469 ( 
.A(n_3213),
.B(n_3219),
.Y(n_3469)
);

NAND2xp5_ASAP7_75t_L g3470 ( 
.A(n_3082),
.B(n_1885),
.Y(n_3470)
);

NAND2xp5_ASAP7_75t_L g3471 ( 
.A(n_3078),
.B(n_1886),
.Y(n_3471)
);

NAND2xp5_ASAP7_75t_L g3472 ( 
.A(n_3078),
.B(n_1887),
.Y(n_3472)
);

O2A1O1Ixp33_ASAP7_75t_L g3473 ( 
.A1(n_3200),
.A2(n_1922),
.B(n_1923),
.C(n_1916),
.Y(n_3473)
);

A2O1A1Ixp33_ASAP7_75t_L g3474 ( 
.A1(n_3127),
.A2(n_1928),
.B(n_1931),
.C(n_1926),
.Y(n_3474)
);

INVx1_ASAP7_75t_L g3475 ( 
.A(n_3276),
.Y(n_3475)
);

INVx2_ASAP7_75t_L g3476 ( 
.A(n_3266),
.Y(n_3476)
);

BUFx5_ASAP7_75t_L g3477 ( 
.A(n_3139),
.Y(n_3477)
);

NAND2xp5_ASAP7_75t_SL g3478 ( 
.A(n_3215),
.B(n_1888),
.Y(n_3478)
);

INVx1_ASAP7_75t_L g3479 ( 
.A(n_3274),
.Y(n_3479)
);

NOR2xp33_ASAP7_75t_L g3480 ( 
.A(n_3188),
.B(n_1889),
.Y(n_3480)
);

INVx1_ASAP7_75t_L g3481 ( 
.A(n_3139),
.Y(n_3481)
);

INVx2_ASAP7_75t_SL g3482 ( 
.A(n_3275),
.Y(n_3482)
);

NAND2xp5_ASAP7_75t_L g3483 ( 
.A(n_3205),
.B(n_1890),
.Y(n_3483)
);

INVx2_ASAP7_75t_L g3484 ( 
.A(n_3277),
.Y(n_3484)
);

INVx1_ASAP7_75t_L g3485 ( 
.A(n_3101),
.Y(n_3485)
);

NAND2xp5_ASAP7_75t_SL g3486 ( 
.A(n_3202),
.B(n_1893),
.Y(n_3486)
);

NAND2xp5_ASAP7_75t_SL g3487 ( 
.A(n_3224),
.B(n_1895),
.Y(n_3487)
);

CKINVDCx5p33_ASAP7_75t_R g3488 ( 
.A(n_3146),
.Y(n_3488)
);

NOR2xp33_ASAP7_75t_L g3489 ( 
.A(n_3196),
.B(n_1898),
.Y(n_3489)
);

INVxp67_ASAP7_75t_SL g3490 ( 
.A(n_3206),
.Y(n_3490)
);

NAND2xp5_ASAP7_75t_SL g3491 ( 
.A(n_3076),
.B(n_1905),
.Y(n_3491)
);

NAND2xp5_ASAP7_75t_L g3492 ( 
.A(n_3133),
.B(n_3138),
.Y(n_3492)
);

NAND2xp5_ASAP7_75t_L g3493 ( 
.A(n_3133),
.B(n_1906),
.Y(n_3493)
);

INVx2_ASAP7_75t_L g3494 ( 
.A(n_3183),
.Y(n_3494)
);

OAI21xp5_ASAP7_75t_L g3495 ( 
.A1(n_3101),
.A2(n_1937),
.B(n_1934),
.Y(n_3495)
);

AOI22xp5_ASAP7_75t_L g3496 ( 
.A1(n_3071),
.A2(n_1909),
.B1(n_1914),
.B2(n_1908),
.Y(n_3496)
);

NAND2xp5_ASAP7_75t_L g3497 ( 
.A(n_3052),
.B(n_1917),
.Y(n_3497)
);

AOI22xp33_ASAP7_75t_L g3498 ( 
.A1(n_3229),
.A2(n_1940),
.B1(n_1942),
.B2(n_1938),
.Y(n_3498)
);

NOR2xp33_ASAP7_75t_L g3499 ( 
.A(n_3226),
.B(n_1919),
.Y(n_3499)
);

AND2x6_ASAP7_75t_SL g3500 ( 
.A(n_3193),
.B(n_1944),
.Y(n_3500)
);

BUFx2_ASAP7_75t_L g3501 ( 
.A(n_3154),
.Y(n_3501)
);

NAND2xp5_ASAP7_75t_SL g3502 ( 
.A(n_3077),
.B(n_1920),
.Y(n_3502)
);

INVx1_ASAP7_75t_L g3503 ( 
.A(n_3048),
.Y(n_3503)
);

NOR2xp33_ASAP7_75t_L g3504 ( 
.A(n_3043),
.B(n_1924),
.Y(n_3504)
);

AOI21xp5_ASAP7_75t_L g3505 ( 
.A1(n_3072),
.A2(n_1962),
.B(n_1957),
.Y(n_3505)
);

NOR2xp33_ASAP7_75t_L g3506 ( 
.A(n_3043),
.B(n_1927),
.Y(n_3506)
);

NOR2xp33_ASAP7_75t_SL g3507 ( 
.A(n_3204),
.B(n_2279),
.Y(n_3507)
);

INVx1_ASAP7_75t_L g3508 ( 
.A(n_3048),
.Y(n_3508)
);

BUFx3_ASAP7_75t_L g3509 ( 
.A(n_3084),
.Y(n_3509)
);

INVx1_ASAP7_75t_L g3510 ( 
.A(n_3048),
.Y(n_3510)
);

AND2x4_ASAP7_75t_SL g3511 ( 
.A(n_3158),
.B(n_2439),
.Y(n_3511)
);

NAND2xp5_ASAP7_75t_SL g3512 ( 
.A(n_3077),
.B(n_1933),
.Y(n_3512)
);

NAND2xp5_ASAP7_75t_SL g3513 ( 
.A(n_3077),
.B(n_1946),
.Y(n_3513)
);

BUFx3_ASAP7_75t_L g3514 ( 
.A(n_3084),
.Y(n_3514)
);

NAND2xp5_ASAP7_75t_L g3515 ( 
.A(n_3153),
.B(n_1948),
.Y(n_3515)
);

BUFx6f_ASAP7_75t_L g3516 ( 
.A(n_3049),
.Y(n_3516)
);

NAND2xp5_ASAP7_75t_L g3517 ( 
.A(n_3153),
.B(n_1953),
.Y(n_3517)
);

AO221x1_ASAP7_75t_L g3518 ( 
.A1(n_3248),
.A2(n_1977),
.B1(n_1979),
.B2(n_1970),
.C(n_1965),
.Y(n_3518)
);

NAND2xp5_ASAP7_75t_L g3519 ( 
.A(n_3153),
.B(n_1956),
.Y(n_3519)
);

NAND2xp5_ASAP7_75t_L g3520 ( 
.A(n_3153),
.B(n_1959),
.Y(n_3520)
);

AOI22xp33_ASAP7_75t_L g3521 ( 
.A1(n_3142),
.A2(n_1988),
.B1(n_1989),
.B2(n_1983),
.Y(n_3521)
);

AOI22xp33_ASAP7_75t_L g3522 ( 
.A1(n_3142),
.A2(n_1998),
.B1(n_2002),
.B2(n_1994),
.Y(n_3522)
);

NAND2xp5_ASAP7_75t_L g3523 ( 
.A(n_3153),
.B(n_1960),
.Y(n_3523)
);

AOI22xp5_ASAP7_75t_L g3524 ( 
.A1(n_3142),
.A2(n_1964),
.B1(n_1967),
.B2(n_1963),
.Y(n_3524)
);

AOI22xp5_ASAP7_75t_L g3525 ( 
.A1(n_3142),
.A2(n_1972),
.B1(n_1973),
.B2(n_1971),
.Y(n_3525)
);

INVx2_ASAP7_75t_SL g3526 ( 
.A(n_3121),
.Y(n_3526)
);

A2O1A1Ixp33_ASAP7_75t_L g3527 ( 
.A1(n_3083),
.A2(n_2025),
.B(n_2028),
.C(n_2020),
.Y(n_3527)
);

INVx2_ASAP7_75t_SL g3528 ( 
.A(n_3121),
.Y(n_3528)
);

AND2x2_ASAP7_75t_L g3529 ( 
.A(n_3083),
.B(n_2439),
.Y(n_3529)
);

INVx2_ASAP7_75t_SL g3530 ( 
.A(n_3121),
.Y(n_3530)
);

NOR2xp33_ASAP7_75t_L g3531 ( 
.A(n_3043),
.B(n_1974),
.Y(n_3531)
);

NAND2xp5_ASAP7_75t_L g3532 ( 
.A(n_3153),
.B(n_1978),
.Y(n_3532)
);

INVx2_ASAP7_75t_SL g3533 ( 
.A(n_3121),
.Y(n_3533)
);

NOR2xp33_ASAP7_75t_L g3534 ( 
.A(n_3043),
.B(n_1980),
.Y(n_3534)
);

NAND2xp5_ASAP7_75t_L g3535 ( 
.A(n_3153),
.B(n_1984),
.Y(n_3535)
);

NOR2xp33_ASAP7_75t_L g3536 ( 
.A(n_3043),
.B(n_1985),
.Y(n_3536)
);

NOR2xp33_ASAP7_75t_L g3537 ( 
.A(n_3043),
.B(n_1992),
.Y(n_3537)
);

AOI22xp5_ASAP7_75t_L g3538 ( 
.A1(n_3142),
.A2(n_1996),
.B1(n_1997),
.B2(n_1993),
.Y(n_3538)
);

BUFx12f_ASAP7_75t_SL g3539 ( 
.A(n_3141),
.Y(n_3539)
);

AOI21xp5_ASAP7_75t_L g3540 ( 
.A1(n_3072),
.A2(n_2031),
.B(n_2030),
.Y(n_3540)
);

NAND2xp5_ASAP7_75t_L g3541 ( 
.A(n_3153),
.B(n_1999),
.Y(n_3541)
);

NAND2xp5_ASAP7_75t_L g3542 ( 
.A(n_3153),
.B(n_2000),
.Y(n_3542)
);

INVx3_ASAP7_75t_L g3543 ( 
.A(n_3049),
.Y(n_3543)
);

INVx2_ASAP7_75t_L g3544 ( 
.A(n_3040),
.Y(n_3544)
);

INVx2_ASAP7_75t_L g3545 ( 
.A(n_3040),
.Y(n_3545)
);

AND2x2_ASAP7_75t_L g3546 ( 
.A(n_3083),
.B(n_2455),
.Y(n_3546)
);

NOR2xp33_ASAP7_75t_L g3547 ( 
.A(n_3043),
.B(n_2003),
.Y(n_3547)
);

INVx1_ASAP7_75t_L g3548 ( 
.A(n_3048),
.Y(n_3548)
);

NAND2xp5_ASAP7_75t_SL g3549 ( 
.A(n_3077),
.B(n_2004),
.Y(n_3549)
);

AOI21xp5_ASAP7_75t_L g3550 ( 
.A1(n_3325),
.A2(n_2038),
.B(n_2037),
.Y(n_3550)
);

OAI21xp5_ASAP7_75t_L g3551 ( 
.A1(n_3299),
.A2(n_2047),
.B(n_2040),
.Y(n_3551)
);

AOI21xp5_ASAP7_75t_L g3552 ( 
.A1(n_3401),
.A2(n_2050),
.B(n_2049),
.Y(n_3552)
);

NAND2xp5_ASAP7_75t_SL g3553 ( 
.A(n_3347),
.B(n_2005),
.Y(n_3553)
);

AOI21xp5_ASAP7_75t_L g3554 ( 
.A1(n_3408),
.A2(n_2057),
.B(n_2055),
.Y(n_3554)
);

AOI21xp5_ASAP7_75t_L g3555 ( 
.A1(n_3353),
.A2(n_2060),
.B(n_2058),
.Y(n_3555)
);

BUFx6f_ASAP7_75t_L g3556 ( 
.A(n_3333),
.Y(n_3556)
);

HB1xp67_ASAP7_75t_L g3557 ( 
.A(n_3539),
.Y(n_3557)
);

OAI22xp5_ASAP7_75t_L g3558 ( 
.A1(n_3311),
.A2(n_3289),
.B1(n_3390),
.B2(n_3404),
.Y(n_3558)
);

O2A1O1Ixp33_ASAP7_75t_L g3559 ( 
.A1(n_3295),
.A2(n_2070),
.B(n_2076),
.C(n_2065),
.Y(n_3559)
);

NAND2xp5_ASAP7_75t_L g3560 ( 
.A(n_3406),
.B(n_2006),
.Y(n_3560)
);

AND2x2_ASAP7_75t_L g3561 ( 
.A(n_3529),
.B(n_2408),
.Y(n_3561)
);

INVx3_ASAP7_75t_L g3562 ( 
.A(n_3328),
.Y(n_3562)
);

NAND2xp5_ASAP7_75t_L g3563 ( 
.A(n_3504),
.B(n_2007),
.Y(n_3563)
);

NOR2xp33_ASAP7_75t_L g3564 ( 
.A(n_3369),
.B(n_2009),
.Y(n_3564)
);

INVx2_ASAP7_75t_L g3565 ( 
.A(n_3292),
.Y(n_3565)
);

INVx2_ASAP7_75t_SL g3566 ( 
.A(n_3469),
.Y(n_3566)
);

AND2x2_ASAP7_75t_L g3567 ( 
.A(n_3546),
.B(n_2440),
.Y(n_3567)
);

A2O1A1Ixp33_ASAP7_75t_L g3568 ( 
.A1(n_3377),
.A2(n_2084),
.B(n_2088),
.C(n_2082),
.Y(n_3568)
);

O2A1O1Ixp33_ASAP7_75t_L g3569 ( 
.A1(n_3297),
.A2(n_2091),
.B(n_2092),
.C(n_2089),
.Y(n_3569)
);

NAND2xp5_ASAP7_75t_L g3570 ( 
.A(n_3506),
.B(n_2010),
.Y(n_3570)
);

AOI21xp5_ASAP7_75t_L g3571 ( 
.A1(n_3298),
.A2(n_2095),
.B(n_2094),
.Y(n_3571)
);

NOR2xp33_ASAP7_75t_L g3572 ( 
.A(n_3283),
.B(n_2014),
.Y(n_3572)
);

INVx2_ASAP7_75t_SL g3573 ( 
.A(n_3344),
.Y(n_3573)
);

INVx3_ASAP7_75t_L g3574 ( 
.A(n_3302),
.Y(n_3574)
);

NAND2xp5_ASAP7_75t_SL g3575 ( 
.A(n_3373),
.B(n_2018),
.Y(n_3575)
);

BUFx6f_ASAP7_75t_L g3576 ( 
.A(n_3333),
.Y(n_3576)
);

NAND2xp5_ASAP7_75t_L g3577 ( 
.A(n_3531),
.B(n_2021),
.Y(n_3577)
);

OAI21x1_ASAP7_75t_SL g3578 ( 
.A1(n_3419),
.A2(n_2124),
.B(n_2120),
.Y(n_3578)
);

O2A1O1Ixp33_ASAP7_75t_SL g3579 ( 
.A1(n_3407),
.A2(n_2130),
.B(n_2131),
.C(n_2129),
.Y(n_3579)
);

NAND2xp5_ASAP7_75t_L g3580 ( 
.A(n_3534),
.B(n_2023),
.Y(n_3580)
);

NAND2xp5_ASAP7_75t_SL g3581 ( 
.A(n_3303),
.B(n_2024),
.Y(n_3581)
);

NAND2xp5_ASAP7_75t_L g3582 ( 
.A(n_3536),
.B(n_2027),
.Y(n_3582)
);

INVx2_ASAP7_75t_L g3583 ( 
.A(n_3544),
.Y(n_3583)
);

NAND2xp5_ASAP7_75t_L g3584 ( 
.A(n_3537),
.B(n_2029),
.Y(n_3584)
);

INVx3_ASAP7_75t_L g3585 ( 
.A(n_3545),
.Y(n_3585)
);

NAND2xp5_ASAP7_75t_SL g3586 ( 
.A(n_3526),
.B(n_2032),
.Y(n_3586)
);

BUFx4f_ASAP7_75t_L g3587 ( 
.A(n_3304),
.Y(n_3587)
);

AOI21xp5_ASAP7_75t_L g3588 ( 
.A1(n_3454),
.A2(n_2172),
.B(n_2168),
.Y(n_3588)
);

NOR2xp33_ASAP7_75t_L g3589 ( 
.A(n_3345),
.B(n_2034),
.Y(n_3589)
);

AND2x4_ASAP7_75t_L g3590 ( 
.A(n_3494),
.B(n_2177),
.Y(n_3590)
);

INVx3_ASAP7_75t_L g3591 ( 
.A(n_3398),
.Y(n_3591)
);

OAI21xp5_ASAP7_75t_L g3592 ( 
.A1(n_3435),
.A2(n_2191),
.B(n_2188),
.Y(n_3592)
);

A2O1A1Ixp33_ASAP7_75t_L g3593 ( 
.A1(n_3378),
.A2(n_3444),
.B(n_3415),
.C(n_3437),
.Y(n_3593)
);

NAND2xp5_ASAP7_75t_L g3594 ( 
.A(n_3547),
.B(n_2039),
.Y(n_3594)
);

AOI21xp5_ASAP7_75t_L g3595 ( 
.A1(n_3368),
.A2(n_2209),
.B(n_2207),
.Y(n_3595)
);

AOI21xp5_ASAP7_75t_L g3596 ( 
.A1(n_3397),
.A2(n_2212),
.B(n_2210),
.Y(n_3596)
);

NAND2xp5_ASAP7_75t_L g3597 ( 
.A(n_3389),
.B(n_2041),
.Y(n_3597)
);

INVx2_ASAP7_75t_L g3598 ( 
.A(n_3314),
.Y(n_3598)
);

O2A1O1Ixp33_ASAP7_75t_SL g3599 ( 
.A1(n_3301),
.A2(n_3334),
.B(n_3527),
.C(n_3381),
.Y(n_3599)
);

NAND2xp5_ASAP7_75t_SL g3600 ( 
.A(n_3528),
.B(n_2042),
.Y(n_3600)
);

NOR2x1_ASAP7_75t_L g3601 ( 
.A(n_3423),
.B(n_2231),
.Y(n_3601)
);

AOI21xp5_ASAP7_75t_L g3602 ( 
.A1(n_3382),
.A2(n_2233),
.B(n_2232),
.Y(n_3602)
);

NAND2xp33_ASAP7_75t_L g3603 ( 
.A(n_3477),
.B(n_3402),
.Y(n_3603)
);

INVx3_ASAP7_75t_L g3604 ( 
.A(n_3399),
.Y(n_3604)
);

INVx1_ASAP7_75t_L g3605 ( 
.A(n_3281),
.Y(n_3605)
);

BUFx2_ASAP7_75t_L g3606 ( 
.A(n_3340),
.Y(n_3606)
);

AND2x2_ASAP7_75t_L g3607 ( 
.A(n_3296),
.B(n_3358),
.Y(n_3607)
);

AOI21xp5_ASAP7_75t_L g3608 ( 
.A1(n_3395),
.A2(n_2274),
.B(n_2265),
.Y(n_3608)
);

CKINVDCx10_ASAP7_75t_R g3609 ( 
.A(n_3410),
.Y(n_3609)
);

AOI21xp5_ASAP7_75t_L g3610 ( 
.A1(n_3400),
.A2(n_2283),
.B(n_2275),
.Y(n_3610)
);

NAND2xp5_ASAP7_75t_SL g3611 ( 
.A(n_3530),
.B(n_2048),
.Y(n_3611)
);

INVx2_ASAP7_75t_SL g3612 ( 
.A(n_3533),
.Y(n_3612)
);

NAND2xp5_ASAP7_75t_L g3613 ( 
.A(n_3320),
.B(n_3305),
.Y(n_3613)
);

AOI21xp5_ASAP7_75t_L g3614 ( 
.A1(n_3284),
.A2(n_2317),
.B(n_2307),
.Y(n_3614)
);

NOR2xp33_ASAP7_75t_L g3615 ( 
.A(n_3317),
.B(n_3350),
.Y(n_3615)
);

AO21x1_ASAP7_75t_L g3616 ( 
.A1(n_3323),
.A2(n_2322),
.B(n_2321),
.Y(n_3616)
);

NAND2xp5_ASAP7_75t_L g3617 ( 
.A(n_3326),
.B(n_3331),
.Y(n_3617)
);

NAND2xp5_ASAP7_75t_L g3618 ( 
.A(n_3346),
.B(n_2063),
.Y(n_3618)
);

NAND2xp5_ASAP7_75t_L g3619 ( 
.A(n_3370),
.B(n_2074),
.Y(n_3619)
);

NAND2xp5_ASAP7_75t_L g3620 ( 
.A(n_3503),
.B(n_3508),
.Y(n_3620)
);

NOR2xp33_ASAP7_75t_L g3621 ( 
.A(n_3313),
.B(n_2077),
.Y(n_3621)
);

NAND2xp5_ASAP7_75t_L g3622 ( 
.A(n_3510),
.B(n_2078),
.Y(n_3622)
);

O2A1O1Ixp33_ASAP7_75t_L g3623 ( 
.A1(n_3474),
.A2(n_2337),
.B(n_2338),
.C(n_2336),
.Y(n_3623)
);

A2O1A1Ixp33_ASAP7_75t_L g3624 ( 
.A1(n_3445),
.A2(n_2353),
.B(n_2359),
.C(n_2352),
.Y(n_3624)
);

CKINVDCx5p33_ASAP7_75t_R g3625 ( 
.A(n_3306),
.Y(n_3625)
);

INVx2_ASAP7_75t_L g3626 ( 
.A(n_3316),
.Y(n_3626)
);

AOI21xp5_ASAP7_75t_L g3627 ( 
.A1(n_3290),
.A2(n_2368),
.B(n_2364),
.Y(n_3627)
);

NAND2xp5_ASAP7_75t_SL g3628 ( 
.A(n_3329),
.B(n_2087),
.Y(n_3628)
);

BUFx12f_ASAP7_75t_L g3629 ( 
.A(n_3361),
.Y(n_3629)
);

AND2x2_ASAP7_75t_L g3630 ( 
.A(n_3363),
.B(n_2090),
.Y(n_3630)
);

INVx1_ASAP7_75t_L g3631 ( 
.A(n_3548),
.Y(n_3631)
);

A2O1A1Ixp33_ASAP7_75t_L g3632 ( 
.A1(n_3388),
.A2(n_3446),
.B(n_3465),
.C(n_3421),
.Y(n_3632)
);

OAI21xp33_ASAP7_75t_L g3633 ( 
.A1(n_3294),
.A2(n_2102),
.B(n_2099),
.Y(n_3633)
);

O2A1O1Ixp33_ASAP7_75t_L g3634 ( 
.A1(n_3332),
.A2(n_2373),
.B(n_2378),
.C(n_2372),
.Y(n_3634)
);

A2O1A1Ixp33_ASAP7_75t_L g3635 ( 
.A1(n_3282),
.A2(n_2397),
.B(n_2399),
.C(n_2381),
.Y(n_3635)
);

NOR2xp33_ASAP7_75t_SL g3636 ( 
.A(n_3488),
.B(n_2104),
.Y(n_3636)
);

AOI22xp5_ASAP7_75t_L g3637 ( 
.A1(n_3336),
.A2(n_2107),
.B1(n_2108),
.B2(n_2106),
.Y(n_3637)
);

AND2x4_ASAP7_75t_L g3638 ( 
.A(n_3420),
.B(n_2403),
.Y(n_3638)
);

BUFx6f_ASAP7_75t_L g3639 ( 
.A(n_3392),
.Y(n_3639)
);

O2A1O1Ixp33_ASAP7_75t_L g3640 ( 
.A1(n_3337),
.A2(n_2418),
.B(n_2421),
.C(n_2414),
.Y(n_3640)
);

AOI22xp33_ASAP7_75t_L g3641 ( 
.A1(n_3518),
.A2(n_2423),
.B1(n_2424),
.B2(n_2422),
.Y(n_3641)
);

NOR2xp33_ASAP7_75t_L g3642 ( 
.A(n_3312),
.B(n_3352),
.Y(n_3642)
);

CKINVDCx20_ASAP7_75t_R g3643 ( 
.A(n_3433),
.Y(n_3643)
);

AOI22xp33_ASAP7_75t_L g3644 ( 
.A1(n_3391),
.A2(n_2438),
.B1(n_2444),
.B2(n_2437),
.Y(n_3644)
);

NAND2xp5_ASAP7_75t_L g3645 ( 
.A(n_3515),
.B(n_3517),
.Y(n_3645)
);

NAND2xp5_ASAP7_75t_L g3646 ( 
.A(n_3519),
.B(n_2114),
.Y(n_3646)
);

NAND2xp5_ASAP7_75t_L g3647 ( 
.A(n_3520),
.B(n_3523),
.Y(n_3647)
);

NAND2xp5_ASAP7_75t_L g3648 ( 
.A(n_3532),
.B(n_2118),
.Y(n_3648)
);

HB1xp67_ASAP7_75t_L g3649 ( 
.A(n_3307),
.Y(n_3649)
);

NAND2xp5_ASAP7_75t_L g3650 ( 
.A(n_3535),
.B(n_2121),
.Y(n_3650)
);

NOR2xp33_ASAP7_75t_L g3651 ( 
.A(n_3489),
.B(n_2122),
.Y(n_3651)
);

INVx2_ASAP7_75t_SL g3652 ( 
.A(n_3392),
.Y(n_3652)
);

NAND2xp5_ASAP7_75t_L g3653 ( 
.A(n_3541),
.B(n_2125),
.Y(n_3653)
);

NAND2xp5_ASAP7_75t_L g3654 ( 
.A(n_3542),
.B(n_2127),
.Y(n_3654)
);

OAI21xp5_ASAP7_75t_L g3655 ( 
.A1(n_3357),
.A2(n_2134),
.B(n_2128),
.Y(n_3655)
);

AOI22xp5_ASAP7_75t_L g3656 ( 
.A1(n_3438),
.A2(n_2136),
.B1(n_2138),
.B2(n_2135),
.Y(n_3656)
);

NAND2xp5_ASAP7_75t_SL g3657 ( 
.A(n_3380),
.B(n_2139),
.Y(n_3657)
);

OAI21xp5_ASAP7_75t_L g3658 ( 
.A1(n_3300),
.A2(n_2146),
.B(n_2142),
.Y(n_3658)
);

NAND2xp5_ASAP7_75t_L g3659 ( 
.A(n_3375),
.B(n_2148),
.Y(n_3659)
);

O2A1O1Ixp33_ASAP7_75t_L g3660 ( 
.A1(n_3426),
.A2(n_2151),
.B(n_2153),
.C(n_2149),
.Y(n_3660)
);

INVxp33_ASAP7_75t_L g3661 ( 
.A(n_3315),
.Y(n_3661)
);

AOI21xp5_ASAP7_75t_L g3662 ( 
.A1(n_3351),
.A2(n_2158),
.B(n_2157),
.Y(n_3662)
);

INVx1_ASAP7_75t_L g3663 ( 
.A(n_3385),
.Y(n_3663)
);

CKINVDCx5p33_ASAP7_75t_R g3664 ( 
.A(n_3509),
.Y(n_3664)
);

NOR2xp33_ASAP7_75t_L g3665 ( 
.A(n_3427),
.B(n_2160),
.Y(n_3665)
);

NAND2x1_ASAP7_75t_L g3666 ( 
.A(n_3450),
.B(n_379),
.Y(n_3666)
);

BUFx3_ASAP7_75t_L g3667 ( 
.A(n_3514),
.Y(n_3667)
);

NAND2xp5_ASAP7_75t_L g3668 ( 
.A(n_3287),
.B(n_2161),
.Y(n_3668)
);

AOI21xp5_ASAP7_75t_L g3669 ( 
.A1(n_3359),
.A2(n_2167),
.B(n_2163),
.Y(n_3669)
);

INVx2_ASAP7_75t_L g3670 ( 
.A(n_3376),
.Y(n_3670)
);

AOI21x1_ASAP7_75t_L g3671 ( 
.A1(n_3411),
.A2(n_3394),
.B(n_3393),
.Y(n_3671)
);

BUFx3_ASAP7_75t_L g3672 ( 
.A(n_3364),
.Y(n_3672)
);

NAND2xp5_ASAP7_75t_SL g3673 ( 
.A(n_3477),
.B(n_2170),
.Y(n_3673)
);

AOI21xp5_ASAP7_75t_L g3674 ( 
.A1(n_3379),
.A2(n_2174),
.B(n_2173),
.Y(n_3674)
);

NAND2xp5_ASAP7_75t_SL g3675 ( 
.A(n_3477),
.B(n_2175),
.Y(n_3675)
);

NAND2xp5_ASAP7_75t_L g3676 ( 
.A(n_3348),
.B(n_2176),
.Y(n_3676)
);

NAND2xp5_ASAP7_75t_L g3677 ( 
.A(n_3403),
.B(n_2179),
.Y(n_3677)
);

O2A1O1Ixp33_ASAP7_75t_L g3678 ( 
.A1(n_3429),
.A2(n_2182),
.B(n_2183),
.C(n_2180),
.Y(n_3678)
);

NOR3xp33_ASAP7_75t_L g3679 ( 
.A(n_3362),
.B(n_2185),
.C(n_2184),
.Y(n_3679)
);

NAND2xp5_ASAP7_75t_SL g3680 ( 
.A(n_3443),
.B(n_3349),
.Y(n_3680)
);

OAI21xp5_ASAP7_75t_L g3681 ( 
.A1(n_3440),
.A2(n_2192),
.B(n_2186),
.Y(n_3681)
);

A2O1A1Ixp33_ASAP7_75t_L g3682 ( 
.A1(n_3455),
.A2(n_2194),
.B(n_2195),
.C(n_2193),
.Y(n_3682)
);

INVx2_ASAP7_75t_L g3683 ( 
.A(n_3384),
.Y(n_3683)
);

AND2x4_ASAP7_75t_L g3684 ( 
.A(n_3461),
.B(n_379),
.Y(n_3684)
);

AOI21xp5_ASAP7_75t_L g3685 ( 
.A1(n_3321),
.A2(n_2197),
.B(n_2196),
.Y(n_3685)
);

NAND2xp5_ASAP7_75t_L g3686 ( 
.A(n_3521),
.B(n_3522),
.Y(n_3686)
);

NAND2x1_ASAP7_75t_L g3687 ( 
.A(n_3279),
.B(n_380),
.Y(n_3687)
);

INVx1_ASAP7_75t_L g3688 ( 
.A(n_3430),
.Y(n_3688)
);

AOI21xp5_ASAP7_75t_L g3689 ( 
.A1(n_3322),
.A2(n_2199),
.B(n_2198),
.Y(n_3689)
);

NAND2xp5_ASAP7_75t_L g3690 ( 
.A(n_3505),
.B(n_2202),
.Y(n_3690)
);

AOI21xp33_ASAP7_75t_L g3691 ( 
.A1(n_3360),
.A2(n_2205),
.B(n_2204),
.Y(n_3691)
);

NAND2xp5_ASAP7_75t_SL g3692 ( 
.A(n_3341),
.B(n_2211),
.Y(n_3692)
);

NAND2xp5_ASAP7_75t_L g3693 ( 
.A(n_3540),
.B(n_2213),
.Y(n_3693)
);

NAND2xp5_ASAP7_75t_L g3694 ( 
.A(n_3327),
.B(n_2215),
.Y(n_3694)
);

CKINVDCx10_ASAP7_75t_R g3695 ( 
.A(n_3410),
.Y(n_3695)
);

OAI321xp33_ASAP7_75t_L g3696 ( 
.A1(n_3495),
.A2(n_2219),
.A3(n_2217),
.B1(n_2220),
.B2(n_2218),
.C(n_2216),
.Y(n_3696)
);

INVxp67_ASAP7_75t_L g3697 ( 
.A(n_3432),
.Y(n_3697)
);

AOI22xp5_ASAP7_75t_L g3698 ( 
.A1(n_3354),
.A2(n_2225),
.B1(n_2229),
.B2(n_2224),
.Y(n_3698)
);

NOR2xp33_ASAP7_75t_L g3699 ( 
.A(n_3291),
.B(n_2230),
.Y(n_3699)
);

NAND2xp5_ASAP7_75t_L g3700 ( 
.A(n_3335),
.B(n_2234),
.Y(n_3700)
);

AOI21xp5_ASAP7_75t_L g3701 ( 
.A1(n_3338),
.A2(n_2237),
.B(n_2235),
.Y(n_3701)
);

A2O1A1Ixp33_ASAP7_75t_L g3702 ( 
.A1(n_3286),
.A2(n_2243),
.B(n_2244),
.C(n_2238),
.Y(n_3702)
);

AOI21xp5_ASAP7_75t_L g3703 ( 
.A1(n_3342),
.A2(n_2247),
.B(n_2245),
.Y(n_3703)
);

NAND2xp5_ASAP7_75t_L g3704 ( 
.A(n_3343),
.B(n_2248),
.Y(n_3704)
);

AOI21xp5_ASAP7_75t_L g3705 ( 
.A1(n_3365),
.A2(n_2252),
.B(n_2250),
.Y(n_3705)
);

AOI21xp5_ASAP7_75t_L g3706 ( 
.A1(n_3366),
.A2(n_2254),
.B(n_2253),
.Y(n_3706)
);

NOR2x1_ASAP7_75t_R g3707 ( 
.A(n_3490),
.B(n_2257),
.Y(n_3707)
);

NAND2xp5_ASAP7_75t_SL g3708 ( 
.A(n_3441),
.B(n_2258),
.Y(n_3708)
);

NOR2xp67_ASAP7_75t_SL g3709 ( 
.A(n_3451),
.B(n_2259),
.Y(n_3709)
);

OAI22xp5_ASAP7_75t_L g3710 ( 
.A1(n_3439),
.A2(n_2261),
.B1(n_2262),
.B2(n_2260),
.Y(n_3710)
);

O2A1O1Ixp33_ASAP7_75t_L g3711 ( 
.A1(n_3417),
.A2(n_2264),
.B(n_2268),
.C(n_2263),
.Y(n_3711)
);

INVx3_ASAP7_75t_L g3712 ( 
.A(n_3516),
.Y(n_3712)
);

AOI22xp5_ASAP7_75t_L g3713 ( 
.A1(n_3355),
.A2(n_2271),
.B1(n_2276),
.B2(n_2270),
.Y(n_3713)
);

NAND2xp5_ASAP7_75t_SL g3714 ( 
.A(n_3468),
.B(n_2285),
.Y(n_3714)
);

BUFx6f_ASAP7_75t_L g3715 ( 
.A(n_3516),
.Y(n_3715)
);

AND2x2_ASAP7_75t_L g3716 ( 
.A(n_3308),
.B(n_2286),
.Y(n_3716)
);

NOR3xp33_ASAP7_75t_L g3717 ( 
.A(n_3310),
.B(n_2291),
.C(n_2290),
.Y(n_3717)
);

OAI22xp5_ASAP7_75t_L g3718 ( 
.A1(n_3449),
.A2(n_2298),
.B1(n_2299),
.B2(n_2296),
.Y(n_3718)
);

AO21x1_ASAP7_75t_L g3719 ( 
.A1(n_3330),
.A2(n_383),
.B(n_381),
.Y(n_3719)
);

INVx1_ASAP7_75t_L g3720 ( 
.A(n_3456),
.Y(n_3720)
);

AOI21xp5_ASAP7_75t_L g3721 ( 
.A1(n_3470),
.A2(n_2301),
.B(n_2300),
.Y(n_3721)
);

AND2x4_ASAP7_75t_L g3722 ( 
.A(n_3482),
.B(n_383),
.Y(n_3722)
);

NAND2xp5_ASAP7_75t_L g3723 ( 
.A(n_3480),
.B(n_2304),
.Y(n_3723)
);

NAND2xp5_ASAP7_75t_SL g3724 ( 
.A(n_3424),
.B(n_2305),
.Y(n_3724)
);

INVx2_ASAP7_75t_SL g3725 ( 
.A(n_3484),
.Y(n_3725)
);

HB1xp67_ASAP7_75t_L g3726 ( 
.A(n_3501),
.Y(n_3726)
);

NOR2xp33_ASAP7_75t_L g3727 ( 
.A(n_3293),
.B(n_2306),
.Y(n_3727)
);

AOI21xp5_ASAP7_75t_L g3728 ( 
.A1(n_3434),
.A2(n_2311),
.B(n_2310),
.Y(n_3728)
);

OAI21xp5_ASAP7_75t_L g3729 ( 
.A1(n_3371),
.A2(n_2313),
.B(n_2312),
.Y(n_3729)
);

AOI21xp5_ASAP7_75t_L g3730 ( 
.A1(n_3288),
.A2(n_2315),
.B(n_2314),
.Y(n_3730)
);

NAND2xp5_ASAP7_75t_SL g3731 ( 
.A(n_3425),
.B(n_2316),
.Y(n_3731)
);

NAND2xp5_ASAP7_75t_L g3732 ( 
.A(n_3524),
.B(n_2332),
.Y(n_3732)
);

NOR2xp33_ASAP7_75t_L g3733 ( 
.A(n_3459),
.B(n_2333),
.Y(n_3733)
);

AOI21xp5_ASAP7_75t_L g3734 ( 
.A1(n_3486),
.A2(n_2347),
.B(n_2345),
.Y(n_3734)
);

NAND2xp5_ASAP7_75t_L g3735 ( 
.A(n_3525),
.B(n_2348),
.Y(n_3735)
);

NAND2xp5_ASAP7_75t_L g3736 ( 
.A(n_3538),
.B(n_2349),
.Y(n_3736)
);

NAND2xp5_ASAP7_75t_L g3737 ( 
.A(n_3453),
.B(n_2350),
.Y(n_3737)
);

NAND2xp5_ASAP7_75t_L g3738 ( 
.A(n_3498),
.B(n_2351),
.Y(n_3738)
);

NAND2xp5_ASAP7_75t_L g3739 ( 
.A(n_3462),
.B(n_2356),
.Y(n_3739)
);

O2A1O1Ixp33_ASAP7_75t_L g3740 ( 
.A1(n_3478),
.A2(n_2366),
.B(n_2370),
.C(n_2361),
.Y(n_3740)
);

INVx2_ASAP7_75t_L g3741 ( 
.A(n_3457),
.Y(n_3741)
);

BUFx6f_ASAP7_75t_L g3742 ( 
.A(n_3448),
.Y(n_3742)
);

AND2x2_ASAP7_75t_L g3743 ( 
.A(n_3447),
.B(n_2376),
.Y(n_3743)
);

AOI21xp5_ASAP7_75t_L g3744 ( 
.A1(n_3418),
.A2(n_2379),
.B(n_2377),
.Y(n_3744)
);

OAI22xp5_ASAP7_75t_L g3745 ( 
.A1(n_3458),
.A2(n_2387),
.B1(n_2388),
.B2(n_2384),
.Y(n_3745)
);

INVx3_ASAP7_75t_L g3746 ( 
.A(n_3356),
.Y(n_3746)
);

AOI21xp5_ASAP7_75t_L g3747 ( 
.A1(n_3452),
.A2(n_2390),
.B(n_2389),
.Y(n_3747)
);

AOI21x1_ASAP7_75t_L g3748 ( 
.A1(n_3502),
.A2(n_385),
.B(n_384),
.Y(n_3748)
);

INVx1_ASAP7_75t_L g3749 ( 
.A(n_3367),
.Y(n_3749)
);

NAND2xp5_ASAP7_75t_L g3750 ( 
.A(n_3374),
.B(n_3481),
.Y(n_3750)
);

AND2x2_ASAP7_75t_L g3751 ( 
.A(n_3499),
.B(n_2391),
.Y(n_3751)
);

AOI21xp5_ASAP7_75t_L g3752 ( 
.A1(n_3428),
.A2(n_2395),
.B(n_2392),
.Y(n_3752)
);

AOI21xp5_ASAP7_75t_L g3753 ( 
.A1(n_3309),
.A2(n_2407),
.B(n_2405),
.Y(n_3753)
);

CKINVDCx5p33_ASAP7_75t_R g3754 ( 
.A(n_3405),
.Y(n_3754)
);

AOI21xp5_ASAP7_75t_L g3755 ( 
.A1(n_3339),
.A2(n_2415),
.B(n_2411),
.Y(n_3755)
);

HB1xp67_ASAP7_75t_L g3756 ( 
.A(n_3412),
.Y(n_3756)
);

AOI21x1_ASAP7_75t_L g3757 ( 
.A1(n_3512),
.A2(n_386),
.B(n_385),
.Y(n_3757)
);

HB1xp67_ASAP7_75t_L g3758 ( 
.A(n_3413),
.Y(n_3758)
);

AOI211xp5_ASAP7_75t_L g3759 ( 
.A1(n_3280),
.A2(n_2426),
.B(n_2430),
.C(n_2425),
.Y(n_3759)
);

BUFx3_ASAP7_75t_L g3760 ( 
.A(n_3476),
.Y(n_3760)
);

NAND2xp5_ASAP7_75t_SL g3761 ( 
.A(n_3507),
.B(n_2431),
.Y(n_3761)
);

AND2x2_ASAP7_75t_L g3762 ( 
.A(n_3318),
.B(n_2433),
.Y(n_3762)
);

INVx1_ASAP7_75t_L g3763 ( 
.A(n_3543),
.Y(n_3763)
);

NOR2xp33_ASAP7_75t_L g3764 ( 
.A(n_3615),
.B(n_3324),
.Y(n_3764)
);

NAND2xp5_ASAP7_75t_SL g3765 ( 
.A(n_3593),
.B(n_3436),
.Y(n_3765)
);

NOR2xp33_ASAP7_75t_L g3766 ( 
.A(n_3558),
.B(n_3487),
.Y(n_3766)
);

NOR2xp33_ASAP7_75t_L g3767 ( 
.A(n_3564),
.B(n_3396),
.Y(n_3767)
);

NAND2xp5_ASAP7_75t_SL g3768 ( 
.A(n_3607),
.B(n_3492),
.Y(n_3768)
);

BUFx6f_ASAP7_75t_L g3769 ( 
.A(n_3556),
.Y(n_3769)
);

A2O1A1Ixp33_ASAP7_75t_SL g3770 ( 
.A1(n_3651),
.A2(n_3485),
.B(n_3473),
.C(n_3497),
.Y(n_3770)
);

HB1xp67_ASAP7_75t_L g3771 ( 
.A(n_3573),
.Y(n_3771)
);

NAND3xp33_ASAP7_75t_SL g3772 ( 
.A(n_3632),
.B(n_3422),
.C(n_3496),
.Y(n_3772)
);

BUFx5_ASAP7_75t_L g3773 ( 
.A(n_3605),
.Y(n_3773)
);

OAI22xp5_ASAP7_75t_L g3774 ( 
.A1(n_3645),
.A2(n_3647),
.B1(n_3642),
.B2(n_3613),
.Y(n_3774)
);

BUFx6f_ASAP7_75t_L g3775 ( 
.A(n_3556),
.Y(n_3775)
);

AND2x6_ASAP7_75t_L g3776 ( 
.A(n_3684),
.B(n_3464),
.Y(n_3776)
);

NAND2xp5_ASAP7_75t_L g3777 ( 
.A(n_3589),
.B(n_3372),
.Y(n_3777)
);

INVx2_ASAP7_75t_L g3778 ( 
.A(n_3574),
.Y(n_3778)
);

BUFx6f_ASAP7_75t_L g3779 ( 
.A(n_3556),
.Y(n_3779)
);

NAND2xp5_ASAP7_75t_L g3780 ( 
.A(n_3572),
.B(n_3387),
.Y(n_3780)
);

NAND2xp5_ASAP7_75t_SL g3781 ( 
.A(n_3697),
.B(n_3285),
.Y(n_3781)
);

AND2x2_ASAP7_75t_SL g3782 ( 
.A(n_3603),
.B(n_3511),
.Y(n_3782)
);

OAI22xp5_ASAP7_75t_L g3783 ( 
.A1(n_3617),
.A2(n_3472),
.B1(n_3471),
.B2(n_3493),
.Y(n_3783)
);

INVx4_ASAP7_75t_L g3784 ( 
.A(n_3664),
.Y(n_3784)
);

NAND2xp5_ASAP7_75t_SL g3785 ( 
.A(n_3566),
.B(n_3463),
.Y(n_3785)
);

BUFx6f_ASAP7_75t_L g3786 ( 
.A(n_3576),
.Y(n_3786)
);

AO21x1_ASAP7_75t_L g3787 ( 
.A1(n_3551),
.A2(n_3588),
.B(n_3592),
.Y(n_3787)
);

NAND2xp5_ASAP7_75t_L g3788 ( 
.A(n_3597),
.B(n_3563),
.Y(n_3788)
);

NOR3xp33_ASAP7_75t_SL g3789 ( 
.A(n_3754),
.B(n_3414),
.C(n_3491),
.Y(n_3789)
);

NAND2xp5_ASAP7_75t_L g3790 ( 
.A(n_3570),
.B(n_3513),
.Y(n_3790)
);

BUFx2_ASAP7_75t_L g3791 ( 
.A(n_3606),
.Y(n_3791)
);

NOR2x1_ASAP7_75t_L g3792 ( 
.A(n_3643),
.B(n_3416),
.Y(n_3792)
);

INVx1_ASAP7_75t_L g3793 ( 
.A(n_3631),
.Y(n_3793)
);

NAND2xp5_ASAP7_75t_SL g3794 ( 
.A(n_3759),
.B(n_3383),
.Y(n_3794)
);

NAND2xp5_ASAP7_75t_SL g3795 ( 
.A(n_3751),
.B(n_3467),
.Y(n_3795)
);

O2A1O1Ixp33_ASAP7_75t_SL g3796 ( 
.A1(n_3624),
.A2(n_3549),
.B(n_3442),
.C(n_3431),
.Y(n_3796)
);

BUFx6f_ASAP7_75t_L g3797 ( 
.A(n_3576),
.Y(n_3797)
);

NAND2xp5_ASAP7_75t_SL g3798 ( 
.A(n_3726),
.B(n_3466),
.Y(n_3798)
);

BUFx2_ASAP7_75t_L g3799 ( 
.A(n_3667),
.Y(n_3799)
);

AND2x2_ASAP7_75t_L g3800 ( 
.A(n_3561),
.B(n_3567),
.Y(n_3800)
);

NOR2xp33_ASAP7_75t_L g3801 ( 
.A(n_3577),
.B(n_3500),
.Y(n_3801)
);

CKINVDCx8_ASAP7_75t_R g3802 ( 
.A(n_3609),
.Y(n_3802)
);

OAI21xp5_ASAP7_75t_L g3803 ( 
.A1(n_3750),
.A2(n_3460),
.B(n_3483),
.Y(n_3803)
);

O2A1O1Ixp5_ASAP7_75t_L g3804 ( 
.A1(n_3621),
.A2(n_3475),
.B(n_3479),
.C(n_3386),
.Y(n_3804)
);

INVx2_ASAP7_75t_SL g3805 ( 
.A(n_3742),
.Y(n_3805)
);

NAND2xp5_ASAP7_75t_L g3806 ( 
.A(n_3580),
.B(n_3582),
.Y(n_3806)
);

A2O1A1Ixp33_ASAP7_75t_L g3807 ( 
.A1(n_3660),
.A2(n_3678),
.B(n_3594),
.C(n_3584),
.Y(n_3807)
);

AND2x2_ASAP7_75t_L g3808 ( 
.A(n_3630),
.B(n_3319),
.Y(n_3808)
);

A2O1A1Ixp33_ASAP7_75t_L g3809 ( 
.A1(n_3727),
.A2(n_2443),
.B(n_2445),
.C(n_2441),
.Y(n_3809)
);

NAND2xp5_ASAP7_75t_SL g3810 ( 
.A(n_3625),
.B(n_2446),
.Y(n_3810)
);

AOI22xp33_ASAP7_75t_L g3811 ( 
.A1(n_3699),
.A2(n_3409),
.B1(n_3416),
.B2(n_2447),
.Y(n_3811)
);

INVx1_ASAP7_75t_L g3812 ( 
.A(n_3663),
.Y(n_3812)
);

INVx1_ASAP7_75t_L g3813 ( 
.A(n_3620),
.Y(n_3813)
);

INVx2_ASAP7_75t_L g3814 ( 
.A(n_3585),
.Y(n_3814)
);

NAND2xp5_ASAP7_75t_L g3815 ( 
.A(n_3560),
.B(n_2451),
.Y(n_3815)
);

INVx6_ASAP7_75t_L g3816 ( 
.A(n_3742),
.Y(n_3816)
);

INVx1_ASAP7_75t_L g3817 ( 
.A(n_3565),
.Y(n_3817)
);

INVx1_ASAP7_75t_L g3818 ( 
.A(n_3583),
.Y(n_3818)
);

A2O1A1Ixp33_ASAP7_75t_L g3819 ( 
.A1(n_3711),
.A2(n_2459),
.B(n_2460),
.C(n_2457),
.Y(n_3819)
);

OAI22xp5_ASAP7_75t_L g3820 ( 
.A1(n_3686),
.A2(n_2468),
.B1(n_2466),
.B2(n_387),
.Y(n_3820)
);

CKINVDCx8_ASAP7_75t_R g3821 ( 
.A(n_3695),
.Y(n_3821)
);

OAI22xp5_ASAP7_75t_SL g3822 ( 
.A1(n_3661),
.A2(n_2),
.B1(n_0),
.B2(n_1),
.Y(n_3822)
);

AOI21xp5_ASAP7_75t_L g3823 ( 
.A1(n_3646),
.A2(n_389),
.B(n_388),
.Y(n_3823)
);

NAND2xp5_ASAP7_75t_L g3824 ( 
.A(n_3723),
.B(n_1),
.Y(n_3824)
);

NOR2xp33_ASAP7_75t_L g3825 ( 
.A(n_3648),
.B(n_390),
.Y(n_3825)
);

INVx1_ASAP7_75t_L g3826 ( 
.A(n_3585),
.Y(n_3826)
);

BUFx2_ASAP7_75t_L g3827 ( 
.A(n_3557),
.Y(n_3827)
);

A2O1A1Ixp33_ASAP7_75t_L g3828 ( 
.A1(n_3740),
.A2(n_4),
.B(n_1),
.C(n_3),
.Y(n_3828)
);

NAND2xp5_ASAP7_75t_L g3829 ( 
.A(n_3650),
.B(n_3),
.Y(n_3829)
);

OR2x6_ASAP7_75t_SL g3830 ( 
.A(n_3732),
.B(n_5),
.Y(n_3830)
);

CKINVDCx20_ASAP7_75t_R g3831 ( 
.A(n_3629),
.Y(n_3831)
);

A2O1A1Ixp33_ASAP7_75t_L g3832 ( 
.A1(n_3559),
.A2(n_7),
.B(n_5),
.C(n_6),
.Y(n_3832)
);

AOI22xp5_ASAP7_75t_L g3833 ( 
.A1(n_3679),
.A2(n_392),
.B1(n_393),
.B2(n_391),
.Y(n_3833)
);

AOI21xp5_ASAP7_75t_L g3834 ( 
.A1(n_3653),
.A2(n_392),
.B(n_391),
.Y(n_3834)
);

INVxp67_ASAP7_75t_L g3835 ( 
.A(n_3649),
.Y(n_3835)
);

AOI21xp5_ASAP7_75t_L g3836 ( 
.A1(n_3654),
.A2(n_394),
.B(n_393),
.Y(n_3836)
);

NAND2xp5_ASAP7_75t_L g3837 ( 
.A(n_3677),
.B(n_6),
.Y(n_3837)
);

AND3x2_ASAP7_75t_L g3838 ( 
.A(n_3636),
.B(n_7),
.C(n_8),
.Y(n_3838)
);

NAND2xp5_ASAP7_75t_L g3839 ( 
.A(n_3694),
.B(n_9),
.Y(n_3839)
);

INVx2_ASAP7_75t_L g3840 ( 
.A(n_3598),
.Y(n_3840)
);

O2A1O1Ixp5_ASAP7_75t_L g3841 ( 
.A1(n_3552),
.A2(n_3655),
.B(n_3675),
.C(n_3673),
.Y(n_3841)
);

INVx2_ASAP7_75t_L g3842 ( 
.A(n_3626),
.Y(n_3842)
);

NAND2x1p5_ASAP7_75t_L g3843 ( 
.A(n_3742),
.B(n_395),
.Y(n_3843)
);

AOI221xp5_ASAP7_75t_L g3844 ( 
.A1(n_3691),
.A2(n_11),
.B1(n_9),
.B2(n_10),
.C(n_12),
.Y(n_3844)
);

CKINVDCx5p33_ASAP7_75t_R g3845 ( 
.A(n_3587),
.Y(n_3845)
);

INVx2_ASAP7_75t_L g3846 ( 
.A(n_3670),
.Y(n_3846)
);

NAND2xp5_ASAP7_75t_SL g3847 ( 
.A(n_3612),
.B(n_396),
.Y(n_3847)
);

A2O1A1Ixp33_ASAP7_75t_L g3848 ( 
.A1(n_3569),
.A2(n_11),
.B(n_9),
.C(n_10),
.Y(n_3848)
);

AOI22xp5_ASAP7_75t_L g3849 ( 
.A1(n_3717),
.A2(n_397),
.B1(n_398),
.B2(n_396),
.Y(n_3849)
);

AND2x2_ASAP7_75t_L g3850 ( 
.A(n_3762),
.B(n_397),
.Y(n_3850)
);

NAND2xp5_ASAP7_75t_L g3851 ( 
.A(n_3700),
.B(n_12),
.Y(n_3851)
);

AOI22xp5_ASAP7_75t_L g3852 ( 
.A1(n_3680),
.A2(n_399),
.B1(n_401),
.B2(n_398),
.Y(n_3852)
);

NAND2xp5_ASAP7_75t_L g3853 ( 
.A(n_3704),
.B(n_12),
.Y(n_3853)
);

INVx2_ASAP7_75t_L g3854 ( 
.A(n_3683),
.Y(n_3854)
);

BUFx6f_ASAP7_75t_L g3855 ( 
.A(n_3639),
.Y(n_3855)
);

NOR2xp33_ASAP7_75t_L g3856 ( 
.A(n_3553),
.B(n_403),
.Y(n_3856)
);

BUFx4f_ASAP7_75t_SL g3857 ( 
.A(n_3639),
.Y(n_3857)
);

BUFx8_ASAP7_75t_SL g3858 ( 
.A(n_3672),
.Y(n_3858)
);

NAND2xp5_ASAP7_75t_SL g3859 ( 
.A(n_3725),
.B(n_404),
.Y(n_3859)
);

INVx3_ASAP7_75t_L g3860 ( 
.A(n_3639),
.Y(n_3860)
);

NOR2xp33_ASAP7_75t_L g3861 ( 
.A(n_3676),
.B(n_405),
.Y(n_3861)
);

AOI21xp5_ASAP7_75t_L g3862 ( 
.A1(n_3724),
.A2(n_3731),
.B(n_3599),
.Y(n_3862)
);

AOI21xp5_ASAP7_75t_L g3863 ( 
.A1(n_3749),
.A2(n_407),
.B(n_406),
.Y(n_3863)
);

AND2x4_ASAP7_75t_L g3864 ( 
.A(n_3760),
.B(n_406),
.Y(n_3864)
);

NOR2xp33_ASAP7_75t_L g3865 ( 
.A(n_3668),
.B(n_407),
.Y(n_3865)
);

NAND2xp5_ASAP7_75t_SL g3866 ( 
.A(n_3715),
.B(n_408),
.Y(n_3866)
);

OAI22x1_ASAP7_75t_L g3867 ( 
.A1(n_3684),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.Y(n_3867)
);

O2A1O1Ixp33_ASAP7_75t_L g3868 ( 
.A1(n_3635),
.A2(n_412),
.B(n_414),
.C(n_411),
.Y(n_3868)
);

BUFx6f_ASAP7_75t_L g3869 ( 
.A(n_3715),
.Y(n_3869)
);

BUFx3_ASAP7_75t_L g3870 ( 
.A(n_3652),
.Y(n_3870)
);

NOR2xp33_ASAP7_75t_L g3871 ( 
.A(n_3735),
.B(n_412),
.Y(n_3871)
);

NOR2xp33_ASAP7_75t_SL g3872 ( 
.A(n_3707),
.B(n_13),
.Y(n_3872)
);

NAND2xp5_ASAP7_75t_L g3873 ( 
.A(n_3638),
.B(n_15),
.Y(n_3873)
);

AOI22xp5_ASAP7_75t_L g3874 ( 
.A1(n_3733),
.A2(n_3716),
.B1(n_3714),
.B2(n_3628),
.Y(n_3874)
);

O2A1O1Ixp33_ASAP7_75t_L g3875 ( 
.A1(n_3682),
.A2(n_416),
.B(n_417),
.C(n_415),
.Y(n_3875)
);

OAI21xp33_ASAP7_75t_L g3876 ( 
.A1(n_3633),
.A2(n_16),
.B(n_17),
.Y(n_3876)
);

INVx2_ASAP7_75t_L g3877 ( 
.A(n_3671),
.Y(n_3877)
);

AND2x2_ASAP7_75t_L g3878 ( 
.A(n_3590),
.B(n_417),
.Y(n_3878)
);

NAND2xp5_ASAP7_75t_L g3879 ( 
.A(n_3638),
.B(n_16),
.Y(n_3879)
);

INVx1_ASAP7_75t_L g3880 ( 
.A(n_3720),
.Y(n_3880)
);

AOI22xp5_ASAP7_75t_L g3881 ( 
.A1(n_3665),
.A2(n_420),
.B1(n_421),
.B2(n_419),
.Y(n_3881)
);

HB1xp67_ASAP7_75t_L g3882 ( 
.A(n_3756),
.Y(n_3882)
);

INVx1_ASAP7_75t_SL g3883 ( 
.A(n_3758),
.Y(n_3883)
);

NOR2xp33_ASAP7_75t_R g3884 ( 
.A(n_3712),
.B(n_422),
.Y(n_3884)
);

BUFx6f_ASAP7_75t_L g3885 ( 
.A(n_3712),
.Y(n_3885)
);

NOR2xp33_ASAP7_75t_L g3886 ( 
.A(n_3736),
.B(n_424),
.Y(n_3886)
);

NAND2xp5_ASAP7_75t_L g3887 ( 
.A(n_3618),
.B(n_17),
.Y(n_3887)
);

O2A1O1Ixp33_ASAP7_75t_L g3888 ( 
.A1(n_3568),
.A2(n_426),
.B(n_427),
.C(n_425),
.Y(n_3888)
);

INVx4_ASAP7_75t_L g3889 ( 
.A(n_3746),
.Y(n_3889)
);

INVx1_ASAP7_75t_SL g3890 ( 
.A(n_3590),
.Y(n_3890)
);

AO21x1_ASAP7_75t_L g3891 ( 
.A1(n_3550),
.A2(n_430),
.B(n_429),
.Y(n_3891)
);

A2O1A1Ixp33_ASAP7_75t_L g3892 ( 
.A1(n_3696),
.A2(n_20),
.B(n_18),
.C(n_19),
.Y(n_3892)
);

AND2x2_ASAP7_75t_L g3893 ( 
.A(n_3681),
.B(n_431),
.Y(n_3893)
);

BUFx2_ASAP7_75t_SL g3894 ( 
.A(n_3746),
.Y(n_3894)
);

NOR2x1_ASAP7_75t_L g3895 ( 
.A(n_3562),
.B(n_432),
.Y(n_3895)
);

O2A1O1Ixp33_ASAP7_75t_L g3896 ( 
.A1(n_3702),
.A2(n_433),
.B(n_434),
.C(n_432),
.Y(n_3896)
);

AOI21xp5_ASAP7_75t_L g3897 ( 
.A1(n_3708),
.A2(n_3575),
.B(n_3571),
.Y(n_3897)
);

BUFx6f_ASAP7_75t_L g3898 ( 
.A(n_3722),
.Y(n_3898)
);

AO32x1_ASAP7_75t_L g3899 ( 
.A1(n_3710),
.A2(n_24),
.A3(n_21),
.B1(n_23),
.B2(n_25),
.Y(n_3899)
);

NAND2xp5_ASAP7_75t_L g3900 ( 
.A(n_3619),
.B(n_21),
.Y(n_3900)
);

AOI21xp5_ASAP7_75t_L g3901 ( 
.A1(n_3581),
.A2(n_436),
.B(n_435),
.Y(n_3901)
);

AOI21xp5_ASAP7_75t_L g3902 ( 
.A1(n_3586),
.A2(n_436),
.B(n_435),
.Y(n_3902)
);

NOR2xp67_ASAP7_75t_SL g3903 ( 
.A(n_3761),
.B(n_23),
.Y(n_3903)
);

NAND2xp5_ASAP7_75t_L g3904 ( 
.A(n_3622),
.B(n_24),
.Y(n_3904)
);

INVx1_ASAP7_75t_L g3905 ( 
.A(n_3591),
.Y(n_3905)
);

AOI22xp33_ASAP7_75t_L g3906 ( 
.A1(n_3616),
.A2(n_28),
.B1(n_26),
.B2(n_27),
.Y(n_3906)
);

INVx1_ASAP7_75t_L g3907 ( 
.A(n_3604),
.Y(n_3907)
);

CKINVDCx5p33_ASAP7_75t_R g3908 ( 
.A(n_3743),
.Y(n_3908)
);

INVx1_ASAP7_75t_SL g3909 ( 
.A(n_3763),
.Y(n_3909)
);

O2A1O1Ixp33_ASAP7_75t_SL g3910 ( 
.A1(n_3657),
.A2(n_28),
.B(n_26),
.C(n_27),
.Y(n_3910)
);

BUFx12f_ASAP7_75t_L g3911 ( 
.A(n_3709),
.Y(n_3911)
);

INVx3_ASAP7_75t_L g3912 ( 
.A(n_3741),
.Y(n_3912)
);

INVx2_ASAP7_75t_L g3913 ( 
.A(n_3578),
.Y(n_3913)
);

AOI21xp5_ASAP7_75t_L g3914 ( 
.A1(n_3600),
.A2(n_438),
.B(n_437),
.Y(n_3914)
);

NAND2xp5_ASAP7_75t_L g3915 ( 
.A(n_3659),
.B(n_29),
.Y(n_3915)
);

CKINVDCx11_ASAP7_75t_R g3916 ( 
.A(n_3718),
.Y(n_3916)
);

OAI21x1_ASAP7_75t_L g3917 ( 
.A1(n_3748),
.A2(n_29),
.B(n_30),
.Y(n_3917)
);

INVx1_ASAP7_75t_L g3918 ( 
.A(n_3757),
.Y(n_3918)
);

HB1xp67_ASAP7_75t_L g3919 ( 
.A(n_3687),
.Y(n_3919)
);

AOI21xp5_ASAP7_75t_L g3920 ( 
.A1(n_3611),
.A2(n_439),
.B(n_437),
.Y(n_3920)
);

NAND2xp5_ASAP7_75t_L g3921 ( 
.A(n_3610),
.B(n_30),
.Y(n_3921)
);

INVx2_ASAP7_75t_L g3922 ( 
.A(n_3690),
.Y(n_3922)
);

BUFx2_ASAP7_75t_L g3923 ( 
.A(n_3601),
.Y(n_3923)
);

NAND2xp5_ASAP7_75t_L g3924 ( 
.A(n_3596),
.B(n_31),
.Y(n_3924)
);

OAI21xp5_ASAP7_75t_L g3925 ( 
.A1(n_3685),
.A2(n_31),
.B(n_32),
.Y(n_3925)
);

INVx2_ASAP7_75t_L g3926 ( 
.A(n_3693),
.Y(n_3926)
);

NAND2xp5_ASAP7_75t_L g3927 ( 
.A(n_3555),
.B(n_31),
.Y(n_3927)
);

BUFx2_ASAP7_75t_L g3928 ( 
.A(n_3739),
.Y(n_3928)
);

NAND2xp5_ASAP7_75t_SL g3929 ( 
.A(n_3656),
.B(n_442),
.Y(n_3929)
);

AOI22xp33_ASAP7_75t_L g3930 ( 
.A1(n_3738),
.A2(n_3729),
.B1(n_3658),
.B2(n_3737),
.Y(n_3930)
);

NAND2xp5_ASAP7_75t_L g3931 ( 
.A(n_3614),
.B(n_33),
.Y(n_3931)
);

AND2x2_ASAP7_75t_L g3932 ( 
.A(n_3637),
.B(n_445),
.Y(n_3932)
);

O2A1O1Ixp33_ASAP7_75t_L g3933 ( 
.A1(n_3634),
.A2(n_448),
.B(n_449),
.C(n_446),
.Y(n_3933)
);

AND2x4_ASAP7_75t_L g3934 ( 
.A(n_3692),
.B(n_448),
.Y(n_3934)
);

NAND2xp5_ASAP7_75t_SL g3935 ( 
.A(n_3713),
.B(n_450),
.Y(n_3935)
);

NAND3xp33_ASAP7_75t_SL g3936 ( 
.A(n_3698),
.B(n_33),
.C(n_34),
.Y(n_3936)
);

NOR2xp33_ASAP7_75t_L g3937 ( 
.A(n_3728),
.B(n_450),
.Y(n_3937)
);

INVx3_ASAP7_75t_L g3938 ( 
.A(n_3666),
.Y(n_3938)
);

OAI22xp5_ASAP7_75t_L g3939 ( 
.A1(n_3641),
.A2(n_454),
.B1(n_455),
.B2(n_453),
.Y(n_3939)
);

BUFx2_ASAP7_75t_L g3940 ( 
.A(n_3719),
.Y(n_3940)
);

NOR2xp33_ASAP7_75t_L g3941 ( 
.A(n_3689),
.B(n_453),
.Y(n_3941)
);

INVx2_ASAP7_75t_L g3942 ( 
.A(n_3745),
.Y(n_3942)
);

BUFx6f_ASAP7_75t_L g3943 ( 
.A(n_3753),
.Y(n_3943)
);

OR2x6_ASAP7_75t_L g3944 ( 
.A(n_3554),
.B(n_455),
.Y(n_3944)
);

INVx1_ASAP7_75t_L g3945 ( 
.A(n_3627),
.Y(n_3945)
);

BUFx2_ASAP7_75t_L g3946 ( 
.A(n_3755),
.Y(n_3946)
);

NAND2xp5_ASAP7_75t_SL g3947 ( 
.A(n_3721),
.B(n_456),
.Y(n_3947)
);

OAI21xp5_ASAP7_75t_L g3948 ( 
.A1(n_3701),
.A2(n_35),
.B(n_36),
.Y(n_3948)
);

INVx4_ASAP7_75t_L g3949 ( 
.A(n_3579),
.Y(n_3949)
);

NOR2xp33_ASAP7_75t_R g3950 ( 
.A(n_3644),
.B(n_457),
.Y(n_3950)
);

INVx3_ASAP7_75t_L g3951 ( 
.A(n_3595),
.Y(n_3951)
);

BUFx6f_ASAP7_75t_L g3952 ( 
.A(n_3640),
.Y(n_3952)
);

INVx3_ASAP7_75t_L g3953 ( 
.A(n_3623),
.Y(n_3953)
);

A2O1A1Ixp33_ASAP7_75t_L g3954 ( 
.A1(n_3703),
.A2(n_37),
.B(n_35),
.C(n_36),
.Y(n_3954)
);

CKINVDCx5p33_ASAP7_75t_R g3955 ( 
.A(n_3744),
.Y(n_3955)
);

NAND3xp33_ASAP7_75t_L g3956 ( 
.A(n_3705),
.B(n_37),
.C(n_38),
.Y(n_3956)
);

O2A1O1Ixp33_ASAP7_75t_L g3957 ( 
.A1(n_3602),
.A2(n_459),
.B(n_460),
.C(n_458),
.Y(n_3957)
);

HB1xp67_ASAP7_75t_L g3958 ( 
.A(n_3752),
.Y(n_3958)
);

AOI21x1_ASAP7_75t_L g3959 ( 
.A1(n_3662),
.A2(n_461),
.B(n_459),
.Y(n_3959)
);

NAND2xp5_ASAP7_75t_L g3960 ( 
.A(n_3706),
.B(n_3608),
.Y(n_3960)
);

NAND2xp5_ASAP7_75t_L g3961 ( 
.A(n_3669),
.B(n_38),
.Y(n_3961)
);

NAND2xp5_ASAP7_75t_L g3962 ( 
.A(n_3674),
.B(n_39),
.Y(n_3962)
);

INVx1_ASAP7_75t_L g3963 ( 
.A(n_3734),
.Y(n_3963)
);

NAND2xp5_ASAP7_75t_L g3964 ( 
.A(n_3747),
.B(n_39),
.Y(n_3964)
);

NAND2xp5_ASAP7_75t_L g3965 ( 
.A(n_3730),
.B(n_39),
.Y(n_3965)
);

INVx4_ASAP7_75t_L g3966 ( 
.A(n_3664),
.Y(n_3966)
);

OAI22xp5_ASAP7_75t_L g3967 ( 
.A1(n_3593),
.A2(n_463),
.B1(n_464),
.B2(n_462),
.Y(n_3967)
);

O2A1O1Ixp33_ASAP7_75t_L g3968 ( 
.A1(n_3593),
.A2(n_466),
.B(n_467),
.C(n_465),
.Y(n_3968)
);

O2A1O1Ixp33_ASAP7_75t_SL g3969 ( 
.A1(n_3593),
.A2(n_42),
.B(n_40),
.C(n_41),
.Y(n_3969)
);

INVx1_ASAP7_75t_L g3970 ( 
.A(n_3688),
.Y(n_3970)
);

AOI21xp5_ASAP7_75t_L g3971 ( 
.A1(n_3593),
.A2(n_468),
.B(n_467),
.Y(n_3971)
);

INVxp67_ASAP7_75t_L g3972 ( 
.A(n_3573),
.Y(n_3972)
);

NAND2xp5_ASAP7_75t_L g3973 ( 
.A(n_3615),
.B(n_41),
.Y(n_3973)
);

NAND2xp5_ASAP7_75t_SL g3974 ( 
.A(n_3593),
.B(n_468),
.Y(n_3974)
);

AOI21xp5_ASAP7_75t_L g3975 ( 
.A1(n_3593),
.A2(n_470),
.B(n_469),
.Y(n_3975)
);

AND2x4_ASAP7_75t_L g3976 ( 
.A(n_3667),
.B(n_471),
.Y(n_3976)
);

NAND2xp5_ASAP7_75t_L g3977 ( 
.A(n_3774),
.B(n_3813),
.Y(n_3977)
);

NAND2xp5_ASAP7_75t_L g3978 ( 
.A(n_3764),
.B(n_43),
.Y(n_3978)
);

INVxp67_ASAP7_75t_L g3979 ( 
.A(n_3771),
.Y(n_3979)
);

AOI21x1_ASAP7_75t_SL g3980 ( 
.A1(n_3893),
.A2(n_43),
.B(n_44),
.Y(n_3980)
);

NAND2xp5_ASAP7_75t_L g3981 ( 
.A(n_3788),
.B(n_43),
.Y(n_3981)
);

A2O1A1Ixp33_ASAP7_75t_L g3982 ( 
.A1(n_3766),
.A2(n_46),
.B(n_44),
.C(n_45),
.Y(n_3982)
);

BUFx2_ASAP7_75t_L g3983 ( 
.A(n_3791),
.Y(n_3983)
);

OA21x2_ASAP7_75t_L g3984 ( 
.A1(n_3877),
.A2(n_44),
.B(n_45),
.Y(n_3984)
);

OAI21x1_ASAP7_75t_L g3985 ( 
.A1(n_3913),
.A2(n_45),
.B(n_47),
.Y(n_3985)
);

NAND2xp5_ASAP7_75t_L g3986 ( 
.A(n_3806),
.B(n_47),
.Y(n_3986)
);

AO31x2_ASAP7_75t_L g3987 ( 
.A1(n_3787),
.A2(n_3940),
.A3(n_3918),
.B(n_3891),
.Y(n_3987)
);

HB1xp67_ASAP7_75t_L g3988 ( 
.A(n_3972),
.Y(n_3988)
);

NOR2xp33_ASAP7_75t_L g3989 ( 
.A(n_3767),
.B(n_472),
.Y(n_3989)
);

INVxp67_ASAP7_75t_SL g3990 ( 
.A(n_3882),
.Y(n_3990)
);

CKINVDCx20_ASAP7_75t_R g3991 ( 
.A(n_3831),
.Y(n_3991)
);

OAI21x1_ASAP7_75t_L g3992 ( 
.A1(n_3862),
.A2(n_48),
.B(n_49),
.Y(n_3992)
);

OAI21xp5_ASAP7_75t_L g3993 ( 
.A1(n_3777),
.A2(n_49),
.B(n_50),
.Y(n_3993)
);

AO31x2_ASAP7_75t_L g3994 ( 
.A1(n_3807),
.A2(n_52),
.A3(n_49),
.B(n_51),
.Y(n_3994)
);

AND2x2_ASAP7_75t_L g3995 ( 
.A(n_3800),
.B(n_3850),
.Y(n_3995)
);

NOR2xp67_ASAP7_75t_L g3996 ( 
.A(n_3784),
.B(n_51),
.Y(n_3996)
);

NAND3xp33_ASAP7_75t_L g3997 ( 
.A(n_3871),
.B(n_52),
.C(n_53),
.Y(n_3997)
);

NOR2x1_ASAP7_75t_SL g3998 ( 
.A(n_3768),
.B(n_473),
.Y(n_3998)
);

AO31x2_ASAP7_75t_L g3999 ( 
.A1(n_3949),
.A2(n_56),
.A3(n_54),
.B(n_55),
.Y(n_3999)
);

A2O1A1Ixp33_ASAP7_75t_L g4000 ( 
.A1(n_3765),
.A2(n_56),
.B(n_54),
.C(n_55),
.Y(n_4000)
);

OAI21x1_ASAP7_75t_L g4001 ( 
.A1(n_3841),
.A2(n_56),
.B(n_57),
.Y(n_4001)
);

INVx3_ASAP7_75t_L g4002 ( 
.A(n_3858),
.Y(n_4002)
);

OAI21xp5_ASAP7_75t_L g4003 ( 
.A1(n_3780),
.A2(n_57),
.B(n_58),
.Y(n_4003)
);

OAI21x1_ASAP7_75t_L g4004 ( 
.A1(n_3917),
.A2(n_59),
.B(n_60),
.Y(n_4004)
);

CKINVDCx5p33_ASAP7_75t_R g4005 ( 
.A(n_3802),
.Y(n_4005)
);

OAI21xp5_ASAP7_75t_L g4006 ( 
.A1(n_3930),
.A2(n_59),
.B(n_60),
.Y(n_4006)
);

NOR4xp25_ASAP7_75t_L g4007 ( 
.A(n_3968),
.B(n_64),
.C(n_62),
.D(n_63),
.Y(n_4007)
);

AOI21xp5_ASAP7_75t_L g4008 ( 
.A1(n_3960),
.A2(n_475),
.B(n_474),
.Y(n_4008)
);

BUFx3_ASAP7_75t_L g4009 ( 
.A(n_3857),
.Y(n_4009)
);

INVx1_ASAP7_75t_L g4010 ( 
.A(n_3793),
.Y(n_4010)
);

NAND2xp5_ASAP7_75t_L g4011 ( 
.A(n_3922),
.B(n_3926),
.Y(n_4011)
);

NAND3xp33_ASAP7_75t_L g4012 ( 
.A(n_3886),
.B(n_62),
.C(n_63),
.Y(n_4012)
);

INVx4_ASAP7_75t_L g4013 ( 
.A(n_3816),
.Y(n_4013)
);

CKINVDCx5p33_ASAP7_75t_R g4014 ( 
.A(n_3821),
.Y(n_4014)
);

OAI22xp5_ASAP7_75t_L g4015 ( 
.A1(n_3874),
.A2(n_64),
.B1(n_62),
.B2(n_63),
.Y(n_4015)
);

AOI21xp5_ASAP7_75t_L g4016 ( 
.A1(n_3790),
.A2(n_475),
.B(n_474),
.Y(n_4016)
);

OAI21xp5_ASAP7_75t_L g4017 ( 
.A1(n_3803),
.A2(n_3783),
.B(n_3772),
.Y(n_4017)
);

O2A1O1Ixp33_ASAP7_75t_L g4018 ( 
.A1(n_3973),
.A2(n_67),
.B(n_65),
.C(n_66),
.Y(n_4018)
);

BUFx2_ASAP7_75t_R g4019 ( 
.A(n_3845),
.Y(n_4019)
);

OA21x2_ASAP7_75t_L g4020 ( 
.A1(n_3971),
.A2(n_3975),
.B(n_3948),
.Y(n_4020)
);

AO22x2_ASAP7_75t_L g4021 ( 
.A1(n_3967),
.A2(n_67),
.B1(n_65),
.B2(n_66),
.Y(n_4021)
);

OR2x6_ASAP7_75t_L g4022 ( 
.A(n_3799),
.B(n_477),
.Y(n_4022)
);

NAND2xp5_ASAP7_75t_L g4023 ( 
.A(n_3801),
.B(n_65),
.Y(n_4023)
);

OAI21x1_ASAP7_75t_L g4024 ( 
.A1(n_3963),
.A2(n_68),
.B(n_69),
.Y(n_4024)
);

AOI21xp5_ASAP7_75t_L g4025 ( 
.A1(n_3897),
.A2(n_479),
.B(n_478),
.Y(n_4025)
);

AND2x4_ASAP7_75t_L g4026 ( 
.A(n_3805),
.B(n_479),
.Y(n_4026)
);

OR2x6_ASAP7_75t_L g4027 ( 
.A(n_3966),
.B(n_480),
.Y(n_4027)
);

OAI21xp5_ASAP7_75t_L g4028 ( 
.A1(n_3825),
.A2(n_68),
.B(n_69),
.Y(n_4028)
);

AOI22xp5_ASAP7_75t_L g4029 ( 
.A1(n_3955),
.A2(n_3856),
.B1(n_3794),
.B2(n_3861),
.Y(n_4029)
);

AOI21xp5_ASAP7_75t_L g4030 ( 
.A1(n_3945),
.A2(n_481),
.B(n_480),
.Y(n_4030)
);

NOR2xp33_ASAP7_75t_L g4031 ( 
.A(n_3928),
.B(n_481),
.Y(n_4031)
);

NAND2xp5_ASAP7_75t_L g4032 ( 
.A(n_3890),
.B(n_68),
.Y(n_4032)
);

NAND2xp33_ASAP7_75t_R g4033 ( 
.A(n_3789),
.B(n_482),
.Y(n_4033)
);

AND2x2_ASAP7_75t_L g4034 ( 
.A(n_3878),
.B(n_69),
.Y(n_4034)
);

INVx5_ASAP7_75t_L g4035 ( 
.A(n_3769),
.Y(n_4035)
);

OAI21x1_ASAP7_75t_L g4036 ( 
.A1(n_3951),
.A2(n_70),
.B(n_71),
.Y(n_4036)
);

INVx2_ASAP7_75t_SL g4037 ( 
.A(n_3885),
.Y(n_4037)
);

OAI21xp5_ASAP7_75t_L g4038 ( 
.A1(n_3815),
.A2(n_70),
.B(n_71),
.Y(n_4038)
);

INVx1_ASAP7_75t_L g4039 ( 
.A(n_3812),
.Y(n_4039)
);

OAI21xp5_ASAP7_75t_L g4040 ( 
.A1(n_3925),
.A2(n_72),
.B(n_73),
.Y(n_4040)
);

AOI21xp5_ASAP7_75t_L g4041 ( 
.A1(n_3796),
.A2(n_483),
.B(n_482),
.Y(n_4041)
);

AND2x4_ASAP7_75t_L g4042 ( 
.A(n_3827),
.B(n_484),
.Y(n_4042)
);

NAND2xp5_ASAP7_75t_L g4043 ( 
.A(n_3776),
.B(n_74),
.Y(n_4043)
);

OAI22xp5_ASAP7_75t_L g4044 ( 
.A1(n_3942),
.A2(n_76),
.B1(n_74),
.B2(n_75),
.Y(n_4044)
);

NAND2xp5_ASAP7_75t_L g4045 ( 
.A(n_3776),
.B(n_3865),
.Y(n_4045)
);

OAI21x1_ASAP7_75t_L g4046 ( 
.A1(n_3959),
.A2(n_75),
.B(n_76),
.Y(n_4046)
);

BUFx2_ASAP7_75t_SL g4047 ( 
.A(n_3870),
.Y(n_4047)
);

NAND2xp5_ASAP7_75t_L g4048 ( 
.A(n_3824),
.B(n_75),
.Y(n_4048)
);

A2O1A1Ixp33_ASAP7_75t_L g4049 ( 
.A1(n_3937),
.A2(n_79),
.B(n_77),
.C(n_78),
.Y(n_4049)
);

BUFx3_ASAP7_75t_L g4050 ( 
.A(n_3769),
.Y(n_4050)
);

OAI22x1_ASAP7_75t_L g4051 ( 
.A1(n_3833),
.A2(n_80),
.B1(n_78),
.B2(n_79),
.Y(n_4051)
);

INVx1_ASAP7_75t_L g4052 ( 
.A(n_3970),
.Y(n_4052)
);

INVxp67_ASAP7_75t_SL g4053 ( 
.A(n_3912),
.Y(n_4053)
);

AO21x2_ASAP7_75t_L g4054 ( 
.A1(n_3974),
.A2(n_81),
.B(n_82),
.Y(n_4054)
);

NAND2xp5_ASAP7_75t_L g4055 ( 
.A(n_3837),
.B(n_3829),
.Y(n_4055)
);

HB1xp67_ASAP7_75t_L g4056 ( 
.A(n_3883),
.Y(n_4056)
);

NOR2xp33_ASAP7_75t_R g4057 ( 
.A(n_3908),
.B(n_485),
.Y(n_4057)
);

NAND2xp5_ASAP7_75t_L g4058 ( 
.A(n_3839),
.B(n_83),
.Y(n_4058)
);

BUFx3_ASAP7_75t_L g4059 ( 
.A(n_3775),
.Y(n_4059)
);

NAND2xp5_ASAP7_75t_L g4060 ( 
.A(n_3851),
.B(n_84),
.Y(n_4060)
);

CKINVDCx11_ASAP7_75t_R g4061 ( 
.A(n_3830),
.Y(n_4061)
);

OAI22xp5_ASAP7_75t_SL g4062 ( 
.A1(n_3822),
.A2(n_86),
.B1(n_84),
.B2(n_85),
.Y(n_4062)
);

INVx2_ASAP7_75t_L g4063 ( 
.A(n_3840),
.Y(n_4063)
);

INVx1_ASAP7_75t_L g4064 ( 
.A(n_3880),
.Y(n_4064)
);

BUFx4_ASAP7_75t_SL g4065 ( 
.A(n_3923),
.Y(n_4065)
);

NAND3xp33_ASAP7_75t_L g4066 ( 
.A(n_3941),
.B(n_84),
.C(n_85),
.Y(n_4066)
);

OR2x2_ASAP7_75t_L g4067 ( 
.A(n_3853),
.B(n_487),
.Y(n_4067)
);

AOI21xp33_ASAP7_75t_L g4068 ( 
.A1(n_3770),
.A2(n_3958),
.B(n_3965),
.Y(n_4068)
);

AND2x2_ASAP7_75t_L g4069 ( 
.A(n_3932),
.B(n_87),
.Y(n_4069)
);

INVx1_ASAP7_75t_L g4070 ( 
.A(n_3817),
.Y(n_4070)
);

AOI21xp5_ASAP7_75t_L g4071 ( 
.A1(n_3946),
.A2(n_489),
.B(n_488),
.Y(n_4071)
);

AO21x2_ASAP7_75t_L g4072 ( 
.A1(n_3863),
.A2(n_87),
.B(n_88),
.Y(n_4072)
);

INVx1_ASAP7_75t_L g4073 ( 
.A(n_3818),
.Y(n_4073)
);

INVx1_ASAP7_75t_L g4074 ( 
.A(n_3842),
.Y(n_4074)
);

OR2x2_ASAP7_75t_L g4075 ( 
.A(n_3887),
.B(n_490),
.Y(n_4075)
);

AO21x2_ASAP7_75t_L g4076 ( 
.A1(n_3947),
.A2(n_88),
.B(n_89),
.Y(n_4076)
);

OAI21x1_ASAP7_75t_L g4077 ( 
.A1(n_3938),
.A2(n_89),
.B(n_90),
.Y(n_4077)
);

INVx1_ASAP7_75t_L g4078 ( 
.A(n_3846),
.Y(n_4078)
);

OAI21xp33_ASAP7_75t_L g4079 ( 
.A1(n_3950),
.A2(n_3876),
.B(n_3809),
.Y(n_4079)
);

AOI21xp5_ASAP7_75t_L g4080 ( 
.A1(n_3943),
.A2(n_493),
.B(n_492),
.Y(n_4080)
);

BUFx6f_ASAP7_75t_SL g4081 ( 
.A(n_3976),
.Y(n_4081)
);

OAI21xp5_ASAP7_75t_L g4082 ( 
.A1(n_3892),
.A2(n_90),
.B(n_91),
.Y(n_4082)
);

INVx1_ASAP7_75t_L g4083 ( 
.A(n_3854),
.Y(n_4083)
);

AND2x2_ASAP7_75t_L g4084 ( 
.A(n_3808),
.B(n_92),
.Y(n_4084)
);

NAND2xp5_ASAP7_75t_L g4085 ( 
.A(n_3900),
.B(n_3904),
.Y(n_4085)
);

OAI22xp5_ASAP7_75t_L g4086 ( 
.A1(n_3811),
.A2(n_95),
.B1(n_93),
.B2(n_94),
.Y(n_4086)
);

INVx1_ASAP7_75t_L g4087 ( 
.A(n_3826),
.Y(n_4087)
);

INVx5_ASAP7_75t_L g4088 ( 
.A(n_3779),
.Y(n_4088)
);

AO21x2_ASAP7_75t_L g4089 ( 
.A1(n_3964),
.A2(n_95),
.B(n_96),
.Y(n_4089)
);

AOI21x1_ASAP7_75t_L g4090 ( 
.A1(n_3919),
.A2(n_96),
.B(n_97),
.Y(n_4090)
);

O2A1O1Ixp5_ASAP7_75t_L g4091 ( 
.A1(n_3935),
.A2(n_98),
.B(n_96),
.C(n_97),
.Y(n_4091)
);

INVx1_ASAP7_75t_SL g4092 ( 
.A(n_3909),
.Y(n_4092)
);

INVx2_ASAP7_75t_L g4093 ( 
.A(n_3778),
.Y(n_4093)
);

NOR2xp67_ASAP7_75t_SL g4094 ( 
.A(n_3911),
.B(n_98),
.Y(n_4094)
);

OAI21x1_ASAP7_75t_L g4095 ( 
.A1(n_3953),
.A2(n_98),
.B(n_100),
.Y(n_4095)
);

AND2x2_ASAP7_75t_L g4096 ( 
.A(n_3898),
.B(n_100),
.Y(n_4096)
);

NAND2xp5_ASAP7_75t_L g4097 ( 
.A(n_3915),
.B(n_101),
.Y(n_4097)
);

AND2x2_ASAP7_75t_L g4098 ( 
.A(n_3898),
.B(n_102),
.Y(n_4098)
);

O2A1O1Ixp33_ASAP7_75t_L g4099 ( 
.A1(n_3929),
.A2(n_104),
.B(n_102),
.C(n_103),
.Y(n_4099)
);

AOI21xp5_ASAP7_75t_L g4100 ( 
.A1(n_3782),
.A2(n_497),
.B(n_495),
.Y(n_4100)
);

A2O1A1Ixp33_ASAP7_75t_L g4101 ( 
.A1(n_3875),
.A2(n_106),
.B(n_104),
.C(n_105),
.Y(n_4101)
);

AOI211x1_ASAP7_75t_L g4102 ( 
.A1(n_3936),
.A2(n_107),
.B(n_105),
.C(n_106),
.Y(n_4102)
);

AND2x2_ASAP7_75t_L g4103 ( 
.A(n_3934),
.B(n_106),
.Y(n_4103)
);

AO31x2_ASAP7_75t_L g4104 ( 
.A1(n_3828),
.A2(n_109),
.A3(n_107),
.B(n_108),
.Y(n_4104)
);

AO31x2_ASAP7_75t_L g4105 ( 
.A1(n_3954),
.A2(n_112),
.A3(n_110),
.B(n_111),
.Y(n_4105)
);

NOR2x1_ASAP7_75t_L g4106 ( 
.A(n_3889),
.B(n_495),
.Y(n_4106)
);

NOR2xp33_ASAP7_75t_SL g4107 ( 
.A(n_3792),
.B(n_110),
.Y(n_4107)
);

AOI21xp5_ASAP7_75t_L g4108 ( 
.A1(n_3795),
.A2(n_498),
.B(n_497),
.Y(n_4108)
);

AOI21xp5_ASAP7_75t_L g4109 ( 
.A1(n_3969),
.A2(n_501),
.B(n_500),
.Y(n_4109)
);

AO31x2_ASAP7_75t_L g4110 ( 
.A1(n_3832),
.A2(n_113),
.A3(n_111),
.B(n_112),
.Y(n_4110)
);

HB1xp67_ASAP7_75t_L g4111 ( 
.A(n_3835),
.Y(n_4111)
);

NAND2xp5_ASAP7_75t_L g4112 ( 
.A(n_3873),
.B(n_112),
.Y(n_4112)
);

AO31x2_ASAP7_75t_L g4113 ( 
.A1(n_3848),
.A2(n_116),
.A3(n_114),
.B(n_115),
.Y(n_4113)
);

OAI21x1_ASAP7_75t_L g4114 ( 
.A1(n_3823),
.A2(n_114),
.B(n_115),
.Y(n_4114)
);

NOR2xp33_ASAP7_75t_L g4115 ( 
.A(n_3916),
.B(n_501),
.Y(n_4115)
);

NAND2xp5_ASAP7_75t_L g4116 ( 
.A(n_3879),
.B(n_3814),
.Y(n_4116)
);

INVx3_ASAP7_75t_L g4117 ( 
.A(n_3779),
.Y(n_4117)
);

AOI221x1_ASAP7_75t_L g4118 ( 
.A1(n_3820),
.A2(n_504),
.B1(n_505),
.B2(n_503),
.C(n_502),
.Y(n_4118)
);

OAI21xp5_ASAP7_75t_L g4119 ( 
.A1(n_3956),
.A2(n_116),
.B(n_117),
.Y(n_4119)
);

BUFx2_ASAP7_75t_L g4120 ( 
.A(n_3860),
.Y(n_4120)
);

INVx1_ASAP7_75t_L g4121 ( 
.A(n_3905),
.Y(n_4121)
);

NOR2xp33_ASAP7_75t_L g4122 ( 
.A(n_3810),
.B(n_502),
.Y(n_4122)
);

OAI21xp5_ASAP7_75t_L g4123 ( 
.A1(n_3819),
.A2(n_117),
.B(n_118),
.Y(n_4123)
);

OAI21x1_ASAP7_75t_L g4124 ( 
.A1(n_3834),
.A2(n_118),
.B(n_119),
.Y(n_4124)
);

OA21x2_ASAP7_75t_L g4125 ( 
.A1(n_3961),
.A2(n_119),
.B(n_120),
.Y(n_4125)
);

NOR4xp25_ASAP7_75t_L g4126 ( 
.A(n_3933),
.B(n_3957),
.C(n_3868),
.D(n_3888),
.Y(n_4126)
);

OAI21x1_ASAP7_75t_L g4127 ( 
.A1(n_3836),
.A2(n_119),
.B(n_120),
.Y(n_4127)
);

NAND3x1_ASAP7_75t_L g4128 ( 
.A(n_3881),
.B(n_121),
.C(n_122),
.Y(n_4128)
);

INVx1_ASAP7_75t_L g4129 ( 
.A(n_3907),
.Y(n_4129)
);

AOI21xp5_ASAP7_75t_L g4130 ( 
.A1(n_3896),
.A2(n_507),
.B(n_506),
.Y(n_4130)
);

INVx4_ASAP7_75t_L g4131 ( 
.A(n_3786),
.Y(n_4131)
);

NOR2xp33_ASAP7_75t_R g4132 ( 
.A(n_3786),
.B(n_508),
.Y(n_4132)
);

NAND2xp5_ASAP7_75t_L g4133 ( 
.A(n_3798),
.B(n_121),
.Y(n_4133)
);

NAND2xp5_ASAP7_75t_L g4134 ( 
.A(n_3952),
.B(n_122),
.Y(n_4134)
);

NAND2xp5_ASAP7_75t_L g4135 ( 
.A(n_3785),
.B(n_124),
.Y(n_4135)
);

OAI21xp5_ASAP7_75t_L g4136 ( 
.A1(n_3804),
.A2(n_124),
.B(n_125),
.Y(n_4136)
);

INVx2_ASAP7_75t_SL g4137 ( 
.A(n_3797),
.Y(n_4137)
);

O2A1O1Ixp5_ASAP7_75t_L g4138 ( 
.A1(n_3903),
.A2(n_128),
.B(n_125),
.C(n_126),
.Y(n_4138)
);

A2O1A1Ixp33_ASAP7_75t_L g4139 ( 
.A1(n_3901),
.A2(n_130),
.B(n_128),
.C(n_129),
.Y(n_4139)
);

INVx1_ASAP7_75t_L g4140 ( 
.A(n_3773),
.Y(n_4140)
);

OAI21xp5_ASAP7_75t_L g4141 ( 
.A1(n_3902),
.A2(n_129),
.B(n_130),
.Y(n_4141)
);

BUFx8_ASAP7_75t_L g4142 ( 
.A(n_4081),
.Y(n_4142)
);

OAI211xp5_ASAP7_75t_L g4143 ( 
.A1(n_4028),
.A2(n_3844),
.B(n_3849),
.C(n_3852),
.Y(n_4143)
);

AOI21xp5_ASAP7_75t_L g4144 ( 
.A1(n_4017),
.A2(n_3899),
.B(n_3927),
.Y(n_4144)
);

OA21x2_ASAP7_75t_L g4145 ( 
.A1(n_4068),
.A2(n_3920),
.B(n_3914),
.Y(n_4145)
);

OAI21x1_ASAP7_75t_L g4146 ( 
.A1(n_4001),
.A2(n_3895),
.B(n_3962),
.Y(n_4146)
);

INVx2_ASAP7_75t_L g4147 ( 
.A(n_4063),
.Y(n_4147)
);

A2O1A1Ixp33_ASAP7_75t_L g4148 ( 
.A1(n_4029),
.A2(n_3924),
.B(n_3921),
.C(n_3931),
.Y(n_4148)
);

INVx1_ASAP7_75t_L g4149 ( 
.A(n_4010),
.Y(n_4149)
);

OAI22xp5_ASAP7_75t_L g4150 ( 
.A1(n_3989),
.A2(n_3906),
.B1(n_3944),
.B2(n_3781),
.Y(n_4150)
);

INVx2_ASAP7_75t_L g4151 ( 
.A(n_4093),
.Y(n_4151)
);

INVx1_ASAP7_75t_L g4152 ( 
.A(n_4039),
.Y(n_4152)
);

AND2x2_ASAP7_75t_L g4153 ( 
.A(n_3995),
.B(n_3867),
.Y(n_4153)
);

AND2x2_ASAP7_75t_L g4154 ( 
.A(n_4069),
.B(n_3843),
.Y(n_4154)
);

OA21x2_ASAP7_75t_L g4155 ( 
.A1(n_4041),
.A2(n_3866),
.B(n_3859),
.Y(n_4155)
);

OAI22xp5_ASAP7_75t_L g4156 ( 
.A1(n_4045),
.A2(n_3894),
.B1(n_3847),
.B2(n_3939),
.Y(n_4156)
);

CKINVDCx20_ASAP7_75t_R g4157 ( 
.A(n_3991),
.Y(n_4157)
);

OAI21x1_ASAP7_75t_L g4158 ( 
.A1(n_4036),
.A2(n_3773),
.B(n_3899),
.Y(n_4158)
);

OAI21x1_ASAP7_75t_L g4159 ( 
.A1(n_4046),
.A2(n_3773),
.B(n_3910),
.Y(n_4159)
);

INVx1_ASAP7_75t_L g4160 ( 
.A(n_4052),
.Y(n_4160)
);

AO21x2_ASAP7_75t_L g4161 ( 
.A1(n_4040),
.A2(n_3884),
.B(n_3864),
.Y(n_4161)
);

OAI21x1_ASAP7_75t_L g4162 ( 
.A1(n_3992),
.A2(n_3838),
.B(n_3855),
.Y(n_4162)
);

AO32x2_ASAP7_75t_L g4163 ( 
.A1(n_4062),
.A2(n_4015),
.A3(n_4044),
.B1(n_4086),
.B2(n_3980),
.Y(n_4163)
);

INVx1_ASAP7_75t_L g4164 ( 
.A(n_4064),
.Y(n_4164)
);

OAI21x1_ASAP7_75t_L g4165 ( 
.A1(n_4024),
.A2(n_3869),
.B(n_3872),
.Y(n_4165)
);

NAND2xp5_ASAP7_75t_L g4166 ( 
.A(n_4055),
.B(n_4085),
.Y(n_4166)
);

OAI22xp5_ASAP7_75t_L g4167 ( 
.A1(n_3978),
.A2(n_133),
.B1(n_131),
.B2(n_132),
.Y(n_4167)
);

CKINVDCx5p33_ASAP7_75t_R g4168 ( 
.A(n_4005),
.Y(n_4168)
);

NAND2xp5_ASAP7_75t_L g4169 ( 
.A(n_4011),
.B(n_509),
.Y(n_4169)
);

INVx2_ASAP7_75t_L g4170 ( 
.A(n_4074),
.Y(n_4170)
);

HB1xp67_ASAP7_75t_L g4171 ( 
.A(n_3990),
.Y(n_4171)
);

AOI22xp33_ASAP7_75t_L g4172 ( 
.A1(n_4079),
.A2(n_137),
.B1(n_135),
.B2(n_136),
.Y(n_4172)
);

OAI22xp5_ASAP7_75t_L g4173 ( 
.A1(n_3977),
.A2(n_139),
.B1(n_135),
.B2(n_138),
.Y(n_4173)
);

AOI22xp33_ASAP7_75t_SL g4174 ( 
.A1(n_4123),
.A2(n_140),
.B1(n_138),
.B2(n_139),
.Y(n_4174)
);

NOR2x1_ASAP7_75t_SL g4175 ( 
.A(n_4140),
.B(n_4072),
.Y(n_4175)
);

INVx1_ASAP7_75t_L g4176 ( 
.A(n_4070),
.Y(n_4176)
);

NAND3xp33_ASAP7_75t_SL g4177 ( 
.A(n_4107),
.B(n_140),
.C(n_141),
.Y(n_4177)
);

HB1xp67_ASAP7_75t_L g4178 ( 
.A(n_4056),
.Y(n_4178)
);

INVx2_ASAP7_75t_L g4179 ( 
.A(n_4078),
.Y(n_4179)
);

BUFx6f_ASAP7_75t_L g4180 ( 
.A(n_4009),
.Y(n_4180)
);

INVx2_ASAP7_75t_L g4181 ( 
.A(n_4083),
.Y(n_4181)
);

INVx1_ASAP7_75t_L g4182 ( 
.A(n_4073),
.Y(n_4182)
);

INVx1_ASAP7_75t_L g4183 ( 
.A(n_4087),
.Y(n_4183)
);

OAI21x1_ASAP7_75t_L g4184 ( 
.A1(n_4025),
.A2(n_140),
.B(n_141),
.Y(n_4184)
);

NAND2xp5_ASAP7_75t_L g4185 ( 
.A(n_3981),
.B(n_510),
.Y(n_4185)
);

O2A1O1Ixp33_ASAP7_75t_SL g4186 ( 
.A1(n_4049),
.A2(n_143),
.B(n_141),
.C(n_142),
.Y(n_4186)
);

INVx1_ASAP7_75t_L g4187 ( 
.A(n_4121),
.Y(n_4187)
);

OAI21x1_ASAP7_75t_L g4188 ( 
.A1(n_4004),
.A2(n_142),
.B(n_143),
.Y(n_4188)
);

AOI21x1_ASAP7_75t_L g4189 ( 
.A1(n_4130),
.A2(n_142),
.B(n_144),
.Y(n_4189)
);

OAI221xp5_ASAP7_75t_L g4190 ( 
.A1(n_4038),
.A2(n_146),
.B1(n_144),
.B2(n_145),
.C(n_147),
.Y(n_4190)
);

INVx1_ASAP7_75t_L g4191 ( 
.A(n_4129),
.Y(n_4191)
);

INVx1_ASAP7_75t_SL g4192 ( 
.A(n_4092),
.Y(n_4192)
);

AO31x2_ASAP7_75t_L g4193 ( 
.A1(n_4118),
.A2(n_147),
.A3(n_145),
.B(n_146),
.Y(n_4193)
);

BUFx12f_ASAP7_75t_L g4194 ( 
.A(n_4014),
.Y(n_4194)
);

INVx1_ASAP7_75t_L g4195 ( 
.A(n_3984),
.Y(n_4195)
);

AND2x2_ASAP7_75t_L g4196 ( 
.A(n_4034),
.B(n_511),
.Y(n_4196)
);

OR2x6_ASAP7_75t_L g4197 ( 
.A(n_4047),
.B(n_511),
.Y(n_4197)
);

NAND2xp5_ASAP7_75t_L g4198 ( 
.A(n_3986),
.B(n_512),
.Y(n_4198)
);

OAI22xp33_ASAP7_75t_L g4199 ( 
.A1(n_3997),
.A2(n_516),
.B1(n_517),
.B2(n_513),
.Y(n_4199)
);

BUFx3_ASAP7_75t_L g4200 ( 
.A(n_4050),
.Y(n_4200)
);

INVx1_ASAP7_75t_L g4201 ( 
.A(n_3994),
.Y(n_4201)
);

INVx3_ASAP7_75t_L g4202 ( 
.A(n_4013),
.Y(n_4202)
);

AO21x1_ASAP7_75t_L g4203 ( 
.A1(n_4006),
.A2(n_145),
.B(n_146),
.Y(n_4203)
);

CKINVDCx5p33_ASAP7_75t_R g4204 ( 
.A(n_4065),
.Y(n_4204)
);

CKINVDCx5p33_ASAP7_75t_R g4205 ( 
.A(n_4019),
.Y(n_4205)
);

BUFx2_ASAP7_75t_L g4206 ( 
.A(n_3983),
.Y(n_4206)
);

NAND2x1p5_ASAP7_75t_L g4207 ( 
.A(n_4035),
.B(n_4088),
.Y(n_4207)
);

OR2x6_ASAP7_75t_L g4208 ( 
.A(n_4027),
.B(n_518),
.Y(n_4208)
);

OAI21x1_ASAP7_75t_L g4209 ( 
.A1(n_4095),
.A2(n_148),
.B(n_150),
.Y(n_4209)
);

OAI22xp5_ASAP7_75t_L g4210 ( 
.A1(n_4128),
.A2(n_152),
.B1(n_150),
.B2(n_151),
.Y(n_4210)
);

AO31x2_ASAP7_75t_L g4211 ( 
.A1(n_4101),
.A2(n_152),
.A3(n_150),
.B(n_151),
.Y(n_4211)
);

AOI21xp5_ASAP7_75t_L g4212 ( 
.A1(n_4020),
.A2(n_519),
.B(n_518),
.Y(n_4212)
);

OAI21x1_ASAP7_75t_L g4213 ( 
.A1(n_3985),
.A2(n_151),
.B(n_153),
.Y(n_4213)
);

AO31x2_ASAP7_75t_L g4214 ( 
.A1(n_4109),
.A2(n_156),
.A3(n_154),
.B(n_155),
.Y(n_4214)
);

OAI21xp5_ASAP7_75t_L g4215 ( 
.A1(n_4141),
.A2(n_154),
.B(n_155),
.Y(n_4215)
);

OAI221xp5_ASAP7_75t_L g4216 ( 
.A1(n_3993),
.A2(n_4003),
.B1(n_4136),
.B2(n_4082),
.C(n_4126),
.Y(n_4216)
);

O2A1O1Ixp33_ASAP7_75t_L g4217 ( 
.A1(n_3982),
.A2(n_157),
.B(n_155),
.C(n_156),
.Y(n_4217)
);

AOI22xp33_ASAP7_75t_L g4218 ( 
.A1(n_4066),
.A2(n_158),
.B1(n_156),
.B2(n_157),
.Y(n_4218)
);

OAI21x1_ASAP7_75t_L g4219 ( 
.A1(n_4114),
.A2(n_4127),
.B(n_4124),
.Y(n_4219)
);

AO21x2_ASAP7_75t_L g4220 ( 
.A1(n_4119),
.A2(n_4007),
.B(n_4008),
.Y(n_4220)
);

INVx1_ASAP7_75t_L g4221 ( 
.A(n_3987),
.Y(n_4221)
);

INVx1_ASAP7_75t_L g4222 ( 
.A(n_3987),
.Y(n_4222)
);

INVx1_ASAP7_75t_L g4223 ( 
.A(n_3999),
.Y(n_4223)
);

OAI21x1_ASAP7_75t_SL g4224 ( 
.A1(n_3998),
.A2(n_157),
.B(n_158),
.Y(n_4224)
);

AOI22xp33_ASAP7_75t_L g4225 ( 
.A1(n_4012),
.A2(n_160),
.B1(n_158),
.B2(n_159),
.Y(n_4225)
);

CKINVDCx11_ASAP7_75t_R g4226 ( 
.A(n_4061),
.Y(n_4226)
);

OAI21x1_ASAP7_75t_SL g4227 ( 
.A1(n_4100),
.A2(n_4090),
.B(n_4071),
.Y(n_4227)
);

INVx1_ASAP7_75t_SL g4228 ( 
.A(n_3988),
.Y(n_4228)
);

AO21x2_ASAP7_75t_L g4229 ( 
.A1(n_4030),
.A2(n_159),
.B(n_161),
.Y(n_4229)
);

AO31x2_ASAP7_75t_L g4230 ( 
.A1(n_4139),
.A2(n_162),
.A3(n_159),
.B(n_161),
.Y(n_4230)
);

BUFx8_ASAP7_75t_L g4231 ( 
.A(n_4084),
.Y(n_4231)
);

NAND2xp5_ASAP7_75t_L g4232 ( 
.A(n_4116),
.B(n_520),
.Y(n_4232)
);

OAI21x1_ASAP7_75t_L g4233 ( 
.A1(n_4077),
.A2(n_162),
.B(n_163),
.Y(n_4233)
);

INVx4_ASAP7_75t_SL g4234 ( 
.A(n_4027),
.Y(n_4234)
);

NOR2xp33_ASAP7_75t_L g4235 ( 
.A(n_3979),
.B(n_4111),
.Y(n_4235)
);

INVxp67_ASAP7_75t_SL g4236 ( 
.A(n_4053),
.Y(n_4236)
);

CKINVDCx5p33_ASAP7_75t_R g4237 ( 
.A(n_4057),
.Y(n_4237)
);

INVx1_ASAP7_75t_L g4238 ( 
.A(n_3999),
.Y(n_4238)
);

INVx1_ASAP7_75t_L g4239 ( 
.A(n_4125),
.Y(n_4239)
);

A2O1A1Ixp33_ASAP7_75t_L g4240 ( 
.A1(n_4099),
.A2(n_522),
.B(n_523),
.C(n_521),
.Y(n_4240)
);

INVx5_ASAP7_75t_SL g4241 ( 
.A(n_4022),
.Y(n_4241)
);

AND2x2_ASAP7_75t_L g4242 ( 
.A(n_4089),
.B(n_4096),
.Y(n_4242)
);

OAI21x1_ASAP7_75t_L g4243 ( 
.A1(n_4080),
.A2(n_164),
.B(n_165),
.Y(n_4243)
);

CKINVDCx16_ASAP7_75t_R g4244 ( 
.A(n_4132),
.Y(n_4244)
);

OR2x2_ASAP7_75t_L g4245 ( 
.A(n_4067),
.B(n_524),
.Y(n_4245)
);

AND2x4_ASAP7_75t_L g4246 ( 
.A(n_4059),
.B(n_524),
.Y(n_4246)
);

INVx1_ASAP7_75t_L g4247 ( 
.A(n_4105),
.Y(n_4247)
);

OAI22xp33_ASAP7_75t_L g4248 ( 
.A1(n_4033),
.A2(n_526),
.B1(n_527),
.B2(n_525),
.Y(n_4248)
);

OAI21xp5_ASAP7_75t_L g4249 ( 
.A1(n_4016),
.A2(n_164),
.B(n_165),
.Y(n_4249)
);

NAND2x1p5_ASAP7_75t_L g4250 ( 
.A(n_4035),
.B(n_526),
.Y(n_4250)
);

OA21x2_ASAP7_75t_L g4251 ( 
.A1(n_4138),
.A2(n_166),
.B(n_167),
.Y(n_4251)
);

OAI21xp5_ASAP7_75t_SL g4252 ( 
.A1(n_4122),
.A2(n_168),
.B(n_169),
.Y(n_4252)
);

INVx1_ASAP7_75t_L g4253 ( 
.A(n_4105),
.Y(n_4253)
);

INVx2_ASAP7_75t_L g4254 ( 
.A(n_4120),
.Y(n_4254)
);

AOI21xp5_ASAP7_75t_L g4255 ( 
.A1(n_4021),
.A2(n_530),
.B(n_529),
.Y(n_4255)
);

CKINVDCx8_ASAP7_75t_R g4256 ( 
.A(n_4042),
.Y(n_4256)
);

INVx3_ASAP7_75t_L g4257 ( 
.A(n_4131),
.Y(n_4257)
);

HB1xp67_ASAP7_75t_L g4258 ( 
.A(n_4171),
.Y(n_4258)
);

AOI22xp33_ASAP7_75t_L g4259 ( 
.A1(n_4216),
.A2(n_4021),
.B1(n_4051),
.B2(n_4115),
.Y(n_4259)
);

AND2x2_ASAP7_75t_L g4260 ( 
.A(n_4242),
.B(n_4098),
.Y(n_4260)
);

HB1xp67_ASAP7_75t_L g4261 ( 
.A(n_4178),
.Y(n_4261)
);

AO31x2_ASAP7_75t_L g4262 ( 
.A1(n_4175),
.A2(n_4000),
.A3(n_4108),
.B(n_4043),
.Y(n_4262)
);

BUFx8_ASAP7_75t_SL g4263 ( 
.A(n_4157),
.Y(n_4263)
);

AO21x2_ASAP7_75t_L g4264 ( 
.A1(n_4144),
.A2(n_4134),
.B(n_4048),
.Y(n_4264)
);

INVx2_ASAP7_75t_L g4265 ( 
.A(n_4170),
.Y(n_4265)
);

NAND2x1p5_ASAP7_75t_L g4266 ( 
.A(n_4228),
.B(n_4002),
.Y(n_4266)
);

BUFx4_ASAP7_75t_R g4267 ( 
.A(n_4200),
.Y(n_4267)
);

OAI21x1_ASAP7_75t_L g4268 ( 
.A1(n_4219),
.A2(n_4091),
.B(n_4106),
.Y(n_4268)
);

AO31x2_ASAP7_75t_L g4269 ( 
.A1(n_4223),
.A2(n_4097),
.A3(n_4058),
.B(n_4060),
.Y(n_4269)
);

INVx4_ASAP7_75t_L g4270 ( 
.A(n_4204),
.Y(n_4270)
);

OAI21x1_ASAP7_75t_L g4271 ( 
.A1(n_4159),
.A2(n_4135),
.B(n_4018),
.Y(n_4271)
);

NAND2xp5_ASAP7_75t_SL g4272 ( 
.A(n_4166),
.B(n_4031),
.Y(n_4272)
);

OA21x2_ASAP7_75t_L g4273 ( 
.A1(n_4212),
.A2(n_4133),
.B(n_4112),
.Y(n_4273)
);

NAND2xp5_ASAP7_75t_L g4274 ( 
.A(n_4236),
.B(n_4075),
.Y(n_4274)
);

BUFx2_ASAP7_75t_SL g4275 ( 
.A(n_4202),
.Y(n_4275)
);

INVx2_ASAP7_75t_L g4276 ( 
.A(n_4179),
.Y(n_4276)
);

AND2x2_ASAP7_75t_L g4277 ( 
.A(n_4254),
.B(n_4103),
.Y(n_4277)
);

AO21x2_ASAP7_75t_L g4278 ( 
.A1(n_4221),
.A2(n_4076),
.B(n_4054),
.Y(n_4278)
);

INVxp67_ASAP7_75t_L g4279 ( 
.A(n_4235),
.Y(n_4279)
);

OAI21x1_ASAP7_75t_SL g4280 ( 
.A1(n_4203),
.A2(n_4023),
.B(n_4032),
.Y(n_4280)
);

NAND2xp5_ASAP7_75t_L g4281 ( 
.A(n_4181),
.B(n_4102),
.Y(n_4281)
);

HB1xp67_ASAP7_75t_L g4282 ( 
.A(n_4239),
.Y(n_4282)
);

NAND3xp33_ASAP7_75t_L g4283 ( 
.A(n_4249),
.B(n_4094),
.C(n_3996),
.Y(n_4283)
);

AOI21x1_ASAP7_75t_L g4284 ( 
.A1(n_4189),
.A2(n_4022),
.B(n_4026),
.Y(n_4284)
);

AND2x4_ASAP7_75t_L g4285 ( 
.A(n_4206),
.B(n_4117),
.Y(n_4285)
);

AOI21xp5_ASAP7_75t_L g4286 ( 
.A1(n_4148),
.A2(n_4137),
.B(n_4037),
.Y(n_4286)
);

OA21x2_ASAP7_75t_L g4287 ( 
.A1(n_4238),
.A2(n_4255),
.B(n_4146),
.Y(n_4287)
);

AOI21xp5_ASAP7_75t_L g4288 ( 
.A1(n_4215),
.A2(n_4104),
.B(n_4110),
.Y(n_4288)
);

AO21x2_ASAP7_75t_L g4289 ( 
.A1(n_4222),
.A2(n_4104),
.B(n_4110),
.Y(n_4289)
);

INVx1_ASAP7_75t_L g4290 ( 
.A(n_4149),
.Y(n_4290)
);

AOI222xp33_ASAP7_75t_L g4291 ( 
.A1(n_4252),
.A2(n_4177),
.B1(n_4143),
.B2(n_4190),
.C1(n_4150),
.C2(n_4210),
.Y(n_4291)
);

INVx1_ASAP7_75t_L g4292 ( 
.A(n_4152),
.Y(n_4292)
);

BUFx2_ASAP7_75t_L g4293 ( 
.A(n_4207),
.Y(n_4293)
);

NAND2xp5_ASAP7_75t_L g4294 ( 
.A(n_4192),
.B(n_4113),
.Y(n_4294)
);

AO31x2_ASAP7_75t_L g4295 ( 
.A1(n_4201),
.A2(n_4113),
.A3(n_170),
.B(n_168),
.Y(n_4295)
);

OR2x6_ASAP7_75t_L g4296 ( 
.A(n_4194),
.B(n_530),
.Y(n_4296)
);

INVx1_ASAP7_75t_L g4297 ( 
.A(n_4160),
.Y(n_4297)
);

OAI21x1_ASAP7_75t_L g4298 ( 
.A1(n_4158),
.A2(n_170),
.B(n_171),
.Y(n_4298)
);

OAI21x1_ASAP7_75t_L g4299 ( 
.A1(n_4227),
.A2(n_171),
.B(n_172),
.Y(n_4299)
);

NAND2xp5_ASAP7_75t_L g4300 ( 
.A(n_4176),
.B(n_531),
.Y(n_4300)
);

OA21x2_ASAP7_75t_L g4301 ( 
.A1(n_4165),
.A2(n_4209),
.B(n_4188),
.Y(n_4301)
);

INVx1_ASAP7_75t_L g4302 ( 
.A(n_4164),
.Y(n_4302)
);

HB1xp67_ASAP7_75t_L g4303 ( 
.A(n_4182),
.Y(n_4303)
);

OA21x2_ASAP7_75t_L g4304 ( 
.A1(n_4233),
.A2(n_172),
.B(n_173),
.Y(n_4304)
);

OAI21x1_ASAP7_75t_SL g4305 ( 
.A1(n_4224),
.A2(n_173),
.B(n_174),
.Y(n_4305)
);

AO21x2_ASAP7_75t_L g4306 ( 
.A1(n_4195),
.A2(n_174),
.B(n_175),
.Y(n_4306)
);

NOR2xp33_ASAP7_75t_L g4307 ( 
.A(n_4256),
.B(n_532),
.Y(n_4307)
);

BUFx6f_ASAP7_75t_L g4308 ( 
.A(n_4180),
.Y(n_4308)
);

INVx3_ASAP7_75t_L g4309 ( 
.A(n_4257),
.Y(n_4309)
);

AO31x2_ASAP7_75t_L g4310 ( 
.A1(n_4247),
.A2(n_180),
.A3(n_177),
.B(n_178),
.Y(n_4310)
);

INVx1_ASAP7_75t_L g4311 ( 
.A(n_4183),
.Y(n_4311)
);

INVx2_ASAP7_75t_SL g4312 ( 
.A(n_4142),
.Y(n_4312)
);

INVx1_ASAP7_75t_L g4313 ( 
.A(n_4187),
.Y(n_4313)
);

INVx1_ASAP7_75t_L g4314 ( 
.A(n_4191),
.Y(n_4314)
);

OAI22xp5_ASAP7_75t_L g4315 ( 
.A1(n_4174),
.A2(n_181),
.B1(n_178),
.B2(n_180),
.Y(n_4315)
);

INVx1_ASAP7_75t_L g4316 ( 
.A(n_4253),
.Y(n_4316)
);

NAND2x1p5_ASAP7_75t_L g4317 ( 
.A(n_4155),
.B(n_535),
.Y(n_4317)
);

INVx2_ASAP7_75t_L g4318 ( 
.A(n_4147),
.Y(n_4318)
);

BUFx8_ASAP7_75t_L g4319 ( 
.A(n_4196),
.Y(n_4319)
);

AO21x2_ASAP7_75t_L g4320 ( 
.A1(n_4184),
.A2(n_180),
.B(n_181),
.Y(n_4320)
);

OAI21x1_ASAP7_75t_L g4321 ( 
.A1(n_4213),
.A2(n_182),
.B(n_183),
.Y(n_4321)
);

NAND2xp5_ASAP7_75t_L g4322 ( 
.A(n_4151),
.B(n_535),
.Y(n_4322)
);

CKINVDCx6p67_ASAP7_75t_R g4323 ( 
.A(n_4244),
.Y(n_4323)
);

NAND2xp5_ASAP7_75t_L g4324 ( 
.A(n_4232),
.B(n_536),
.Y(n_4324)
);

AOI21xp5_ASAP7_75t_L g4325 ( 
.A1(n_4145),
.A2(n_185),
.B(n_186),
.Y(n_4325)
);

NOR2xp33_ASAP7_75t_L g4326 ( 
.A(n_4168),
.B(n_4237),
.Y(n_4326)
);

INVx2_ASAP7_75t_L g4327 ( 
.A(n_4169),
.Y(n_4327)
);

NAND2xp5_ASAP7_75t_L g4328 ( 
.A(n_4220),
.B(n_537),
.Y(n_4328)
);

AO31x2_ASAP7_75t_L g4329 ( 
.A1(n_4240),
.A2(n_187),
.A3(n_185),
.B(n_186),
.Y(n_4329)
);

OAI21xp5_ASAP7_75t_L g4330 ( 
.A1(n_4217),
.A2(n_185),
.B(n_186),
.Y(n_4330)
);

INVxp67_ASAP7_75t_SL g4331 ( 
.A(n_4162),
.Y(n_4331)
);

NAND2xp5_ASAP7_75t_L g4332 ( 
.A(n_4153),
.B(n_538),
.Y(n_4332)
);

INVx2_ASAP7_75t_L g4333 ( 
.A(n_4243),
.Y(n_4333)
);

BUFx2_ASAP7_75t_L g4334 ( 
.A(n_4234),
.Y(n_4334)
);

NAND2xp5_ASAP7_75t_L g4335 ( 
.A(n_4185),
.B(n_538),
.Y(n_4335)
);

OAI21x1_ASAP7_75t_L g4336 ( 
.A1(n_4251),
.A2(n_187),
.B(n_188),
.Y(n_4336)
);

INVx1_ASAP7_75t_L g4337 ( 
.A(n_4214),
.Y(n_4337)
);

INVx1_ASAP7_75t_L g4338 ( 
.A(n_4214),
.Y(n_4338)
);

OAI21x1_ASAP7_75t_L g4339 ( 
.A1(n_4156),
.A2(n_187),
.B(n_188),
.Y(n_4339)
);

AND2x2_ASAP7_75t_L g4340 ( 
.A(n_4154),
.B(n_540),
.Y(n_4340)
);

INVx1_ASAP7_75t_L g4341 ( 
.A(n_4230),
.Y(n_4341)
);

AND2x2_ASAP7_75t_L g4342 ( 
.A(n_4161),
.B(n_542),
.Y(n_4342)
);

AOI21xp5_ASAP7_75t_L g4343 ( 
.A1(n_4186),
.A2(n_189),
.B(n_190),
.Y(n_4343)
);

INVx1_ASAP7_75t_L g4344 ( 
.A(n_4230),
.Y(n_4344)
);

OA21x2_ASAP7_75t_L g4345 ( 
.A1(n_4198),
.A2(n_189),
.B(n_190),
.Y(n_4345)
);

INVx1_ASAP7_75t_L g4346 ( 
.A(n_4193),
.Y(n_4346)
);

INVx1_ASAP7_75t_L g4347 ( 
.A(n_4193),
.Y(n_4347)
);

OAI21x1_ASAP7_75t_L g4348 ( 
.A1(n_4173),
.A2(n_191),
.B(n_192),
.Y(n_4348)
);

AOI22xp33_ASAP7_75t_L g4349 ( 
.A1(n_4199),
.A2(n_194),
.B1(n_192),
.B2(n_193),
.Y(n_4349)
);

INVx1_ASAP7_75t_L g4350 ( 
.A(n_4211),
.Y(n_4350)
);

OAI21xp5_ASAP7_75t_L g4351 ( 
.A1(n_4218),
.A2(n_4225),
.B(n_4172),
.Y(n_4351)
);

O2A1O1Ixp33_ASAP7_75t_L g4352 ( 
.A1(n_4248),
.A2(n_195),
.B(n_192),
.C(n_193),
.Y(n_4352)
);

BUFx6f_ASAP7_75t_L g4353 ( 
.A(n_4246),
.Y(n_4353)
);

BUFx6f_ASAP7_75t_L g4354 ( 
.A(n_4226),
.Y(n_4354)
);

INVx2_ASAP7_75t_L g4355 ( 
.A(n_4229),
.Y(n_4355)
);

AOI222xp33_ASAP7_75t_L g4356 ( 
.A1(n_4167),
.A2(n_4241),
.B1(n_4163),
.B2(n_4231),
.C1(n_4205),
.C2(n_4208),
.Y(n_4356)
);

NAND2xp5_ASAP7_75t_L g4357 ( 
.A(n_4245),
.B(n_543),
.Y(n_4357)
);

INVx1_ASAP7_75t_L g4358 ( 
.A(n_4197),
.Y(n_4358)
);

AOI22xp5_ASAP7_75t_L g4359 ( 
.A1(n_4291),
.A2(n_4208),
.B1(n_4241),
.B2(n_4197),
.Y(n_4359)
);

OR2x2_ASAP7_75t_L g4360 ( 
.A(n_4258),
.B(n_4250),
.Y(n_4360)
);

INVx2_ASAP7_75t_L g4361 ( 
.A(n_4290),
.Y(n_4361)
);

INVx1_ASAP7_75t_L g4362 ( 
.A(n_4292),
.Y(n_4362)
);

OR2x2_ASAP7_75t_L g4363 ( 
.A(n_4261),
.B(n_543),
.Y(n_4363)
);

HB1xp67_ASAP7_75t_L g4364 ( 
.A(n_4282),
.Y(n_4364)
);

AND2x2_ASAP7_75t_L g4365 ( 
.A(n_4279),
.B(n_546),
.Y(n_4365)
);

INVx1_ASAP7_75t_L g4366 ( 
.A(n_4297),
.Y(n_4366)
);

AND2x2_ASAP7_75t_L g4367 ( 
.A(n_4266),
.B(n_547),
.Y(n_4367)
);

HB1xp67_ASAP7_75t_L g4368 ( 
.A(n_4294),
.Y(n_4368)
);

AOI22xp33_ASAP7_75t_L g4369 ( 
.A1(n_4330),
.A2(n_549),
.B1(n_550),
.B2(n_548),
.Y(n_4369)
);

OR2x2_ASAP7_75t_L g4370 ( 
.A(n_4274),
.B(n_549),
.Y(n_4370)
);

INVx1_ASAP7_75t_L g4371 ( 
.A(n_4302),
.Y(n_4371)
);

INVx4_ASAP7_75t_L g4372 ( 
.A(n_4267),
.Y(n_4372)
);

INVx1_ASAP7_75t_L g4373 ( 
.A(n_4311),
.Y(n_4373)
);

OR2x2_ASAP7_75t_L g4374 ( 
.A(n_4313),
.B(n_550),
.Y(n_4374)
);

INVx2_ASAP7_75t_L g4375 ( 
.A(n_4314),
.Y(n_4375)
);

AND2x2_ASAP7_75t_L g4376 ( 
.A(n_4277),
.B(n_551),
.Y(n_4376)
);

INVx2_ASAP7_75t_L g4377 ( 
.A(n_4265),
.Y(n_4377)
);

INVx2_ASAP7_75t_L g4378 ( 
.A(n_4276),
.Y(n_4378)
);

AND2x2_ASAP7_75t_L g4379 ( 
.A(n_4285),
.B(n_4358),
.Y(n_4379)
);

NAND2xp5_ASAP7_75t_L g4380 ( 
.A(n_4264),
.B(n_554),
.Y(n_4380)
);

INVx1_ASAP7_75t_L g4381 ( 
.A(n_4316),
.Y(n_4381)
);

BUFx3_ASAP7_75t_L g4382 ( 
.A(n_4263),
.Y(n_4382)
);

NAND2xp5_ASAP7_75t_L g4383 ( 
.A(n_4327),
.B(n_554),
.Y(n_4383)
);

INVx2_ASAP7_75t_L g4384 ( 
.A(n_4318),
.Y(n_4384)
);

INVx1_ASAP7_75t_L g4385 ( 
.A(n_4341),
.Y(n_4385)
);

AND2x4_ASAP7_75t_L g4386 ( 
.A(n_4293),
.B(n_555),
.Y(n_4386)
);

INVx2_ASAP7_75t_L g4387 ( 
.A(n_4287),
.Y(n_4387)
);

CKINVDCx5p33_ASAP7_75t_R g4388 ( 
.A(n_4323),
.Y(n_4388)
);

INVx3_ASAP7_75t_L g4389 ( 
.A(n_4309),
.Y(n_4389)
);

CKINVDCx5p33_ASAP7_75t_R g4390 ( 
.A(n_4354),
.Y(n_4390)
);

INVx2_ASAP7_75t_L g4391 ( 
.A(n_4333),
.Y(n_4391)
);

INVx1_ASAP7_75t_L g4392 ( 
.A(n_4344),
.Y(n_4392)
);

INVx2_ASAP7_75t_L g4393 ( 
.A(n_4355),
.Y(n_4393)
);

AND2x2_ASAP7_75t_L g4394 ( 
.A(n_4334),
.B(n_555),
.Y(n_4394)
);

INVx4_ASAP7_75t_L g4395 ( 
.A(n_4308),
.Y(n_4395)
);

OA21x2_ASAP7_75t_L g4396 ( 
.A1(n_4328),
.A2(n_557),
.B(n_556),
.Y(n_4396)
);

NOR2xp67_ASAP7_75t_SL g4397 ( 
.A(n_4283),
.B(n_196),
.Y(n_4397)
);

INVx2_ASAP7_75t_L g4398 ( 
.A(n_4278),
.Y(n_4398)
);

INVx1_ASAP7_75t_L g4399 ( 
.A(n_4350),
.Y(n_4399)
);

INVx2_ASAP7_75t_L g4400 ( 
.A(n_4269),
.Y(n_4400)
);

NOR2xp33_ASAP7_75t_L g4401 ( 
.A(n_4272),
.B(n_556),
.Y(n_4401)
);

INVx2_ASAP7_75t_L g4402 ( 
.A(n_4269),
.Y(n_4402)
);

INVx3_ASAP7_75t_L g4403 ( 
.A(n_4308),
.Y(n_4403)
);

OA21x2_ASAP7_75t_L g4404 ( 
.A1(n_4298),
.A2(n_559),
.B(n_558),
.Y(n_4404)
);

INVx1_ASAP7_75t_L g4405 ( 
.A(n_4337),
.Y(n_4405)
);

INVx1_ASAP7_75t_L g4406 ( 
.A(n_4338),
.Y(n_4406)
);

INVx1_ASAP7_75t_L g4407 ( 
.A(n_4289),
.Y(n_4407)
);

INVx2_ASAP7_75t_SL g4408 ( 
.A(n_4354),
.Y(n_4408)
);

INVx1_ASAP7_75t_L g4409 ( 
.A(n_4346),
.Y(n_4409)
);

INVx2_ASAP7_75t_L g4410 ( 
.A(n_4301),
.Y(n_4410)
);

HB1xp67_ASAP7_75t_L g4411 ( 
.A(n_4347),
.Y(n_4411)
);

HB1xp67_ASAP7_75t_L g4412 ( 
.A(n_4331),
.Y(n_4412)
);

AND2x2_ASAP7_75t_L g4413 ( 
.A(n_4275),
.B(n_560),
.Y(n_4413)
);

OR2x2_ASAP7_75t_L g4414 ( 
.A(n_4273),
.B(n_4300),
.Y(n_4414)
);

INVx1_ASAP7_75t_L g4415 ( 
.A(n_4295),
.Y(n_4415)
);

NOR2x1_ASAP7_75t_R g4416 ( 
.A(n_4270),
.B(n_197),
.Y(n_4416)
);

INVx1_ASAP7_75t_L g4417 ( 
.A(n_4295),
.Y(n_4417)
);

AND2x4_ASAP7_75t_L g4418 ( 
.A(n_4312),
.B(n_561),
.Y(n_4418)
);

INVx3_ASAP7_75t_L g4419 ( 
.A(n_4353),
.Y(n_4419)
);

AND2x2_ASAP7_75t_L g4420 ( 
.A(n_4340),
.B(n_561),
.Y(n_4420)
);

INVx2_ASAP7_75t_L g4421 ( 
.A(n_4317),
.Y(n_4421)
);

NOR2xp33_ASAP7_75t_L g4422 ( 
.A(n_4324),
.B(n_562),
.Y(n_4422)
);

HB1xp67_ASAP7_75t_L g4423 ( 
.A(n_4271),
.Y(n_4423)
);

INVx1_ASAP7_75t_L g4424 ( 
.A(n_4310),
.Y(n_4424)
);

INVx1_ASAP7_75t_L g4425 ( 
.A(n_4322),
.Y(n_4425)
);

BUFx2_ASAP7_75t_L g4426 ( 
.A(n_4342),
.Y(n_4426)
);

AO21x2_ASAP7_75t_L g4427 ( 
.A1(n_4325),
.A2(n_198),
.B(n_199),
.Y(n_4427)
);

INVx2_ASAP7_75t_L g4428 ( 
.A(n_4268),
.Y(n_4428)
);

INVx1_ASAP7_75t_L g4429 ( 
.A(n_4336),
.Y(n_4429)
);

AND2x2_ASAP7_75t_L g4430 ( 
.A(n_4332),
.B(n_563),
.Y(n_4430)
);

BUFx2_ASAP7_75t_L g4431 ( 
.A(n_4262),
.Y(n_4431)
);

INVx1_ASAP7_75t_L g4432 ( 
.A(n_4345),
.Y(n_4432)
);

INVx2_ASAP7_75t_L g4433 ( 
.A(n_4299),
.Y(n_4433)
);

BUFx3_ASAP7_75t_L g4434 ( 
.A(n_4319),
.Y(n_4434)
);

NAND2xp5_ASAP7_75t_L g4435 ( 
.A(n_4259),
.B(n_563),
.Y(n_4435)
);

NOR2xp33_ASAP7_75t_L g4436 ( 
.A(n_4335),
.B(n_564),
.Y(n_4436)
);

BUFx6f_ASAP7_75t_L g4437 ( 
.A(n_4296),
.Y(n_4437)
);

NAND2xp5_ASAP7_75t_L g4438 ( 
.A(n_4288),
.B(n_565),
.Y(n_4438)
);

INVx3_ASAP7_75t_L g4439 ( 
.A(n_4284),
.Y(n_4439)
);

INVx2_ASAP7_75t_L g4440 ( 
.A(n_4306),
.Y(n_4440)
);

INVxp67_ASAP7_75t_SL g4441 ( 
.A(n_4281),
.Y(n_4441)
);

BUFx6f_ASAP7_75t_L g4442 ( 
.A(n_4326),
.Y(n_4442)
);

INVx2_ASAP7_75t_L g4443 ( 
.A(n_4321),
.Y(n_4443)
);

INVx3_ASAP7_75t_L g4444 ( 
.A(n_4339),
.Y(n_4444)
);

INVx2_ASAP7_75t_SL g4445 ( 
.A(n_4357),
.Y(n_4445)
);

INVx2_ASAP7_75t_L g4446 ( 
.A(n_4304),
.Y(n_4446)
);

OAI22xp5_ASAP7_75t_L g4447 ( 
.A1(n_4349),
.A2(n_201),
.B1(n_199),
.B2(n_200),
.Y(n_4447)
);

NAND2xp5_ASAP7_75t_L g4448 ( 
.A(n_4356),
.B(n_566),
.Y(n_4448)
);

HB1xp67_ASAP7_75t_L g4449 ( 
.A(n_4320),
.Y(n_4449)
);

BUFx6f_ASAP7_75t_L g4450 ( 
.A(n_4307),
.Y(n_4450)
);

INVx1_ASAP7_75t_L g4451 ( 
.A(n_4329),
.Y(n_4451)
);

AND2x2_ASAP7_75t_L g4452 ( 
.A(n_4286),
.B(n_567),
.Y(n_4452)
);

INVx2_ASAP7_75t_L g4453 ( 
.A(n_4305),
.Y(n_4453)
);

AND2x4_ASAP7_75t_L g4454 ( 
.A(n_4348),
.B(n_569),
.Y(n_4454)
);

INVx2_ASAP7_75t_L g4455 ( 
.A(n_4280),
.Y(n_4455)
);

CKINVDCx6p67_ASAP7_75t_R g4456 ( 
.A(n_4352),
.Y(n_4456)
);

INVx1_ASAP7_75t_L g4457 ( 
.A(n_4343),
.Y(n_4457)
);

INVx2_ASAP7_75t_SL g4458 ( 
.A(n_4315),
.Y(n_4458)
);

NOR2xp33_ASAP7_75t_L g4459 ( 
.A(n_4351),
.B(n_571),
.Y(n_4459)
);

INVx1_ASAP7_75t_L g4460 ( 
.A(n_4303),
.Y(n_4460)
);

HB1xp67_ASAP7_75t_L g4461 ( 
.A(n_4258),
.Y(n_4461)
);

AND2x2_ASAP7_75t_L g4462 ( 
.A(n_4260),
.B(n_572),
.Y(n_4462)
);

BUFx2_ASAP7_75t_L g4463 ( 
.A(n_4261),
.Y(n_4463)
);

OAI22xp5_ASAP7_75t_L g4464 ( 
.A1(n_4456),
.A2(n_204),
.B1(n_202),
.B2(n_203),
.Y(n_4464)
);

AOI22xp33_ASAP7_75t_L g4465 ( 
.A1(n_4459),
.A2(n_575),
.B1(n_576),
.B2(n_574),
.Y(n_4465)
);

OAI22xp5_ASAP7_75t_L g4466 ( 
.A1(n_4369),
.A2(n_204),
.B1(n_202),
.B2(n_203),
.Y(n_4466)
);

NAND2xp5_ASAP7_75t_L g4467 ( 
.A(n_4441),
.B(n_575),
.Y(n_4467)
);

AOI221xp5_ASAP7_75t_L g4468 ( 
.A1(n_4438),
.A2(n_206),
.B1(n_203),
.B2(n_205),
.C(n_207),
.Y(n_4468)
);

INVx1_ASAP7_75t_L g4469 ( 
.A(n_4366),
.Y(n_4469)
);

AOI21xp5_ASAP7_75t_L g4470 ( 
.A1(n_4457),
.A2(n_205),
.B(n_206),
.Y(n_4470)
);

OAI22xp5_ASAP7_75t_L g4471 ( 
.A1(n_4359),
.A2(n_207),
.B1(n_205),
.B2(n_206),
.Y(n_4471)
);

AOI22xp33_ASAP7_75t_L g4472 ( 
.A1(n_4397),
.A2(n_579),
.B1(n_581),
.B2(n_578),
.Y(n_4472)
);

INVx2_ASAP7_75t_L g4473 ( 
.A(n_4463),
.Y(n_4473)
);

OA21x2_ASAP7_75t_L g4474 ( 
.A1(n_4410),
.A2(n_208),
.B(n_210),
.Y(n_4474)
);

AND2x2_ASAP7_75t_L g4475 ( 
.A(n_4426),
.B(n_211),
.Y(n_4475)
);

OAI22xp5_ASAP7_75t_L g4476 ( 
.A1(n_4435),
.A2(n_213),
.B1(n_211),
.B2(n_212),
.Y(n_4476)
);

OAI33xp33_ASAP7_75t_L g4477 ( 
.A1(n_4432),
.A2(n_4380),
.A3(n_4414),
.B1(n_4448),
.B2(n_4451),
.B3(n_4425),
.Y(n_4477)
);

OAI22xp5_ASAP7_75t_L g4478 ( 
.A1(n_4458),
.A2(n_214),
.B1(n_212),
.B2(n_213),
.Y(n_4478)
);

AOI21xp5_ASAP7_75t_L g4479 ( 
.A1(n_4449),
.A2(n_212),
.B(n_213),
.Y(n_4479)
);

NOR2xp33_ASAP7_75t_L g4480 ( 
.A(n_4442),
.B(n_585),
.Y(n_4480)
);

INVxp67_ASAP7_75t_L g4481 ( 
.A(n_4461),
.Y(n_4481)
);

OAI221xp5_ASAP7_75t_L g4482 ( 
.A1(n_4401),
.A2(n_217),
.B1(n_215),
.B2(n_216),
.C(n_218),
.Y(n_4482)
);

OAI21x1_ASAP7_75t_L g4483 ( 
.A1(n_4387),
.A2(n_215),
.B(n_216),
.Y(n_4483)
);

INVx1_ASAP7_75t_L g4484 ( 
.A(n_4371),
.Y(n_4484)
);

OAI21xp5_ASAP7_75t_L g4485 ( 
.A1(n_4422),
.A2(n_586),
.B(n_585),
.Y(n_4485)
);

OAI21x1_ASAP7_75t_L g4486 ( 
.A1(n_4439),
.A2(n_4398),
.B(n_4400),
.Y(n_4486)
);

OAI221xp5_ASAP7_75t_L g4487 ( 
.A1(n_4436),
.A2(n_218),
.B1(n_215),
.B2(n_217),
.C(n_219),
.Y(n_4487)
);

AOI22xp5_ASAP7_75t_L g4488 ( 
.A1(n_4455),
.A2(n_588),
.B1(n_589),
.B2(n_587),
.Y(n_4488)
);

AND2x2_ASAP7_75t_L g4489 ( 
.A(n_4379),
.B(n_4368),
.Y(n_4489)
);

INVx1_ASAP7_75t_L g4490 ( 
.A(n_4373),
.Y(n_4490)
);

OR2x2_ASAP7_75t_L g4491 ( 
.A(n_4364),
.B(n_224),
.Y(n_4491)
);

OAI22xp5_ASAP7_75t_L g4492 ( 
.A1(n_4453),
.A2(n_226),
.B1(n_224),
.B2(n_225),
.Y(n_4492)
);

INVx2_ASAP7_75t_L g4493 ( 
.A(n_4361),
.Y(n_4493)
);

INVx2_ASAP7_75t_L g4494 ( 
.A(n_4375),
.Y(n_4494)
);

OAI321xp33_ASAP7_75t_L g4495 ( 
.A1(n_4431),
.A2(n_227),
.A3(n_229),
.B1(n_225),
.B2(n_226),
.C(n_228),
.Y(n_4495)
);

AOI21xp5_ASAP7_75t_L g4496 ( 
.A1(n_4440),
.A2(n_225),
.B(n_226),
.Y(n_4496)
);

OAI22xp33_ASAP7_75t_L g4497 ( 
.A1(n_4396),
.A2(n_591),
.B1(n_592),
.B2(n_590),
.Y(n_4497)
);

AOI22xp5_ASAP7_75t_L g4498 ( 
.A1(n_4421),
.A2(n_593),
.B1(n_594),
.B2(n_592),
.Y(n_4498)
);

AOI221x1_ASAP7_75t_L g4499 ( 
.A1(n_4383),
.A2(n_229),
.B1(n_227),
.B2(n_228),
.C(n_230),
.Y(n_4499)
);

OAI21x1_ASAP7_75t_L g4500 ( 
.A1(n_4402),
.A2(n_228),
.B(n_230),
.Y(n_4500)
);

INVx1_ASAP7_75t_L g4501 ( 
.A(n_4381),
.Y(n_4501)
);

AOI22xp33_ASAP7_75t_L g4502 ( 
.A1(n_4450),
.A2(n_594),
.B1(n_595),
.B2(n_593),
.Y(n_4502)
);

BUFx6f_ASAP7_75t_L g4503 ( 
.A(n_4434),
.Y(n_4503)
);

AND2x2_ASAP7_75t_L g4504 ( 
.A(n_4460),
.B(n_232),
.Y(n_4504)
);

AOI211xp5_ASAP7_75t_L g4505 ( 
.A1(n_4416),
.A2(n_234),
.B(n_232),
.C(n_233),
.Y(n_4505)
);

AOI22xp33_ASAP7_75t_L g4506 ( 
.A1(n_4450),
.A2(n_596),
.B1(n_597),
.B2(n_595),
.Y(n_4506)
);

AOI22xp5_ASAP7_75t_L g4507 ( 
.A1(n_4427),
.A2(n_598),
.B1(n_599),
.B2(n_597),
.Y(n_4507)
);

OAI21xp33_ASAP7_75t_L g4508 ( 
.A1(n_4452),
.A2(n_233),
.B(n_234),
.Y(n_4508)
);

INVx1_ASAP7_75t_L g4509 ( 
.A(n_4409),
.Y(n_4509)
);

AOI21xp5_ASAP7_75t_L g4510 ( 
.A1(n_4423),
.A2(n_237),
.B(n_239),
.Y(n_4510)
);

AOI22xp33_ASAP7_75t_L g4511 ( 
.A1(n_4454),
.A2(n_601),
.B1(n_602),
.B2(n_600),
.Y(n_4511)
);

INVx1_ASAP7_75t_L g4512 ( 
.A(n_4405),
.Y(n_4512)
);

NAND2xp5_ASAP7_75t_L g4513 ( 
.A(n_4377),
.B(n_602),
.Y(n_4513)
);

AND2x2_ASAP7_75t_L g4514 ( 
.A(n_4389),
.B(n_237),
.Y(n_4514)
);

BUFx8_ASAP7_75t_L g4515 ( 
.A(n_4394),
.Y(n_4515)
);

OAI22xp33_ASAP7_75t_L g4516 ( 
.A1(n_4370),
.A2(n_4444),
.B1(n_4445),
.B2(n_4447),
.Y(n_4516)
);

INVx1_ASAP7_75t_L g4517 ( 
.A(n_4406),
.Y(n_4517)
);

INVx1_ASAP7_75t_L g4518 ( 
.A(n_4385),
.Y(n_4518)
);

OAI22xp5_ASAP7_75t_L g4519 ( 
.A1(n_4360),
.A2(n_241),
.B1(n_239),
.B2(n_240),
.Y(n_4519)
);

OA21x2_ASAP7_75t_L g4520 ( 
.A1(n_4407),
.A2(n_239),
.B(n_240),
.Y(n_4520)
);

AND2x4_ASAP7_75t_L g4521 ( 
.A(n_4429),
.B(n_242),
.Y(n_4521)
);

NAND2xp5_ASAP7_75t_L g4522 ( 
.A(n_4378),
.B(n_603),
.Y(n_4522)
);

BUFx4f_ASAP7_75t_SL g4523 ( 
.A(n_4408),
.Y(n_4523)
);

AOI22xp33_ASAP7_75t_L g4524 ( 
.A1(n_4437),
.A2(n_4430),
.B1(n_4433),
.B2(n_4443),
.Y(n_4524)
);

INVx2_ASAP7_75t_L g4525 ( 
.A(n_4384),
.Y(n_4525)
);

BUFx3_ASAP7_75t_L g4526 ( 
.A(n_4390),
.Y(n_4526)
);

AND2x2_ASAP7_75t_L g4527 ( 
.A(n_4419),
.B(n_243),
.Y(n_4527)
);

OAI22xp5_ASAP7_75t_L g4528 ( 
.A1(n_4403),
.A2(n_246),
.B1(n_244),
.B2(n_245),
.Y(n_4528)
);

OAI21x1_ASAP7_75t_L g4529 ( 
.A1(n_4428),
.A2(n_244),
.B(n_245),
.Y(n_4529)
);

NAND2xp5_ASAP7_75t_L g4530 ( 
.A(n_4393),
.B(n_604),
.Y(n_4530)
);

AOI22xp33_ASAP7_75t_L g4531 ( 
.A1(n_4367),
.A2(n_607),
.B1(n_608),
.B2(n_606),
.Y(n_4531)
);

BUFx2_ASAP7_75t_L g4532 ( 
.A(n_4412),
.Y(n_4532)
);

AOI22xp33_ASAP7_75t_L g4533 ( 
.A1(n_4404),
.A2(n_608),
.B1(n_609),
.B2(n_606),
.Y(n_4533)
);

AOI22xp33_ASAP7_75t_L g4534 ( 
.A1(n_4446),
.A2(n_4462),
.B1(n_4386),
.B2(n_4420),
.Y(n_4534)
);

INVx1_ASAP7_75t_L g4535 ( 
.A(n_4392),
.Y(n_4535)
);

INVx1_ASAP7_75t_L g4536 ( 
.A(n_4399),
.Y(n_4536)
);

NAND2xp5_ASAP7_75t_L g4537 ( 
.A(n_4415),
.B(n_609),
.Y(n_4537)
);

OAI221xp5_ASAP7_75t_L g4538 ( 
.A1(n_4374),
.A2(n_250),
.B1(n_248),
.B2(n_249),
.C(n_251),
.Y(n_4538)
);

AOI211xp5_ASAP7_75t_L g4539 ( 
.A1(n_4413),
.A2(n_251),
.B(n_249),
.C(n_250),
.Y(n_4539)
);

INVx1_ASAP7_75t_L g4540 ( 
.A(n_4411),
.Y(n_4540)
);

NAND2xp5_ASAP7_75t_L g4541 ( 
.A(n_4417),
.B(n_4424),
.Y(n_4541)
);

INVx1_ASAP7_75t_SL g4542 ( 
.A(n_4388),
.Y(n_4542)
);

OAI22xp33_ASAP7_75t_L g4543 ( 
.A1(n_4363),
.A2(n_612),
.B1(n_613),
.B2(n_611),
.Y(n_4543)
);

INVx1_ASAP7_75t_L g4544 ( 
.A(n_4391),
.Y(n_4544)
);

NAND3xp33_ASAP7_75t_L g4545 ( 
.A(n_4365),
.B(n_615),
.C(n_614),
.Y(n_4545)
);

INVxp67_ASAP7_75t_L g4546 ( 
.A(n_4376),
.Y(n_4546)
);

NAND2xp5_ASAP7_75t_L g4547 ( 
.A(n_4395),
.B(n_616),
.Y(n_4547)
);

OA21x2_ASAP7_75t_L g4548 ( 
.A1(n_4418),
.A2(n_252),
.B(n_253),
.Y(n_4548)
);

AND2x2_ASAP7_75t_L g4549 ( 
.A(n_4463),
.B(n_253),
.Y(n_4549)
);

INVx2_ASAP7_75t_L g4550 ( 
.A(n_4463),
.Y(n_4550)
);

INVx1_ASAP7_75t_L g4551 ( 
.A(n_4362),
.Y(n_4551)
);

BUFx2_ASAP7_75t_L g4552 ( 
.A(n_4463),
.Y(n_4552)
);

OAI221xp5_ASAP7_75t_L g4553 ( 
.A1(n_4459),
.A2(n_256),
.B1(n_254),
.B2(n_255),
.C(n_257),
.Y(n_4553)
);

AND2x2_ASAP7_75t_L g4554 ( 
.A(n_4463),
.B(n_254),
.Y(n_4554)
);

AOI22xp33_ASAP7_75t_SL g4555 ( 
.A1(n_4459),
.A2(n_617),
.B1(n_618),
.B2(n_616),
.Y(n_4555)
);

BUFx2_ASAP7_75t_SL g4556 ( 
.A(n_4372),
.Y(n_4556)
);

AOI22xp33_ASAP7_75t_L g4557 ( 
.A1(n_4456),
.A2(n_618),
.B1(n_619),
.B2(n_617),
.Y(n_4557)
);

INVx2_ASAP7_75t_L g4558 ( 
.A(n_4463),
.Y(n_4558)
);

AOI22xp33_ASAP7_75t_L g4559 ( 
.A1(n_4456),
.A2(n_621),
.B1(n_622),
.B2(n_620),
.Y(n_4559)
);

INVx1_ASAP7_75t_SL g4560 ( 
.A(n_4382),
.Y(n_4560)
);

CKINVDCx5p33_ASAP7_75t_R g4561 ( 
.A(n_4382),
.Y(n_4561)
);

CKINVDCx5p33_ASAP7_75t_R g4562 ( 
.A(n_4382),
.Y(n_4562)
);

OAI22xp5_ASAP7_75t_L g4563 ( 
.A1(n_4456),
.A2(n_262),
.B1(n_259),
.B2(n_261),
.Y(n_4563)
);

AND2x2_ASAP7_75t_L g4564 ( 
.A(n_4463),
.B(n_259),
.Y(n_4564)
);

OAI22xp5_ASAP7_75t_L g4565 ( 
.A1(n_4456),
.A2(n_263),
.B1(n_261),
.B2(n_262),
.Y(n_4565)
);

NAND2xp5_ASAP7_75t_L g4566 ( 
.A(n_4441),
.B(n_620),
.Y(n_4566)
);

OAI22xp33_ASAP7_75t_L g4567 ( 
.A1(n_4456),
.A2(n_623),
.B1(n_624),
.B2(n_622),
.Y(n_4567)
);

AOI221xp5_ASAP7_75t_L g4568 ( 
.A1(n_4459),
.A2(n_265),
.B1(n_263),
.B2(n_264),
.C(n_266),
.Y(n_4568)
);

OAI221xp5_ASAP7_75t_L g4569 ( 
.A1(n_4459),
.A2(n_266),
.B1(n_264),
.B2(n_265),
.C(n_267),
.Y(n_4569)
);

OAI221xp5_ASAP7_75t_L g4570 ( 
.A1(n_4459),
.A2(n_266),
.B1(n_264),
.B2(n_265),
.C(n_267),
.Y(n_4570)
);

OAI21x1_ASAP7_75t_L g4571 ( 
.A1(n_4387),
.A2(n_267),
.B(n_268),
.Y(n_4571)
);

OAI221xp5_ASAP7_75t_SL g4572 ( 
.A1(n_4456),
.A2(n_270),
.B1(n_268),
.B2(n_269),
.C(n_271),
.Y(n_4572)
);

INVx1_ASAP7_75t_L g4573 ( 
.A(n_4362),
.Y(n_4573)
);

AND2x2_ASAP7_75t_L g4574 ( 
.A(n_4463),
.B(n_269),
.Y(n_4574)
);

INVx1_ASAP7_75t_SL g4575 ( 
.A(n_4382),
.Y(n_4575)
);

OAI22xp33_ASAP7_75t_L g4576 ( 
.A1(n_4456),
.A2(n_625),
.B1(n_626),
.B2(n_623),
.Y(n_4576)
);

INVx1_ASAP7_75t_L g4577 ( 
.A(n_4362),
.Y(n_4577)
);

AND2x4_ASAP7_75t_L g4578 ( 
.A(n_4552),
.B(n_625),
.Y(n_4578)
);

INVx2_ASAP7_75t_L g4579 ( 
.A(n_4532),
.Y(n_4579)
);

INVx1_ASAP7_75t_L g4580 ( 
.A(n_4509),
.Y(n_4580)
);

HB1xp67_ASAP7_75t_L g4581 ( 
.A(n_4540),
.Y(n_4581)
);

OR2x6_ASAP7_75t_SL g4582 ( 
.A(n_4561),
.B(n_269),
.Y(n_4582)
);

NAND2xp5_ASAP7_75t_L g4583 ( 
.A(n_4481),
.B(n_627),
.Y(n_4583)
);

INVx1_ASAP7_75t_L g4584 ( 
.A(n_4512),
.Y(n_4584)
);

INVx1_ASAP7_75t_L g4585 ( 
.A(n_4517),
.Y(n_4585)
);

NAND2xp5_ASAP7_75t_L g4586 ( 
.A(n_4473),
.B(n_628),
.Y(n_4586)
);

OR2x2_ASAP7_75t_L g4587 ( 
.A(n_4550),
.B(n_271),
.Y(n_4587)
);

INVx2_ASAP7_75t_L g4588 ( 
.A(n_4486),
.Y(n_4588)
);

INVx1_ASAP7_75t_L g4589 ( 
.A(n_4518),
.Y(n_4589)
);

OR2x2_ASAP7_75t_L g4590 ( 
.A(n_4558),
.B(n_272),
.Y(n_4590)
);

INVx1_ASAP7_75t_L g4591 ( 
.A(n_4535),
.Y(n_4591)
);

AND2x4_ASAP7_75t_L g4592 ( 
.A(n_4521),
.B(n_629),
.Y(n_4592)
);

AND2x4_ASAP7_75t_L g4593 ( 
.A(n_4521),
.B(n_629),
.Y(n_4593)
);

INVx1_ASAP7_75t_L g4594 ( 
.A(n_4536),
.Y(n_4594)
);

AND2x2_ASAP7_75t_L g4595 ( 
.A(n_4524),
.B(n_274),
.Y(n_4595)
);

AND2x2_ASAP7_75t_L g4596 ( 
.A(n_4556),
.B(n_275),
.Y(n_4596)
);

INVx1_ASAP7_75t_SL g4597 ( 
.A(n_4542),
.Y(n_4597)
);

AND2x2_ASAP7_75t_L g4598 ( 
.A(n_4546),
.B(n_276),
.Y(n_4598)
);

NAND2xp5_ASAP7_75t_L g4599 ( 
.A(n_4469),
.B(n_630),
.Y(n_4599)
);

INVx4_ASAP7_75t_L g4600 ( 
.A(n_4503),
.Y(n_4600)
);

INVx2_ASAP7_75t_L g4601 ( 
.A(n_4544),
.Y(n_4601)
);

NAND2xp5_ASAP7_75t_L g4602 ( 
.A(n_4484),
.B(n_631),
.Y(n_4602)
);

INVx1_ASAP7_75t_L g4603 ( 
.A(n_4541),
.Y(n_4603)
);

INVxp67_ASAP7_75t_SL g4604 ( 
.A(n_4467),
.Y(n_4604)
);

NOR2xp33_ASAP7_75t_L g4605 ( 
.A(n_4503),
.B(n_632),
.Y(n_4605)
);

AND2x4_ASAP7_75t_L g4606 ( 
.A(n_4490),
.B(n_632),
.Y(n_4606)
);

INVx1_ASAP7_75t_L g4607 ( 
.A(n_4501),
.Y(n_4607)
);

INVx1_ASAP7_75t_L g4608 ( 
.A(n_4551),
.Y(n_4608)
);

BUFx3_ASAP7_75t_L g4609 ( 
.A(n_4526),
.Y(n_4609)
);

NAND2xp5_ASAP7_75t_L g4610 ( 
.A(n_4573),
.B(n_4577),
.Y(n_4610)
);

NAND2xp5_ASAP7_75t_L g4611 ( 
.A(n_4525),
.B(n_633),
.Y(n_4611)
);

INVx1_ASAP7_75t_SL g4612 ( 
.A(n_4523),
.Y(n_4612)
);

INVx2_ASAP7_75t_L g4613 ( 
.A(n_4493),
.Y(n_4613)
);

NAND2xp5_ASAP7_75t_L g4614 ( 
.A(n_4494),
.B(n_634),
.Y(n_4614)
);

CKINVDCx11_ASAP7_75t_R g4615 ( 
.A(n_4560),
.Y(n_4615)
);

AND2x2_ASAP7_75t_L g4616 ( 
.A(n_4534),
.B(n_4475),
.Y(n_4616)
);

INVxp67_ASAP7_75t_SL g4617 ( 
.A(n_4566),
.Y(n_4617)
);

AND2x2_ASAP7_75t_L g4618 ( 
.A(n_4549),
.B(n_277),
.Y(n_4618)
);

HB1xp67_ASAP7_75t_L g4619 ( 
.A(n_4474),
.Y(n_4619)
);

INVx2_ASAP7_75t_L g4620 ( 
.A(n_4491),
.Y(n_4620)
);

NAND2xp5_ASAP7_75t_L g4621 ( 
.A(n_4516),
.B(n_635),
.Y(n_4621)
);

AND2x2_ASAP7_75t_L g4622 ( 
.A(n_4554),
.B(n_278),
.Y(n_4622)
);

AND2x4_ASAP7_75t_L g4623 ( 
.A(n_4504),
.B(n_635),
.Y(n_4623)
);

INVx1_ASAP7_75t_L g4624 ( 
.A(n_4520),
.Y(n_4624)
);

INVx1_ASAP7_75t_L g4625 ( 
.A(n_4520),
.Y(n_4625)
);

AND2x2_ASAP7_75t_L g4626 ( 
.A(n_4564),
.B(n_4574),
.Y(n_4626)
);

AND2x2_ASAP7_75t_L g4627 ( 
.A(n_4575),
.B(n_278),
.Y(n_4627)
);

HB1xp67_ASAP7_75t_L g4628 ( 
.A(n_4474),
.Y(n_4628)
);

INVx2_ASAP7_75t_L g4629 ( 
.A(n_4513),
.Y(n_4629)
);

INVxp67_ASAP7_75t_L g4630 ( 
.A(n_4548),
.Y(n_4630)
);

NAND2xp5_ASAP7_75t_L g4631 ( 
.A(n_4537),
.B(n_637),
.Y(n_4631)
);

NAND2xp5_ASAP7_75t_L g4632 ( 
.A(n_4530),
.B(n_638),
.Y(n_4632)
);

CKINVDCx20_ASAP7_75t_R g4633 ( 
.A(n_4562),
.Y(n_4633)
);

INVx1_ASAP7_75t_L g4634 ( 
.A(n_4522),
.Y(n_4634)
);

NOR2xp33_ASAP7_75t_L g4635 ( 
.A(n_4477),
.B(n_638),
.Y(n_4635)
);

INVx2_ASAP7_75t_L g4636 ( 
.A(n_4514),
.Y(n_4636)
);

INVx1_ASAP7_75t_L g4637 ( 
.A(n_4500),
.Y(n_4637)
);

AND2x4_ASAP7_75t_L g4638 ( 
.A(n_4527),
.B(n_639),
.Y(n_4638)
);

AND2x2_ASAP7_75t_L g4639 ( 
.A(n_4548),
.B(n_279),
.Y(n_4639)
);

AND2x2_ASAP7_75t_L g4640 ( 
.A(n_4480),
.B(n_279),
.Y(n_4640)
);

INVx1_ASAP7_75t_L g4641 ( 
.A(n_4529),
.Y(n_4641)
);

INVx2_ASAP7_75t_L g4642 ( 
.A(n_4483),
.Y(n_4642)
);

NAND2xp5_ASAP7_75t_L g4643 ( 
.A(n_4479),
.B(n_640),
.Y(n_4643)
);

AND2x2_ASAP7_75t_L g4644 ( 
.A(n_4547),
.B(n_279),
.Y(n_4644)
);

INVx1_ASAP7_75t_L g4645 ( 
.A(n_4571),
.Y(n_4645)
);

INVx2_ASAP7_75t_SL g4646 ( 
.A(n_4515),
.Y(n_4646)
);

NAND2xp5_ASAP7_75t_L g4647 ( 
.A(n_4510),
.B(n_641),
.Y(n_4647)
);

NAND2xp5_ASAP7_75t_L g4648 ( 
.A(n_4496),
.B(n_641),
.Y(n_4648)
);

NAND2xp5_ASAP7_75t_L g4649 ( 
.A(n_4497),
.B(n_642),
.Y(n_4649)
);

INVx3_ASAP7_75t_L g4650 ( 
.A(n_4545),
.Y(n_4650)
);

AND2x2_ASAP7_75t_L g4651 ( 
.A(n_4485),
.B(n_280),
.Y(n_4651)
);

INVx1_ASAP7_75t_L g4652 ( 
.A(n_4507),
.Y(n_4652)
);

OR2x2_ASAP7_75t_L g4653 ( 
.A(n_4508),
.B(n_281),
.Y(n_4653)
);

AND2x4_ASAP7_75t_SL g4654 ( 
.A(n_4498),
.B(n_4531),
.Y(n_4654)
);

AND2x2_ASAP7_75t_L g4655 ( 
.A(n_4539),
.B(n_281),
.Y(n_4655)
);

AND2x4_ASAP7_75t_L g4656 ( 
.A(n_4470),
.B(n_642),
.Y(n_4656)
);

AOI22xp33_ASAP7_75t_SL g4657 ( 
.A1(n_4553),
.A2(n_4570),
.B1(n_4569),
.B2(n_4471),
.Y(n_4657)
);

NAND2xp5_ASAP7_75t_L g4658 ( 
.A(n_4476),
.B(n_643),
.Y(n_4658)
);

INVx1_ASAP7_75t_L g4659 ( 
.A(n_4519),
.Y(n_4659)
);

CKINVDCx20_ASAP7_75t_R g4660 ( 
.A(n_4464),
.Y(n_4660)
);

AOI22xp33_ASAP7_75t_L g4661 ( 
.A1(n_4568),
.A2(n_644),
.B1(n_645),
.B2(n_643),
.Y(n_4661)
);

NAND2xp5_ASAP7_75t_L g4662 ( 
.A(n_4468),
.B(n_644),
.Y(n_4662)
);

HB1xp67_ASAP7_75t_L g4663 ( 
.A(n_4538),
.Y(n_4663)
);

INVx2_ASAP7_75t_L g4664 ( 
.A(n_4482),
.Y(n_4664)
);

INVx2_ASAP7_75t_L g4665 ( 
.A(n_4488),
.Y(n_4665)
);

NAND2xp5_ASAP7_75t_L g4666 ( 
.A(n_4543),
.B(n_646),
.Y(n_4666)
);

INVx2_ASAP7_75t_L g4667 ( 
.A(n_4487),
.Y(n_4667)
);

AND2x4_ASAP7_75t_L g4668 ( 
.A(n_4499),
.B(n_647),
.Y(n_4668)
);

AND2x4_ASAP7_75t_L g4669 ( 
.A(n_4533),
.B(n_647),
.Y(n_4669)
);

HB1xp67_ASAP7_75t_L g4670 ( 
.A(n_4563),
.Y(n_4670)
);

NAND2xp5_ASAP7_75t_L g4671 ( 
.A(n_4555),
.B(n_648),
.Y(n_4671)
);

NAND2x1_ASAP7_75t_L g4672 ( 
.A(n_4495),
.B(n_284),
.Y(n_4672)
);

INVx1_ASAP7_75t_L g4673 ( 
.A(n_4492),
.Y(n_4673)
);

OR2x2_ASAP7_75t_L g4674 ( 
.A(n_4565),
.B(n_284),
.Y(n_4674)
);

AND2x2_ASAP7_75t_L g4675 ( 
.A(n_4505),
.B(n_285),
.Y(n_4675)
);

AND2x2_ASAP7_75t_L g4676 ( 
.A(n_4511),
.B(n_285),
.Y(n_4676)
);

INVx2_ASAP7_75t_L g4677 ( 
.A(n_4478),
.Y(n_4677)
);

OAI222xp33_ASAP7_75t_L g4678 ( 
.A1(n_4572),
.A2(n_4465),
.B1(n_4576),
.B2(n_4567),
.C1(n_4557),
.C2(n_4559),
.Y(n_4678)
);

INVx1_ASAP7_75t_L g4679 ( 
.A(n_4528),
.Y(n_4679)
);

AND2x2_ASAP7_75t_L g4680 ( 
.A(n_4502),
.B(n_286),
.Y(n_4680)
);

BUFx3_ASAP7_75t_L g4681 ( 
.A(n_4466),
.Y(n_4681)
);

AND2x4_ASAP7_75t_L g4682 ( 
.A(n_4506),
.B(n_650),
.Y(n_4682)
);

AND2x2_ASAP7_75t_L g4683 ( 
.A(n_4472),
.B(n_287),
.Y(n_4683)
);

AND2x2_ASAP7_75t_L g4684 ( 
.A(n_4489),
.B(n_287),
.Y(n_4684)
);

INVx1_ASAP7_75t_L g4685 ( 
.A(n_4509),
.Y(n_4685)
);

INVx1_ASAP7_75t_L g4686 ( 
.A(n_4509),
.Y(n_4686)
);

AND2x2_ASAP7_75t_L g4687 ( 
.A(n_4489),
.B(n_288),
.Y(n_4687)
);

AND2x2_ASAP7_75t_L g4688 ( 
.A(n_4489),
.B(n_288),
.Y(n_4688)
);

INVx1_ASAP7_75t_L g4689 ( 
.A(n_4509),
.Y(n_4689)
);

INVxp67_ASAP7_75t_L g4690 ( 
.A(n_4552),
.Y(n_4690)
);

OR2x6_ASAP7_75t_L g4691 ( 
.A(n_4556),
.B(n_653),
.Y(n_4691)
);

NAND2xp5_ASAP7_75t_L g4692 ( 
.A(n_4481),
.B(n_653),
.Y(n_4692)
);

INVx2_ASAP7_75t_SL g4693 ( 
.A(n_4503),
.Y(n_4693)
);

AND2x2_ASAP7_75t_L g4694 ( 
.A(n_4489),
.B(n_289),
.Y(n_4694)
);

AND2x2_ASAP7_75t_L g4695 ( 
.A(n_4489),
.B(n_289),
.Y(n_4695)
);

NAND2xp5_ASAP7_75t_L g4696 ( 
.A(n_4481),
.B(n_654),
.Y(n_4696)
);

HB1xp67_ASAP7_75t_L g4697 ( 
.A(n_4532),
.Y(n_4697)
);

INVx3_ASAP7_75t_L g4698 ( 
.A(n_4503),
.Y(n_4698)
);

BUFx3_ASAP7_75t_L g4699 ( 
.A(n_4526),
.Y(n_4699)
);

NAND2xp5_ASAP7_75t_L g4700 ( 
.A(n_4481),
.B(n_654),
.Y(n_4700)
);

INVx1_ASAP7_75t_L g4701 ( 
.A(n_4509),
.Y(n_4701)
);

AND2x2_ASAP7_75t_L g4702 ( 
.A(n_4489),
.B(n_291),
.Y(n_4702)
);

INVx1_ASAP7_75t_L g4703 ( 
.A(n_4509),
.Y(n_4703)
);

AND2x2_ASAP7_75t_L g4704 ( 
.A(n_4489),
.B(n_292),
.Y(n_4704)
);

INVx2_ASAP7_75t_L g4705 ( 
.A(n_4532),
.Y(n_4705)
);

INVx1_ASAP7_75t_L g4706 ( 
.A(n_4509),
.Y(n_4706)
);

INVx1_ASAP7_75t_L g4707 ( 
.A(n_4509),
.Y(n_4707)
);

INVx1_ASAP7_75t_L g4708 ( 
.A(n_4509),
.Y(n_4708)
);

INVx2_ASAP7_75t_L g4709 ( 
.A(n_4532),
.Y(n_4709)
);

INVx2_ASAP7_75t_L g4710 ( 
.A(n_4588),
.Y(n_4710)
);

INVx1_ASAP7_75t_L g4711 ( 
.A(n_4580),
.Y(n_4711)
);

NAND2xp5_ASAP7_75t_L g4712 ( 
.A(n_4604),
.B(n_655),
.Y(n_4712)
);

INVx1_ASAP7_75t_L g4713 ( 
.A(n_4584),
.Y(n_4713)
);

BUFx2_ASAP7_75t_L g4714 ( 
.A(n_4697),
.Y(n_4714)
);

AND2x2_ASAP7_75t_L g4715 ( 
.A(n_4617),
.B(n_292),
.Y(n_4715)
);

AND2x4_ASAP7_75t_L g4716 ( 
.A(n_4690),
.B(n_4693),
.Y(n_4716)
);

INVx1_ASAP7_75t_L g4717 ( 
.A(n_4585),
.Y(n_4717)
);

NAND2xp5_ASAP7_75t_L g4718 ( 
.A(n_4629),
.B(n_656),
.Y(n_4718)
);

NAND2xp5_ASAP7_75t_L g4719 ( 
.A(n_4642),
.B(n_657),
.Y(n_4719)
);

NAND2xp5_ASAP7_75t_L g4720 ( 
.A(n_4641),
.B(n_657),
.Y(n_4720)
);

HB1xp67_ASAP7_75t_L g4721 ( 
.A(n_4619),
.Y(n_4721)
);

NOR2xp33_ASAP7_75t_L g4722 ( 
.A(n_4600),
.B(n_658),
.Y(n_4722)
);

OAI221xp5_ASAP7_75t_L g4723 ( 
.A1(n_4657),
.A2(n_295),
.B1(n_293),
.B2(n_294),
.C(n_296),
.Y(n_4723)
);

HB1xp67_ASAP7_75t_L g4724 ( 
.A(n_4628),
.Y(n_4724)
);

AND2x2_ASAP7_75t_L g4725 ( 
.A(n_4579),
.B(n_4705),
.Y(n_4725)
);

OAI21xp5_ASAP7_75t_L g4726 ( 
.A1(n_4663),
.A2(n_293),
.B(n_294),
.Y(n_4726)
);

AND2x2_ASAP7_75t_L g4727 ( 
.A(n_4709),
.B(n_295),
.Y(n_4727)
);

AND2x2_ASAP7_75t_L g4728 ( 
.A(n_4620),
.B(n_296),
.Y(n_4728)
);

AND2x2_ASAP7_75t_L g4729 ( 
.A(n_4636),
.B(n_297),
.Y(n_4729)
);

NAND2xp5_ASAP7_75t_L g4730 ( 
.A(n_4645),
.B(n_4634),
.Y(n_4730)
);

AOI22xp33_ASAP7_75t_L g4731 ( 
.A1(n_4667),
.A2(n_661),
.B1(n_662),
.B2(n_659),
.Y(n_4731)
);

INVx1_ASAP7_75t_L g4732 ( 
.A(n_4589),
.Y(n_4732)
);

INVxp33_ASAP7_75t_SL g4733 ( 
.A(n_4615),
.Y(n_4733)
);

INVx1_ASAP7_75t_SL g4734 ( 
.A(n_4612),
.Y(n_4734)
);

INVx1_ASAP7_75t_L g4735 ( 
.A(n_4591),
.Y(n_4735)
);

INVxp67_ASAP7_75t_L g4736 ( 
.A(n_4582),
.Y(n_4736)
);

INVx2_ASAP7_75t_L g4737 ( 
.A(n_4613),
.Y(n_4737)
);

OAI221xp5_ASAP7_75t_SL g4738 ( 
.A1(n_4661),
.A2(n_301),
.B1(n_299),
.B2(n_300),
.C(n_302),
.Y(n_4738)
);

OR2x2_ASAP7_75t_L g4739 ( 
.A(n_4637),
.B(n_300),
.Y(n_4739)
);

AND2x2_ASAP7_75t_L g4740 ( 
.A(n_4616),
.B(n_301),
.Y(n_4740)
);

INVx1_ASAP7_75t_L g4741 ( 
.A(n_4594),
.Y(n_4741)
);

INVx1_ASAP7_75t_L g4742 ( 
.A(n_4607),
.Y(n_4742)
);

INVx1_ASAP7_75t_L g4743 ( 
.A(n_4608),
.Y(n_4743)
);

AND2x2_ASAP7_75t_L g4744 ( 
.A(n_4626),
.B(n_301),
.Y(n_4744)
);

NAND2xp5_ASAP7_75t_L g4745 ( 
.A(n_4650),
.B(n_663),
.Y(n_4745)
);

AOI22xp33_ASAP7_75t_L g4746 ( 
.A1(n_4664),
.A2(n_665),
.B1(n_666),
.B2(n_664),
.Y(n_4746)
);

OR2x2_ASAP7_75t_L g4747 ( 
.A(n_4624),
.B(n_302),
.Y(n_4747)
);

HB1xp67_ASAP7_75t_L g4748 ( 
.A(n_4625),
.Y(n_4748)
);

INVx1_ASAP7_75t_L g4749 ( 
.A(n_4685),
.Y(n_4749)
);

INVx1_ASAP7_75t_L g4750 ( 
.A(n_4686),
.Y(n_4750)
);

NAND2xp5_ASAP7_75t_L g4751 ( 
.A(n_4581),
.B(n_666),
.Y(n_4751)
);

INVx2_ASAP7_75t_L g4752 ( 
.A(n_4601),
.Y(n_4752)
);

OR2x2_ASAP7_75t_L g4753 ( 
.A(n_4610),
.B(n_303),
.Y(n_4753)
);

INVx1_ASAP7_75t_L g4754 ( 
.A(n_4689),
.Y(n_4754)
);

NAND2xp5_ASAP7_75t_L g4755 ( 
.A(n_4652),
.B(n_667),
.Y(n_4755)
);

AND2x2_ASAP7_75t_L g4756 ( 
.A(n_4698),
.B(n_303),
.Y(n_4756)
);

INVx1_ASAP7_75t_L g4757 ( 
.A(n_4701),
.Y(n_4757)
);

NOR2xp67_ASAP7_75t_L g4758 ( 
.A(n_4646),
.B(n_304),
.Y(n_4758)
);

OR2x2_ASAP7_75t_L g4759 ( 
.A(n_4587),
.B(n_4590),
.Y(n_4759)
);

NAND3xp33_ASAP7_75t_L g4760 ( 
.A(n_4672),
.B(n_4647),
.C(n_4662),
.Y(n_4760)
);

AND2x2_ASAP7_75t_L g4761 ( 
.A(n_4684),
.B(n_304),
.Y(n_4761)
);

AND2x2_ASAP7_75t_L g4762 ( 
.A(n_4687),
.B(n_305),
.Y(n_4762)
);

OR2x2_ASAP7_75t_L g4763 ( 
.A(n_4603),
.B(n_305),
.Y(n_4763)
);

NOR2x1_ASAP7_75t_L g4764 ( 
.A(n_4609),
.B(n_4699),
.Y(n_4764)
);

AND2x2_ASAP7_75t_L g4765 ( 
.A(n_4688),
.B(n_305),
.Y(n_4765)
);

AND2x2_ASAP7_75t_L g4766 ( 
.A(n_4694),
.B(n_306),
.Y(n_4766)
);

HB1xp67_ASAP7_75t_L g4767 ( 
.A(n_4703),
.Y(n_4767)
);

HB1xp67_ASAP7_75t_L g4768 ( 
.A(n_4706),
.Y(n_4768)
);

AND2x2_ASAP7_75t_L g4769 ( 
.A(n_4695),
.B(n_306),
.Y(n_4769)
);

OR2x6_ASAP7_75t_L g4770 ( 
.A(n_4691),
.B(n_668),
.Y(n_4770)
);

INVx1_ASAP7_75t_L g4771 ( 
.A(n_4707),
.Y(n_4771)
);

INVx1_ASAP7_75t_L g4772 ( 
.A(n_4708),
.Y(n_4772)
);

NAND2xp5_ASAP7_75t_SL g4773 ( 
.A(n_4597),
.B(n_308),
.Y(n_4773)
);

NAND2xp5_ASAP7_75t_L g4774 ( 
.A(n_4639),
.B(n_668),
.Y(n_4774)
);

INVx2_ASAP7_75t_L g4775 ( 
.A(n_4606),
.Y(n_4775)
);

INVx1_ASAP7_75t_L g4776 ( 
.A(n_4611),
.Y(n_4776)
);

NAND3xp33_ASAP7_75t_L g4777 ( 
.A(n_4643),
.B(n_309),
.C(n_311),
.Y(n_4777)
);

OR2x2_ASAP7_75t_L g4778 ( 
.A(n_4586),
.B(n_309),
.Y(n_4778)
);

OR2x2_ASAP7_75t_L g4779 ( 
.A(n_4673),
.B(n_311),
.Y(n_4779)
);

OR2x2_ASAP7_75t_L g4780 ( 
.A(n_4599),
.B(n_312),
.Y(n_4780)
);

INVx2_ASAP7_75t_L g4781 ( 
.A(n_4592),
.Y(n_4781)
);

OR2x2_ASAP7_75t_L g4782 ( 
.A(n_4602),
.B(n_312),
.Y(n_4782)
);

INVx2_ASAP7_75t_L g4783 ( 
.A(n_4593),
.Y(n_4783)
);

AND2x4_ASAP7_75t_SL g4784 ( 
.A(n_4633),
.B(n_313),
.Y(n_4784)
);

INVxp67_ASAP7_75t_L g4785 ( 
.A(n_4670),
.Y(n_4785)
);

INVx2_ASAP7_75t_L g4786 ( 
.A(n_4596),
.Y(n_4786)
);

NOR3xp33_ASAP7_75t_L g4787 ( 
.A(n_4678),
.B(n_314),
.C(n_315),
.Y(n_4787)
);

INVx1_ASAP7_75t_L g4788 ( 
.A(n_4614),
.Y(n_4788)
);

NAND2xp5_ASAP7_75t_L g4789 ( 
.A(n_4665),
.B(n_670),
.Y(n_4789)
);

AND2x2_ASAP7_75t_L g4790 ( 
.A(n_4702),
.B(n_4704),
.Y(n_4790)
);

INVxp67_ASAP7_75t_SL g4791 ( 
.A(n_4621),
.Y(n_4791)
);

INVxp67_ASAP7_75t_SL g4792 ( 
.A(n_4677),
.Y(n_4792)
);

INVx2_ASAP7_75t_L g4793 ( 
.A(n_4598),
.Y(n_4793)
);

NAND2xp5_ASAP7_75t_L g4794 ( 
.A(n_4595),
.B(n_672),
.Y(n_4794)
);

OR2x2_ASAP7_75t_L g4795 ( 
.A(n_4583),
.B(n_315),
.Y(n_4795)
);

NOR2x1_ASAP7_75t_L g4796 ( 
.A(n_4692),
.B(n_4696),
.Y(n_4796)
);

OR2x2_ASAP7_75t_L g4797 ( 
.A(n_4700),
.B(n_316),
.Y(n_4797)
);

INVx2_ASAP7_75t_L g4798 ( 
.A(n_4638),
.Y(n_4798)
);

NAND2xp5_ASAP7_75t_L g4799 ( 
.A(n_4659),
.B(n_673),
.Y(n_4799)
);

INVx1_ASAP7_75t_L g4800 ( 
.A(n_4631),
.Y(n_4800)
);

NAND2xp5_ASAP7_75t_L g4801 ( 
.A(n_4679),
.B(n_674),
.Y(n_4801)
);

AND2x2_ASAP7_75t_L g4802 ( 
.A(n_4644),
.B(n_316),
.Y(n_4802)
);

AND2x4_ASAP7_75t_L g4803 ( 
.A(n_4656),
.B(n_316),
.Y(n_4803)
);

AND2x2_ASAP7_75t_L g4804 ( 
.A(n_4618),
.B(n_317),
.Y(n_4804)
);

AOI211xp5_ASAP7_75t_L g4805 ( 
.A1(n_4655),
.A2(n_319),
.B(n_320),
.C(n_318),
.Y(n_4805)
);

NAND2xp5_ASAP7_75t_SL g4806 ( 
.A(n_4668),
.B(n_317),
.Y(n_4806)
);

AND2x2_ASAP7_75t_L g4807 ( 
.A(n_4622),
.B(n_317),
.Y(n_4807)
);

INVx1_ASAP7_75t_L g4808 ( 
.A(n_4632),
.Y(n_4808)
);

INVx1_ASAP7_75t_L g4809 ( 
.A(n_4648),
.Y(n_4809)
);

AND2x2_ASAP7_75t_L g4810 ( 
.A(n_4623),
.B(n_319),
.Y(n_4810)
);

OR2x2_ASAP7_75t_L g4811 ( 
.A(n_4681),
.B(n_319),
.Y(n_4811)
);

OAI221xp5_ASAP7_75t_SL g4812 ( 
.A1(n_4649),
.A2(n_322),
.B1(n_320),
.B2(n_321),
.C(n_323),
.Y(n_4812)
);

INVxp67_ASAP7_75t_L g4813 ( 
.A(n_4605),
.Y(n_4813)
);

OR2x2_ASAP7_75t_L g4814 ( 
.A(n_4653),
.B(n_4674),
.Y(n_4814)
);

INVx1_ASAP7_75t_L g4815 ( 
.A(n_4627),
.Y(n_4815)
);

AOI221xp5_ASAP7_75t_L g4816 ( 
.A1(n_4675),
.A2(n_323),
.B1(n_321),
.B2(n_322),
.C(n_324),
.Y(n_4816)
);

NAND2xp5_ASAP7_75t_L g4817 ( 
.A(n_4651),
.B(n_674),
.Y(n_4817)
);

INVx1_ASAP7_75t_L g4818 ( 
.A(n_4658),
.Y(n_4818)
);

OAI21xp5_ASAP7_75t_SL g4819 ( 
.A1(n_4654),
.A2(n_323),
.B(n_324),
.Y(n_4819)
);

INVx1_ASAP7_75t_L g4820 ( 
.A(n_4666),
.Y(n_4820)
);

INVx4_ASAP7_75t_L g4821 ( 
.A(n_4640),
.Y(n_4821)
);

OR2x6_ASAP7_75t_L g4822 ( 
.A(n_4671),
.B(n_4682),
.Y(n_4822)
);

AND2x2_ASAP7_75t_L g4823 ( 
.A(n_4680),
.B(n_329),
.Y(n_4823)
);

NOR2xp33_ASAP7_75t_L g4824 ( 
.A(n_4676),
.B(n_675),
.Y(n_4824)
);

INVx1_ASAP7_75t_L g4825 ( 
.A(n_4683),
.Y(n_4825)
);

INVx2_ASAP7_75t_L g4826 ( 
.A(n_4669),
.Y(n_4826)
);

INVx1_ASAP7_75t_L g4827 ( 
.A(n_4580),
.Y(n_4827)
);

INVx1_ASAP7_75t_L g4828 ( 
.A(n_4580),
.Y(n_4828)
);

NAND2x1p5_ASAP7_75t_L g4829 ( 
.A(n_4578),
.B(n_330),
.Y(n_4829)
);

NAND2x1p5_ASAP7_75t_L g4830 ( 
.A(n_4578),
.B(n_330),
.Y(n_4830)
);

INVx1_ASAP7_75t_L g4831 ( 
.A(n_4580),
.Y(n_4831)
);

NAND2xp5_ASAP7_75t_L g4832 ( 
.A(n_4604),
.B(n_676),
.Y(n_4832)
);

INVx2_ASAP7_75t_L g4833 ( 
.A(n_4588),
.Y(n_4833)
);

INVx2_ASAP7_75t_L g4834 ( 
.A(n_4588),
.Y(n_4834)
);

INVx2_ASAP7_75t_L g4835 ( 
.A(n_4588),
.Y(n_4835)
);

AND2x4_ASAP7_75t_L g4836 ( 
.A(n_4690),
.B(n_331),
.Y(n_4836)
);

AND2x2_ASAP7_75t_L g4837 ( 
.A(n_4604),
.B(n_331),
.Y(n_4837)
);

NAND2xp5_ASAP7_75t_SL g4838 ( 
.A(n_4597),
.B(n_332),
.Y(n_4838)
);

HB1xp67_ASAP7_75t_L g4839 ( 
.A(n_4619),
.Y(n_4839)
);

NAND2xp5_ASAP7_75t_L g4840 ( 
.A(n_4604),
.B(n_677),
.Y(n_4840)
);

NAND2xp5_ASAP7_75t_L g4841 ( 
.A(n_4604),
.B(n_678),
.Y(n_4841)
);

AND2x2_ASAP7_75t_L g4842 ( 
.A(n_4604),
.B(n_333),
.Y(n_4842)
);

NAND2xp5_ASAP7_75t_L g4843 ( 
.A(n_4604),
.B(n_678),
.Y(n_4843)
);

AND2x2_ASAP7_75t_L g4844 ( 
.A(n_4604),
.B(n_335),
.Y(n_4844)
);

AND2x2_ASAP7_75t_L g4845 ( 
.A(n_4604),
.B(n_335),
.Y(n_4845)
);

AND2x2_ASAP7_75t_L g4846 ( 
.A(n_4604),
.B(n_336),
.Y(n_4846)
);

INVxp67_ASAP7_75t_L g4847 ( 
.A(n_4582),
.Y(n_4847)
);

INVx1_ASAP7_75t_L g4848 ( 
.A(n_4580),
.Y(n_4848)
);

INVx2_ASAP7_75t_L g4849 ( 
.A(n_4588),
.Y(n_4849)
);

NAND2xp33_ASAP7_75t_SL g4850 ( 
.A(n_4660),
.B(n_337),
.Y(n_4850)
);

AND2x2_ASAP7_75t_L g4851 ( 
.A(n_4604),
.B(n_337),
.Y(n_4851)
);

AND2x2_ASAP7_75t_L g4852 ( 
.A(n_4604),
.B(n_338),
.Y(n_4852)
);

NAND2xp33_ASAP7_75t_SL g4853 ( 
.A(n_4660),
.B(n_338),
.Y(n_4853)
);

NOR3xp33_ASAP7_75t_L g4854 ( 
.A(n_4635),
.B(n_339),
.C(n_340),
.Y(n_4854)
);

NOR2xp33_ASAP7_75t_L g4855 ( 
.A(n_4600),
.B(n_679),
.Y(n_4855)
);

AOI22xp33_ASAP7_75t_L g4856 ( 
.A1(n_4663),
.A2(n_682),
.B1(n_683),
.B2(n_681),
.Y(n_4856)
);

INVx1_ASAP7_75t_L g4857 ( 
.A(n_4580),
.Y(n_4857)
);

INVx2_ASAP7_75t_L g4858 ( 
.A(n_4588),
.Y(n_4858)
);

NAND2xp5_ASAP7_75t_L g4859 ( 
.A(n_4604),
.B(n_681),
.Y(n_4859)
);

NAND2xp5_ASAP7_75t_L g4860 ( 
.A(n_4604),
.B(n_682),
.Y(n_4860)
);

INVx1_ASAP7_75t_L g4861 ( 
.A(n_4580),
.Y(n_4861)
);

OA21x2_ASAP7_75t_L g4862 ( 
.A1(n_4630),
.A2(n_340),
.B(n_341),
.Y(n_4862)
);

AND2x2_ASAP7_75t_L g4863 ( 
.A(n_4604),
.B(n_341),
.Y(n_4863)
);

OR2x2_ASAP7_75t_L g4864 ( 
.A(n_4604),
.B(n_342),
.Y(n_4864)
);

OAI21xp5_ASAP7_75t_SL g4865 ( 
.A1(n_4678),
.A2(n_343),
.B(n_344),
.Y(n_4865)
);

AND2x2_ASAP7_75t_L g4866 ( 
.A(n_4604),
.B(n_343),
.Y(n_4866)
);

NOR2x1_ASAP7_75t_L g4867 ( 
.A(n_4600),
.B(n_343),
.Y(n_4867)
);

AND2x2_ASAP7_75t_L g4868 ( 
.A(n_4604),
.B(n_344),
.Y(n_4868)
);

INVx2_ASAP7_75t_L g4869 ( 
.A(n_4588),
.Y(n_4869)
);

INVx1_ASAP7_75t_L g4870 ( 
.A(n_4580),
.Y(n_4870)
);

NAND2xp5_ASAP7_75t_L g4871 ( 
.A(n_4604),
.B(n_684),
.Y(n_4871)
);

INVxp67_ASAP7_75t_SL g4872 ( 
.A(n_4736),
.Y(n_4872)
);

AOI21xp5_ASAP7_75t_SL g4873 ( 
.A1(n_4806),
.A2(n_345),
.B(n_346),
.Y(n_4873)
);

INVx1_ASAP7_75t_L g4874 ( 
.A(n_4767),
.Y(n_4874)
);

NAND2xp5_ASAP7_75t_L g4875 ( 
.A(n_4791),
.B(n_346),
.Y(n_4875)
);

O2A1O1Ixp33_ASAP7_75t_L g4876 ( 
.A1(n_4865),
.A2(n_349),
.B(n_347),
.C(n_348),
.Y(n_4876)
);

BUFx2_ASAP7_75t_SL g4877 ( 
.A(n_4758),
.Y(n_4877)
);

OAI321xp33_ASAP7_75t_L g4878 ( 
.A1(n_4723),
.A2(n_372),
.A3(n_355),
.B1(n_363),
.B2(n_347),
.C(n_349),
.Y(n_4878)
);

INVx1_ASAP7_75t_L g4879 ( 
.A(n_4768),
.Y(n_4879)
);

AND2x2_ASAP7_75t_L g4880 ( 
.A(n_4764),
.B(n_348),
.Y(n_4880)
);

NAND3xp33_ASAP7_75t_L g4881 ( 
.A(n_4787),
.B(n_350),
.C(n_351),
.Y(n_4881)
);

AND2x4_ASAP7_75t_L g4882 ( 
.A(n_4716),
.B(n_350),
.Y(n_4882)
);

INVx1_ASAP7_75t_L g4883 ( 
.A(n_4748),
.Y(n_4883)
);

HB1xp67_ASAP7_75t_L g4884 ( 
.A(n_4721),
.Y(n_4884)
);

AOI22xp33_ASAP7_75t_L g4885 ( 
.A1(n_4854),
.A2(n_353),
.B1(n_351),
.B2(n_352),
.Y(n_4885)
);

NOR2xp33_ASAP7_75t_L g4886 ( 
.A(n_4733),
.B(n_352),
.Y(n_4886)
);

HB1xp67_ASAP7_75t_L g4887 ( 
.A(n_4724),
.Y(n_4887)
);

INVx1_ASAP7_75t_L g4888 ( 
.A(n_4839),
.Y(n_4888)
);

INVx2_ASAP7_75t_L g4889 ( 
.A(n_4714),
.Y(n_4889)
);

NAND2xp5_ASAP7_75t_L g4890 ( 
.A(n_4820),
.B(n_4792),
.Y(n_4890)
);

BUFx3_ASAP7_75t_L g4891 ( 
.A(n_4784),
.Y(n_4891)
);

AOI33xp33_ASAP7_75t_L g4892 ( 
.A1(n_4805),
.A2(n_354),
.A3(n_356),
.B1(n_352),
.B2(n_353),
.B3(n_355),
.Y(n_4892)
);

NAND2xp5_ASAP7_75t_L g4893 ( 
.A(n_4818),
.B(n_353),
.Y(n_4893)
);

AND2x2_ASAP7_75t_L g4894 ( 
.A(n_4725),
.B(n_354),
.Y(n_4894)
);

OAI221xp5_ASAP7_75t_L g4895 ( 
.A1(n_4819),
.A2(n_357),
.B1(n_355),
.B2(n_356),
.C(n_358),
.Y(n_4895)
);

NOR3xp33_ASAP7_75t_SL g4896 ( 
.A(n_4812),
.B(n_4853),
.C(n_4850),
.Y(n_4896)
);

OAI221xp5_ASAP7_75t_L g4897 ( 
.A1(n_4726),
.A2(n_359),
.B1(n_357),
.B2(n_358),
.C(n_360),
.Y(n_4897)
);

OAI221xp5_ASAP7_75t_L g4898 ( 
.A1(n_4847),
.A2(n_360),
.B1(n_357),
.B2(n_359),
.C(n_361),
.Y(n_4898)
);

AOI21xp5_ASAP7_75t_SL g4899 ( 
.A1(n_4770),
.A2(n_4838),
.B(n_4773),
.Y(n_4899)
);

INVx3_ASAP7_75t_L g4900 ( 
.A(n_4821),
.Y(n_4900)
);

AOI31xp33_ASAP7_75t_L g4901 ( 
.A1(n_4867),
.A2(n_364),
.A3(n_362),
.B(n_363),
.Y(n_4901)
);

AOI22xp5_ASAP7_75t_L g4902 ( 
.A1(n_4785),
.A2(n_364),
.B1(n_362),
.B2(n_363),
.Y(n_4902)
);

INVx1_ASAP7_75t_L g4903 ( 
.A(n_4711),
.Y(n_4903)
);

INVx3_ASAP7_75t_L g4904 ( 
.A(n_4734),
.Y(n_4904)
);

OAI211xp5_ASAP7_75t_SL g4905 ( 
.A1(n_4816),
.A2(n_367),
.B(n_365),
.C(n_366),
.Y(n_4905)
);

INVx1_ASAP7_75t_L g4906 ( 
.A(n_4713),
.Y(n_4906)
);

NOR2x1_ASAP7_75t_L g4907 ( 
.A(n_4862),
.B(n_366),
.Y(n_4907)
);

AOI22xp5_ASAP7_75t_L g4908 ( 
.A1(n_4760),
.A2(n_370),
.B1(n_367),
.B2(n_369),
.Y(n_4908)
);

INVx3_ASAP7_75t_L g4909 ( 
.A(n_4781),
.Y(n_4909)
);

AND2x2_ASAP7_75t_L g4910 ( 
.A(n_4809),
.B(n_369),
.Y(n_4910)
);

INVx1_ASAP7_75t_L g4911 ( 
.A(n_4717),
.Y(n_4911)
);

A2O1A1Ixp33_ASAP7_75t_SL g4912 ( 
.A1(n_4722),
.A2(n_372),
.B(n_370),
.C(n_371),
.Y(n_4912)
);

INVxp67_ASAP7_75t_SL g4913 ( 
.A(n_4811),
.Y(n_4913)
);

INVx5_ASAP7_75t_L g4914 ( 
.A(n_4770),
.Y(n_4914)
);

HB1xp67_ASAP7_75t_L g4915 ( 
.A(n_4786),
.Y(n_4915)
);

AND2x2_ASAP7_75t_L g4916 ( 
.A(n_4800),
.B(n_373),
.Y(n_4916)
);

INVx1_ASAP7_75t_L g4917 ( 
.A(n_4732),
.Y(n_4917)
);

INVx1_ASAP7_75t_L g4918 ( 
.A(n_4735),
.Y(n_4918)
);

OAI33xp33_ASAP7_75t_L g4919 ( 
.A1(n_4730),
.A2(n_376),
.A3(n_375),
.B1(n_374),
.B2(n_377),
.B3(n_684),
.Y(n_4919)
);

INVx1_ASAP7_75t_L g4920 ( 
.A(n_4741),
.Y(n_4920)
);

BUFx2_ASAP7_75t_L g4921 ( 
.A(n_4815),
.Y(n_4921)
);

BUFx2_ASAP7_75t_L g4922 ( 
.A(n_4759),
.Y(n_4922)
);

INVx1_ASAP7_75t_L g4923 ( 
.A(n_4742),
.Y(n_4923)
);

OAI33xp33_ASAP7_75t_L g4924 ( 
.A1(n_4745),
.A2(n_689),
.A3(n_692),
.B1(n_686),
.B2(n_688),
.B3(n_690),
.Y(n_4924)
);

INVx1_ASAP7_75t_L g4925 ( 
.A(n_4743),
.Y(n_4925)
);

INVx2_ASAP7_75t_L g4926 ( 
.A(n_4793),
.Y(n_4926)
);

OAI221xp5_ASAP7_75t_L g4927 ( 
.A1(n_4777),
.A2(n_692),
.B1(n_688),
.B2(n_689),
.C(n_693),
.Y(n_4927)
);

AOI33xp33_ASAP7_75t_L g4928 ( 
.A1(n_4856),
.A2(n_696),
.A3(n_698),
.B1(n_694),
.B2(n_695),
.B3(n_697),
.Y(n_4928)
);

AND2x2_ASAP7_75t_L g4929 ( 
.A(n_4808),
.B(n_697),
.Y(n_4929)
);

NAND2xp5_ASAP7_75t_L g4930 ( 
.A(n_4776),
.B(n_698),
.Y(n_4930)
);

NAND3xp33_ASAP7_75t_L g4931 ( 
.A(n_4738),
.B(n_699),
.C(n_700),
.Y(n_4931)
);

AO21x2_ASAP7_75t_L g4932 ( 
.A1(n_4751),
.A2(n_699),
.B(n_701),
.Y(n_4932)
);

INVx5_ASAP7_75t_L g4933 ( 
.A(n_4715),
.Y(n_4933)
);

AOI22xp33_ASAP7_75t_L g4934 ( 
.A1(n_4824),
.A2(n_707),
.B1(n_705),
.B2(n_706),
.Y(n_4934)
);

AOI22xp33_ASAP7_75t_L g4935 ( 
.A1(n_4825),
.A2(n_707),
.B1(n_705),
.B2(n_706),
.Y(n_4935)
);

BUFx2_ASAP7_75t_L g4936 ( 
.A(n_4829),
.Y(n_4936)
);

AND2x2_ASAP7_75t_L g4937 ( 
.A(n_4788),
.B(n_708),
.Y(n_4937)
);

INVx1_ASAP7_75t_L g4938 ( 
.A(n_4749),
.Y(n_4938)
);

INVxp67_ASAP7_75t_L g4939 ( 
.A(n_4747),
.Y(n_4939)
);

INVx1_ASAP7_75t_L g4940 ( 
.A(n_4750),
.Y(n_4940)
);

OAI221xp5_ASAP7_75t_SL g4941 ( 
.A1(n_4731),
.A2(n_4746),
.B1(n_4822),
.B2(n_4814),
.C(n_4712),
.Y(n_4941)
);

OAI221xp5_ASAP7_75t_L g4942 ( 
.A1(n_4813),
.A2(n_712),
.B1(n_710),
.B2(n_711),
.C(n_713),
.Y(n_4942)
);

INVx5_ASAP7_75t_L g4943 ( 
.A(n_4837),
.Y(n_4943)
);

INVx1_ASAP7_75t_L g4944 ( 
.A(n_4754),
.Y(n_4944)
);

INVx1_ASAP7_75t_L g4945 ( 
.A(n_4757),
.Y(n_4945)
);

INVx1_ASAP7_75t_L g4946 ( 
.A(n_4771),
.Y(n_4946)
);

INVxp67_ASAP7_75t_L g4947 ( 
.A(n_4739),
.Y(n_4947)
);

INVx2_ASAP7_75t_L g4948 ( 
.A(n_4737),
.Y(n_4948)
);

OR2x2_ASAP7_75t_L g4949 ( 
.A(n_4753),
.B(n_713),
.Y(n_4949)
);

OAI211xp5_ASAP7_75t_L g4950 ( 
.A1(n_4720),
.A2(n_716),
.B(n_714),
.C(n_715),
.Y(n_4950)
);

INVx1_ASAP7_75t_L g4951 ( 
.A(n_4772),
.Y(n_4951)
);

INVx2_ASAP7_75t_L g4952 ( 
.A(n_4710),
.Y(n_4952)
);

INVx2_ASAP7_75t_L g4953 ( 
.A(n_4833),
.Y(n_4953)
);

AND2x2_ASAP7_75t_L g4954 ( 
.A(n_4775),
.B(n_717),
.Y(n_4954)
);

AND2x2_ASAP7_75t_L g4955 ( 
.A(n_4790),
.B(n_720),
.Y(n_4955)
);

NAND4xp25_ASAP7_75t_L g4956 ( 
.A(n_4796),
.B(n_725),
.C(n_726),
.D(n_724),
.Y(n_4956)
);

INVx1_ASAP7_75t_L g4957 ( 
.A(n_4827),
.Y(n_4957)
);

AND2x2_ASAP7_75t_L g4958 ( 
.A(n_4798),
.B(n_721),
.Y(n_4958)
);

AOI221xp5_ASAP7_75t_L g4959 ( 
.A1(n_4755),
.A2(n_726),
.B1(n_724),
.B2(n_725),
.C(n_728),
.Y(n_4959)
);

OAI221xp5_ASAP7_75t_L g4960 ( 
.A1(n_4822),
.A2(n_730),
.B1(n_728),
.B2(n_729),
.C(n_731),
.Y(n_4960)
);

BUFx2_ASAP7_75t_L g4961 ( 
.A(n_4830),
.Y(n_4961)
);

AOI22xp5_ASAP7_75t_L g4962 ( 
.A1(n_4855),
.A2(n_732),
.B1(n_730),
.B2(n_731),
.Y(n_4962)
);

AND2x2_ASAP7_75t_L g4963 ( 
.A(n_4783),
.B(n_4826),
.Y(n_4963)
);

INVx1_ASAP7_75t_L g4964 ( 
.A(n_4828),
.Y(n_4964)
);

INVx1_ASAP7_75t_L g4965 ( 
.A(n_4831),
.Y(n_4965)
);

OAI22xp5_ASAP7_75t_L g4966 ( 
.A1(n_4719),
.A2(n_4801),
.B1(n_4799),
.B2(n_4832),
.Y(n_4966)
);

INVx4_ASAP7_75t_L g4967 ( 
.A(n_4836),
.Y(n_4967)
);

NAND3xp33_ASAP7_75t_L g4968 ( 
.A(n_4840),
.B(n_4843),
.C(n_4841),
.Y(n_4968)
);

INVx1_ASAP7_75t_L g4969 ( 
.A(n_4848),
.Y(n_4969)
);

AND2x2_ASAP7_75t_L g4970 ( 
.A(n_4727),
.B(n_735),
.Y(n_4970)
);

AOI211xp5_ASAP7_75t_L g4971 ( 
.A1(n_4871),
.A2(n_738),
.B(n_736),
.C(n_737),
.Y(n_4971)
);

INVx1_ASAP7_75t_L g4972 ( 
.A(n_4857),
.Y(n_4972)
);

NAND2xp5_ASAP7_75t_L g4973 ( 
.A(n_4842),
.B(n_738),
.Y(n_4973)
);

INVx1_ASAP7_75t_L g4974 ( 
.A(n_4861),
.Y(n_4974)
);

NOR3xp33_ASAP7_75t_SL g4975 ( 
.A(n_4789),
.B(n_742),
.C(n_743),
.Y(n_4975)
);

OAI33xp33_ASAP7_75t_L g4976 ( 
.A1(n_4859),
.A2(n_747),
.A3(n_749),
.B1(n_745),
.B2(n_746),
.B3(n_748),
.Y(n_4976)
);

INVx2_ASAP7_75t_L g4977 ( 
.A(n_4834),
.Y(n_4977)
);

OAI31xp33_ASAP7_75t_L g4978 ( 
.A1(n_4740),
.A2(n_1619),
.A3(n_1620),
.B(n_1618),
.Y(n_4978)
);

INVx1_ASAP7_75t_L g4979 ( 
.A(n_4870),
.Y(n_4979)
);

OAI221xp5_ASAP7_75t_L g4980 ( 
.A1(n_4860),
.A2(n_752),
.B1(n_750),
.B2(n_751),
.C(n_753),
.Y(n_4980)
);

NAND2xp5_ASAP7_75t_L g4981 ( 
.A(n_4844),
.B(n_750),
.Y(n_4981)
);

NOR2x1_ASAP7_75t_SL g4982 ( 
.A(n_4864),
.B(n_1620),
.Y(n_4982)
);

INVx2_ASAP7_75t_L g4983 ( 
.A(n_4835),
.Y(n_4983)
);

AND2x2_ASAP7_75t_L g4984 ( 
.A(n_4752),
.B(n_752),
.Y(n_4984)
);

INVxp67_ASAP7_75t_L g4985 ( 
.A(n_4779),
.Y(n_4985)
);

INVxp67_ASAP7_75t_L g4986 ( 
.A(n_4763),
.Y(n_4986)
);

NAND2xp5_ASAP7_75t_L g4987 ( 
.A(n_4845),
.B(n_757),
.Y(n_4987)
);

INVx1_ASAP7_75t_L g4988 ( 
.A(n_4728),
.Y(n_4988)
);

AND2x2_ASAP7_75t_L g4989 ( 
.A(n_4846),
.B(n_758),
.Y(n_4989)
);

INVx2_ASAP7_75t_L g4990 ( 
.A(n_4904),
.Y(n_4990)
);

INVx1_ASAP7_75t_L g4991 ( 
.A(n_4922),
.Y(n_4991)
);

AND2x2_ASAP7_75t_L g4992 ( 
.A(n_4872),
.B(n_4744),
.Y(n_4992)
);

AND2x2_ASAP7_75t_L g4993 ( 
.A(n_4933),
.B(n_4943),
.Y(n_4993)
);

INVx1_ASAP7_75t_L g4994 ( 
.A(n_4884),
.Y(n_4994)
);

AND2x2_ASAP7_75t_L g4995 ( 
.A(n_4933),
.B(n_4851),
.Y(n_4995)
);

AND2x2_ASAP7_75t_L g4996 ( 
.A(n_4943),
.B(n_4852),
.Y(n_4996)
);

INVx1_ASAP7_75t_SL g4997 ( 
.A(n_4877),
.Y(n_4997)
);

INVx1_ASAP7_75t_L g4998 ( 
.A(n_4887),
.Y(n_4998)
);

NAND3xp33_ASAP7_75t_L g4999 ( 
.A(n_4881),
.B(n_4896),
.C(n_4876),
.Y(n_4999)
);

NAND2xp5_ASAP7_75t_L g5000 ( 
.A(n_4907),
.B(n_4863),
.Y(n_5000)
);

NAND2xp5_ASAP7_75t_SL g5001 ( 
.A(n_4914),
.B(n_4866),
.Y(n_5001)
);

AOI211x1_ASAP7_75t_SL g5002 ( 
.A1(n_4931),
.A2(n_4905),
.B(n_4956),
.C(n_4889),
.Y(n_5002)
);

NAND2xp5_ASAP7_75t_L g5003 ( 
.A(n_4913),
.B(n_4868),
.Y(n_5003)
);

NAND4xp25_ASAP7_75t_SL g5004 ( 
.A(n_4899),
.B(n_4817),
.C(n_4794),
.D(n_4774),
.Y(n_5004)
);

AND2x2_ASAP7_75t_L g5005 ( 
.A(n_4900),
.B(n_4802),
.Y(n_5005)
);

INVx3_ASAP7_75t_L g5006 ( 
.A(n_4967),
.Y(n_5006)
);

AND2x2_ASAP7_75t_L g5007 ( 
.A(n_4936),
.B(n_4803),
.Y(n_5007)
);

NAND2xp5_ASAP7_75t_L g5008 ( 
.A(n_4914),
.B(n_4718),
.Y(n_5008)
);

AND2x2_ASAP7_75t_L g5009 ( 
.A(n_4961),
.B(n_4804),
.Y(n_5009)
);

INVxp67_ASAP7_75t_L g5010 ( 
.A(n_4982),
.Y(n_5010)
);

OR2x2_ASAP7_75t_L g5011 ( 
.A(n_4921),
.B(n_4780),
.Y(n_5011)
);

AND2x2_ASAP7_75t_L g5012 ( 
.A(n_4963),
.B(n_4807),
.Y(n_5012)
);

INVx1_ASAP7_75t_SL g5013 ( 
.A(n_4891),
.Y(n_5013)
);

NAND2x1p5_ASAP7_75t_L g5014 ( 
.A(n_4882),
.B(n_4756),
.Y(n_5014)
);

NAND5xp2_ASAP7_75t_L g5015 ( 
.A(n_4941),
.B(n_4823),
.C(n_4762),
.D(n_4766),
.E(n_4765),
.Y(n_5015)
);

NAND2xp5_ASAP7_75t_L g5016 ( 
.A(n_4988),
.B(n_4729),
.Y(n_5016)
);

AND2x2_ASAP7_75t_L g5017 ( 
.A(n_4909),
.B(n_4761),
.Y(n_5017)
);

OR2x2_ASAP7_75t_L g5018 ( 
.A(n_4890),
.B(n_4985),
.Y(n_5018)
);

INVx1_ASAP7_75t_L g5019 ( 
.A(n_4883),
.Y(n_5019)
);

OR2x2_ASAP7_75t_L g5020 ( 
.A(n_4915),
.B(n_4782),
.Y(n_5020)
);

NAND2xp5_ASAP7_75t_L g5021 ( 
.A(n_4880),
.B(n_4769),
.Y(n_5021)
);

OR2x2_ASAP7_75t_L g5022 ( 
.A(n_4939),
.B(n_4778),
.Y(n_5022)
);

AND2x4_ASAP7_75t_SL g5023 ( 
.A(n_4975),
.B(n_4810),
.Y(n_5023)
);

INVx1_ASAP7_75t_L g5024 ( 
.A(n_4903),
.Y(n_5024)
);

AND2x2_ASAP7_75t_L g5025 ( 
.A(n_4986),
.B(n_4795),
.Y(n_5025)
);

OR2x2_ASAP7_75t_L g5026 ( 
.A(n_4947),
.B(n_4797),
.Y(n_5026)
);

OR2x2_ASAP7_75t_L g5027 ( 
.A(n_4926),
.B(n_4849),
.Y(n_5027)
);

INVx1_ASAP7_75t_L g5028 ( 
.A(n_4906),
.Y(n_5028)
);

OAI21xp5_ASAP7_75t_L g5029 ( 
.A1(n_4901),
.A2(n_4869),
.B(n_4858),
.Y(n_5029)
);

AND2x2_ASAP7_75t_L g5030 ( 
.A(n_4894),
.B(n_759),
.Y(n_5030)
);

NAND2xp5_ASAP7_75t_L g5031 ( 
.A(n_4932),
.B(n_759),
.Y(n_5031)
);

INVx1_ASAP7_75t_L g5032 ( 
.A(n_4911),
.Y(n_5032)
);

OR2x2_ASAP7_75t_L g5033 ( 
.A(n_4888),
.B(n_1613),
.Y(n_5033)
);

INVx1_ASAP7_75t_L g5034 ( 
.A(n_4917),
.Y(n_5034)
);

AND2x2_ASAP7_75t_L g5035 ( 
.A(n_4955),
.B(n_760),
.Y(n_5035)
);

NAND2xp5_ASAP7_75t_SL g5036 ( 
.A(n_4968),
.B(n_760),
.Y(n_5036)
);

INVx1_ASAP7_75t_L g5037 ( 
.A(n_4918),
.Y(n_5037)
);

AND2x2_ASAP7_75t_L g5038 ( 
.A(n_4929),
.B(n_761),
.Y(n_5038)
);

NAND2xp5_ASAP7_75t_L g5039 ( 
.A(n_4966),
.B(n_762),
.Y(n_5039)
);

AND2x2_ASAP7_75t_L g5040 ( 
.A(n_4937),
.B(n_763),
.Y(n_5040)
);

AOI221x1_ASAP7_75t_L g5041 ( 
.A1(n_4873),
.A2(n_766),
.B1(n_764),
.B2(n_765),
.C(n_767),
.Y(n_5041)
);

AND2x2_ASAP7_75t_L g5042 ( 
.A(n_4910),
.B(n_765),
.Y(n_5042)
);

AND2x2_ASAP7_75t_L g5043 ( 
.A(n_4916),
.B(n_766),
.Y(n_5043)
);

NAND4xp25_ASAP7_75t_L g5044 ( 
.A(n_4892),
.B(n_772),
.C(n_767),
.D(n_771),
.Y(n_5044)
);

INVx1_ASAP7_75t_L g5045 ( 
.A(n_4920),
.Y(n_5045)
);

INVx1_ASAP7_75t_L g5046 ( 
.A(n_4923),
.Y(n_5046)
);

AOI22xp33_ASAP7_75t_L g5047 ( 
.A1(n_4895),
.A2(n_1628),
.B1(n_1627),
.B2(n_775),
.Y(n_5047)
);

INVx1_ASAP7_75t_L g5048 ( 
.A(n_4925),
.Y(n_5048)
);

INVx1_ASAP7_75t_L g5049 ( 
.A(n_4938),
.Y(n_5049)
);

NAND5xp2_ASAP7_75t_L g5050 ( 
.A(n_4971),
.B(n_777),
.C(n_774),
.D(n_776),
.E(n_778),
.Y(n_5050)
);

NAND2xp5_ASAP7_75t_L g5051 ( 
.A(n_4874),
.B(n_777),
.Y(n_5051)
);

AND2x2_ASAP7_75t_L g5052 ( 
.A(n_4954),
.B(n_778),
.Y(n_5052)
);

AND2x2_ASAP7_75t_L g5053 ( 
.A(n_4958),
.B(n_779),
.Y(n_5053)
);

NAND2xp5_ASAP7_75t_L g5054 ( 
.A(n_4879),
.B(n_780),
.Y(n_5054)
);

AND2x2_ASAP7_75t_L g5055 ( 
.A(n_4989),
.B(n_780),
.Y(n_5055)
);

INVx1_ASAP7_75t_L g5056 ( 
.A(n_4940),
.Y(n_5056)
);

HB1xp67_ASAP7_75t_SL g5057 ( 
.A(n_4886),
.Y(n_5057)
);

INVx2_ASAP7_75t_L g5058 ( 
.A(n_4948),
.Y(n_5058)
);

INVx1_ASAP7_75t_L g5059 ( 
.A(n_4944),
.Y(n_5059)
);

AND2x2_ASAP7_75t_L g5060 ( 
.A(n_4970),
.B(n_782),
.Y(n_5060)
);

INVx2_ASAP7_75t_L g5061 ( 
.A(n_4952),
.Y(n_5061)
);

INVx2_ASAP7_75t_L g5062 ( 
.A(n_4953),
.Y(n_5062)
);

INVx2_ASAP7_75t_L g5063 ( 
.A(n_4977),
.Y(n_5063)
);

INVx3_ASAP7_75t_R g5064 ( 
.A(n_4949),
.Y(n_5064)
);

NAND2x1_ASAP7_75t_L g5065 ( 
.A(n_4983),
.B(n_783),
.Y(n_5065)
);

INVx1_ASAP7_75t_L g5066 ( 
.A(n_4945),
.Y(n_5066)
);

INVx1_ASAP7_75t_L g5067 ( 
.A(n_4946),
.Y(n_5067)
);

INVx1_ASAP7_75t_L g5068 ( 
.A(n_4951),
.Y(n_5068)
);

INVx1_ASAP7_75t_L g5069 ( 
.A(n_4957),
.Y(n_5069)
);

BUFx12f_ASAP7_75t_L g5070 ( 
.A(n_4984),
.Y(n_5070)
);

OR2x2_ASAP7_75t_L g5071 ( 
.A(n_4893),
.B(n_1626),
.Y(n_5071)
);

INVx1_ASAP7_75t_L g5072 ( 
.A(n_4964),
.Y(n_5072)
);

OR2x2_ASAP7_75t_L g5073 ( 
.A(n_4930),
.B(n_1626),
.Y(n_5073)
);

OAI22xp5_ASAP7_75t_L g5074 ( 
.A1(n_4999),
.A2(n_4897),
.B1(n_4885),
.B2(n_4908),
.Y(n_5074)
);

AND3x2_ASAP7_75t_L g5075 ( 
.A(n_4993),
.B(n_4978),
.C(n_4959),
.Y(n_5075)
);

AND2x2_ASAP7_75t_L g5076 ( 
.A(n_4997),
.B(n_4965),
.Y(n_5076)
);

INVx1_ASAP7_75t_L g5077 ( 
.A(n_4994),
.Y(n_5077)
);

NAND2xp5_ASAP7_75t_L g5078 ( 
.A(n_4995),
.B(n_4902),
.Y(n_5078)
);

NAND2xp5_ASAP7_75t_L g5079 ( 
.A(n_4996),
.B(n_4875),
.Y(n_5079)
);

INVx1_ASAP7_75t_L g5080 ( 
.A(n_4998),
.Y(n_5080)
);

INVx1_ASAP7_75t_L g5081 ( 
.A(n_5020),
.Y(n_5081)
);

AND2x2_ASAP7_75t_L g5082 ( 
.A(n_5013),
.B(n_4969),
.Y(n_5082)
);

INVx1_ASAP7_75t_L g5083 ( 
.A(n_5016),
.Y(n_5083)
);

NAND2xp5_ASAP7_75t_L g5084 ( 
.A(n_4992),
.B(n_4972),
.Y(n_5084)
);

NAND4xp25_ASAP7_75t_L g5085 ( 
.A(n_5002),
.B(n_4898),
.C(n_4912),
.D(n_4928),
.Y(n_5085)
);

NOR3xp33_ASAP7_75t_L g5086 ( 
.A(n_5004),
.B(n_4878),
.C(n_4980),
.Y(n_5086)
);

AND2x2_ASAP7_75t_L g5087 ( 
.A(n_5009),
.B(n_4974),
.Y(n_5087)
);

INVx2_ASAP7_75t_L g5088 ( 
.A(n_5006),
.Y(n_5088)
);

INVx1_ASAP7_75t_L g5089 ( 
.A(n_4991),
.Y(n_5089)
);

NAND2x1p5_ASAP7_75t_L g5090 ( 
.A(n_5065),
.B(n_4962),
.Y(n_5090)
);

AND2x2_ASAP7_75t_L g5091 ( 
.A(n_5007),
.B(n_4979),
.Y(n_5091)
);

AND2x2_ASAP7_75t_L g5092 ( 
.A(n_5005),
.B(n_5012),
.Y(n_5092)
);

BUFx3_ASAP7_75t_L g5093 ( 
.A(n_5070),
.Y(n_5093)
);

NOR2xp33_ASAP7_75t_L g5094 ( 
.A(n_5057),
.B(n_4973),
.Y(n_5094)
);

HB1xp67_ASAP7_75t_L g5095 ( 
.A(n_5010),
.Y(n_5095)
);

INVx2_ASAP7_75t_L g5096 ( 
.A(n_5014),
.Y(n_5096)
);

INVx2_ASAP7_75t_SL g5097 ( 
.A(n_5017),
.Y(n_5097)
);

CKINVDCx14_ASAP7_75t_R g5098 ( 
.A(n_5055),
.Y(n_5098)
);

INVx1_ASAP7_75t_L g5099 ( 
.A(n_5033),
.Y(n_5099)
);

INVx2_ASAP7_75t_L g5100 ( 
.A(n_4990),
.Y(n_5100)
);

OR2x2_ASAP7_75t_L g5101 ( 
.A(n_5000),
.B(n_4981),
.Y(n_5101)
);

INVx3_ASAP7_75t_L g5102 ( 
.A(n_5011),
.Y(n_5102)
);

OR2x2_ASAP7_75t_L g5103 ( 
.A(n_5003),
.B(n_4987),
.Y(n_5103)
);

OR2x2_ASAP7_75t_L g5104 ( 
.A(n_5015),
.B(n_4960),
.Y(n_5104)
);

AOI22xp33_ASAP7_75t_L g5105 ( 
.A1(n_5044),
.A2(n_4976),
.B1(n_4924),
.B2(n_4919),
.Y(n_5105)
);

OR2x2_ASAP7_75t_L g5106 ( 
.A(n_5026),
.B(n_4950),
.Y(n_5106)
);

AND2x2_ASAP7_75t_L g5107 ( 
.A(n_5025),
.B(n_4934),
.Y(n_5107)
);

INVx2_ASAP7_75t_SL g5108 ( 
.A(n_5001),
.Y(n_5108)
);

OR2x2_ASAP7_75t_L g5109 ( 
.A(n_5022),
.B(n_4942),
.Y(n_5109)
);

NAND2xp5_ASAP7_75t_SL g5110 ( 
.A(n_5023),
.B(n_4935),
.Y(n_5110)
);

OR2x2_ASAP7_75t_L g5111 ( 
.A(n_5021),
.B(n_4927),
.Y(n_5111)
);

NAND2xp5_ASAP7_75t_L g5112 ( 
.A(n_5039),
.B(n_784),
.Y(n_5112)
);

OR2x2_ASAP7_75t_L g5113 ( 
.A(n_5018),
.B(n_784),
.Y(n_5113)
);

NAND2x1_ASAP7_75t_L g5114 ( 
.A(n_5029),
.B(n_785),
.Y(n_5114)
);

INVx1_ASAP7_75t_L g5115 ( 
.A(n_5024),
.Y(n_5115)
);

AND2x2_ASAP7_75t_L g5116 ( 
.A(n_5008),
.B(n_786),
.Y(n_5116)
);

INVx2_ASAP7_75t_L g5117 ( 
.A(n_5027),
.Y(n_5117)
);

AND2x2_ASAP7_75t_L g5118 ( 
.A(n_5030),
.B(n_787),
.Y(n_5118)
);

INVx2_ASAP7_75t_SL g5119 ( 
.A(n_5060),
.Y(n_5119)
);

INVx1_ASAP7_75t_L g5120 ( 
.A(n_5028),
.Y(n_5120)
);

OR2x2_ASAP7_75t_L g5121 ( 
.A(n_5019),
.B(n_789),
.Y(n_5121)
);

OR2x2_ASAP7_75t_L g5122 ( 
.A(n_5058),
.B(n_789),
.Y(n_5122)
);

INVx2_ASAP7_75t_L g5123 ( 
.A(n_5061),
.Y(n_5123)
);

AND2x2_ASAP7_75t_L g5124 ( 
.A(n_5035),
.B(n_791),
.Y(n_5124)
);

AND2x2_ASAP7_75t_L g5125 ( 
.A(n_5052),
.B(n_791),
.Y(n_5125)
);

OR2x2_ASAP7_75t_L g5126 ( 
.A(n_5062),
.B(n_792),
.Y(n_5126)
);

INVx2_ASAP7_75t_L g5127 ( 
.A(n_5063),
.Y(n_5127)
);

INVx1_ASAP7_75t_L g5128 ( 
.A(n_5032),
.Y(n_5128)
);

OR2x2_ASAP7_75t_L g5129 ( 
.A(n_5051),
.B(n_793),
.Y(n_5129)
);

INVx1_ASAP7_75t_SL g5130 ( 
.A(n_5042),
.Y(n_5130)
);

OR2x2_ASAP7_75t_L g5131 ( 
.A(n_5054),
.B(n_794),
.Y(n_5131)
);

INVxp67_ASAP7_75t_L g5132 ( 
.A(n_5036),
.Y(n_5132)
);

HB1xp67_ASAP7_75t_L g5133 ( 
.A(n_5064),
.Y(n_5133)
);

INVx1_ASAP7_75t_L g5134 ( 
.A(n_5034),
.Y(n_5134)
);

INVx1_ASAP7_75t_L g5135 ( 
.A(n_5037),
.Y(n_5135)
);

OR2x2_ASAP7_75t_L g5136 ( 
.A(n_5073),
.B(n_5031),
.Y(n_5136)
);

INVx1_ASAP7_75t_SL g5137 ( 
.A(n_5043),
.Y(n_5137)
);

AND2x2_ASAP7_75t_L g5138 ( 
.A(n_5053),
.B(n_795),
.Y(n_5138)
);

AND2x2_ASAP7_75t_L g5139 ( 
.A(n_5038),
.B(n_795),
.Y(n_5139)
);

INVx1_ASAP7_75t_L g5140 ( 
.A(n_5045),
.Y(n_5140)
);

INVx1_ASAP7_75t_L g5141 ( 
.A(n_5046),
.Y(n_5141)
);

AND2x2_ASAP7_75t_L g5142 ( 
.A(n_5040),
.B(n_797),
.Y(n_5142)
);

INVx1_ASAP7_75t_L g5143 ( 
.A(n_5048),
.Y(n_5143)
);

INVx2_ASAP7_75t_L g5144 ( 
.A(n_5071),
.Y(n_5144)
);

INVx2_ASAP7_75t_L g5145 ( 
.A(n_5049),
.Y(n_5145)
);

NAND2xp5_ASAP7_75t_L g5146 ( 
.A(n_5041),
.B(n_798),
.Y(n_5146)
);

HB1xp67_ASAP7_75t_L g5147 ( 
.A(n_5056),
.Y(n_5147)
);

INVx1_ASAP7_75t_L g5148 ( 
.A(n_5059),
.Y(n_5148)
);

AND2x2_ASAP7_75t_L g5149 ( 
.A(n_5066),
.B(n_799),
.Y(n_5149)
);

AND2x2_ASAP7_75t_L g5150 ( 
.A(n_5067),
.B(n_801),
.Y(n_5150)
);

OAI31xp33_ASAP7_75t_L g5151 ( 
.A1(n_5050),
.A2(n_804),
.A3(n_801),
.B(n_803),
.Y(n_5151)
);

OR2x2_ASAP7_75t_L g5152 ( 
.A(n_5068),
.B(n_803),
.Y(n_5152)
);

NAND2xp5_ASAP7_75t_L g5153 ( 
.A(n_5069),
.B(n_805),
.Y(n_5153)
);

AND2x2_ASAP7_75t_L g5154 ( 
.A(n_5072),
.B(n_806),
.Y(n_5154)
);

AND2x2_ASAP7_75t_SL g5155 ( 
.A(n_5047),
.B(n_807),
.Y(n_5155)
);

INVx1_ASAP7_75t_SL g5156 ( 
.A(n_5133),
.Y(n_5156)
);

NAND2xp5_ASAP7_75t_L g5157 ( 
.A(n_5095),
.B(n_807),
.Y(n_5157)
);

HB1xp67_ASAP7_75t_L g5158 ( 
.A(n_5098),
.Y(n_5158)
);

INVxp67_ASAP7_75t_L g5159 ( 
.A(n_5094),
.Y(n_5159)
);

INVx1_ASAP7_75t_L g5160 ( 
.A(n_5102),
.Y(n_5160)
);

OR2x2_ASAP7_75t_L g5161 ( 
.A(n_5106),
.B(n_809),
.Y(n_5161)
);

NOR2x1_ASAP7_75t_L g5162 ( 
.A(n_5085),
.B(n_809),
.Y(n_5162)
);

OAI22xp5_ASAP7_75t_L g5163 ( 
.A1(n_5105),
.A2(n_812),
.B1(n_813),
.B2(n_811),
.Y(n_5163)
);

INVx1_ASAP7_75t_L g5164 ( 
.A(n_5122),
.Y(n_5164)
);

INVx1_ASAP7_75t_L g5165 ( 
.A(n_5126),
.Y(n_5165)
);

NAND2xp5_ASAP7_75t_L g5166 ( 
.A(n_5075),
.B(n_814),
.Y(n_5166)
);

INVx3_ASAP7_75t_L g5167 ( 
.A(n_5088),
.Y(n_5167)
);

AOI22xp33_ASAP7_75t_L g5168 ( 
.A1(n_5086),
.A2(n_817),
.B1(n_815),
.B2(n_816),
.Y(n_5168)
);

OR2x6_ASAP7_75t_L g5169 ( 
.A(n_5108),
.B(n_818),
.Y(n_5169)
);

OAI222xp33_ASAP7_75t_L g5170 ( 
.A1(n_5104),
.A2(n_1613),
.B1(n_1605),
.B2(n_822),
.C1(n_823),
.C2(n_820),
.Y(n_5170)
);

AND2x2_ASAP7_75t_SL g5171 ( 
.A(n_5155),
.B(n_821),
.Y(n_5171)
);

NOR2xp33_ASAP7_75t_SL g5172 ( 
.A(n_5132),
.B(n_1608),
.Y(n_5172)
);

NAND2xp5_ASAP7_75t_L g5173 ( 
.A(n_5092),
.B(n_821),
.Y(n_5173)
);

NAND2xp5_ASAP7_75t_L g5174 ( 
.A(n_5130),
.B(n_5137),
.Y(n_5174)
);

NAND2xp5_ASAP7_75t_L g5175 ( 
.A(n_5097),
.B(n_824),
.Y(n_5175)
);

INVx1_ASAP7_75t_SL g5176 ( 
.A(n_5082),
.Y(n_5176)
);

INVx1_ASAP7_75t_L g5177 ( 
.A(n_5081),
.Y(n_5177)
);

INVx1_ASAP7_75t_SL g5178 ( 
.A(n_5076),
.Y(n_5178)
);

AND2x4_ASAP7_75t_L g5179 ( 
.A(n_5096),
.B(n_825),
.Y(n_5179)
);

INVx1_ASAP7_75t_L g5180 ( 
.A(n_5149),
.Y(n_5180)
);

INVx1_ASAP7_75t_L g5181 ( 
.A(n_5150),
.Y(n_5181)
);

INVx1_ASAP7_75t_L g5182 ( 
.A(n_5154),
.Y(n_5182)
);

AND2x2_ASAP7_75t_L g5183 ( 
.A(n_5091),
.B(n_1612),
.Y(n_5183)
);

INVx1_ASAP7_75t_L g5184 ( 
.A(n_5147),
.Y(n_5184)
);

INVxp67_ASAP7_75t_SL g5185 ( 
.A(n_5090),
.Y(n_5185)
);

NAND2xp5_ASAP7_75t_L g5186 ( 
.A(n_5119),
.B(n_826),
.Y(n_5186)
);

NOR2xp67_ASAP7_75t_L g5187 ( 
.A(n_5099),
.B(n_1623),
.Y(n_5187)
);

AND2x2_ASAP7_75t_L g5188 ( 
.A(n_5087),
.B(n_1627),
.Y(n_5188)
);

NOR2xp33_ASAP7_75t_L g5189 ( 
.A(n_5110),
.B(n_1628),
.Y(n_5189)
);

INVx1_ASAP7_75t_SL g5190 ( 
.A(n_5113),
.Y(n_5190)
);

OAI22xp5_ASAP7_75t_L g5191 ( 
.A1(n_5074),
.A2(n_828),
.B1(n_829),
.B2(n_827),
.Y(n_5191)
);

OAI21xp5_ASAP7_75t_L g5192 ( 
.A1(n_5114),
.A2(n_832),
.B(n_833),
.Y(n_5192)
);

INVx2_ASAP7_75t_L g5193 ( 
.A(n_5100),
.Y(n_5193)
);

OR2x2_ASAP7_75t_L g5194 ( 
.A(n_5078),
.B(n_5079),
.Y(n_5194)
);

AND2x4_ASAP7_75t_L g5195 ( 
.A(n_5117),
.B(n_833),
.Y(n_5195)
);

AOI21xp33_ASAP7_75t_L g5196 ( 
.A1(n_5109),
.A2(n_834),
.B(n_835),
.Y(n_5196)
);

AOI222xp33_ASAP7_75t_L g5197 ( 
.A1(n_5107),
.A2(n_837),
.B1(n_839),
.B2(n_841),
.C1(n_836),
.C2(n_838),
.Y(n_5197)
);

OR2x2_ASAP7_75t_L g5198 ( 
.A(n_5101),
.B(n_834),
.Y(n_5198)
);

NAND2x1p5_ASAP7_75t_L g5199 ( 
.A(n_5125),
.B(n_841),
.Y(n_5199)
);

AND2x2_ASAP7_75t_L g5200 ( 
.A(n_5116),
.B(n_1615),
.Y(n_5200)
);

INVx2_ASAP7_75t_L g5201 ( 
.A(n_5138),
.Y(n_5201)
);

OAI22xp5_ASAP7_75t_L g5202 ( 
.A1(n_5111),
.A2(n_844),
.B1(n_845),
.B2(n_843),
.Y(n_5202)
);

AND2x2_ASAP7_75t_L g5203 ( 
.A(n_5144),
.B(n_1615),
.Y(n_5203)
);

NAND2x1p5_ASAP7_75t_L g5204 ( 
.A(n_5139),
.B(n_843),
.Y(n_5204)
);

INVx1_ASAP7_75t_L g5205 ( 
.A(n_5152),
.Y(n_5205)
);

INVx3_ASAP7_75t_L g5206 ( 
.A(n_5123),
.Y(n_5206)
);

INVx1_ASAP7_75t_L g5207 ( 
.A(n_5121),
.Y(n_5207)
);

INVx2_ASAP7_75t_L g5208 ( 
.A(n_5142),
.Y(n_5208)
);

OAI21xp5_ASAP7_75t_L g5209 ( 
.A1(n_5146),
.A2(n_844),
.B(n_847),
.Y(n_5209)
);

NAND2x2_ASAP7_75t_L g5210 ( 
.A(n_5103),
.B(n_849),
.Y(n_5210)
);

NAND2xp5_ASAP7_75t_L g5211 ( 
.A(n_5089),
.B(n_849),
.Y(n_5211)
);

AOI221xp5_ASAP7_75t_L g5212 ( 
.A1(n_5077),
.A2(n_852),
.B1(n_850),
.B2(n_851),
.C(n_853),
.Y(n_5212)
);

INVx1_ASAP7_75t_L g5213 ( 
.A(n_5084),
.Y(n_5213)
);

NAND2xp5_ASAP7_75t_L g5214 ( 
.A(n_5080),
.B(n_851),
.Y(n_5214)
);

AND2x2_ASAP7_75t_L g5215 ( 
.A(n_5083),
.B(n_1607),
.Y(n_5215)
);

NAND3xp33_ASAP7_75t_L g5216 ( 
.A(n_5151),
.B(n_854),
.C(n_855),
.Y(n_5216)
);

OR2x2_ASAP7_75t_L g5217 ( 
.A(n_5136),
.B(n_855),
.Y(n_5217)
);

INVx2_ASAP7_75t_L g5218 ( 
.A(n_5124),
.Y(n_5218)
);

AO22x1_ASAP7_75t_L g5219 ( 
.A1(n_5145),
.A2(n_858),
.B1(n_856),
.B2(n_857),
.Y(n_5219)
);

INVx2_ASAP7_75t_L g5220 ( 
.A(n_5118),
.Y(n_5220)
);

AND2x2_ASAP7_75t_L g5221 ( 
.A(n_5127),
.B(n_1614),
.Y(n_5221)
);

NAND2xp5_ASAP7_75t_L g5222 ( 
.A(n_5112),
.B(n_857),
.Y(n_5222)
);

INVxp67_ASAP7_75t_L g5223 ( 
.A(n_5129),
.Y(n_5223)
);

INVx3_ASAP7_75t_L g5224 ( 
.A(n_5131),
.Y(n_5224)
);

NAND2xp5_ASAP7_75t_L g5225 ( 
.A(n_5153),
.B(n_858),
.Y(n_5225)
);

NAND2xp5_ASAP7_75t_L g5226 ( 
.A(n_5115),
.B(n_860),
.Y(n_5226)
);

INVx1_ASAP7_75t_L g5227 ( 
.A(n_5120),
.Y(n_5227)
);

OAI211xp5_ASAP7_75t_L g5228 ( 
.A1(n_5128),
.A2(n_5135),
.B(n_5140),
.C(n_5134),
.Y(n_5228)
);

AOI211xp5_ASAP7_75t_L g5229 ( 
.A1(n_5141),
.A2(n_863),
.B(n_861),
.C(n_862),
.Y(n_5229)
);

AOI32xp33_ASAP7_75t_L g5230 ( 
.A1(n_5143),
.A2(n_863),
.A3(n_861),
.B1(n_862),
.B2(n_864),
.Y(n_5230)
);

INVx1_ASAP7_75t_L g5231 ( 
.A(n_5148),
.Y(n_5231)
);

NAND2xp5_ASAP7_75t_L g5232 ( 
.A(n_5133),
.B(n_865),
.Y(n_5232)
);

NAND2xp5_ASAP7_75t_L g5233 ( 
.A(n_5133),
.B(n_866),
.Y(n_5233)
);

INVx2_ASAP7_75t_L g5234 ( 
.A(n_5093),
.Y(n_5234)
);

AOI222xp33_ASAP7_75t_L g5235 ( 
.A1(n_5163),
.A2(n_888),
.B1(n_873),
.B2(n_894),
.C1(n_880),
.C2(n_868),
.Y(n_5235)
);

OR2x2_ASAP7_75t_L g5236 ( 
.A(n_5156),
.B(n_869),
.Y(n_5236)
);

INVx1_ASAP7_75t_L g5237 ( 
.A(n_5158),
.Y(n_5237)
);

OR2x2_ASAP7_75t_L g5238 ( 
.A(n_5178),
.B(n_870),
.Y(n_5238)
);

AND2x4_ASAP7_75t_L g5239 ( 
.A(n_5185),
.B(n_873),
.Y(n_5239)
);

OAI22xp5_ASAP7_75t_L g5240 ( 
.A1(n_5216),
.A2(n_876),
.B1(n_874),
.B2(n_875),
.Y(n_5240)
);

OR2x2_ASAP7_75t_L g5241 ( 
.A(n_5176),
.B(n_875),
.Y(n_5241)
);

OAI22xp5_ASAP7_75t_L g5242 ( 
.A1(n_5168),
.A2(n_879),
.B1(n_877),
.B2(n_878),
.Y(n_5242)
);

INVx2_ASAP7_75t_L g5243 ( 
.A(n_5234),
.Y(n_5243)
);

INVx1_ASAP7_75t_L g5244 ( 
.A(n_5174),
.Y(n_5244)
);

INVx1_ASAP7_75t_L g5245 ( 
.A(n_5187),
.Y(n_5245)
);

AOI21xp5_ASAP7_75t_L g5246 ( 
.A1(n_5209),
.A2(n_880),
.B(n_882),
.Y(n_5246)
);

NAND4xp25_ASAP7_75t_L g5247 ( 
.A(n_5159),
.B(n_884),
.C(n_882),
.D(n_883),
.Y(n_5247)
);

INVx1_ASAP7_75t_L g5248 ( 
.A(n_5232),
.Y(n_5248)
);

HB1xp67_ASAP7_75t_L g5249 ( 
.A(n_5169),
.Y(n_5249)
);

INVx1_ASAP7_75t_L g5250 ( 
.A(n_5233),
.Y(n_5250)
);

NAND2xp5_ASAP7_75t_L g5251 ( 
.A(n_5167),
.B(n_885),
.Y(n_5251)
);

OAI22xp5_ASAP7_75t_L g5252 ( 
.A1(n_5210),
.A2(n_5194),
.B1(n_5189),
.B2(n_5160),
.Y(n_5252)
);

AOI21xp5_ASAP7_75t_L g5253 ( 
.A1(n_5192),
.A2(n_885),
.B(n_886),
.Y(n_5253)
);

A2O1A1Ixp33_ASAP7_75t_SL g5254 ( 
.A1(n_5223),
.A2(n_888),
.B(n_886),
.C(n_887),
.Y(n_5254)
);

NAND2xp5_ASAP7_75t_L g5255 ( 
.A(n_5183),
.B(n_889),
.Y(n_5255)
);

AOI21xp33_ASAP7_75t_L g5256 ( 
.A1(n_5190),
.A2(n_1608),
.B(n_1606),
.Y(n_5256)
);

OR2x2_ASAP7_75t_L g5257 ( 
.A(n_5161),
.B(n_5169),
.Y(n_5257)
);

OAI21xp5_ASAP7_75t_L g5258 ( 
.A1(n_5170),
.A2(n_891),
.B(n_893),
.Y(n_5258)
);

INVx1_ASAP7_75t_SL g5259 ( 
.A(n_5188),
.Y(n_5259)
);

AND2x2_ASAP7_75t_L g5260 ( 
.A(n_5201),
.B(n_891),
.Y(n_5260)
);

AO21x1_ASAP7_75t_L g5261 ( 
.A1(n_5191),
.A2(n_897),
.B(n_895),
.Y(n_5261)
);

NAND2xp5_ASAP7_75t_SL g5262 ( 
.A(n_5172),
.B(n_893),
.Y(n_5262)
);

INVx1_ASAP7_75t_L g5263 ( 
.A(n_5203),
.Y(n_5263)
);

A2O1A1Ixp33_ASAP7_75t_SL g5264 ( 
.A1(n_5224),
.A2(n_5184),
.B(n_5206),
.C(n_5193),
.Y(n_5264)
);

OAI221xp5_ASAP7_75t_SL g5265 ( 
.A1(n_5230),
.A2(n_917),
.B1(n_923),
.B2(n_906),
.C(n_899),
.Y(n_5265)
);

INVx1_ASAP7_75t_SL g5266 ( 
.A(n_5199),
.Y(n_5266)
);

AOI22xp33_ASAP7_75t_L g5267 ( 
.A1(n_5208),
.A2(n_902),
.B1(n_900),
.B2(n_901),
.Y(n_5267)
);

NAND3xp33_ASAP7_75t_L g5268 ( 
.A(n_5197),
.B(n_903),
.C(n_904),
.Y(n_5268)
);

AOI22xp5_ASAP7_75t_L g5269 ( 
.A1(n_5180),
.A2(n_905),
.B1(n_903),
.B2(n_904),
.Y(n_5269)
);

INVx1_ASAP7_75t_L g5270 ( 
.A(n_5218),
.Y(n_5270)
);

OAI321xp33_ASAP7_75t_L g5271 ( 
.A1(n_5177),
.A2(n_908),
.A3(n_911),
.B1(n_905),
.B2(n_907),
.C(n_910),
.Y(n_5271)
);

INVx1_ASAP7_75t_L g5272 ( 
.A(n_5220),
.Y(n_5272)
);

OAI21xp5_ASAP7_75t_L g5273 ( 
.A1(n_5196),
.A2(n_914),
.B(n_916),
.Y(n_5273)
);

NAND2xp5_ASAP7_75t_L g5274 ( 
.A(n_5179),
.B(n_916),
.Y(n_5274)
);

NOR5xp2_ASAP7_75t_L g5275 ( 
.A(n_5228),
.B(n_920),
.C(n_918),
.D(n_919),
.E(n_921),
.Y(n_5275)
);

INVx2_ASAP7_75t_L g5276 ( 
.A(n_5204),
.Y(n_5276)
);

AND2x2_ASAP7_75t_L g5277 ( 
.A(n_5181),
.B(n_919),
.Y(n_5277)
);

AND2x2_ASAP7_75t_L g5278 ( 
.A(n_5182),
.B(n_920),
.Y(n_5278)
);

NAND2xp5_ASAP7_75t_L g5279 ( 
.A(n_5195),
.B(n_922),
.Y(n_5279)
);

OR2x2_ASAP7_75t_L g5280 ( 
.A(n_5157),
.B(n_5198),
.Y(n_5280)
);

INVxp67_ASAP7_75t_L g5281 ( 
.A(n_5200),
.Y(n_5281)
);

INVx1_ASAP7_75t_L g5282 ( 
.A(n_5175),
.Y(n_5282)
);

NAND2xp5_ASAP7_75t_L g5283 ( 
.A(n_5221),
.B(n_928),
.Y(n_5283)
);

INVx1_ASAP7_75t_L g5284 ( 
.A(n_5186),
.Y(n_5284)
);

OAI21xp5_ASAP7_75t_L g5285 ( 
.A1(n_5212),
.A2(n_929),
.B(n_930),
.Y(n_5285)
);

AND2x2_ASAP7_75t_L g5286 ( 
.A(n_5205),
.B(n_933),
.Y(n_5286)
);

INVxp67_ASAP7_75t_L g5287 ( 
.A(n_5173),
.Y(n_5287)
);

AOI22xp5_ASAP7_75t_L g5288 ( 
.A1(n_5213),
.A2(n_937),
.B1(n_934),
.B2(n_936),
.Y(n_5288)
);

AOI211xp5_ASAP7_75t_L g5289 ( 
.A1(n_5202),
.A2(n_942),
.B(n_938),
.C(n_941),
.Y(n_5289)
);

NOR2xp33_ASAP7_75t_SL g5290 ( 
.A(n_5207),
.B(n_938),
.Y(n_5290)
);

AND2x2_ASAP7_75t_L g5291 ( 
.A(n_5164),
.B(n_943),
.Y(n_5291)
);

AO22x1_ASAP7_75t_L g5292 ( 
.A1(n_5165),
.A2(n_948),
.B1(n_945),
.B2(n_947),
.Y(n_5292)
);

AOI31xp33_ASAP7_75t_L g5293 ( 
.A1(n_5229),
.A2(n_954),
.A3(n_949),
.B(n_953),
.Y(n_5293)
);

AOI211xp5_ASAP7_75t_L g5294 ( 
.A1(n_5219),
.A2(n_957),
.B(n_955),
.C(n_956),
.Y(n_5294)
);

INVx1_ASAP7_75t_L g5295 ( 
.A(n_5217),
.Y(n_5295)
);

INVx1_ASAP7_75t_L g5296 ( 
.A(n_5215),
.Y(n_5296)
);

OAI322xp33_ASAP7_75t_L g5297 ( 
.A1(n_5227),
.A2(n_965),
.A3(n_964),
.B1(n_962),
.B2(n_959),
.C1(n_961),
.C2(n_963),
.Y(n_5297)
);

OAI22xp33_ASAP7_75t_L g5298 ( 
.A1(n_5211),
.A2(n_965),
.B1(n_961),
.B2(n_962),
.Y(n_5298)
);

AOI221xp5_ASAP7_75t_L g5299 ( 
.A1(n_5231),
.A2(n_981),
.B1(n_988),
.B2(n_974),
.C(n_966),
.Y(n_5299)
);

OR2x2_ASAP7_75t_L g5300 ( 
.A(n_5214),
.B(n_966),
.Y(n_5300)
);

O2A1O1Ixp33_ASAP7_75t_L g5301 ( 
.A1(n_5226),
.A2(n_1610),
.B(n_1611),
.C(n_1609),
.Y(n_5301)
);

INVx2_ASAP7_75t_L g5302 ( 
.A(n_5222),
.Y(n_5302)
);

AOI222xp33_ASAP7_75t_L g5303 ( 
.A1(n_5225),
.A2(n_991),
.B1(n_975),
.B2(n_1001),
.C1(n_984),
.C2(n_967),
.Y(n_5303)
);

OR2x2_ASAP7_75t_L g5304 ( 
.A(n_5156),
.B(n_967),
.Y(n_5304)
);

AND2x2_ASAP7_75t_L g5305 ( 
.A(n_5158),
.B(n_969),
.Y(n_5305)
);

INVx1_ASAP7_75t_L g5306 ( 
.A(n_5158),
.Y(n_5306)
);

INVx1_ASAP7_75t_L g5307 ( 
.A(n_5158),
.Y(n_5307)
);

INVx1_ASAP7_75t_L g5308 ( 
.A(n_5158),
.Y(n_5308)
);

INVx2_ASAP7_75t_L g5309 ( 
.A(n_5158),
.Y(n_5309)
);

NAND2xp5_ASAP7_75t_L g5310 ( 
.A(n_5158),
.B(n_970),
.Y(n_5310)
);

OAI22xp33_ASAP7_75t_L g5311 ( 
.A1(n_5216),
.A2(n_972),
.B1(n_970),
.B2(n_971),
.Y(n_5311)
);

AOI21xp33_ASAP7_75t_L g5312 ( 
.A1(n_5158),
.A2(n_1599),
.B(n_1598),
.Y(n_5312)
);

OAI21xp5_ASAP7_75t_SL g5313 ( 
.A1(n_5166),
.A2(n_1600),
.B(n_1599),
.Y(n_5313)
);

AND2x2_ASAP7_75t_L g5314 ( 
.A(n_5158),
.B(n_974),
.Y(n_5314)
);

INVx1_ASAP7_75t_L g5315 ( 
.A(n_5158),
.Y(n_5315)
);

AOI21xp33_ASAP7_75t_L g5316 ( 
.A1(n_5158),
.A2(n_1604),
.B(n_1602),
.Y(n_5316)
);

OAI221xp5_ASAP7_75t_L g5317 ( 
.A1(n_5166),
.A2(n_979),
.B1(n_977),
.B2(n_978),
.C(n_980),
.Y(n_5317)
);

INVx1_ASAP7_75t_L g5318 ( 
.A(n_5158),
.Y(n_5318)
);

INVxp67_ASAP7_75t_SL g5319 ( 
.A(n_5158),
.Y(n_5319)
);

AOI22xp5_ASAP7_75t_L g5320 ( 
.A1(n_5156),
.A2(n_990),
.B1(n_987),
.B2(n_989),
.Y(n_5320)
);

AOI21xp5_ASAP7_75t_L g5321 ( 
.A1(n_5166),
.A2(n_992),
.B(n_994),
.Y(n_5321)
);

AOI22xp33_ASAP7_75t_L g5322 ( 
.A1(n_5162),
.A2(n_996),
.B1(n_994),
.B2(n_995),
.Y(n_5322)
);

INVx2_ASAP7_75t_SL g5323 ( 
.A(n_5158),
.Y(n_5323)
);

NAND2xp5_ASAP7_75t_SL g5324 ( 
.A(n_5171),
.B(n_995),
.Y(n_5324)
);

INVx1_ASAP7_75t_L g5325 ( 
.A(n_5158),
.Y(n_5325)
);

INVx1_ASAP7_75t_L g5326 ( 
.A(n_5158),
.Y(n_5326)
);

INVxp67_ASAP7_75t_L g5327 ( 
.A(n_5158),
.Y(n_5327)
);

OAI22xp5_ASAP7_75t_L g5328 ( 
.A1(n_5216),
.A2(n_999),
.B1(n_997),
.B2(n_998),
.Y(n_5328)
);

OAI22xp33_ASAP7_75t_SL g5329 ( 
.A1(n_5166),
.A2(n_1003),
.B1(n_998),
.B2(n_1002),
.Y(n_5329)
);

AOI22xp5_ASAP7_75t_L g5330 ( 
.A1(n_5156),
.A2(n_1004),
.B1(n_1002),
.B2(n_1003),
.Y(n_5330)
);

AND2x2_ASAP7_75t_L g5331 ( 
.A(n_5158),
.B(n_1006),
.Y(n_5331)
);

OAI21xp33_ASAP7_75t_L g5332 ( 
.A1(n_5156),
.A2(n_1007),
.B(n_1008),
.Y(n_5332)
);

INVx2_ASAP7_75t_L g5333 ( 
.A(n_5158),
.Y(n_5333)
);

OAI22xp33_ASAP7_75t_L g5334 ( 
.A1(n_5216),
.A2(n_1011),
.B1(n_1009),
.B2(n_1010),
.Y(n_5334)
);

INVxp67_ASAP7_75t_L g5335 ( 
.A(n_5158),
.Y(n_5335)
);

AOI21xp33_ASAP7_75t_L g5336 ( 
.A1(n_5158),
.A2(n_1624),
.B(n_1013),
.Y(n_5336)
);

INVx1_ASAP7_75t_L g5337 ( 
.A(n_5158),
.Y(n_5337)
);

INVxp67_ASAP7_75t_SL g5338 ( 
.A(n_5158),
.Y(n_5338)
);

AOI22xp33_ASAP7_75t_L g5339 ( 
.A1(n_5162),
.A2(n_1017),
.B1(n_1015),
.B2(n_1016),
.Y(n_5339)
);

AND2x2_ASAP7_75t_SL g5340 ( 
.A(n_5171),
.B(n_1017),
.Y(n_5340)
);

BUFx2_ASAP7_75t_L g5341 ( 
.A(n_5158),
.Y(n_5341)
);

XOR2x2_ASAP7_75t_L g5342 ( 
.A(n_5216),
.B(n_1021),
.Y(n_5342)
);

HB1xp67_ASAP7_75t_L g5343 ( 
.A(n_5249),
.Y(n_5343)
);

NAND2xp5_ASAP7_75t_L g5344 ( 
.A(n_5319),
.B(n_5338),
.Y(n_5344)
);

AOI21xp33_ASAP7_75t_L g5345 ( 
.A1(n_5264),
.A2(n_1025),
.B(n_1026),
.Y(n_5345)
);

OAI21xp5_ASAP7_75t_L g5346 ( 
.A1(n_5268),
.A2(n_1029),
.B(n_1027),
.Y(n_5346)
);

NAND3xp33_ASAP7_75t_L g5347 ( 
.A(n_5245),
.B(n_1030),
.C(n_1031),
.Y(n_5347)
);

OAI321xp33_ASAP7_75t_L g5348 ( 
.A1(n_5327),
.A2(n_1034),
.A3(n_1036),
.B1(n_1032),
.B2(n_1033),
.C(n_1035),
.Y(n_5348)
);

O2A1O1Ixp33_ASAP7_75t_L g5349 ( 
.A1(n_5254),
.A2(n_1037),
.B(n_1034),
.C(n_1035),
.Y(n_5349)
);

INVx1_ASAP7_75t_L g5350 ( 
.A(n_5341),
.Y(n_5350)
);

INVxp67_ASAP7_75t_L g5351 ( 
.A(n_5290),
.Y(n_5351)
);

INVx1_ASAP7_75t_L g5352 ( 
.A(n_5305),
.Y(n_5352)
);

INVx1_ASAP7_75t_L g5353 ( 
.A(n_5314),
.Y(n_5353)
);

INVx1_ASAP7_75t_L g5354 ( 
.A(n_5331),
.Y(n_5354)
);

INVx1_ASAP7_75t_L g5355 ( 
.A(n_5237),
.Y(n_5355)
);

AOI22xp5_ASAP7_75t_SL g5356 ( 
.A1(n_5292),
.A2(n_1042),
.B1(n_1038),
.B2(n_1041),
.Y(n_5356)
);

OAI22xp5_ASAP7_75t_L g5357 ( 
.A1(n_5335),
.A2(n_5322),
.B1(n_5339),
.B2(n_5323),
.Y(n_5357)
);

NAND2xp5_ASAP7_75t_L g5358 ( 
.A(n_5340),
.B(n_1043),
.Y(n_5358)
);

HB1xp67_ASAP7_75t_L g5359 ( 
.A(n_5257),
.Y(n_5359)
);

NAND2xp5_ASAP7_75t_L g5360 ( 
.A(n_5309),
.B(n_1045),
.Y(n_5360)
);

OAI22xp5_ASAP7_75t_L g5361 ( 
.A1(n_5333),
.A2(n_1050),
.B1(n_1047),
.B2(n_1049),
.Y(n_5361)
);

OAI22xp5_ASAP7_75t_L g5362 ( 
.A1(n_5306),
.A2(n_1050),
.B1(n_1047),
.B2(n_1049),
.Y(n_5362)
);

OR2x2_ASAP7_75t_L g5363 ( 
.A(n_5307),
.B(n_5308),
.Y(n_5363)
);

INVx1_ASAP7_75t_L g5364 ( 
.A(n_5315),
.Y(n_5364)
);

INVx1_ASAP7_75t_L g5365 ( 
.A(n_5318),
.Y(n_5365)
);

NAND2xp5_ASAP7_75t_L g5366 ( 
.A(n_5325),
.B(n_1054),
.Y(n_5366)
);

NAND2xp5_ASAP7_75t_L g5367 ( 
.A(n_5326),
.B(n_1055),
.Y(n_5367)
);

INVx1_ASAP7_75t_L g5368 ( 
.A(n_5337),
.Y(n_5368)
);

NOR2xp33_ASAP7_75t_L g5369 ( 
.A(n_5266),
.B(n_1056),
.Y(n_5369)
);

INVx1_ASAP7_75t_L g5370 ( 
.A(n_5236),
.Y(n_5370)
);

AOI22xp5_ASAP7_75t_SL g5371 ( 
.A1(n_5329),
.A2(n_1060),
.B1(n_1058),
.B2(n_1059),
.Y(n_5371)
);

INVx1_ASAP7_75t_L g5372 ( 
.A(n_5304),
.Y(n_5372)
);

O2A1O1Ixp33_ASAP7_75t_L g5373 ( 
.A1(n_5258),
.A2(n_1062),
.B(n_1059),
.C(n_1060),
.Y(n_5373)
);

OAI22xp5_ASAP7_75t_L g5374 ( 
.A1(n_5265),
.A2(n_5259),
.B1(n_5281),
.B2(n_5244),
.Y(n_5374)
);

NAND2xp5_ASAP7_75t_L g5375 ( 
.A(n_5239),
.B(n_1063),
.Y(n_5375)
);

OA21x2_ASAP7_75t_L g5376 ( 
.A1(n_5321),
.A2(n_1065),
.B(n_1066),
.Y(n_5376)
);

OAI22xp5_ASAP7_75t_L g5377 ( 
.A1(n_5320),
.A2(n_1067),
.B1(n_1065),
.B2(n_1066),
.Y(n_5377)
);

INVx1_ASAP7_75t_L g5378 ( 
.A(n_5310),
.Y(n_5378)
);

OAI21xp33_ASAP7_75t_L g5379 ( 
.A1(n_5243),
.A2(n_1068),
.B(n_1069),
.Y(n_5379)
);

INVx2_ASAP7_75t_L g5380 ( 
.A(n_5239),
.Y(n_5380)
);

INVx2_ASAP7_75t_L g5381 ( 
.A(n_5276),
.Y(n_5381)
);

INVx1_ASAP7_75t_SL g5382 ( 
.A(n_5324),
.Y(n_5382)
);

INVx1_ASAP7_75t_SL g5383 ( 
.A(n_5238),
.Y(n_5383)
);

OAI22xp5_ASAP7_75t_L g5384 ( 
.A1(n_5330),
.A2(n_1073),
.B1(n_1071),
.B2(n_1072),
.Y(n_5384)
);

AND2x2_ASAP7_75t_L g5385 ( 
.A(n_5296),
.B(n_1072),
.Y(n_5385)
);

AOI21xp33_ASAP7_75t_L g5386 ( 
.A1(n_5252),
.A2(n_1073),
.B(n_1074),
.Y(n_5386)
);

OAI32xp33_ASAP7_75t_L g5387 ( 
.A1(n_5270),
.A2(n_1093),
.A3(n_1101),
.B1(n_1083),
.B2(n_1075),
.Y(n_5387)
);

AOI222xp33_ASAP7_75t_L g5388 ( 
.A1(n_5285),
.A2(n_1078),
.B1(n_1080),
.B2(n_1076),
.C1(n_1077),
.C2(n_1079),
.Y(n_5388)
);

AOI222xp33_ASAP7_75t_L g5389 ( 
.A1(n_5273),
.A2(n_1081),
.B1(n_1084),
.B2(n_1077),
.C1(n_1079),
.C2(n_1082),
.Y(n_5389)
);

INVx3_ASAP7_75t_L g5390 ( 
.A(n_5241),
.Y(n_5390)
);

NAND2xp5_ASAP7_75t_L g5391 ( 
.A(n_5294),
.B(n_1084),
.Y(n_5391)
);

AOI221xp5_ASAP7_75t_L g5392 ( 
.A1(n_5311),
.A2(n_1596),
.B1(n_1597),
.B2(n_1595),
.C(n_1594),
.Y(n_5392)
);

OAI21xp33_ASAP7_75t_L g5393 ( 
.A1(n_5263),
.A2(n_1086),
.B(n_1087),
.Y(n_5393)
);

AOI22xp5_ASAP7_75t_L g5394 ( 
.A1(n_5342),
.A2(n_1090),
.B1(n_1087),
.B2(n_1089),
.Y(n_5394)
);

A2O1A1Ixp33_ASAP7_75t_L g5395 ( 
.A1(n_5275),
.A2(n_1093),
.B(n_1090),
.C(n_1091),
.Y(n_5395)
);

NAND2xp5_ASAP7_75t_SL g5396 ( 
.A(n_5261),
.B(n_1091),
.Y(n_5396)
);

AOI221xp5_ASAP7_75t_L g5397 ( 
.A1(n_5334),
.A2(n_1587),
.B1(n_1588),
.B2(n_1586),
.C(n_1585),
.Y(n_5397)
);

AOI22xp5_ASAP7_75t_L g5398 ( 
.A1(n_5240),
.A2(n_1590),
.B1(n_1592),
.B2(n_1589),
.Y(n_5398)
);

INVx1_ASAP7_75t_L g5399 ( 
.A(n_5286),
.Y(n_5399)
);

AOI22xp33_ASAP7_75t_SL g5400 ( 
.A1(n_5328),
.A2(n_1097),
.B1(n_1094),
.B2(n_1096),
.Y(n_5400)
);

AOI21xp5_ASAP7_75t_L g5401 ( 
.A1(n_5246),
.A2(n_1098),
.B(n_1099),
.Y(n_5401)
);

NAND3xp33_ASAP7_75t_L g5402 ( 
.A(n_5303),
.B(n_1098),
.C(n_1100),
.Y(n_5402)
);

AOI22xp33_ASAP7_75t_L g5403 ( 
.A1(n_5302),
.A2(n_5250),
.B1(n_5248),
.B2(n_5272),
.Y(n_5403)
);

INVx3_ASAP7_75t_L g5404 ( 
.A(n_5291),
.Y(n_5404)
);

INVx1_ASAP7_75t_L g5405 ( 
.A(n_5274),
.Y(n_5405)
);

AOI21xp5_ASAP7_75t_L g5406 ( 
.A1(n_5301),
.A2(n_1101),
.B(n_1102),
.Y(n_5406)
);

AOI21xp5_ASAP7_75t_L g5407 ( 
.A1(n_5253),
.A2(n_1102),
.B(n_1103),
.Y(n_5407)
);

INVx1_ASAP7_75t_L g5408 ( 
.A(n_5277),
.Y(n_5408)
);

INVxp67_ASAP7_75t_L g5409 ( 
.A(n_5262),
.Y(n_5409)
);

INVx1_ASAP7_75t_L g5410 ( 
.A(n_5278),
.Y(n_5410)
);

OAI221xp5_ASAP7_75t_L g5411 ( 
.A1(n_5313),
.A2(n_1592),
.B1(n_1593),
.B2(n_1587),
.C(n_1585),
.Y(n_5411)
);

NAND3xp33_ASAP7_75t_SL g5412 ( 
.A(n_5235),
.B(n_1108),
.C(n_1109),
.Y(n_5412)
);

OAI21xp5_ASAP7_75t_L g5413 ( 
.A1(n_5293),
.A2(n_1111),
.B(n_1110),
.Y(n_5413)
);

INVx1_ASAP7_75t_L g5414 ( 
.A(n_5255),
.Y(n_5414)
);

INVx1_ASAP7_75t_L g5415 ( 
.A(n_5260),
.Y(n_5415)
);

OAI32xp33_ASAP7_75t_L g5416 ( 
.A1(n_5295),
.A2(n_1126),
.A3(n_1134),
.B1(n_1118),
.B2(n_1114),
.Y(n_5416)
);

INVx2_ASAP7_75t_L g5417 ( 
.A(n_5280),
.Y(n_5417)
);

INVx2_ASAP7_75t_SL g5418 ( 
.A(n_5251),
.Y(n_5418)
);

INVx1_ASAP7_75t_L g5419 ( 
.A(n_5279),
.Y(n_5419)
);

INVx1_ASAP7_75t_SL g5420 ( 
.A(n_5300),
.Y(n_5420)
);

INVx1_ASAP7_75t_L g5421 ( 
.A(n_5283),
.Y(n_5421)
);

NAND2xp5_ASAP7_75t_SL g5422 ( 
.A(n_5271),
.B(n_1116),
.Y(n_5422)
);

OAI21xp33_ASAP7_75t_L g5423 ( 
.A1(n_5287),
.A2(n_1119),
.B(n_1120),
.Y(n_5423)
);

AOI221xp5_ASAP7_75t_L g5424 ( 
.A1(n_5357),
.A2(n_5297),
.B1(n_5312),
.B2(n_5336),
.C(n_5316),
.Y(n_5424)
);

AOI221xp5_ASAP7_75t_L g5425 ( 
.A1(n_5386),
.A2(n_5242),
.B1(n_5256),
.B2(n_5317),
.C(n_5298),
.Y(n_5425)
);

NAND2xp5_ASAP7_75t_L g5426 ( 
.A(n_5356),
.B(n_5332),
.Y(n_5426)
);

INVx1_ASAP7_75t_L g5427 ( 
.A(n_5343),
.Y(n_5427)
);

OAI221xp5_ASAP7_75t_SL g5428 ( 
.A1(n_5344),
.A2(n_5282),
.B1(n_5284),
.B2(n_5299),
.C(n_5267),
.Y(n_5428)
);

OAI22xp5_ASAP7_75t_L g5429 ( 
.A1(n_5350),
.A2(n_5289),
.B1(n_5288),
.B2(n_5269),
.Y(n_5429)
);

AOI222xp33_ASAP7_75t_L g5430 ( 
.A1(n_5396),
.A2(n_5412),
.B1(n_5382),
.B2(n_5351),
.C1(n_5402),
.C2(n_5374),
.Y(n_5430)
);

NAND2xp5_ASAP7_75t_L g5431 ( 
.A(n_5404),
.B(n_5247),
.Y(n_5431)
);

NAND2xp5_ASAP7_75t_L g5432 ( 
.A(n_5404),
.B(n_1120),
.Y(n_5432)
);

NAND2xp5_ASAP7_75t_L g5433 ( 
.A(n_5371),
.B(n_1124),
.Y(n_5433)
);

OAI221xp5_ASAP7_75t_L g5434 ( 
.A1(n_5346),
.A2(n_1127),
.B1(n_1124),
.B2(n_1126),
.C(n_1129),
.Y(n_5434)
);

OAI221xp5_ASAP7_75t_L g5435 ( 
.A1(n_5409),
.A2(n_1131),
.B1(n_1129),
.B2(n_1130),
.C(n_1132),
.Y(n_5435)
);

A2O1A1Ixp33_ASAP7_75t_L g5436 ( 
.A1(n_5395),
.A2(n_5406),
.B(n_5373),
.C(n_5348),
.Y(n_5436)
);

AOI21xp5_ASAP7_75t_L g5437 ( 
.A1(n_5422),
.A2(n_5407),
.B(n_5401),
.Y(n_5437)
);

OAI221xp5_ASAP7_75t_L g5438 ( 
.A1(n_5403),
.A2(n_1138),
.B1(n_1136),
.B2(n_1137),
.C(n_1139),
.Y(n_5438)
);

OAI221xp5_ASAP7_75t_L g5439 ( 
.A1(n_5355),
.A2(n_1140),
.B1(n_1138),
.B2(n_1139),
.C(n_1141),
.Y(n_5439)
);

AOI22xp5_ASAP7_75t_L g5440 ( 
.A1(n_5352),
.A2(n_1142),
.B1(n_1140),
.B2(n_1141),
.Y(n_5440)
);

OAI321xp33_ASAP7_75t_L g5441 ( 
.A1(n_5364),
.A2(n_5368),
.A3(n_5365),
.B1(n_5363),
.B2(n_5381),
.C(n_5354),
.Y(n_5441)
);

AOI22xp5_ASAP7_75t_L g5442 ( 
.A1(n_5353),
.A2(n_1146),
.B1(n_1144),
.B2(n_1145),
.Y(n_5442)
);

OAI211xp5_ASAP7_75t_L g5443 ( 
.A1(n_5388),
.A2(n_1147),
.B(n_1145),
.C(n_1146),
.Y(n_5443)
);

OAI21xp33_ASAP7_75t_L g5444 ( 
.A1(n_5417),
.A2(n_1148),
.B(n_1149),
.Y(n_5444)
);

AOI31xp33_ASAP7_75t_L g5445 ( 
.A1(n_5413),
.A2(n_1150),
.A3(n_1148),
.B(n_1149),
.Y(n_5445)
);

NAND2xp5_ASAP7_75t_SL g5446 ( 
.A(n_5390),
.B(n_1152),
.Y(n_5446)
);

NOR2xp67_ASAP7_75t_L g5447 ( 
.A(n_5390),
.B(n_1153),
.Y(n_5447)
);

NAND3x1_ASAP7_75t_L g5448 ( 
.A(n_5358),
.B(n_1157),
.C(n_1158),
.Y(n_5448)
);

OAI22xp5_ASAP7_75t_L g5449 ( 
.A1(n_5394),
.A2(n_1159),
.B1(n_1157),
.B2(n_1158),
.Y(n_5449)
);

AOI21xp33_ASAP7_75t_L g5450 ( 
.A1(n_5383),
.A2(n_5372),
.B(n_5370),
.Y(n_5450)
);

INVx1_ASAP7_75t_L g5451 ( 
.A(n_5375),
.Y(n_5451)
);

OAI21xp5_ASAP7_75t_SL g5452 ( 
.A1(n_5420),
.A2(n_1161),
.B(n_1162),
.Y(n_5452)
);

O2A1O1Ixp33_ASAP7_75t_SL g5453 ( 
.A1(n_5391),
.A2(n_1164),
.B(n_1162),
.C(n_1163),
.Y(n_5453)
);

AOI22xp5_ASAP7_75t_L g5454 ( 
.A1(n_5369),
.A2(n_1166),
.B1(n_1163),
.B2(n_1165),
.Y(n_5454)
);

AOI21xp33_ASAP7_75t_SL g5455 ( 
.A1(n_5376),
.A2(n_1169),
.B(n_1168),
.Y(n_5455)
);

OAI221xp5_ASAP7_75t_L g5456 ( 
.A1(n_5400),
.A2(n_1170),
.B1(n_1167),
.B2(n_1169),
.C(n_1171),
.Y(n_5456)
);

NAND3xp33_ASAP7_75t_L g5457 ( 
.A(n_5389),
.B(n_1172),
.C(n_1173),
.Y(n_5457)
);

INVx2_ASAP7_75t_L g5458 ( 
.A(n_5385),
.Y(n_5458)
);

OAI221xp5_ASAP7_75t_L g5459 ( 
.A1(n_5399),
.A2(n_5410),
.B1(n_5408),
.B2(n_5360),
.C(n_5415),
.Y(n_5459)
);

NAND3xp33_ASAP7_75t_L g5460 ( 
.A(n_5392),
.B(n_1174),
.C(n_1175),
.Y(n_5460)
);

XNOR2x1_ASAP7_75t_L g5461 ( 
.A(n_5377),
.B(n_1175),
.Y(n_5461)
);

NOR2xp33_ASAP7_75t_L g5462 ( 
.A(n_5393),
.B(n_5411),
.Y(n_5462)
);

OAI21xp5_ASAP7_75t_L g5463 ( 
.A1(n_5366),
.A2(n_1174),
.B(n_1176),
.Y(n_5463)
);

INVx1_ASAP7_75t_L g5464 ( 
.A(n_5367),
.Y(n_5464)
);

OAI21xp5_ASAP7_75t_L g5465 ( 
.A1(n_5347),
.A2(n_1177),
.B(n_1179),
.Y(n_5465)
);

AOI211xp5_ASAP7_75t_L g5466 ( 
.A1(n_5384),
.A2(n_5416),
.B(n_5387),
.C(n_5378),
.Y(n_5466)
);

AOI21xp5_ASAP7_75t_L g5467 ( 
.A1(n_5418),
.A2(n_1181),
.B(n_1182),
.Y(n_5467)
);

AOI222xp33_ASAP7_75t_L g5468 ( 
.A1(n_5397),
.A2(n_1186),
.B1(n_1188),
.B2(n_1183),
.C1(n_1185),
.C2(n_1187),
.Y(n_5468)
);

INVx1_ASAP7_75t_L g5469 ( 
.A(n_5361),
.Y(n_5469)
);

AOI211xp5_ASAP7_75t_SL g5470 ( 
.A1(n_5405),
.A2(n_1194),
.B(n_1192),
.C(n_1193),
.Y(n_5470)
);

AOI21xp5_ASAP7_75t_L g5471 ( 
.A1(n_5414),
.A2(n_1195),
.B(n_1198),
.Y(n_5471)
);

AOI211xp5_ASAP7_75t_L g5472 ( 
.A1(n_5419),
.A2(n_5421),
.B(n_5379),
.C(n_5423),
.Y(n_5472)
);

INVx1_ASAP7_75t_L g5473 ( 
.A(n_5362),
.Y(n_5473)
);

AOI21xp5_ASAP7_75t_SL g5474 ( 
.A1(n_5398),
.A2(n_1203),
.B(n_1207),
.Y(n_5474)
);

OAI221xp5_ASAP7_75t_L g5475 ( 
.A1(n_5345),
.A2(n_1210),
.B1(n_1208),
.B2(n_1209),
.C(n_1212),
.Y(n_5475)
);

NOR3xp33_ASAP7_75t_SL g5476 ( 
.A(n_5357),
.B(n_1212),
.C(n_1213),
.Y(n_5476)
);

OAI211xp5_ASAP7_75t_L g5477 ( 
.A1(n_5345),
.A2(n_1216),
.B(n_1214),
.C(n_1215),
.Y(n_5477)
);

NAND2xp5_ASAP7_75t_L g5478 ( 
.A(n_5356),
.B(n_1217),
.Y(n_5478)
);

AND2x2_ASAP7_75t_L g5479 ( 
.A(n_5359),
.B(n_1218),
.Y(n_5479)
);

OAI221xp5_ASAP7_75t_SL g5480 ( 
.A1(n_5344),
.A2(n_1598),
.B1(n_1601),
.B2(n_1584),
.C(n_1583),
.Y(n_5480)
);

NAND2xp5_ASAP7_75t_L g5481 ( 
.A(n_5356),
.B(n_1222),
.Y(n_5481)
);

NAND2xp5_ASAP7_75t_L g5482 ( 
.A(n_5356),
.B(n_1223),
.Y(n_5482)
);

NAND2xp5_ASAP7_75t_L g5483 ( 
.A(n_5356),
.B(n_1223),
.Y(n_5483)
);

NAND3xp33_ASAP7_75t_L g5484 ( 
.A(n_5345),
.B(n_1224),
.C(n_1227),
.Y(n_5484)
);

NAND2xp5_ASAP7_75t_SL g5485 ( 
.A(n_5356),
.B(n_1227),
.Y(n_5485)
);

NAND3xp33_ASAP7_75t_L g5486 ( 
.A(n_5345),
.B(n_1228),
.C(n_1229),
.Y(n_5486)
);

NAND3xp33_ASAP7_75t_L g5487 ( 
.A(n_5345),
.B(n_1228),
.C(n_1229),
.Y(n_5487)
);

OAI22xp5_ASAP7_75t_L g5488 ( 
.A1(n_5350),
.A2(n_1233),
.B1(n_1230),
.B2(n_1231),
.Y(n_5488)
);

OAI21xp5_ASAP7_75t_SL g5489 ( 
.A1(n_5345),
.A2(n_1234),
.B(n_1235),
.Y(n_5489)
);

OAI221xp5_ASAP7_75t_SL g5490 ( 
.A1(n_5344),
.A2(n_1582),
.B1(n_1239),
.B2(n_1236),
.C(n_1238),
.Y(n_5490)
);

A2O1A1Ixp33_ASAP7_75t_L g5491 ( 
.A1(n_5349),
.A2(n_1246),
.B(n_1253),
.C(n_1238),
.Y(n_5491)
);

NOR2xp33_ASAP7_75t_L g5492 ( 
.A(n_5380),
.B(n_1239),
.Y(n_5492)
);

OAI32xp33_ASAP7_75t_L g5493 ( 
.A1(n_5345),
.A2(n_1243),
.A3(n_1245),
.B1(n_1241),
.B2(n_1244),
.Y(n_5493)
);

OAI21xp5_ASAP7_75t_L g5494 ( 
.A1(n_5345),
.A2(n_1250),
.B(n_1251),
.Y(n_5494)
);

NAND2xp5_ASAP7_75t_L g5495 ( 
.A(n_5356),
.B(n_1253),
.Y(n_5495)
);

OAI21xp33_ASAP7_75t_SL g5496 ( 
.A1(n_5345),
.A2(n_1254),
.B(n_1255),
.Y(n_5496)
);

OAI221xp5_ASAP7_75t_L g5497 ( 
.A1(n_5345),
.A2(n_1259),
.B1(n_1257),
.B2(n_1258),
.C(n_1260),
.Y(n_5497)
);

NAND3xp33_ASAP7_75t_L g5498 ( 
.A(n_5345),
.B(n_1261),
.C(n_1262),
.Y(n_5498)
);

NAND2xp5_ASAP7_75t_L g5499 ( 
.A(n_5356),
.B(n_1261),
.Y(n_5499)
);

OAI221xp5_ASAP7_75t_L g5500 ( 
.A1(n_5345),
.A2(n_1266),
.B1(n_1264),
.B2(n_1265),
.C(n_1267),
.Y(n_5500)
);

NAND2xp5_ASAP7_75t_SL g5501 ( 
.A(n_5356),
.B(n_1267),
.Y(n_5501)
);

OAI221xp5_ASAP7_75t_L g5502 ( 
.A1(n_5345),
.A2(n_1270),
.B1(n_1268),
.B2(n_1269),
.C(n_1271),
.Y(n_5502)
);

AOI21xp5_ASAP7_75t_L g5503 ( 
.A1(n_5345),
.A2(n_1268),
.B(n_1269),
.Y(n_5503)
);

NAND2xp5_ASAP7_75t_L g5504 ( 
.A(n_5356),
.B(n_1271),
.Y(n_5504)
);

NAND2xp5_ASAP7_75t_SL g5505 ( 
.A(n_5356),
.B(n_1272),
.Y(n_5505)
);

NOR2x1_ASAP7_75t_L g5506 ( 
.A(n_5447),
.B(n_1272),
.Y(n_5506)
);

INVx1_ASAP7_75t_L g5507 ( 
.A(n_5479),
.Y(n_5507)
);

AOI322xp5_ASAP7_75t_L g5508 ( 
.A1(n_5476),
.A2(n_1280),
.A3(n_1279),
.B1(n_1277),
.B2(n_1274),
.C1(n_1276),
.C2(n_1278),
.Y(n_5508)
);

NOR3xp33_ASAP7_75t_SL g5509 ( 
.A(n_5441),
.B(n_1277),
.C(n_1278),
.Y(n_5509)
);

AOI221xp5_ASAP7_75t_L g5510 ( 
.A1(n_5424),
.A2(n_1285),
.B1(n_1287),
.B2(n_1282),
.C(n_1286),
.Y(n_5510)
);

OAI221xp5_ASAP7_75t_SL g5511 ( 
.A1(n_5427),
.A2(n_1287),
.B1(n_1281),
.B2(n_1286),
.C(n_1288),
.Y(n_5511)
);

OR2x2_ASAP7_75t_L g5512 ( 
.A(n_5426),
.B(n_1289),
.Y(n_5512)
);

NAND2xp5_ASAP7_75t_SL g5513 ( 
.A(n_5455),
.B(n_1289),
.Y(n_5513)
);

AND2x2_ASAP7_75t_L g5514 ( 
.A(n_5458),
.B(n_1290),
.Y(n_5514)
);

OAI211xp5_ASAP7_75t_L g5515 ( 
.A1(n_5430),
.A2(n_1293),
.B(n_1291),
.C(n_1292),
.Y(n_5515)
);

NOR2xp33_ASAP7_75t_L g5516 ( 
.A(n_5496),
.B(n_1291),
.Y(n_5516)
);

AOI21xp33_ASAP7_75t_SL g5517 ( 
.A1(n_5485),
.A2(n_5505),
.B(n_5501),
.Y(n_5517)
);

AOI22xp5_ASAP7_75t_L g5518 ( 
.A1(n_5462),
.A2(n_1296),
.B1(n_1294),
.B2(n_1295),
.Y(n_5518)
);

AOI222xp33_ASAP7_75t_L g5519 ( 
.A1(n_5429),
.A2(n_1297),
.B1(n_1300),
.B2(n_1295),
.C1(n_1296),
.C2(n_1298),
.Y(n_5519)
);

O2A1O1Ixp33_ASAP7_75t_SL g5520 ( 
.A1(n_5491),
.A2(n_1303),
.B(n_1301),
.C(n_1302),
.Y(n_5520)
);

INVxp67_ASAP7_75t_L g5521 ( 
.A(n_5492),
.Y(n_5521)
);

OAI321xp33_ASAP7_75t_L g5522 ( 
.A1(n_5428),
.A2(n_1306),
.A3(n_1308),
.B1(n_1304),
.B2(n_1305),
.C(n_1307),
.Y(n_5522)
);

NAND2xp5_ASAP7_75t_L g5523 ( 
.A(n_5470),
.B(n_1308),
.Y(n_5523)
);

OAI221xp5_ASAP7_75t_SL g5524 ( 
.A1(n_5466),
.A2(n_1312),
.B1(n_1310),
.B2(n_1311),
.C(n_1313),
.Y(n_5524)
);

AOI22xp5_ASAP7_75t_L g5525 ( 
.A1(n_5473),
.A2(n_1315),
.B1(n_1312),
.B2(n_1314),
.Y(n_5525)
);

NAND2x1_ASAP7_75t_L g5526 ( 
.A(n_5474),
.B(n_1315),
.Y(n_5526)
);

NAND4xp25_ASAP7_75t_L g5527 ( 
.A(n_5472),
.B(n_5450),
.C(n_5431),
.D(n_5437),
.Y(n_5527)
);

AOI22xp33_ASAP7_75t_L g5528 ( 
.A1(n_5469),
.A2(n_1321),
.B1(n_1316),
.B2(n_1320),
.Y(n_5528)
);

INVx1_ASAP7_75t_L g5529 ( 
.A(n_5432),
.Y(n_5529)
);

INVx2_ASAP7_75t_L g5530 ( 
.A(n_5448),
.Y(n_5530)
);

NOR2xp33_ASAP7_75t_L g5531 ( 
.A(n_5477),
.B(n_1321),
.Y(n_5531)
);

AOI21xp5_ASAP7_75t_L g5532 ( 
.A1(n_5446),
.A2(n_1322),
.B(n_1323),
.Y(n_5532)
);

OAI21xp5_ASAP7_75t_SL g5533 ( 
.A1(n_5489),
.A2(n_1322),
.B(n_1324),
.Y(n_5533)
);

AOI322xp5_ASAP7_75t_L g5534 ( 
.A1(n_5425),
.A2(n_1330),
.A3(n_1329),
.B1(n_1327),
.B2(n_1325),
.C1(n_1326),
.C2(n_1328),
.Y(n_5534)
);

INVx1_ASAP7_75t_L g5535 ( 
.A(n_5478),
.Y(n_5535)
);

OAI322xp33_ASAP7_75t_L g5536 ( 
.A1(n_5459),
.A2(n_1332),
.A3(n_1331),
.B1(n_1329),
.B2(n_1326),
.C1(n_1327),
.C2(n_1330),
.Y(n_5536)
);

INVx1_ASAP7_75t_L g5537 ( 
.A(n_5481),
.Y(n_5537)
);

OAI22xp5_ASAP7_75t_L g5538 ( 
.A1(n_5436),
.A2(n_5484),
.B1(n_5487),
.B2(n_5486),
.Y(n_5538)
);

AND2x2_ASAP7_75t_L g5539 ( 
.A(n_5465),
.B(n_1333),
.Y(n_5539)
);

AOI221xp5_ASAP7_75t_L g5540 ( 
.A1(n_5493),
.A2(n_1336),
.B1(n_1338),
.B2(n_1335),
.C(n_1337),
.Y(n_5540)
);

OAI32xp33_ASAP7_75t_L g5541 ( 
.A1(n_5433),
.A2(n_1339),
.A3(n_1334),
.B1(n_1337),
.B2(n_1340),
.Y(n_5541)
);

NOR2xp33_ASAP7_75t_L g5542 ( 
.A(n_5452),
.B(n_1339),
.Y(n_5542)
);

OAI32xp33_ASAP7_75t_L g5543 ( 
.A1(n_5482),
.A2(n_1347),
.A3(n_1344),
.B1(n_1345),
.B2(n_1348),
.Y(n_5543)
);

NOR2xp33_ASAP7_75t_L g5544 ( 
.A(n_5483),
.B(n_1344),
.Y(n_5544)
);

INVx1_ASAP7_75t_L g5545 ( 
.A(n_5495),
.Y(n_5545)
);

AOI21xp5_ASAP7_75t_L g5546 ( 
.A1(n_5453),
.A2(n_1350),
.B(n_1353),
.Y(n_5546)
);

INVx1_ASAP7_75t_L g5547 ( 
.A(n_5499),
.Y(n_5547)
);

AOI211xp5_ASAP7_75t_L g5548 ( 
.A1(n_5443),
.A2(n_1355),
.B(n_1350),
.C(n_1354),
.Y(n_5548)
);

AOI221xp5_ASAP7_75t_L g5549 ( 
.A1(n_5457),
.A2(n_5494),
.B1(n_5503),
.B2(n_5498),
.C(n_5445),
.Y(n_5549)
);

AOI221xp5_ASAP7_75t_L g5550 ( 
.A1(n_5475),
.A2(n_1357),
.B1(n_1359),
.B2(n_1356),
.C(n_1358),
.Y(n_5550)
);

INVx1_ASAP7_75t_L g5551 ( 
.A(n_5504),
.Y(n_5551)
);

AOI22xp33_ASAP7_75t_L g5552 ( 
.A1(n_5464),
.A2(n_1357),
.B1(n_1354),
.B2(n_1356),
.Y(n_5552)
);

AND2x2_ASAP7_75t_L g5553 ( 
.A(n_5451),
.B(n_1360),
.Y(n_5553)
);

INVx1_ASAP7_75t_SL g5554 ( 
.A(n_5461),
.Y(n_5554)
);

AOI22xp33_ASAP7_75t_L g5555 ( 
.A1(n_5460),
.A2(n_1364),
.B1(n_1362),
.B2(n_1363),
.Y(n_5555)
);

NAND2xp5_ASAP7_75t_L g5556 ( 
.A(n_5467),
.B(n_1365),
.Y(n_5556)
);

AOI211xp5_ASAP7_75t_L g5557 ( 
.A1(n_5524),
.A2(n_5500),
.B(n_5502),
.C(n_5497),
.Y(n_5557)
);

INVx2_ASAP7_75t_L g5558 ( 
.A(n_5506),
.Y(n_5558)
);

AOI211xp5_ASAP7_75t_SL g5559 ( 
.A1(n_5522),
.A2(n_5480),
.B(n_5490),
.C(n_5438),
.Y(n_5559)
);

AOI211xp5_ASAP7_75t_L g5560 ( 
.A1(n_5517),
.A2(n_5456),
.B(n_5434),
.C(n_5449),
.Y(n_5560)
);

OAI21xp33_ASAP7_75t_L g5561 ( 
.A1(n_5527),
.A2(n_5444),
.B(n_5468),
.Y(n_5561)
);

AOI21xp5_ASAP7_75t_L g5562 ( 
.A1(n_5513),
.A2(n_5471),
.B(n_5463),
.Y(n_5562)
);

INVxp33_ASAP7_75t_L g5563 ( 
.A(n_5526),
.Y(n_5563)
);

OAI22xp5_ASAP7_75t_L g5564 ( 
.A1(n_5555),
.A2(n_5528),
.B1(n_5525),
.B2(n_5512),
.Y(n_5564)
);

INVx2_ASAP7_75t_L g5565 ( 
.A(n_5530),
.Y(n_5565)
);

INVxp33_ASAP7_75t_SL g5566 ( 
.A(n_5538),
.Y(n_5566)
);

INVx1_ASAP7_75t_L g5567 ( 
.A(n_5514),
.Y(n_5567)
);

AOI211xp5_ASAP7_75t_L g5568 ( 
.A1(n_5515),
.A2(n_5435),
.B(n_5439),
.C(n_5488),
.Y(n_5568)
);

CKINVDCx5p33_ASAP7_75t_R g5569 ( 
.A(n_5509),
.Y(n_5569)
);

NAND4xp25_ASAP7_75t_L g5570 ( 
.A(n_5549),
.B(n_5454),
.C(n_5442),
.D(n_5440),
.Y(n_5570)
);

OAI22xp33_ASAP7_75t_L g5571 ( 
.A1(n_5523),
.A2(n_1367),
.B1(n_1369),
.B2(n_1366),
.Y(n_5571)
);

OAI21xp33_ASAP7_75t_L g5572 ( 
.A1(n_5554),
.A2(n_1370),
.B(n_1371),
.Y(n_5572)
);

INVx1_ASAP7_75t_L g5573 ( 
.A(n_5507),
.Y(n_5573)
);

NAND2xp5_ASAP7_75t_L g5574 ( 
.A(n_5508),
.B(n_5546),
.Y(n_5574)
);

INVx1_ASAP7_75t_L g5575 ( 
.A(n_5556),
.Y(n_5575)
);

OAI21xp33_ASAP7_75t_SL g5576 ( 
.A1(n_5535),
.A2(n_1372),
.B(n_1375),
.Y(n_5576)
);

AOI21xp5_ASAP7_75t_L g5577 ( 
.A1(n_5520),
.A2(n_5532),
.B(n_5516),
.Y(n_5577)
);

OAI22xp5_ASAP7_75t_L g5578 ( 
.A1(n_5548),
.A2(n_1380),
.B1(n_1377),
.B2(n_1379),
.Y(n_5578)
);

NAND5xp2_ASAP7_75t_L g5579 ( 
.A(n_5537),
.B(n_1581),
.C(n_1383),
.D(n_1381),
.E(n_1382),
.Y(n_5579)
);

OAI221xp5_ASAP7_75t_SL g5580 ( 
.A1(n_5533),
.A2(n_1386),
.B1(n_1384),
.B2(n_1385),
.C(n_1387),
.Y(n_5580)
);

NAND3xp33_ASAP7_75t_L g5581 ( 
.A(n_5510),
.B(n_1386),
.C(n_1388),
.Y(n_5581)
);

INVx2_ASAP7_75t_L g5582 ( 
.A(n_5553),
.Y(n_5582)
);

INVx1_ASAP7_75t_L g5583 ( 
.A(n_5539),
.Y(n_5583)
);

AOI22xp33_ASAP7_75t_L g5584 ( 
.A1(n_5545),
.A2(n_1392),
.B1(n_1389),
.B2(n_1391),
.Y(n_5584)
);

NOR2x1_ASAP7_75t_L g5585 ( 
.A(n_5536),
.B(n_1392),
.Y(n_5585)
);

BUFx6f_ASAP7_75t_L g5586 ( 
.A(n_5529),
.Y(n_5586)
);

AOI211xp5_ASAP7_75t_L g5587 ( 
.A1(n_5543),
.A2(n_1396),
.B(n_1394),
.C(n_1395),
.Y(n_5587)
);

NAND2xp5_ASAP7_75t_SL g5588 ( 
.A(n_5519),
.B(n_1397),
.Y(n_5588)
);

AOI211xp5_ASAP7_75t_L g5589 ( 
.A1(n_5563),
.A2(n_5541),
.B(n_5551),
.C(n_5547),
.Y(n_5589)
);

NOR2xp67_ASAP7_75t_L g5590 ( 
.A(n_5576),
.B(n_5521),
.Y(n_5590)
);

AOI211xp5_ASAP7_75t_SL g5591 ( 
.A1(n_5561),
.A2(n_5531),
.B(n_5511),
.C(n_5544),
.Y(n_5591)
);

NAND2xp5_ASAP7_75t_L g5592 ( 
.A(n_5558),
.B(n_5534),
.Y(n_5592)
);

AOI22xp5_ASAP7_75t_L g5593 ( 
.A1(n_5566),
.A2(n_5542),
.B1(n_5540),
.B2(n_5550),
.Y(n_5593)
);

OAI22xp33_ASAP7_75t_L g5594 ( 
.A1(n_5559),
.A2(n_5518),
.B1(n_5552),
.B2(n_1400),
.Y(n_5594)
);

NAND2xp5_ASAP7_75t_L g5595 ( 
.A(n_5569),
.B(n_1398),
.Y(n_5595)
);

O2A1O1Ixp33_ASAP7_75t_L g5596 ( 
.A1(n_5588),
.A2(n_1405),
.B(n_1403),
.C(n_1404),
.Y(n_5596)
);

A2O1A1Ixp33_ASAP7_75t_L g5597 ( 
.A1(n_5562),
.A2(n_5577),
.B(n_5572),
.C(n_5565),
.Y(n_5597)
);

NAND2xp5_ASAP7_75t_L g5598 ( 
.A(n_5587),
.B(n_1406),
.Y(n_5598)
);

INVx1_ASAP7_75t_L g5599 ( 
.A(n_5567),
.Y(n_5599)
);

XOR2xp5_ASAP7_75t_L g5600 ( 
.A(n_5570),
.B(n_1406),
.Y(n_5600)
);

NAND2xp5_ASAP7_75t_L g5601 ( 
.A(n_5585),
.B(n_1407),
.Y(n_5601)
);

INVx2_ASAP7_75t_L g5602 ( 
.A(n_5586),
.Y(n_5602)
);

AOI21xp33_ASAP7_75t_SL g5603 ( 
.A1(n_5571),
.A2(n_1409),
.B(n_1410),
.Y(n_5603)
);

NOR2xp33_ASAP7_75t_L g5604 ( 
.A(n_5579),
.B(n_1410),
.Y(n_5604)
);

AO22x2_ASAP7_75t_L g5605 ( 
.A1(n_5600),
.A2(n_5573),
.B1(n_5582),
.B2(n_5583),
.Y(n_5605)
);

INVx1_ASAP7_75t_L g5606 ( 
.A(n_5601),
.Y(n_5606)
);

HB1xp67_ASAP7_75t_L g5607 ( 
.A(n_5590),
.Y(n_5607)
);

NAND4xp25_ASAP7_75t_L g5608 ( 
.A(n_5591),
.B(n_5560),
.C(n_5557),
.D(n_5568),
.Y(n_5608)
);

INVx1_ASAP7_75t_L g5609 ( 
.A(n_5595),
.Y(n_5609)
);

AOI22xp5_ASAP7_75t_L g5610 ( 
.A1(n_5604),
.A2(n_5564),
.B1(n_5574),
.B2(n_5578),
.Y(n_5610)
);

OR2x2_ASAP7_75t_L g5611 ( 
.A(n_5602),
.B(n_5580),
.Y(n_5611)
);

INVx1_ASAP7_75t_L g5612 ( 
.A(n_5598),
.Y(n_5612)
);

INVx1_ASAP7_75t_L g5613 ( 
.A(n_5592),
.Y(n_5613)
);

OAI22xp5_ASAP7_75t_SL g5614 ( 
.A1(n_5593),
.A2(n_5575),
.B1(n_5581),
.B2(n_5584),
.Y(n_5614)
);

XNOR2xp5_ASAP7_75t_L g5615 ( 
.A(n_5610),
.B(n_5589),
.Y(n_5615)
);

INVx1_ASAP7_75t_L g5616 ( 
.A(n_5607),
.Y(n_5616)
);

NOR3xp33_ASAP7_75t_L g5617 ( 
.A(n_5608),
.B(n_5597),
.C(n_5614),
.Y(n_5617)
);

NOR3xp33_ASAP7_75t_L g5618 ( 
.A(n_5613),
.B(n_5599),
.C(n_5594),
.Y(n_5618)
);

INVx1_ASAP7_75t_L g5619 ( 
.A(n_5605),
.Y(n_5619)
);

INVx1_ASAP7_75t_L g5620 ( 
.A(n_5605),
.Y(n_5620)
);

NOR2x1_ASAP7_75t_L g5621 ( 
.A(n_5611),
.B(n_5596),
.Y(n_5621)
);

NOR2xp67_ASAP7_75t_SL g5622 ( 
.A(n_5606),
.B(n_5603),
.Y(n_5622)
);

AOI221xp5_ASAP7_75t_L g5623 ( 
.A1(n_5619),
.A2(n_5620),
.B1(n_5617),
.B2(n_5618),
.C(n_5616),
.Y(n_5623)
);

OA22x2_ASAP7_75t_L g5624 ( 
.A1(n_5615),
.A2(n_5609),
.B1(n_5612),
.B2(n_1412),
.Y(n_5624)
);

NOR3xp33_ASAP7_75t_L g5625 ( 
.A(n_5621),
.B(n_1415),
.C(n_1416),
.Y(n_5625)
);

AND4x1_ASAP7_75t_L g5626 ( 
.A(n_5622),
.B(n_1420),
.C(n_1418),
.D(n_1419),
.Y(n_5626)
);

INVx3_ASAP7_75t_L g5627 ( 
.A(n_5626),
.Y(n_5627)
);

INVx1_ASAP7_75t_L g5628 ( 
.A(n_5624),
.Y(n_5628)
);

INVx2_ASAP7_75t_L g5629 ( 
.A(n_5627),
.Y(n_5629)
);

AOI22xp33_ASAP7_75t_L g5630 ( 
.A1(n_5629),
.A2(n_5623),
.B1(n_5628),
.B2(n_5625),
.Y(n_5630)
);

INVx1_ASAP7_75t_L g5631 ( 
.A(n_5630),
.Y(n_5631)
);

NOR2xp67_ASAP7_75t_L g5632 ( 
.A(n_5631),
.B(n_1422),
.Y(n_5632)
);

AOI22xp33_ASAP7_75t_L g5633 ( 
.A1(n_5632),
.A2(n_1427),
.B1(n_1425),
.B2(n_1426),
.Y(n_5633)
);

AOI21xp33_ASAP7_75t_SL g5634 ( 
.A1(n_5633),
.A2(n_1429),
.B(n_1430),
.Y(n_5634)
);

AOI21xp5_ASAP7_75t_L g5635 ( 
.A1(n_5634),
.A2(n_1431),
.B(n_1432),
.Y(n_5635)
);

AOI22xp5_ASAP7_75t_L g5636 ( 
.A1(n_5635),
.A2(n_1434),
.B1(n_1432),
.B2(n_1433),
.Y(n_5636)
);

OAI21xp5_ASAP7_75t_L g5637 ( 
.A1(n_5636),
.A2(n_1435),
.B(n_1436),
.Y(n_5637)
);

AOI211xp5_ASAP7_75t_L g5638 ( 
.A1(n_5637),
.A2(n_1440),
.B(n_1438),
.C(n_1439),
.Y(n_5638)
);

AOI211xp5_ASAP7_75t_L g5639 ( 
.A1(n_5638),
.A2(n_1443),
.B(n_1441),
.C(n_1442),
.Y(n_5639)
);


endmodule