module fake_jpeg_3259_n_220 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_220);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_220;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_39),
.Y(n_53)
);

CKINVDCx14_ASAP7_75t_R g54 ( 
.A(n_16),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_29),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_0),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_9),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_46),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_26),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_13),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_4),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_13),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_43),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_16),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_23),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_25),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_35),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_30),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

INVx4_ASAP7_75t_SL g76 ( 
.A(n_66),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_79),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_80),
.A2(n_55),
.B1(n_52),
.B2(n_72),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_0),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_81),
.B(n_62),
.Y(n_85)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_76),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_78),
.A2(n_71),
.B1(n_70),
.B2(n_67),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_83),
.A2(n_80),
.B1(n_77),
.B2(n_74),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_81),
.B(n_56),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_84),
.B(n_87),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_88),
.Y(n_96)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_86),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_82),
.B(n_56),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_82),
.B(n_57),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_79),
.B(n_57),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_89),
.B(n_75),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_76),
.A2(n_67),
.B1(n_70),
.B2(n_71),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_93),
.A2(n_79),
.B1(n_78),
.B2(n_75),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_94),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_94),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_99),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_98),
.A2(n_106),
.B1(n_95),
.B2(n_59),
.Y(n_125)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_95),
.Y(n_100)
);

INVx2_ASAP7_75t_SL g121 ( 
.A(n_100),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_102),
.Y(n_132)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_95),
.Y(n_103)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_103),
.Y(n_119)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_105),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_83),
.A2(n_77),
.B1(n_69),
.B2(n_72),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_87),
.A2(n_88),
.B1(n_89),
.B2(n_92),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_107),
.A2(n_90),
.B1(n_59),
.B2(n_69),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_84),
.B(n_60),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_108),
.B(n_110),
.Y(n_123)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_95),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_109),
.Y(n_117)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_92),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_111),
.B(n_113),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_90),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_85),
.B(n_60),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_61),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_97),
.A2(n_95),
.B1(n_80),
.B2(n_53),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_115),
.A2(n_126),
.B1(n_3),
.B2(n_4),
.Y(n_152)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_120),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_96),
.B(n_104),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_122),
.B(n_124),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_110),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_125),
.A2(n_64),
.B1(n_58),
.B2(n_42),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_105),
.A2(n_90),
.B(n_74),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_127),
.A2(n_130),
.B(n_131),
.Y(n_143)
);

AND2x6_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_50),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_128),
.B(n_133),
.Y(n_136)
);

OAI21xp33_ASAP7_75t_L g130 ( 
.A1(n_107),
.A2(n_73),
.B(n_63),
.Y(n_130)
);

O2A1O1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_106),
.A2(n_73),
.B(n_63),
.C(n_53),
.Y(n_131)
);

AND2x6_ASAP7_75t_L g134 ( 
.A(n_112),
.B(n_48),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_134),
.B(n_45),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_109),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_135),
.B(n_100),
.Y(n_142)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_118),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_137),
.B(n_138),
.Y(n_159)
);

HB1xp67_ASAP7_75t_L g138 ( 
.A(n_121),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_132),
.A2(n_101),
.B1(n_113),
.B2(n_111),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_139),
.A2(n_144),
.B1(n_146),
.B2(n_156),
.Y(n_165)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_121),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_140),
.B(n_145),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_116),
.B(n_103),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_141),
.B(n_131),
.Y(n_160)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_142),
.Y(n_162)
);

OAI22x1_ASAP7_75t_L g144 ( 
.A1(n_120),
.A2(n_58),
.B1(n_54),
.B2(n_68),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_129),
.B(n_1),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_147),
.B(n_149),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_130),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_148),
.A2(n_152),
.B1(n_6),
.B2(n_8),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_115),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_123),
.B(n_2),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_151),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g153 ( 
.A(n_117),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_153),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_117),
.Y(n_154)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_154),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_119),
.B(n_5),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_155),
.A2(n_9),
.B(n_10),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_125),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_143),
.A2(n_134),
.B(n_128),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_158),
.B(n_164),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_160),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_152),
.A2(n_119),
.B1(n_7),
.B2(n_8),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_161),
.A2(n_163),
.B1(n_171),
.B2(n_157),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_141),
.B(n_40),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_166),
.B(n_174),
.C(n_176),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_143),
.A2(n_136),
.B(n_149),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g182 ( 
.A(n_170),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_150),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_156),
.B(n_38),
.Y(n_174)
);

OA22x2_ASAP7_75t_L g175 ( 
.A1(n_139),
.A2(n_11),
.B1(n_12),
.B2(n_14),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_175),
.A2(n_15),
.B1(n_17),
.B2(n_18),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_155),
.A2(n_14),
.B(n_15),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_176),
.A2(n_164),
.B(n_168),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_154),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_177),
.Y(n_190)
);

BUFx12_ASAP7_75t_L g178 ( 
.A(n_172),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_178),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_179),
.A2(n_187),
.B1(n_17),
.B2(n_20),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_165),
.A2(n_157),
.B1(n_155),
.B2(n_144),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_183),
.A2(n_167),
.B1(n_175),
.B2(n_174),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_184),
.B(n_185),
.Y(n_193)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_159),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_186),
.B(n_190),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_166),
.B(n_37),
.C(n_34),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_188),
.B(n_189),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_160),
.B(n_33),
.C(n_32),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_180),
.A2(n_165),
.B1(n_162),
.B2(n_169),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_191),
.A2(n_192),
.B1(n_194),
.B2(n_195),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_180),
.A2(n_175),
.B1(n_173),
.B2(n_19),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_182),
.A2(n_173),
.B1(n_18),
.B2(n_19),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_196),
.B(n_197),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_183),
.A2(n_28),
.B(n_20),
.Y(n_197)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_199),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_200),
.B(n_189),
.C(n_181),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_201),
.B(n_203),
.C(n_205),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_200),
.B(n_193),
.C(n_198),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_191),
.B(n_185),
.C(n_188),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_192),
.B(n_179),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_206),
.B(n_197),
.C(n_195),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_204),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_209),
.B(n_202),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_210),
.B(n_211),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_207),
.A2(n_196),
.B1(n_178),
.B2(n_23),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_213),
.B(n_202),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_214),
.B(n_212),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_215),
.B(n_208),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_216),
.B(n_178),
.C(n_22),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_217),
.B(n_21),
.C(n_22),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_218),
.B(n_21),
.C(n_24),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_219),
.B(n_24),
.Y(n_220)
);


endmodule